

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
         n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
         n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
         n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
         n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
         n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797,
         n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807,
         n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817,
         n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827,
         n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
         n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
         n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857,
         n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867,
         n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
         n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887,
         n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897,
         n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907,
         n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917,
         n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
         n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
         n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957,
         n6958, n6959;

  NOR2_X1 U3553 ( .A1(n5981), .A2(n3775), .ZN(n4713) );
  CLKBUF_X2 U3554 ( .A(n3776), .Z(n5189) );
  BUF_X2 U3555 ( .A(n3778), .Z(n3111) );
  AND2_X2 U3557 ( .A1(n3776), .A2(n3778), .ZN(n5273) );
  NAND2_X2 U3558 ( .A1(n4214), .A2(n4190), .ZN(n3778) );
  CLKBUF_X2 U3559 ( .A(n3353), .Z(n5109) );
  CLKBUF_X2 U3560 ( .A(n3275), .Z(n5135) );
  CLKBUF_X2 U3561 ( .A(n3303), .Z(n5129) );
  CLKBUF_X2 U3562 ( .A(n3302), .Z(n5110) );
  CLKBUF_X2 U3563 ( .A(n3313), .Z(n5137) );
  CLKBUF_X2 U3564 ( .A(n3351), .Z(n3311) );
  CLKBUF_X2 U3565 ( .A(n3352), .Z(n5136) );
  CLKBUF_X2 U3566 ( .A(n3276), .Z(n5075) );
  CLKBUF_X2 U3567 ( .A(n3312), .Z(n5112) );
  NOR2_X1 U3568 ( .A1(n6009), .A2(n4190), .ZN(n3256) );
  INV_X2 U3569 ( .A(n4190), .ZN(n4121) );
  CLKBUF_X2 U3570 ( .A(n3305), .Z(n5130) );
  CLKBUF_X2 U3571 ( .A(n3304), .Z(n5104) );
  AND2_X1 U3572 ( .A1(n3242), .A2(n5161), .ZN(n3195) );
  AND4_X1 U3573 ( .A1(n3145), .A2(n3144), .A3(n3143), .A4(n3142), .ZN(n3109)
         );
  NAND2_X2 U3574 ( .A1(n3109), .A2(n3110), .ZN(n4031) );
  INV_X1 U3575 ( .A(n5257), .ZN(n5731) );
  INV_X1 U3576 ( .A(n3778), .ZN(n5197) );
  INV_X1 U3577 ( .A(n5979), .ZN(n5967) );
  OR2_X1 U3578 ( .A1(n5195), .A2(n5192), .ZN(n5200) );
  NOR2_X1 U3579 ( .A1(n3255), .A2(n4214), .ZN(n4420) );
  INV_X2 U3580 ( .A(n5731), .ZN(n5822) );
  INV_X2 U3581 ( .A(n5731), .ZN(n5698) );
  OR3_X1 U3582 ( .A1(n3954), .A2(n6229), .A3(n3762), .ZN(n5934) );
  AND2_X1 U3583 ( .A1(n5934), .A2(n3857), .ZN(n5986) );
  OAI21_X1 U3584 ( .B1(n5343), .B2(n5342), .A(n5341), .ZN(n5347) );
  INV_X1 U3585 ( .A(n5986), .ZN(n5977) );
  NAND2_X2 U3586 ( .A1(n4875), .A2(n6111), .ZN(n5623) );
  AOI22_X1 U3587 ( .A1(n3353), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3179) );
  AOI21_X1 U3588 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n5565) );
  AND2_X1 U3589 ( .A1(n5429), .A2(n5428), .ZN(n5995) );
  OR2_X1 U3590 ( .A1(n4884), .A2(n5624), .ZN(n4907) );
  INV_X1 U3591 ( .A(n5731), .ZN(n5568) );
  NAND2_X1 U3592 ( .A1(n4653), .A2(n4652), .ZN(n5257) );
  XNOR2_X1 U3593 ( .A(n4537), .B(n3492), .ZN(n4527) );
  NOR2_X1 U3594 ( .A1(n5455), .A2(n4921), .ZN(n3834) );
  NAND2_X1 U3595 ( .A1(n4043), .A2(n4042), .ZN(n3391) );
  AOI222_X2 U3596 ( .A1(n4125), .A2(STATE2_REG_2__SCAN_IN), .B1(n4136), .B2(
        n6359), .C1(n6433), .C2(n6944), .ZN(n6952) );
  NAND2_X1 U3597 ( .A1(n3376), .A2(n3375), .ZN(n4043) );
  CLKBUF_X1 U3599 ( .A(n4047), .Z(n4767) );
  NAND2_X1 U3600 ( .A1(n3794), .A2(n3793), .ZN(n4428) );
  NOR2_X1 U3601 ( .A1(n4707), .A2(n4423), .ZN(n3793) );
  AND2_X1 U3602 ( .A1(n3788), .A2(n3787), .ZN(n4707) );
  NOR2_X1 U3603 ( .A1(n4187), .A2(n4169), .ZN(n3754) );
  OR2_X1 U3604 ( .A1(n4032), .A2(n5159), .ZN(n4199) );
  AND2_X1 U3605 ( .A1(n3234), .A2(n3237), .ZN(n3106) );
  NAND3_X1 U3606 ( .A1(n3197), .A2(n3196), .A3(n3195), .ZN(n3259) );
  NAND2_X1 U3607 ( .A1(n3942), .A2(n3253), .ZN(n4187) );
  INV_X1 U3608 ( .A(n3783), .ZN(n3912) );
  CLKBUF_X1 U3609 ( .A(n4030), .Z(n5383) );
  BUF_X2 U3610 ( .A(n3256), .Z(n4806) );
  INV_X1 U3611 ( .A(n5161), .ZN(n4030) );
  BUF_X2 U3612 ( .A(n3252), .Z(n4216) );
  OR2_X1 U3613 ( .A1(n3319), .A2(n3318), .ZN(n4655) );
  OR2_X2 U3614 ( .A1(n3194), .A2(n3193), .ZN(n5161) );
  BUF_X2 U3615 ( .A(n3230), .Z(n4349) );
  INV_X1 U3616 ( .A(n4031), .ZN(n3368) );
  OR2_X2 U3617 ( .A1(n3159), .A2(n3158), .ZN(n3225) );
  AND4_X1 U3618 ( .A1(n3149), .A2(n3148), .A3(n3147), .A4(n3146), .ZN(n3110)
         );
  INV_X2 U3619 ( .A(n5617), .ZN(n6137) );
  BUF_X2 U3620 ( .A(n3214), .Z(n5128) );
  INV_X2 U3621 ( .A(n3211), .ZN(n3310) );
  AND2_X2 U3622 ( .A1(n3129), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3987)
         );
  NAND2_X1 U3623 ( .A1(n6538), .A2(STATE_REG_1__SCAN_IN), .ZN(n6589) );
  AND2_X1 U3624 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3107) );
  AND2_X1 U3625 ( .A1(n4633), .A2(n5189), .ZN(n5981) );
  BUF_X2 U3626 ( .A(n3184), .Z(n3276) );
  NAND2_X1 U3627 ( .A1(n3235), .A2(n3106), .ZN(n3104) );
  AND2_X2 U3628 ( .A1(n3104), .A2(n3105), .ZN(n3284) );
  OR2_X1 U3629 ( .A1(n3236), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3105)
         );
  NAND3_X1 U3630 ( .A1(n5569), .A2(n3107), .A3(n5822), .ZN(n5560) );
  CLKBUF_X1 U3631 ( .A(n5260), .Z(n3108) );
  NAND2_X1 U3632 ( .A1(n3235), .A2(n3234), .ZN(n3338) );
  OR2_X4 U3633 ( .A1(n5488), .A2(n5173), .ZN(n5420) );
  AND2_X2 U3634 ( .A1(n6009), .A2(n4190), .ZN(n3776) );
  AOI211_X2 U3635 ( .C1(n5391), .C2(n5216), .A(n5215), .B(n5214), .ZN(n5217)
         );
  NAND2_X2 U3636 ( .A1(n3284), .A2(n3285), .ZN(n3337) );
  NOR2_X4 U3637 ( .A1(n4845), .A2(n4846), .ZN(n4844) );
  NAND2_X2 U3638 ( .A1(n5236), .A2(n5235), .ZN(n5539) );
  NOR2_X2 U3639 ( .A1(n4110), .A2(n4148), .ZN(n4147) );
  AND2_X4 U3640 ( .A1(n5059), .A2(n5491), .ZN(n5492) );
  NAND2_X2 U3641 ( .A1(n3283), .A2(n3117), .ZN(n3369) );
  AND2_X2 U3642 ( .A1(n3987), .A2(n4056), .ZN(n3346) );
  AND2_X4 U3643 ( .A1(n3987), .A2(n4050), .ZN(n3352) );
  XNOR2_X2 U3644 ( .A(n3371), .B(n3370), .ZN(n3372) );
  AND2_X2 U3645 ( .A1(n4055), .A2(n4009), .ZN(n4052) );
  AND2_X2 U3646 ( .A1(n3986), .A2(n4055), .ZN(n3303) );
  NAND2_X1 U3647 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  INV_X1 U3648 ( .A(n3778), .ZN(n3222) );
  NAND2_X1 U3649 ( .A1(n3459), .A2(n3458), .ZN(n3487) );
  INV_X1 U3650 ( .A(n3461), .ZN(n3458) );
  NAND2_X1 U3651 ( .A1(n4349), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4651) );
  NAND3_X1 U3652 ( .A1(n3225), .A2(n6009), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3732) );
  OR2_X1 U3653 ( .A1(n4249), .A2(n4189), .ZN(n4422) );
  OR2_X1 U3654 ( .A1(n5102), .A2(n5284), .ZN(n5127) );
  NAND2_X1 U3655 ( .A1(n4189), .A2(n4518), .ZN(n5750) );
  OR2_X1 U3656 ( .A1(n3715), .A2(n3719), .ZN(n3717) );
  AND2_X1 U3657 ( .A1(n3717), .A2(n3702), .ZN(n3710) );
  NAND2_X1 U3658 ( .A1(n3437), .A2(n3436), .ZN(n3446) );
  NAND2_X1 U3659 ( .A1(n3490), .A2(n3489), .ZN(n4537) );
  OR2_X1 U3660 ( .A1(n3400), .A2(n4121), .ZN(n3234) );
  OR2_X1 U3661 ( .A1(n3410), .A2(n3409), .ZN(n4229) );
  INV_X1 U3662 ( .A(n3732), .ZN(n3743) );
  AND2_X1 U3663 ( .A1(n5051), .A2(n5053), .ZN(n5099) );
  INV_X1 U3664 ( .A(n5091), .ZN(n5152) );
  INV_X1 U3665 ( .A(n3609), .ZN(n3623) );
  NOR2_X1 U3666 ( .A1(n3938), .A2(n3947), .ZN(n3971) );
  NAND2_X1 U3667 ( .A1(n4354), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3609) );
  NAND2_X1 U3668 ( .A1(n3171), .A2(n3170), .ZN(n4192) );
  AND4_X1 U3669 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3171)
         );
  NOR2_X1 U3670 ( .A1(n3169), .A2(n3168), .ZN(n3170) );
  OR2_X1 U3671 ( .A1(n6521), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4097) );
  INV_X1 U3672 ( .A(n4192), .ZN(n3252) );
  AOI21_X1 U3673 ( .B1(n6621), .B2(n6527), .A(n6605), .ZN(n4119) );
  NAND2_X1 U3674 ( .A1(n4250), .A2(n3946), .ZN(n4249) );
  INV_X1 U3675 ( .A(n5096), .ZN(n3766) );
  NAND2_X1 U3676 ( .A1(n3867), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3900)
         );
  NAND2_X1 U3677 ( .A1(n3493), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3510)
         );
  AND2_X1 U3678 ( .A1(n3811), .A2(n3810), .ZN(n4703) );
  NAND2_X1 U3679 ( .A1(n3382), .A2(n6765), .ZN(n3381) );
  NAND2_X1 U3681 ( .A1(n3753), .A2(n3752), .ZN(n4189) );
  OR3_X1 U3682 ( .A1(n4558), .A2(n6354), .A3(n5738), .ZN(n4141) );
  OR2_X1 U3683 ( .A1(n5755), .A2(n5213), .ZN(n5289) );
  AND2_X1 U3684 ( .A1(n5310), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3857) );
  CLKBUF_X1 U3685 ( .A(n4209), .Z(n5738) );
  NAND2_X1 U3686 ( .A1(n4037), .A2(n4214), .ZN(n3242) );
  NAND2_X1 U3687 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n4487), .ZN(n3719) );
  NAND2_X1 U3688 ( .A1(n3706), .A2(n3705), .ZN(n3711) );
  INV_X1 U3689 ( .A(n3310), .ZN(n3202) );
  OR2_X1 U3690 ( .A1(n3477), .A2(n3476), .ZN(n4541) );
  AOI22_X1 U3691 ( .A1(n3302), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3166) );
  OR2_X1 U3692 ( .A1(n3435), .A2(n3434), .ZN(n4242) );
  OR2_X1 U3693 ( .A1(n3282), .A2(n3281), .ZN(n4212) );
  INV_X1 U3694 ( .A(n4212), .ZN(n3325) );
  AOI22_X1 U3695 ( .A1(n3353), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U3696 ( .A1(n3267), .A2(n3119), .ZN(n3335) );
  INV_X1 U3697 ( .A(n4097), .ZN(n3340) );
  AND2_X2 U3698 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4049) );
  OR2_X1 U3699 ( .A1(n5219), .A2(n5125), .ZN(n5156) );
  AND2_X1 U3700 ( .A1(n5401), .A2(n5099), .ZN(n5218) );
  AND2_X1 U3701 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n3764), .ZN(n5013)
         );
  INV_X1 U3702 ( .A(n3900), .ZN(n3764) );
  NAND2_X1 U3703 ( .A1(n3661), .A2(n3660), .ZN(n3698) );
  INV_X1 U3704 ( .A(n5440), .ZN(n3661) );
  NAND2_X1 U3705 ( .A1(n3611), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3612)
         );
  INV_X1 U3706 ( .A(n3610), .ZN(n3611) );
  AND3_X1 U3707 ( .A1(n3945), .A2(n3996), .A3(n3994), .ZN(n4250) );
  INV_X1 U3708 ( .A(n6238), .ZN(n4549) );
  OR2_X1 U3709 ( .A1(n3300), .A2(n3299), .ZN(n4211) );
  NAND2_X1 U3710 ( .A1(n3287), .A2(n3286), .ZN(n3288) );
  AOI221_X1 U3711 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3738), .C1(
        n3984), .C2(n3738), .A(n3708), .ZN(n3758) );
  INV_X1 U3712 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3131) );
  AND2_X2 U3713 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4009) );
  AND2_X2 U3714 ( .A1(n3703), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4055)
         );
  OR2_X1 U3715 ( .A1(n4152), .A2(n3339), .ZN(n4291) );
  INV_X2 U3716 ( .A(n3225), .ZN(n3230) );
  INV_X1 U3717 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U3718 ( .A1(n3412), .A2(n3411), .ZN(n3415) );
  NAND2_X1 U3719 ( .A1(n4047), .A2(n6765), .ZN(n3412) );
  INV_X1 U3720 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U3721 ( .A1(n3958), .A2(n3933), .ZN(n3954) );
  BUF_X1 U3722 ( .A(n3760), .Z(n3966) );
  NOR2_X1 U3723 ( .A1(n3860), .A2(n5879), .ZN(n5435) );
  AND2_X1 U3724 ( .A1(n5050), .A2(n5049), .ZN(n5053) );
  AND2_X1 U3725 ( .A1(n3826), .A2(n3825), .ZN(n5521) );
  NAND2_X1 U3726 ( .A1(n4209), .A2(n3623), .ZN(n3376) );
  NAND2_X1 U3727 ( .A1(n3765), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5096)
         );
  INV_X1 U3728 ( .A(n5094), .ZN(n3765) );
  AND2_X1 U3729 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n4985), .ZN(n5045)
         );
  NAND2_X1 U3730 ( .A1(n5045), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5094)
         );
  NAND2_X1 U3731 ( .A1(n5015), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5021)
         );
  AND2_X1 U3732 ( .A1(n4998), .A2(n4997), .ZN(n5263) );
  NOR2_X1 U3733 ( .A1(n3763), .A2(n3690), .ZN(n3867) );
  AOI21_X1 U3734 ( .B1(n3885), .B2(n5148), .A(n3884), .ZN(n5491) );
  AND2_X1 U3735 ( .A1(n3676), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3677)
         );
  NAND2_X1 U3736 ( .A1(n3677), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3763)
         );
  AND2_X1 U3737 ( .A1(n3656), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3676)
         );
  NAND2_X1 U3738 ( .A1(n5517), .A2(n3594), .ZN(n4929) );
  NAND2_X1 U3739 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n3575), .ZN(n3610)
         );
  OR2_X1 U3740 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  NAND2_X1 U3741 ( .A1(n3593), .A2(n3592), .ZN(n5517) );
  INV_X1 U3742 ( .A(n5520), .ZN(n3592) );
  INV_X1 U3743 ( .A(n5519), .ZN(n3593) );
  NAND2_X1 U3744 ( .A1(n3556), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3557)
         );
  NOR2_X1 U3745 ( .A1(n6891), .A2(n3557), .ZN(n3575) );
  NOR2_X1 U3746 ( .A1(n3540), .A2(n3539), .ZN(n3556) );
  NAND2_X1 U3747 ( .A1(n3524), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3540)
         );
  AND2_X1 U3748 ( .A1(n3509), .A2(n3508), .ZN(n4484) );
  AOI21_X1 U3749 ( .B1(n4527), .B2(n3623), .A(n3496), .ZN(n4397) );
  NAND2_X1 U3750 ( .A1(n3486), .A2(n3485), .ZN(n4334) );
  INV_X1 U3751 ( .A(n3463), .ZN(n3464) );
  AND3_X1 U3752 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .ZN(n3440) );
  AND2_X1 U3753 ( .A1(n5667), .A2(n5331), .ZN(n5353) );
  NOR2_X2 U3754 ( .A1(n5420), .A2(n5182), .ZN(n5475) );
  NAND2_X1 U3755 ( .A1(n5548), .A2(n4939), .ZN(n5234) );
  INV_X1 U3756 ( .A(n5556), .ZN(n5558) );
  NAND2_X1 U3757 ( .A1(n5819), .A2(n4913), .ZN(n5821) );
  OR2_X1 U3758 ( .A1(n5822), .A2(n6914), .ZN(n5605) );
  NOR2_X1 U3759 ( .A1(n4890), .A2(n4889), .ZN(n5705) );
  OR2_X1 U3760 ( .A1(n5522), .A2(n5521), .ZN(n5524) );
  AND2_X1 U3761 ( .A1(n4885), .A2(n4907), .ZN(n5626) );
  NAND2_X1 U3762 ( .A1(n4857), .A2(n4856), .ZN(n5522) );
  NAND2_X1 U3763 ( .A1(n6245), .A2(n4892), .ZN(n5708) );
  NAND2_X1 U3764 ( .A1(n4870), .A2(n3113), .ZN(n6113) );
  NAND2_X1 U3765 ( .A1(n3813), .A2(n3812), .ZN(n4752) );
  INV_X1 U3766 ( .A(n4737), .ZN(n3813) );
  NAND2_X1 U3767 ( .A1(n4198), .A2(n4518), .ZN(n4258) );
  INV_X1 U3768 ( .A(n4711), .ZN(n3794) );
  BUF_X1 U3769 ( .A(n3382), .Z(n6436) );
  AND2_X1 U3771 ( .A1(n3639), .A2(n3638), .ZN(n3998) );
  NOR2_X2 U3772 ( .A1(n3131), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3986)
         );
  INV_X1 U3773 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3703) );
  INV_X1 U3774 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4058) );
  AND3_X1 U3775 ( .A1(n3979), .A2(n4422), .A3(n3978), .ZN(n4491) );
  AND2_X1 U3776 ( .A1(n4265), .A2(n6434), .ZN(n4270) );
  OR3_X1 U3777 ( .A1(n4558), .A2(n3415), .A3(n5738), .ZN(n4156) );
  NAND2_X1 U3778 ( .A1(n3399), .A2(n3398), .ZN(n6325) );
  INV_X1 U3779 ( .A(n4386), .ZN(n4380) );
  AND2_X1 U3780 ( .A1(n6257), .A2(n4767), .ZN(n6437) );
  INV_X1 U3781 ( .A(n6318), .ZN(n6353) );
  AND2_X1 U3782 ( .A1(n4558), .A2(n5738), .ZN(n6254) );
  BUF_X1 U3783 ( .A(n3368), .Z(n4354) );
  INV_X1 U3784 ( .A(n4214), .ZN(n4140) );
  INV_X1 U3785 ( .A(n4119), .ZN(n4120) );
  OR2_X1 U3786 ( .A1(n4558), .A2(n4264), .ZN(n6356) );
  OAI21_X1 U3787 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6397), .A(n4764), 
        .ZN(n6438) );
  OR2_X1 U3788 ( .A1(n4187), .A2(n6618), .ZN(n5747) );
  AND2_X1 U3789 ( .A1(n6708), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4515) );
  INV_X1 U3790 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6397) );
  INV_X1 U3791 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6765) );
  INV_X1 U3792 ( .A(n5753), .ZN(n5945) );
  AND2_X1 U3793 ( .A1(n4809), .A2(n3852), .ZN(n5969) );
  AND2_X1 U3794 ( .A1(n5934), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5952) );
  AND2_X1 U3795 ( .A1(n5980), .A2(n5189), .ZN(n5965) );
  INV_X1 U3796 ( .A(n5969), .ZN(n5994) );
  INV_X1 U3797 ( .A(n5952), .ZN(n5989) );
  AND2_X1 U3798 ( .A1(n4809), .A2(n3854), .ZN(n5979) );
  INV_X1 U3799 ( .A(n5965), .ZN(n5929) );
  INV_X1 U3800 ( .A(n5516), .ZN(n5480) );
  INV_X1 U3801 ( .A(n5565), .ZN(n5533) );
  INV_X1 U3802 ( .A(n5796), .ZN(n6003) );
  AND2_X1 U3803 ( .A1(n5382), .A2(n5160), .ZN(n6002) );
  AND2_X1 U3804 ( .A1(n5382), .A2(n5163), .ZN(n6006) );
  INV_X1 U3805 ( .A(n5535), .ZN(n4336) );
  INV_X1 U3806 ( .A(n6025), .ZN(n6029) );
  INV_X1 U3807 ( .A(n6057), .ZN(n6102) );
  OR2_X1 U3808 ( .A1(n5750), .A2(n5747), .ZN(n6108) );
  OR3_X1 U3809 ( .A1(n5750), .A2(READY_N), .A3(n4201), .ZN(n6104) );
  XNOR2_X1 U3810 ( .A(n3769), .B(n3768), .ZN(n5310) );
  INV_X1 U3811 ( .A(n6140), .ZN(n6117) );
  OR2_X1 U3812 ( .A1(n6130), .A2(n4603), .ZN(n6140) );
  OR2_X1 U3813 ( .A1(n6529), .A2(n6439), .ZN(n5617) );
  INV_X1 U3814 ( .A(n6121), .ZN(n6135) );
  XNOR2_X1 U3815 ( .A(n5305), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5360)
         );
  NAND2_X1 U3816 ( .A1(n3114), .A2(n5303), .ZN(n5304) );
  AND2_X1 U3817 ( .A1(n5661), .A2(n5330), .ZN(n5646) );
  CLKBUF_X1 U3818 ( .A(n5588), .Z(n5589) );
  NOR2_X1 U3819 ( .A1(n5851), .A2(n5326), .ZN(n6143) );
  NOR2_X1 U3820 ( .A1(n5705), .A2(n6143), .ZN(n5687) );
  OR2_X1 U3821 ( .A1(n4258), .A2(n5748), .ZN(n6245) );
  INV_X1 U3822 ( .A(n6207), .ZN(n6247) );
  INV_X1 U3823 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4487) );
  CLKBUF_X1 U3824 ( .A(n4010), .Z(n4011) );
  INV_X1 U3826 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6253) );
  INV_X1 U3827 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6708) );
  NAND2_X1 U3828 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4189), .ZN(n4521) );
  CLKBUF_X1 U3829 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n6699) );
  INV_X1 U3831 ( .A(n4521), .ZN(n6605) );
  INV_X1 U3832 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3984) );
  AND2_X1 U3833 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3396), .ZN(n6383)
         );
  NAND2_X1 U3834 ( .A1(n4142), .A2(n6318), .ZN(n6485) );
  NAND2_X1 U3835 ( .A1(n4515), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6520) );
  NOR2_X1 U3836 ( .A1(n6629), .A2(n5859), .ZN(n6599) );
  INV_X1 U3837 ( .A(n6589), .ZN(n6629) );
  INV_X1 U3838 ( .A(n3777), .ZN(n3783) );
  AND2_X2 U3839 ( .A1(n4049), .A2(n4009), .ZN(n3305) );
  NOR2_X1 U3840 ( .A1(n5822), .A2(n5315), .ZN(n3112) );
  NOR2_X1 U3841 ( .A1(n4869), .A2(n4868), .ZN(n3113) );
  AND2_X1 U3842 ( .A1(n5538), .A2(n5351), .ZN(n3114) );
  NAND2_X1 U3843 ( .A1(n5822), .A2(n5709), .ZN(n3115) );
  NAND2_X1 U3844 ( .A1(n4929), .A2(n4928), .ZN(n4927) );
  AND2_X1 U3845 ( .A1(n4018), .A2(n3245), .ZN(n3116) );
  OR2_X1 U3846 ( .A1(n4651), .A2(n3325), .ZN(n3117) );
  NAND2_X1 U3847 ( .A1(n4335), .A2(n4334), .ZN(n4333) );
  OR2_X1 U3848 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5155) );
  AND2_X1 U3849 ( .A1(n5591), .A2(n5986), .ZN(n3118) );
  AOI21_X1 U3850 ( .B1(n3395), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3342), 
        .ZN(n3343) );
  OR2_X1 U3851 ( .A1(n3266), .A2(n6699), .ZN(n3119) );
  INV_X1 U3852 ( .A(n3385), .ZN(n3881) );
  AND4_X1 U3853 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3120)
         );
  XNOR2_X1 U3854 ( .A(n3269), .B(n3268), .ZN(n3991) );
  OR2_X1 U3855 ( .A1(n5994), .A2(n3922), .ZN(n3121) );
  AND2_X2 U3856 ( .A1(n6121), .A2(n4098), .ZN(n6130) );
  INV_X1 U3857 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4225) );
  AND2_X1 U3858 ( .A1(n3210), .A2(n3209), .ZN(n3122) );
  AND3_X1 U3859 ( .A1(n3122), .A2(n3213), .A3(n3212), .ZN(n3123) );
  NAND2_X1 U3860 ( .A1(n3220), .A2(n3230), .ZN(n3721) );
  OR2_X1 U3861 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3124)
         );
  INV_X1 U3862 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5557) );
  AND2_X1 U3863 ( .A1(n4216), .A2(n4214), .ZN(n3125) );
  OR2_X1 U3864 ( .A1(n3721), .A2(n6009), .ZN(n3126) );
  NAND2_X1 U3865 ( .A1(n5382), .A2(n4040), .ZN(n5796) );
  AND3_X1 U3866 ( .A1(n3924), .A2(n3923), .A3(n3121), .ZN(n3127) );
  OR2_X1 U3867 ( .A1(n6402), .A2(n6401), .ZN(n3128) );
  NOR2_X2 U3868 ( .A1(n3698), .A2(n3697), .ZN(n5059) );
  INV_X1 U3869 ( .A(n3415), .ZN(n6354) );
  AND2_X2 U3870 ( .A1(n4009), .A2(n4050), .ZN(n3313) );
  AND2_X2 U3871 ( .A1(n3987), .A2(n4049), .ZN(n3302) );
  AND2_X1 U3872 ( .A1(n6606), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3245) );
  NOR2_X1 U3873 ( .A1(n4806), .A2(n3714), .ZN(n3731) );
  NOR2_X1 U3874 ( .A1(n3713), .A2(n3755), .ZN(n3737) );
  OR2_X1 U3875 ( .A1(n3243), .A2(n6618), .ZN(n3246) );
  INV_X1 U3876 ( .A(n3371), .ZN(n3330) );
  INV_X1 U3877 ( .A(n3710), .ZN(n3706) );
  AND2_X1 U3878 ( .A1(n3711), .A2(n3707), .ZN(n3742) );
  NOR2_X1 U3879 ( .A1(n3359), .A2(n3358), .ZN(n4204) );
  AND3_X1 U3880 ( .A1(n3247), .A2(n3246), .A3(n3116), .ZN(n3250) );
  NOR2_X1 U3881 ( .A1(n3742), .A2(n3741), .ZN(n3740) );
  INV_X1 U3882 ( .A(n4052), .ZN(n3289) );
  INV_X1 U3883 ( .A(n5506), .ZN(n3660) );
  AND2_X1 U3884 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  INV_X1 U3885 ( .A(n3337), .ZN(n3269) );
  NAND2_X1 U3886 ( .A1(n4169), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3400) );
  NOR2_X2 U3888 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4075) );
  AOI21_X1 U3889 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6320), .A(n3740), 
        .ZN(n3738) );
  OR2_X1 U3890 ( .A1(n5426), .A2(n3696), .ZN(n3697) );
  NOR2_X1 U3891 ( .A1(n3732), .A2(n4650), .ZN(n3745) );
  BUF_X1 U3892 ( .A(n4537), .Z(n4653) );
  AND2_X1 U3893 ( .A1(n5189), .A2(n5197), .ZN(n5176) );
  OR2_X1 U3894 ( .A1(n3457), .A2(n3456), .ZN(n4245) );
  OR2_X1 U3895 ( .A1(n6318), .A2(n4650), .ZN(n4094) );
  NAND2_X1 U3897 ( .A1(n3400), .A2(n4651), .ZN(n3750) );
  INV_X1 U3898 ( .A(n3966), .ZN(n3972) );
  NOR2_X1 U3899 ( .A1(n5021), .A2(n5422), .ZN(n4985) );
  INV_X1 U3900 ( .A(n5273), .ZN(n3833) );
  INV_X1 U3901 ( .A(n4703), .ZN(n3812) );
  INV_X1 U3902 ( .A(n3881), .ZN(n5149) );
  INV_X1 U3903 ( .A(n5024), .ZN(n5306) );
  NAND2_X1 U3904 ( .A1(n3766), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5102)
         );
  AND2_X1 U3905 ( .A1(n3998), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5091) );
  INV_X1 U3907 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3539) );
  AND2_X1 U3908 ( .A1(n3822), .A2(n3821), .ZN(n4856) );
  NAND2_X1 U3909 ( .A1(n4226), .A2(n4225), .ZN(n6123) );
  NAND2_X1 U3910 ( .A1(n3773), .A2(n3772), .ZN(n3775) );
  AND2_X1 U3911 ( .A1(n3337), .A2(n3288), .ZN(n3382) );
  XNOR2_X1 U3912 ( .A(n3394), .B(n6325), .ZN(n4047) );
  NAND2_X1 U3913 ( .A1(n3416), .A2(n3367), .ZN(n4208) );
  NOR2_X1 U3914 ( .A1(n4122), .A2(n6353), .ZN(n6947) );
  AND2_X1 U3915 ( .A1(n5013), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5015)
         );
  OAI21_X1 U3916 ( .B1(n5878), .B2(n6571), .A(n3861), .ZN(n3862) );
  INV_X1 U3917 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6891) );
  INV_X1 U3918 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4738) );
  AND2_X1 U3919 ( .A1(n3479), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3493)
         );
  AND2_X1 U3920 ( .A1(n5934), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4809) );
  NAND2_X1 U3921 ( .A1(n5200), .A2(n3111), .ZN(n5341) );
  AND2_X1 U3922 ( .A1(n5059), .A2(n5052), .ZN(n5054) );
  NAND2_X1 U3923 ( .A1(n3912), .A2(n3111), .ZN(n5345) );
  NOR2_X1 U3924 ( .A1(n3699), .A2(n5157), .ZN(n5308) );
  INV_X1 U3925 ( .A(n5263), .ZN(n5264) );
  NOR2_X1 U3926 ( .A1(n6758), .A2(n3612), .ZN(n3656) );
  NOR2_X1 U3927 ( .A1(n3510), .A2(n4738), .ZN(n3524) );
  AND2_X1 U3928 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3464), .ZN(n3479)
         );
  INV_X1 U3929 ( .A(n6130), .ZN(n5616) );
  AOI21_X1 U3930 ( .B1(n5588), .B2(n5586), .A(n5585), .ZN(n5700) );
  AND2_X1 U3931 ( .A1(n3839), .A2(n3838), .ZN(n5507) );
  CLKBUF_X1 U3932 ( .A(n4723), .Z(n4724) );
  NAND2_X1 U3933 ( .A1(n5708), .A2(n6231), .ZN(n5326) );
  OR2_X1 U3934 ( .A1(n4258), .A2(n4249), .ZN(n5711) );
  NOR2_X1 U3935 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4119), .ZN(n4764) );
  CLKBUF_X1 U3936 ( .A(n4009), .Z(n4020) );
  INV_X1 U3937 ( .A(n6313), .ZN(n4356) );
  OR2_X1 U3938 ( .A1(n4767), .A2(n6439), .ZN(n6400) );
  OR2_X1 U3939 ( .A1(n6434), .A2(n4377), .ZN(n4386) );
  AND2_X1 U3940 ( .A1(n4770), .A2(n6390), .ZN(n4800) );
  NAND2_X1 U3941 ( .A1(n6601), .A2(n4120), .ZN(n4355) );
  INV_X1 U3942 ( .A(n6947), .ZN(n4477) );
  NAND2_X1 U3943 ( .A1(n6397), .A2(n6442), .ZN(n6439) );
  OR2_X1 U3944 ( .A1(n6356), .A2(n4118), .ZN(n6950) );
  INV_X1 U3945 ( .A(n5155), .ZN(n5148) );
  NOR2_X1 U3946 ( .A1(n6439), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3955) );
  INV_X2 U3947 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6442) );
  AND2_X1 U3948 ( .A1(n5407), .A2(n5211), .ZN(n5391) );
  NOR2_X1 U3949 ( .A1(n3118), .A2(n3862), .ZN(n3863) );
  NOR2_X1 U3950 ( .A1(n5967), .A2(n3858), .ZN(n5893) );
  NOR2_X1 U3951 ( .A1(n5310), .A2(n6708), .ZN(n3770) );
  INV_X1 U3952 ( .A(n5971), .ZN(n5953) );
  NAND2_X1 U3953 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3440), .ZN(n3463)
         );
  OR2_X1 U3954 ( .A1(n5979), .A2(n5985), .ZN(n5395) );
  BUF_X1 U3955 ( .A(n5195), .Z(n5279) );
  NOR2_X1 U3956 ( .A1(n4752), .A2(n4751), .ZN(n4849) );
  NOR2_X1 U3957 ( .A1(n4428), .A2(n3800), .ZN(n4552) );
  INV_X1 U3958 ( .A(n5525), .ZN(n5479) );
  NAND2_X1 U3959 ( .A1(n5429), .A2(n3696), .ZN(n3700) );
  AND2_X1 U3960 ( .A1(n5382), .A2(n4041), .ZN(n5535) );
  INV_X1 U3961 ( .A(n6055), .ZN(n6045) );
  INV_X1 U3962 ( .A(n6108), .ZN(n6101) );
  OR2_X1 U3963 ( .A1(n4187), .A2(n5344), .ZN(n4201) );
  INV_X1 U3964 ( .A(n5501), .ZN(n5595) );
  NAND2_X1 U3965 ( .A1(n5364), .A2(n5304), .ZN(n5305) );
  INV_X1 U3966 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5313) );
  AND2_X1 U3967 ( .A1(n5677), .A2(n5317), .ZN(n5661) );
  AOI21_X1 U3968 ( .B1(n5822), .B2(n5684), .A(n5575), .ZN(n5569) );
  AND2_X1 U3969 ( .A1(n5433), .A2(n5432), .ZN(n5832) );
  INV_X1 U3970 ( .A(n5687), .ZN(n6155) );
  NAND2_X1 U3971 ( .A1(n4697), .A2(n4696), .ZN(n4867) );
  OR2_X1 U3972 ( .A1(n4898), .A2(n4251), .ZN(n6232) );
  INV_X1 U3973 ( .A(n6196), .ZN(n6240) );
  INV_X1 U3974 ( .A(n4764), .ZN(n4353) );
  AND2_X1 U3975 ( .A1(n4270), .A2(n6318), .ZN(n4447) );
  AND3_X1 U3976 ( .A1(n6254), .A2(n6434), .A3(n6318), .ZN(n6280) );
  NOR2_X1 U3977 ( .A1(n4156), .A2(n6353), .ZN(n6313) );
  OAI21_X1 U3978 ( .B1(n4160), .B2(n4159), .A(n4158), .ZN(n4360) );
  NOR2_X1 U3979 ( .A1(n4156), .A2(n6318), .ZN(n6349) );
  NAND2_X2 U3980 ( .A1(n3381), .A2(n3380), .ZN(n6318) );
  NOR2_X2 U3981 ( .A1(n4386), .A2(n6353), .ZN(n6426) );
  INV_X1 U3982 ( .A(n4625), .ZN(n4688) );
  INV_X1 U3983 ( .A(n6467), .ZN(n6475) );
  INV_X1 U3984 ( .A(n6520), .ZN(n4518) );
  INV_X1 U3985 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6538) );
  OR2_X1 U3986 ( .A1(n5750), .A2(n3948), .ZN(n3958) );
  AOI21_X1 U3987 ( .B1(n5803), .B2(n5945), .A(n5774), .ZN(n5777) );
  NAND2_X1 U3988 ( .A1(n5934), .A2(n3770), .ZN(n5753) );
  NAND2_X1 U3989 ( .A1(n5202), .A2(n5201), .ZN(n5376) );
  INV_X1 U3990 ( .A(n5995), .ZN(n5504) );
  NAND2_X1 U3991 ( .A1(n5525), .A2(n5383), .ZN(n5516) );
  OAI21_X1 U3992 ( .B1(n5402), .B2(n5401), .A(n5400), .ZN(n5542) );
  NAND2_X1 U3993 ( .A1(n3700), .A2(n3699), .ZN(n5501) );
  INV_X1 U3994 ( .A(n4662), .ZN(n4745) );
  INV_X1 U3995 ( .A(n6047), .ZN(n6039) );
  OR2_X1 U3996 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6527), .ZN(n6626) );
  OR3_X1 U3997 ( .A1(n5750), .A2(n5749), .A3(n6536), .ZN(n6055) );
  INV_X1 U3998 ( .A(n6106), .ZN(n6057) );
  OR2_X2 U3999 ( .A1(n5750), .A2(n4504), .ZN(n6121) );
  AOI211_X1 U4000 ( .C1(n5350), .C2(n6247), .A(n5349), .B(n5348), .ZN(n5359)
         );
  OR2_X1 U4001 ( .A1(n4258), .A2(n4257), .ZN(n6207) );
  OR2_X1 U4002 ( .A1(n4258), .A2(n4203), .ZN(n6196) );
  AND2_X1 U4003 ( .A1(n6244), .A2(n6249), .ZN(n6238) );
  INV_X1 U4004 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6320) );
  NOR2_X1 U4005 ( .A1(n6601), .A2(n3982), .ZN(n6609) );
  NOR2_X1 U4006 ( .A1(n4288), .A2(n4287), .ZN(n4451) );
  NAND2_X1 U4007 ( .A1(n4270), .A2(n6353), .ZN(n4595) );
  NOR2_X1 U4008 ( .A1(n4564), .A2(n4563), .ZN(n4600) );
  NAND3_X1 U4009 ( .A1(n6254), .A2(n6353), .A3(n6434), .ZN(n6317) );
  OR2_X1 U4010 ( .A1(n6356), .A2(n6355), .ZN(n6429) );
  NAND2_X1 U4011 ( .A1(n4380), .A2(n6353), .ZN(n4625) );
  NAND2_X1 U4012 ( .A1(n4760), .A2(n6254), .ZN(n6481) );
  AND2_X1 U4013 ( .A1(n4135), .A2(n4382), .ZN(n6518) );
  AND3_X1 U4014 ( .A1(n4315), .A2(n4624), .A3(n4314), .ZN(n4482) );
  CLKBUF_X1 U4015 ( .A(n6585), .Z(n6592) );
  OR2_X1 U4016 ( .A1(n3927), .A2(n3926), .ZN(U2806) );
  INV_X1 U4017 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3129) );
  INV_X1 U4018 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3130) );
  NOR2_X2 U4019 ( .A1(n3130), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4056)
         );
  AOI22_X1 U4020 ( .A1(n4052), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3135) );
  AND2_X2 U4021 ( .A1(n3986), .A2(n4056), .ZN(n3214) );
  AOI22_X1 U4022 ( .A1(n3214), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3134) );
  NOR2_X4 U4023 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4050) );
  AND2_X2 U4024 ( .A1(n4050), .A2(n4075), .ZN(n3304) );
  AOI22_X1 U4025 ( .A1(n3303), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3133) );
  AND2_X2 U4026 ( .A1(n3986), .A2(n4049), .ZN(n3270) );
  AOI22_X1 U4027 ( .A1(n3270), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3132) );
  NAND4_X1 U4028 ( .A1(n3135), .A2(n3134), .A3(n3133), .A4(n3132), .ZN(n3141)
         );
  AND2_X2 U4029 ( .A1(n4055), .A2(n4075), .ZN(n3351) );
  AOI22_X1 U4030 ( .A1(n3351), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3139) );
  AND2_X2 U4031 ( .A1(n4056), .A2(n4075), .ZN(n3275) );
  AND2_X2 U4032 ( .A1(n4056), .A2(n4009), .ZN(n3211) );
  AOI22_X1 U4033 ( .A1(n3275), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3211), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3138) );
  AND2_X2 U4034 ( .A1(n4055), .A2(n3987), .ZN(n3353) );
  AND2_X2 U4035 ( .A1(n4075), .A2(n4049), .ZN(n3184) );
  AOI22_X1 U4036 ( .A1(n3353), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3137) );
  AND2_X2 U4037 ( .A1(n3986), .A2(n4050), .ZN(n3312) );
  AOI22_X1 U4038 ( .A1(n3312), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3136) );
  NAND4_X1 U4039 ( .A1(n3139), .A2(n3138), .A3(n3137), .A4(n3136), .ZN(n3140)
         );
  OR2_X2 U4040 ( .A1(n3141), .A2(n3140), .ZN(n3173) );
  INV_X2 U4041 ( .A(n3173), .ZN(n5162) );
  AOI22_X1 U4042 ( .A1(n4052), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4043 ( .A1(n3214), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4044 ( .A1(n3303), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3143) );
  AOI22_X1 U4045 ( .A1(n3270), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4046 ( .A1(n3351), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4047 ( .A1(n3275), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3211), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3148) );
  AOI22_X1 U4048 ( .A1(n3312), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3146) );
  NAND2_X2 U4049 ( .A1(n5162), .A2(n4031), .ZN(n3226) );
  AOI22_X1 U4050 ( .A1(n4052), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U4051 ( .A1(n3214), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4052 ( .A1(n3303), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4053 ( .A1(n3270), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3150) );
  NAND4_X1 U4054 ( .A1(n3153), .A2(n3152), .A3(n3151), .A4(n3150), .ZN(n3159)
         );
  AOI22_X1 U4055 ( .A1(n3351), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3157) );
  AOI22_X1 U4056 ( .A1(n3275), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3211), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4057 ( .A1(n3353), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3155) );
  AOI22_X1 U4058 ( .A1(n3312), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3154) );
  NAND4_X1 U4059 ( .A1(n3157), .A2(n3156), .A3(n3155), .A4(n3154), .ZN(n3158)
         );
  NAND2_X2 U4060 ( .A1(n3226), .A2(n3230), .ZN(n3219) );
  AOI22_X1 U4061 ( .A1(n3214), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3163) );
  AOI22_X1 U4062 ( .A1(n3353), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4063 ( .A1(n3351), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3161) );
  AOI22_X1 U4064 ( .A1(n4052), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3160) );
  AOI22_X1 U4065 ( .A1(n3211), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3184), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4066 ( .A1(n3303), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4067 ( .A1(n3165), .A2(n3164), .ZN(n3169) );
  AOI22_X1 U4068 ( .A1(n3312), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4069 ( .A1(n3167), .A2(n3166), .ZN(n3168) );
  NAND2_X1 U4070 ( .A1(n3226), .A2(n3252), .ZN(n3172) );
  MUX2_X2 U4071 ( .A(n3219), .B(n3172), .S(n4031), .Z(n3197) );
  NAND2_X1 U4072 ( .A1(n3219), .A2(n4192), .ZN(n3196) );
  BUF_X2 U4073 ( .A(n3173), .Z(n3220) );
  NAND2_X2 U4074 ( .A1(n3220), .A2(n3368), .ZN(n4037) );
  AOI22_X1 U4075 ( .A1(n4052), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3177) );
  AOI22_X1 U4076 ( .A1(n3214), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4077 ( .A1(n3303), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4078 ( .A1(n3270), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3174) );
  NAND4_X1 U4079 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3183)
         );
  AOI22_X1 U4080 ( .A1(n3275), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3211), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4081 ( .A1(n3351), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4082 ( .A1(n3312), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3178) );
  NAND4_X1 U4083 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3182)
         );
  OR2_X2 U4084 ( .A1(n3183), .A2(n3182), .ZN(n4214) );
  AOI22_X1 U4085 ( .A1(n3275), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4086 ( .A1(n3351), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4087 ( .A1(n3353), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3186) );
  AOI22_X1 U4088 ( .A1(n3312), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3185) );
  NAND4_X1 U4089 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3194)
         );
  AOI22_X1 U4090 ( .A1(n4052), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4091 ( .A1(n3214), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4092 ( .A1(n3303), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3190) );
  AOI22_X1 U4093 ( .A1(n3270), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3189) );
  NAND4_X1 U4094 ( .A1(n3192), .A2(n3191), .A3(n3190), .A4(n3189), .ZN(n3193)
         );
  AOI22_X1 U4095 ( .A1(n4052), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4096 ( .A1(n3303), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4097 ( .A1(n3270), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4098 ( .A1(n3184), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3198) );
  NAND4_X1 U4099 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3208)
         );
  AOI22_X1 U4100 ( .A1(n3346), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3202), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4101 ( .A1(n3275), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4102 ( .A1(n3351), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4103 ( .A1(n3214), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U4104 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3207)
         );
  OR2_X4 U4105 ( .A1(n3208), .A2(n3207), .ZN(n6009) );
  AOI22_X1 U4106 ( .A1(n3312), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3313), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4107 ( .A1(n3351), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4108 ( .A1(n3275), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3211), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3213) );
  AOI22_X1 U4109 ( .A1(n3353), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3276), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4110 ( .A1(n4052), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3346), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4111 ( .A1(n3214), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3302), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U4112 ( .A1(n3303), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3216) );
  AOI22_X1 U4113 ( .A1(n3270), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3215) );
  NAND2_X4 U4114 ( .A1(n3123), .A2(n3120), .ZN(n4190) );
  NAND2_X1 U4115 ( .A1(n3259), .A2(n4806), .ZN(n3238) );
  NOR2_X2 U4116 ( .A1(n3219), .A2(n4030), .ZN(n3942) );
  NAND2_X2 U4117 ( .A1(n4121), .A2(n6009), .ZN(n6618) );
  INV_X1 U4118 ( .A(n3721), .ZN(n3221) );
  OAI21_X1 U4119 ( .B1(n3942), .B2(n6618), .A(n3223), .ZN(n3224) );
  INV_X1 U4120 ( .A(n3224), .ZN(n3251) );
  OAI211_X1 U4121 ( .C1(n4037), .C2(n3225), .A(n5161), .B(n3226), .ZN(n3227)
         );
  INV_X1 U4122 ( .A(n3227), .ZN(n3240) );
  NAND2_X1 U4123 ( .A1(n3240), .A2(n3125), .ZN(n3938) );
  NAND2_X1 U4124 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n3228) );
  OAI21_X1 U4125 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n3228), .ZN(n3848) );
  INV_X1 U4126 ( .A(n3848), .ZN(n3229) );
  NOR2_X1 U4127 ( .A1(n4190), .A2(n3229), .ZN(n3254) );
  INV_X1 U4128 ( .A(n4037), .ZN(n3639) );
  OR2_X2 U4129 ( .A1(n3639), .A2(n4349), .ZN(n3239) );
  OAI21_X1 U4130 ( .B1(n3254), .B2(n3220), .A(n3239), .ZN(n3231) );
  NOR2_X1 U4131 ( .A1(n3938), .A2(n3231), .ZN(n3232) );
  NAND3_X1 U4132 ( .A1(n3238), .A2(n3251), .A3(n3232), .ZN(n3233) );
  NAND2_X1 U4133 ( .A1(n3233), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3235) );
  INV_X4 U4134 ( .A(n6009), .ZN(n4169) );
  INV_X1 U4135 ( .A(n4515), .ZN(n3262) );
  NAND2_X1 U4136 ( .A1(n6708), .A2(n6397), .ZN(n6521) );
  MUX2_X1 U4137 ( .A(n3262), .B(n3340), .S(n4487), .Z(n3236) );
  INV_X1 U4138 ( .A(n3236), .ZN(n3237) );
  NAND3_X1 U4139 ( .A1(n3240), .A2(n4214), .A3(n3239), .ZN(n3241) );
  NAND2_X1 U4140 ( .A1(n3241), .A2(n4190), .ZN(n3247) );
  INV_X1 U4141 ( .A(n3242), .ZN(n3243) );
  NOR2_X1 U4142 ( .A1(n4031), .A2(n4214), .ZN(n3244) );
  AND2_X1 U4143 ( .A1(n3225), .A2(n5161), .ZN(n3638) );
  NAND4_X1 U4144 ( .A1(n4169), .A2(n3244), .A3(n3638), .A4(n4216), .ZN(n4018)
         );
  INV_X1 U4145 ( .A(n6521), .ZN(n6606) );
  MUX2_X1 U4146 ( .A(n3721), .B(n4192), .S(n6009), .Z(n3249) );
  INV_X1 U4147 ( .A(n4806), .ZN(n3248) );
  NAND2_X1 U4148 ( .A1(n3249), .A2(n3248), .ZN(n3939) );
  NAND4_X1 U4149 ( .A1(n3996), .A2(n3251), .A3(n3250), .A4(n3939), .ZN(n3285)
         );
  NAND2_X1 U4150 ( .A1(n3252), .A2(n5162), .ZN(n3255) );
  NOR2_X1 U4151 ( .A1(n3255), .A2(n4140), .ZN(n3253) );
  INV_X1 U4152 ( .A(n3254), .ZN(n3258) );
  NAND2_X1 U4153 ( .A1(n4420), .A2(n3256), .ZN(n4032) );
  NAND2_X1 U4154 ( .A1(n4031), .A2(n5161), .ZN(n5159) );
  INV_X1 U4155 ( .A(n4199), .ZN(n3257) );
  AOI21_X1 U4156 ( .B1(n3754), .B2(n3258), .A(n3257), .ZN(n3260) );
  NOR2_X2 U4157 ( .A1(n3259), .A2(n3126), .ZN(n3760) );
  NAND2_X2 U4158 ( .A1(n4121), .A2(n3760), .ZN(n3969) );
  NAND2_X1 U4159 ( .A1(n3260), .A2(n3969), .ZN(n3261) );
  NAND2_X1 U4160 ( .A1(n3261), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3264) );
  XNOR2_X1 U4161 ( .A(n4378), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6321)
         );
  AOI22_X1 U4162 ( .A1(n3340), .A2(n6321), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3262), .ZN(n3265) );
  NAND2_X1 U4163 ( .A1(n3338), .A2(n6699), .ZN(n3263) );
  NAND3_X1 U4164 ( .A1(n3264), .A2(n3265), .A3(n3263), .ZN(n3334) );
  INV_X1 U4165 ( .A(n3264), .ZN(n3267) );
  INV_X1 U4166 ( .A(n3265), .ZN(n3266) );
  NAND2_X1 U4167 ( .A1(n3334), .A2(n3335), .ZN(n3268) );
  NAND2_X1 U4168 ( .A1(n3991), .A2(n6765), .ZN(n3283) );
  INV_X2 U4169 ( .A(n3289), .ZN(n5111) );
  CLKBUF_X1 U4170 ( .A(n3346), .Z(n3294) );
  AOI22_X1 U4171 ( .A1(n5111), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4172 ( .A1(n5128), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4173 ( .A1(n5129), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3272) );
  INV_X1 U4174 ( .A(n3270), .ZN(n4057) );
  INV_X2 U4175 ( .A(n4057), .ZN(n5028) );
  AOI22_X1 U4176 ( .A1(n5028), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3271) );
  NAND4_X1 U4177 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3282)
         );
  INV_X1 U4178 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6691) );
  INV_X2 U4179 ( .A(n3310), .ZN(n5076) );
  AOI22_X1 U4180 ( .A1(n5135), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4181 ( .A1(n3311), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4182 ( .A1(n5109), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4183 ( .A1(n5112), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3277) );
  NAND4_X1 U4184 ( .A1(n3280), .A2(n3279), .A3(n3278), .A4(n3277), .ZN(n3281)
         );
  INV_X1 U4185 ( .A(n3284), .ZN(n3287) );
  INV_X1 U4186 ( .A(n3285), .ZN(n3286) );
  AOI22_X1 U4187 ( .A1(n5135), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4188 ( .A1(n5128), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4189 ( .A1(n5111), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4190 ( .A1(n5112), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3290) );
  NAND4_X1 U4191 ( .A1(n3293), .A2(n3292), .A3(n3291), .A4(n3290), .ZN(n3300)
         );
  AOI22_X1 U4192 ( .A1(n3294), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3353), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4193 ( .A1(n3311), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3352), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4194 ( .A1(n5129), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4195 ( .A1(n5028), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3295) );
  NAND4_X1 U4196 ( .A1(n3298), .A2(n3297), .A3(n3296), .A4(n3295), .ZN(n3299)
         );
  CLKBUF_X1 U4197 ( .A(n3346), .Z(n3301) );
  AOI22_X1 U4198 ( .A1(n5111), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4199 ( .A1(n3214), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4200 ( .A1(n5129), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4201 ( .A1(n5028), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3306) );
  NAND4_X1 U4202 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3319)
         );
  AOI22_X1 U4203 ( .A1(n5135), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4204 ( .A1(n3311), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4205 ( .A1(n3353), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4206 ( .A1(n5112), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U4207 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  XNOR2_X1 U4208 ( .A(n4211), .B(n4655), .ZN(n3320) );
  NOR2_X1 U4209 ( .A1(n3320), .A2(n4651), .ZN(n3377) );
  INV_X1 U4210 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6747) );
  AOI21_X1 U4211 ( .B1(n4349), .B2(n4655), .A(n6765), .ZN(n3322) );
  NAND2_X1 U4212 ( .A1(n4169), .A2(n4211), .ZN(n3321) );
  OAI211_X1 U4213 ( .C1(n3732), .C2(n6747), .A(n3322), .B(n3321), .ZN(n3379)
         );
  INV_X1 U4214 ( .A(n4651), .ZN(n3323) );
  AOI22_X1 U4215 ( .A1(n3377), .A2(n3379), .B1(n3323), .B2(n4655), .ZN(n3324)
         );
  NAND2_X2 U4216 ( .A1(n3381), .A2(n3324), .ZN(n3371) );
  NAND2_X1 U4217 ( .A1(n3369), .A2(n3371), .ZN(n3329) );
  INV_X1 U4218 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4301) );
  OR2_X1 U4219 ( .A1(n3400), .A2(n3325), .ZN(n3327) );
  OR2_X1 U4220 ( .A1(n4651), .A2(n4655), .ZN(n3326) );
  OAI211_X1 U4221 ( .C1(n4301), .C2(n3732), .A(n3327), .B(n3326), .ZN(n3370)
         );
  INV_X1 U4222 ( .A(n3370), .ZN(n3328) );
  NAND2_X1 U4223 ( .A1(n3329), .A2(n3328), .ZN(n3333) );
  INV_X1 U4224 ( .A(n3369), .ZN(n3331) );
  NAND2_X1 U4225 ( .A1(n3331), .A2(n3330), .ZN(n3332) );
  NAND2_X1 U4226 ( .A1(n3333), .A2(n3332), .ZN(n3365) );
  INV_X1 U4227 ( .A(n3365), .ZN(n3363) );
  INV_X1 U4228 ( .A(n3334), .ZN(n3336) );
  OAI21_X2 U4229 ( .B1(n3337), .B2(n3336), .A(n3335), .ZN(n3345) );
  AND2_X1 U4230 ( .A1(n4378), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4152)
         );
  NOR2_X1 U4231 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4378), .ZN(n4619)
         );
  NAND2_X1 U4232 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4619), .ZN(n6431) );
  OAI21_X1 U4233 ( .B1(n4495), .B2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n6431), 
        .ZN(n3339) );
  NAND2_X1 U4234 ( .A1(n3340), .A2(n4291), .ZN(n3341) );
  OAI21_X1 U4235 ( .B1(n4515), .B2(n4495), .A(n3341), .ZN(n3342) );
  INV_X1 U4236 ( .A(n3343), .ZN(n3344) );
  NAND2_X1 U4237 ( .A1(n3345), .A2(n3344), .ZN(n3394) );
  OAI21_X1 U4238 ( .B1(n3345), .B2(n3344), .A(n3394), .ZN(n4010) );
  AOI22_X1 U4239 ( .A1(n5111), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3350) );
  AOI22_X1 U4240 ( .A1(n5128), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3349) );
  INV_X1 U4241 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6855) );
  AOI22_X1 U4242 ( .A1(n5129), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4243 ( .A1(n5028), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3347) );
  NAND4_X1 U4244 ( .A1(n3350), .A2(n3349), .A3(n3348), .A4(n3347), .ZN(n3359)
         );
  AOI22_X1 U4245 ( .A1(n5135), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4246 ( .A1(n3311), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4247 ( .A1(n5109), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3355) );
  AOI22_X1 U4248 ( .A1(n5112), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3354) );
  NAND4_X1 U4249 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3358)
         );
  OAI22_X1 U4250 ( .A1(n4010), .A2(STATE2_REG_0__SCAN_IN), .B1(n4204), .B2(
        n4651), .ZN(n3362) );
  INV_X1 U4251 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4341) );
  OAI22_X1 U4252 ( .A1(n3400), .A2(n4204), .B1(n3732), .B2(n4341), .ZN(n3360)
         );
  INV_X1 U4253 ( .A(n3360), .ZN(n3361) );
  XNOR2_X1 U4254 ( .A(n3362), .B(n3361), .ZN(n3364) );
  NAND2_X1 U4255 ( .A1(n3363), .A2(n3364), .ZN(n3413) );
  BUF_X2 U4256 ( .A(n3413), .Z(n3416) );
  INV_X1 U4257 ( .A(n3364), .ZN(n3366) );
  NAND2_X1 U4258 ( .A1(n3366), .A2(n3365), .ZN(n3367) );
  NAND2_X1 U4259 ( .A1(n6442), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5024) );
  OAI21_X2 U4260 ( .B1(n4208), .B2(n3609), .A(n5024), .ZN(n4107) );
  XNOR2_X2 U4261 ( .A(n3369), .B(n3372), .ZN(n4209) );
  NOR2_X1 U4262 ( .A1(n5159), .A2(n6442), .ZN(n3438) );
  NAND2_X1 U4263 ( .A1(n3438), .A2(n6699), .ZN(n3374) );
  NOR2_X2 U4264 ( .A1(n5161), .A2(n6442), .ZN(n3385) );
  AOI22_X1 U4265 ( .A1(n3385), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6442), .ZN(n3373) );
  AND2_X1 U4266 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  INV_X1 U4267 ( .A(n3377), .ZN(n3378) );
  XNOR2_X1 U4268 ( .A(n3379), .B(n3378), .ZN(n3380) );
  AOI21_X1 U4269 ( .B1(n6318), .B2(n4354), .A(n6442), .ZN(n4039) );
  INV_X1 U4270 ( .A(n6436), .ZN(n4831) );
  AOI22_X1 U4271 ( .A1(n3385), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6442), .ZN(n3384) );
  NAND2_X1 U4272 ( .A1(n3438), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3383) );
  OAI211_X1 U4273 ( .C1(n4831), .C2(n3609), .A(n3384), .B(n3383), .ZN(n4038)
         );
  MUX2_X1 U4274 ( .A(n5148), .B(n4039), .S(n4038), .Z(n4042) );
  NAND2_X1 U4275 ( .A1(n3438), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3389) );
  INV_X1 U4276 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U4277 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3418) );
  OAI21_X1 U4278 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3418), .ZN(n6129) );
  NAND2_X1 U4279 ( .A1(n5148), .A2(n6129), .ZN(n3386) );
  OAI21_X1 U4280 ( .B1(n5024), .B2(n5460), .A(n3386), .ZN(n3387) );
  AOI21_X1 U4281 ( .B1(n3385), .B2(EAX_REG_2__SCAN_IN), .A(n3387), .ZN(n3388)
         );
  AND2_X1 U4282 ( .A1(n3389), .A2(n3388), .ZN(n4104) );
  NOR2_X1 U4283 ( .A1(n3391), .A2(n4104), .ZN(n3390) );
  OR2_X1 U4284 ( .A1(n4107), .A2(n3390), .ZN(n3393) );
  NAND2_X1 U4285 ( .A1(n3391), .A2(n4104), .ZN(n3392) );
  AND2_X2 U4286 ( .A1(n3393), .A2(n3392), .ZN(n4108) );
  NAND2_X1 U4287 ( .A1(n3395), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3399) );
  NAND3_X1 U4288 ( .A1(n6320), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6362) );
  INV_X1 U4289 ( .A(n6362), .ZN(n3396) );
  NAND3_X1 U4290 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4312) );
  INV_X1 U4291 ( .A(n4312), .ZN(n4125) );
  NAND2_X1 U4292 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4125), .ZN(n4180) );
  OAI21_X1 U4293 ( .B1(n6383), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n4180), 
        .ZN(n4761) );
  OAI22_X1 U4294 ( .A1(n4761), .A2(n4097), .B1(n4515), .B2(n6320), .ZN(n3397)
         );
  INV_X1 U4295 ( .A(n3397), .ZN(n3398) );
  AOI22_X1 U4296 ( .A1(n5111), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4297 ( .A1(n5128), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4298 ( .A1(n5129), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4299 ( .A1(n5028), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3401) );
  NAND4_X1 U4300 ( .A1(n3404), .A2(n3403), .A3(n3402), .A4(n3401), .ZN(n3410)
         );
  AOI22_X1 U4301 ( .A1(n5135), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3408) );
  AOI22_X1 U4302 ( .A1(n3311), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3407) );
  AOI22_X1 U4303 ( .A1(n5109), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4304 ( .A1(n5112), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3405) );
  NAND4_X1 U4305 ( .A1(n3408), .A2(n3407), .A3(n3406), .A4(n3405), .ZN(n3409)
         );
  AOI22_X1 U4306 ( .A1(n3750), .A2(n4229), .B1(n3743), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3411) );
  INV_X1 U4307 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4308 ( .A1(n3415), .A2(n3414), .ZN(n3445) );
  NAND2_X1 U4309 ( .A1(n3416), .A2(n6354), .ZN(n3417) );
  NAND2_X1 U4310 ( .A1(n3445), .A2(n3417), .ZN(n4231) );
  INV_X1 U4311 ( .A(n3438), .ZN(n3423) );
  INV_X1 U4312 ( .A(n3418), .ZN(n3420) );
  INV_X1 U4313 ( .A(n3440), .ZN(n3419) );
  OAI21_X1 U4314 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3420), .A(n3419), 
        .ZN(n4812) );
  AOI22_X1 U4315 ( .A1(n5148), .A2(n4812), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3422) );
  NAND2_X1 U4316 ( .A1(n5149), .A2(EAX_REG_3__SCAN_IN), .ZN(n3421) );
  OAI211_X1 U4317 ( .C1(n3423), .C2(n4058), .A(n3422), .B(n3421), .ZN(n3424)
         );
  INV_X1 U4318 ( .A(n3424), .ZN(n3425) );
  OAI21_X1 U4319 ( .B1(n4231), .B2(n3609), .A(n3425), .ZN(n4111) );
  NAND2_X1 U4320 ( .A1(n4108), .A2(n4111), .ZN(n4110) );
  AOI22_X1 U4321 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3301), .B1(n5111), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4322 ( .A1(n5128), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4323 ( .A1(n5129), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4324 ( .A1(n5028), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4325 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3435)
         );
  AOI22_X1 U4326 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5135), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4327 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3311), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4328 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5109), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4329 ( .A1(n5112), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3430) );
  NAND4_X1 U4330 ( .A1(n3433), .A2(n3432), .A3(n3431), .A4(n3430), .ZN(n3434)
         );
  NAND2_X1 U4331 ( .A1(n3750), .A2(n4242), .ZN(n3437) );
  NAND2_X1 U4332 ( .A1(n3743), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3436) );
  XNOR2_X1 U4333 ( .A(n3445), .B(n3446), .ZN(n4235) );
  NAND2_X1 U4334 ( .A1(n3438), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3443) );
  INV_X1 U4335 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6794) );
  AOI21_X1 U4336 ( .B1(n6794), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3439) );
  AOI21_X1 U4337 ( .B1(n5149), .B2(EAX_REG_4__SCAN_IN), .A(n3439), .ZN(n3442)
         );
  OAI21_X1 U4338 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3440), .A(n3463), 
        .ZN(n5978) );
  NOR2_X1 U4339 ( .A1(n5978), .A2(n5155), .ZN(n3441) );
  AOI21_X1 U4340 ( .B1(n3443), .B2(n3442), .A(n3441), .ZN(n3444) );
  AOI21_X1 U4341 ( .B1(n4235), .B2(n3623), .A(n3444), .ZN(n4148) );
  INV_X1 U4342 ( .A(n3445), .ZN(n3447) );
  NAND2_X1 U4343 ( .A1(n3447), .A2(n3446), .ZN(n3460) );
  INV_X1 U4344 ( .A(n3460), .ZN(n3459) );
  AOI22_X1 U4345 ( .A1(n5111), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4346 ( .A1(n5128), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4347 ( .A1(n5129), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4348 ( .A1(n5028), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4349 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4350 ( .A1(n5135), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4351 ( .A1(n3311), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4352 ( .A1(n5109), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4353 ( .A1(n5112), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4354 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  AOI22_X1 U4355 ( .A1(n3750), .A2(n4245), .B1(n3743), .B2(
        INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U4356 ( .A1(n3460), .A2(n3461), .ZN(n3462) );
  NAND2_X1 U4357 ( .A1(n3487), .A2(n3462), .ZN(n4248) );
  NOR2_X1 U4358 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3464), .ZN(n3465)
         );
  NOR2_X1 U4359 ( .A1(n3479), .A2(n3465), .ZN(n5956) );
  INV_X1 U4360 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4718) );
  OAI22_X1 U4361 ( .A1(n5956), .A2(n5155), .B1(n5024), .B2(n4718), .ZN(n3466)
         );
  AOI21_X1 U4362 ( .B1(n5149), .B2(EAX_REG_5__SCAN_IN), .A(n3466), .ZN(n3467)
         );
  OAI21_X1 U4363 ( .B1(n4248), .B2(n3609), .A(n3467), .ZN(n4282) );
  AND2_X2 U4364 ( .A1(n4147), .A2(n4282), .ZN(n4335) );
  AOI22_X1 U4365 ( .A1(n5111), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3471) );
  AOI22_X1 U4366 ( .A1(n5128), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3470) );
  AOI22_X1 U4367 ( .A1(n5129), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3469) );
  INV_X1 U4368 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U4369 ( .A1(n5028), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3468) );
  NAND4_X1 U4370 ( .A1(n3471), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3477)
         );
  AOI22_X1 U4371 ( .A1(n5135), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4372 ( .A1(n3311), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4373 ( .A1(n5109), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4374 ( .A1(n5112), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4375 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3476)
         );
  AOI22_X1 U4376 ( .A1(n3750), .A2(n4541), .B1(n3743), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U4377 ( .A1(n3487), .A2(n3488), .ZN(n4539) );
  NAND2_X1 U4378 ( .A1(n4539), .A2(n3623), .ZN(n3486) );
  INV_X1 U4379 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3478) );
  INV_X1 U4380 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4726) );
  OAI22_X1 U4381 ( .A1(n3881), .A2(n3478), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4726), .ZN(n3484) );
  INV_X1 U4382 ( .A(n3493), .ZN(n3482) );
  INV_X1 U4383 ( .A(n3479), .ZN(n3480) );
  NAND2_X1 U4384 ( .A1(n3480), .A2(n4726), .ZN(n3481) );
  NAND2_X1 U4385 ( .A1(n3482), .A2(n3481), .ZN(n5951) );
  AND2_X1 U4386 ( .A1(n5951), .A2(n5148), .ZN(n3483) );
  AOI21_X1 U4387 ( .B1(n3484), .B2(n5155), .A(n3483), .ZN(n3485) );
  INV_X1 U4388 ( .A(n3487), .ZN(n3490) );
  INV_X1 U4389 ( .A(n3488), .ZN(n3489) );
  INV_X1 U4390 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4310) );
  NAND2_X1 U4391 ( .A1(n3750), .A2(n4655), .ZN(n3491) );
  OAI21_X1 U4392 ( .B1(n4310), .B2(n3732), .A(n3491), .ZN(n3492) );
  INV_X1 U4393 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3495) );
  OAI21_X1 U4394 ( .B1(n3493), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3510), 
        .ZN(n5931) );
  AOI22_X1 U4395 ( .A1(n5931), .A2(n5148), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3494) );
  OAI21_X1 U4396 ( .B1(n3881), .B2(n3495), .A(n3494), .ZN(n3496) );
  OR2_X2 U4397 ( .A1(n4333), .A2(n4397), .ZN(n4483) );
  AOI22_X1 U4398 ( .A1(n5149), .A2(EAX_REG_8__SCAN_IN), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4399 ( .A1(n5128), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4400 ( .A1(n3301), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4401 ( .A1(n5112), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4402 ( .A1(n5028), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4403 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3506)
         );
  AOI22_X1 U4404 ( .A1(n5135), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4405 ( .A1(n5110), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4406 ( .A1(n5111), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4407 ( .A1(n5136), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4408 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3505)
         );
  OR2_X1 U4409 ( .A1(n3506), .A2(n3505), .ZN(n3507) );
  XNOR2_X1 U4410 ( .A(n3510), .B(n4738), .ZN(n4733) );
  AOI22_X1 U4411 ( .A1(n3623), .A2(n3507), .B1(n5148), .B2(n4733), .ZN(n3508)
         );
  NOR2_X2 U4412 ( .A1(n4483), .A2(n4484), .ZN(n4675) );
  XOR2_X1 U4413 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3524), .Z(n5923) );
  AOI22_X1 U4414 ( .A1(n3294), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4415 ( .A1(n5111), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5135), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4416 ( .A1(n3311), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4417 ( .A1(n5028), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4418 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3520)
         );
  AOI22_X1 U4419 ( .A1(n5128), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4420 ( .A1(n5109), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4421 ( .A1(n5076), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4422 ( .A1(n5112), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3515) );
  NAND4_X1 U4423 ( .A1(n3518), .A2(n3517), .A3(n3516), .A4(n3515), .ZN(n3519)
         );
  OR2_X1 U4424 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  AOI22_X1 U4425 ( .A1(n3623), .A2(n3521), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3523) );
  NAND2_X1 U4426 ( .A1(n3385), .A2(EAX_REG_9__SCAN_IN), .ZN(n3522) );
  OAI211_X1 U4427 ( .C1(n5923), .C2(n5155), .A(n3523), .B(n3522), .ZN(n4674)
         );
  NAND2_X1 U4428 ( .A1(n4675), .A2(n4674), .ZN(n4673) );
  XNOR2_X1 U4429 ( .A(n3540), .B(n3539), .ZN(n4824) );
  AOI22_X1 U4430 ( .A1(n3294), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4431 ( .A1(n3311), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4432 ( .A1(n5104), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3526) );
  AOI22_X1 U4433 ( .A1(n5112), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3525) );
  NAND4_X1 U4434 ( .A1(n3528), .A2(n3527), .A3(n3526), .A4(n3525), .ZN(n3534)
         );
  AOI22_X1 U4435 ( .A1(n5128), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3532) );
  AOI22_X1 U4436 ( .A1(n5111), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4437 ( .A1(n5129), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4438 ( .A1(n5135), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3529) );
  NAND4_X1 U4439 ( .A1(n3532), .A2(n3531), .A3(n3530), .A4(n3529), .ZN(n3533)
         );
  OAI21_X1 U4440 ( .B1(n3534), .B2(n3533), .A(n3623), .ZN(n3537) );
  NAND2_X1 U4441 ( .A1(n5149), .A2(EAX_REG_10__SCAN_IN), .ZN(n3536) );
  NAND2_X1 U4442 ( .A1(n5306), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3535)
         );
  NAND3_X1 U4443 ( .A1(n3537), .A2(n3536), .A3(n3535), .ZN(n3538) );
  AOI21_X1 U4444 ( .B1(n4824), .B2(n5148), .A(n3538), .ZN(n4747) );
  OR2_X2 U4445 ( .A1(n4673), .A2(n4747), .ZN(n4845) );
  XOR2_X1 U4446 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3556), .Z(n6116) );
  INV_X1 U4447 ( .A(n6116), .ZN(n3555) );
  AOI22_X1 U4448 ( .A1(n5135), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4449 ( .A1(n5129), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4450 ( .A1(n5104), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4451 ( .A1(n5136), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4452 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3550)
         );
  AOI22_X1 U4453 ( .A1(n5128), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4454 ( .A1(n5111), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3547) );
  AOI22_X1 U4455 ( .A1(n5112), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4456 ( .A1(n5028), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3545) );
  NAND4_X1 U4457 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3549)
         );
  OAI21_X1 U4458 ( .B1(n3550), .B2(n3549), .A(n3623), .ZN(n3553) );
  NAND2_X1 U4459 ( .A1(n5149), .A2(EAX_REG_11__SCAN_IN), .ZN(n3552) );
  NAND2_X1 U4460 ( .A1(n5306), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3551)
         );
  NAND3_X1 U4461 ( .A1(n3553), .A2(n3552), .A3(n3551), .ZN(n3554) );
  AOI21_X1 U4462 ( .B1(n3555), .B2(n5148), .A(n3554), .ZN(n4846) );
  NAND2_X1 U4463 ( .A1(n3557), .A2(n6891), .ZN(n3559) );
  INV_X1 U4464 ( .A(n3575), .ZN(n3558) );
  NAND2_X1 U4465 ( .A1(n3559), .A2(n3558), .ZN(n4879) );
  AOI22_X1 U4466 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3311), .B1(n5136), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4467 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n5110), .B1(n5104), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4468 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5076), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4469 ( .A1(n5028), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3560) );
  NAND4_X1 U4470 ( .A1(n3563), .A2(n3562), .A3(n3561), .A4(n3560), .ZN(n3569)
         );
  AOI22_X1 U4471 ( .A1(n5128), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4472 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5111), .B1(n3294), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4473 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5135), .B1(n5112), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4474 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5109), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3564) );
  NAND4_X1 U4475 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3568)
         );
  OAI21_X1 U4476 ( .B1(n3569), .B2(n3568), .A(n3623), .ZN(n3572) );
  NAND2_X1 U4477 ( .A1(n3385), .A2(EAX_REG_12__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4478 ( .A1(n5306), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3570)
         );
  NAND3_X1 U4479 ( .A1(n3572), .A2(n3571), .A3(n3570), .ZN(n3573) );
  AOI21_X1 U4480 ( .B1(n4879), .B2(n5148), .A(n3573), .ZN(n4854) );
  INV_X1 U4481 ( .A(n4854), .ZN(n3574) );
  AND2_X2 U4482 ( .A1(n4844), .A2(n3574), .ZN(n3579) );
  NAND2_X1 U4483 ( .A1(n5149), .A2(EAX_REG_13__SCAN_IN), .ZN(n3577) );
  OAI21_X1 U4484 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3575), .A(n3610), 
        .ZN(n5901) );
  AOI22_X1 U4485 ( .A1(n5148), .A2(n5901), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U4486 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  NAND2_X1 U4487 ( .A1(n3579), .A2(n3578), .ZN(n3594) );
  NAND2_X1 U4488 ( .A1(n3580), .A2(n3594), .ZN(n5519) );
  AOI22_X1 U4489 ( .A1(n5111), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4490 ( .A1(n5135), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5112), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4491 ( .A1(n5129), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4492 ( .A1(n5109), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3581) );
  NAND4_X1 U4493 ( .A1(n3584), .A2(n3583), .A3(n3582), .A4(n3581), .ZN(n3590)
         );
  AOI22_X1 U4494 ( .A1(n3311), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3588) );
  AOI22_X1 U4495 ( .A1(n5128), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3587) );
  AOI22_X1 U4496 ( .A1(n5076), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4497 ( .A1(n5028), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3585) );
  NAND4_X1 U4498 ( .A1(n3588), .A2(n3587), .A3(n3586), .A4(n3585), .ZN(n3589)
         );
  OR2_X1 U4499 ( .A1(n3590), .A2(n3589), .ZN(n3591) );
  NAND2_X1 U4500 ( .A1(n3623), .A2(n3591), .ZN(n5520) );
  AOI22_X1 U4501 ( .A1(n5129), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4502 ( .A1(n5111), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4503 ( .A1(n5112), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4504 ( .A1(n5135), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4505 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3604)
         );
  AOI22_X1 U4506 ( .A1(n5109), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4507 ( .A1(n5110), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4508 ( .A1(n5136), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4509 ( .A1(n5128), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3599) );
  NAND4_X1 U4510 ( .A1(n3602), .A2(n3601), .A3(n3600), .A4(n3599), .ZN(n3603)
         );
  NOR2_X1 U4511 ( .A1(n3604), .A2(n3603), .ZN(n3608) );
  XNOR2_X1 U4512 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3610), .ZN(n5890)
         );
  INV_X1 U4513 ( .A(n5890), .ZN(n3605) );
  AOI22_X1 U4514 ( .A1(n5306), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n5148), 
        .B2(n3605), .ZN(n3607) );
  NAND2_X1 U4515 ( .A1(n5149), .A2(EAX_REG_14__SCAN_IN), .ZN(n3606) );
  OAI211_X1 U4516 ( .C1(n3609), .C2(n3608), .A(n3607), .B(n3606), .ZN(n4928)
         );
  INV_X1 U4517 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6758) );
  NAND2_X1 U4518 ( .A1(n3612), .A2(n6758), .ZN(n3614) );
  INV_X1 U4519 ( .A(n3656), .ZN(n3613) );
  NAND2_X1 U4520 ( .A1(n3614), .A2(n3613), .ZN(n5451) );
  AOI22_X1 U4521 ( .A1(n5128), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4522 ( .A1(n5111), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4523 ( .A1(n5028), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3616) );
  AOI22_X1 U4524 ( .A1(n5135), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3615) );
  NAND4_X1 U4525 ( .A1(n3618), .A2(n3617), .A3(n3616), .A4(n3615), .ZN(n3625)
         );
  AOI22_X1 U4526 ( .A1(n5129), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3622) );
  AOI22_X1 U4527 ( .A1(n5076), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5112), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4528 ( .A1(n3311), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4529 ( .A1(n5104), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3619) );
  NAND4_X1 U4530 ( .A1(n3622), .A2(n3621), .A3(n3620), .A4(n3619), .ZN(n3624)
         );
  OAI21_X1 U4531 ( .B1(n3625), .B2(n3624), .A(n3623), .ZN(n3628) );
  NAND2_X1 U4532 ( .A1(n5149), .A2(EAX_REG_15__SCAN_IN), .ZN(n3627) );
  NAND2_X1 U4533 ( .A1(n5306), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3626)
         );
  NAND3_X1 U4534 ( .A1(n3628), .A2(n3627), .A3(n3626), .ZN(n3629) );
  AOI21_X1 U4535 ( .B1(n5451), .B2(n5148), .A(n3629), .ZN(n5449) );
  NOR2_X2 U4536 ( .A1(n4927), .A2(n5449), .ZN(n5439) );
  XNOR2_X1 U4537 ( .A(n5597), .B(n3656), .ZN(n5600) );
  AOI22_X1 U4538 ( .A1(n3385), .A2(EAX_REG_16__SCAN_IN), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4539 ( .A1(n5129), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4540 ( .A1(n3311), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3632) );
  AOI22_X1 U4541 ( .A1(n5111), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4542 ( .A1(n5112), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3630) );
  NAND4_X1 U4543 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3641)
         );
  AOI22_X1 U4544 ( .A1(n3301), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4545 ( .A1(n5135), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4546 ( .A1(n5128), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4547 ( .A1(n5110), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4548 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3640)
         );
  OAI21_X1 U4549 ( .B1(n3641), .B2(n3640), .A(n5091), .ZN(n3642) );
  OAI211_X1 U4550 ( .C1(n5600), .C2(n5155), .A(n3643), .B(n3642), .ZN(n5441)
         );
  NAND2_X1 U4551 ( .A1(n5439), .A2(n5441), .ZN(n5440) );
  AOI22_X1 U4552 ( .A1(n5128), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4553 ( .A1(n5111), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4554 ( .A1(n5112), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4555 ( .A1(n5109), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3644) );
  NAND4_X1 U4556 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3653)
         );
  AOI22_X1 U4557 ( .A1(n5135), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4558 ( .A1(n5129), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4559 ( .A1(n3311), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4560 ( .A1(n5110), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3648) );
  NAND4_X1 U4561 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3652)
         );
  NOR2_X1 U4562 ( .A1(n3653), .A2(n3652), .ZN(n3655) );
  AOI22_X1 U4563 ( .A1(n5149), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6442), .ZN(n3654) );
  OAI21_X1 U4564 ( .B1(n5152), .B2(n3655), .A(n3654), .ZN(n3659) );
  INV_X1 U4565 ( .A(n3676), .ZN(n3657) );
  XNOR2_X1 U4566 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .B(n3657), .ZN(n5881)
         );
  NOR2_X1 U4567 ( .A1(n5881), .A2(n5155), .ZN(n3658) );
  AOI21_X1 U4568 ( .B1(n3659), .B2(n5155), .A(n3658), .ZN(n5506) );
  AOI22_X1 U4569 ( .A1(n3294), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4570 ( .A1(n5135), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3664) );
  AOI22_X1 U4571 ( .A1(n5028), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4572 ( .A1(n5110), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3662) );
  NAND4_X1 U4573 ( .A1(n3665), .A2(n3664), .A3(n3663), .A4(n3662), .ZN(n3671)
         );
  AOI22_X1 U4574 ( .A1(n5128), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4575 ( .A1(n5112), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4576 ( .A1(n5111), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4577 ( .A1(n5076), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3666) );
  NAND4_X1 U4578 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3670)
         );
  NOR2_X1 U4579 ( .A1(n3671), .A2(n3670), .ZN(n3675) );
  NAND2_X1 U4580 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3672)
         );
  NAND2_X1 U4581 ( .A1(n5155), .A2(n3672), .ZN(n3673) );
  AOI21_X1 U4582 ( .B1(n5149), .B2(EAX_REG_18__SCAN_IN), .A(n3673), .ZN(n3674)
         );
  OAI21_X1 U4583 ( .B1(n5152), .B2(n3675), .A(n3674), .ZN(n3679) );
  OAI21_X1 U4584 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3677), .A(n3763), 
        .ZN(n5828) );
  OR2_X1 U4585 ( .A1(n5155), .A2(n5828), .ZN(n3678) );
  NAND2_X1 U4586 ( .A1(n3679), .A2(n3678), .ZN(n5426) );
  OR2_X1 U4587 ( .A1(n5427), .A2(n5426), .ZN(n5429) );
  AOI22_X1 U4588 ( .A1(n5111), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4589 ( .A1(n5128), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4590 ( .A1(n5129), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4591 ( .A1(n5028), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3680) );
  NAND4_X1 U4592 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3689)
         );
  AOI22_X1 U4593 ( .A1(n5135), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4594 ( .A1(n3351), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4595 ( .A1(n5109), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4596 ( .A1(n5112), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4597 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3688)
         );
  NOR2_X1 U4598 ( .A1(n3689), .A2(n3688), .ZN(n3693) );
  INV_X1 U4599 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3690) );
  AOI21_X1 U4600 ( .B1(n3690), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3691) );
  AOI21_X1 U4601 ( .B1(n5149), .B2(EAX_REG_19__SCAN_IN), .A(n3691), .ZN(n3692)
         );
  OAI21_X1 U4602 ( .B1(n5152), .B2(n3693), .A(n3692), .ZN(n3695) );
  XNOR2_X1 U4603 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n3763), .ZN(n5591)
         );
  NAND2_X1 U4604 ( .A1(n5591), .A2(n5148), .ZN(n3694) );
  NAND2_X1 U4605 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  INV_X1 U4606 ( .A(n5059), .ZN(n3699) );
  NAND2_X1 U4607 ( .A1(n4378), .A2(n6699), .ZN(n3702) );
  NAND2_X1 U4608 ( .A1(n3129), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4609 ( .A1(n3702), .A2(n3701), .ZN(n3715) );
  NAND2_X1 U4610 ( .A1(n4495), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4611 ( .A1(n4027), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3704) );
  NAND2_X1 U4612 ( .A1(n3707), .A2(n3704), .ZN(n3709) );
  INV_X1 U4613 ( .A(n3709), .ZN(n3705) );
  XNOR2_X1 U4614 ( .A(n4058), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3741)
         );
  NOR2_X1 U4615 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6253), .ZN(n3708)
         );
  NAND2_X1 U4616 ( .A1(n3220), .A2(n4190), .ZN(n4650) );
  NAND2_X1 U4617 ( .A1(n3758), .A2(n3745), .ZN(n3753) );
  INV_X1 U4618 ( .A(n3750), .ZN(n3713) );
  NAND2_X1 U4619 ( .A1(n3710), .A2(n3709), .ZN(n3712) );
  NAND2_X1 U4620 ( .A1(n3712), .A2(n3711), .ZN(n3755) );
  AND2_X1 U4621 ( .A1(n4121), .A2(n3220), .ZN(n3714) );
  INV_X1 U4622 ( .A(n3731), .ZN(n3736) );
  AOI21_X1 U4623 ( .B1(n3750), .B2(n4190), .A(n5162), .ZN(n3729) );
  NAND2_X1 U4624 ( .A1(n3715), .A2(n3719), .ZN(n3716) );
  NAND2_X1 U4625 ( .A1(n3717), .A2(n3716), .ZN(n3756) );
  INV_X1 U4626 ( .A(n3756), .ZN(n3718) );
  NAND2_X1 U4627 ( .A1(n3718), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3728) );
  INV_X1 U4628 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4007) );
  INV_X1 U4629 ( .A(n3719), .ZN(n3720) );
  AOI21_X1 U4630 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n4007), .A(n3720), 
        .ZN(n3724) );
  INV_X1 U4631 ( .A(n3724), .ZN(n3722) );
  OAI21_X1 U4632 ( .B1(n3221), .B2(n3722), .A(n6009), .ZN(n3723) );
  AOI22_X1 U4633 ( .A1(n3731), .A2(n3723), .B1(n3729), .B2(n3728), .ZN(n3725)
         );
  NAND3_X1 U4634 ( .A1(n3724), .A2(n3725), .A3(n3750), .ZN(n3727) );
  OAI21_X1 U4635 ( .B1(n3725), .B2(n3756), .A(n3745), .ZN(n3726) );
  OAI211_X1 U4636 ( .C1(n3729), .C2(n3728), .A(n3727), .B(n3726), .ZN(n3735)
         );
  INV_X1 U4637 ( .A(n3755), .ZN(n3733) );
  INV_X1 U4638 ( .A(n3737), .ZN(n3730) );
  OAI211_X1 U4639 ( .C1(n3733), .C2(n3732), .A(n3731), .B(n3730), .ZN(n3734)
         );
  AOI22_X1 U4640 ( .A1(n3737), .A2(n3736), .B1(n3735), .B2(n3734), .ZN(n3748)
         );
  AND3_X1 U4641 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3738), .A3(n3984), 
        .ZN(n3739) );
  AOI211_X1 U4642 ( .C1(n3742), .C2(n3741), .A(n3740), .B(n3739), .ZN(n3744)
         );
  NOR2_X1 U4643 ( .A1(n3743), .A2(n3744), .ZN(n3747) );
  INV_X1 U4644 ( .A(n3744), .ZN(n3757) );
  AOI22_X1 U4645 ( .A1(n3745), .A2(n3757), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6765), .ZN(n3746) );
  OAI21_X1 U4646 ( .B1(n3748), .B2(n3747), .A(n3746), .ZN(n3749) );
  AOI21_X1 U4647 ( .B1(n3750), .B2(n3758), .A(n3749), .ZN(n3751) );
  INV_X1 U4648 ( .A(n3751), .ZN(n3752) );
  INV_X1 U4649 ( .A(n3754), .ZN(n3948) );
  NOR3_X1 U4650 ( .A1(n3757), .A2(n3756), .A3(n3755), .ZN(n3759) );
  NOR2_X1 U4651 ( .A1(n3759), .A2(n3758), .ZN(n3970) );
  NOR2_X1 U4652 ( .A1(n3972), .A2(n6520), .ZN(n3761) );
  NAND2_X1 U4653 ( .A1(n3970), .A2(n3761), .ZN(n3933) );
  AND2_X2 U4654 ( .A1(n3955), .A2(n6765), .ZN(n6229) );
  AND2_X1 U4655 ( .A1(n6765), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4090) );
  AND2_X1 U4656 ( .A1(n4090), .A2(n5148), .ZN(n6522) );
  NAND2_X1 U4657 ( .A1(n6442), .A2(n6708), .ZN(n6621) );
  NOR3_X1 U4658 ( .A1(n6765), .A2(n6397), .A3(n6621), .ZN(n4517) );
  OR2_X1 U4659 ( .A1(n6522), .A2(n4517), .ZN(n3762) );
  INV_X1 U4660 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5422) );
  INV_X1 U4661 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5284) );
  INV_X1 U4662 ( .A(n5127), .ZN(n3767) );
  NAND2_X1 U4663 ( .A1(n3767), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n3769)
         );
  INV_X1 U4664 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n3768) );
  NAND2_X1 U4665 ( .A1(n4809), .A2(EBX_REG_31__SCAN_IN), .ZN(n5387) );
  NOR2_X1 U4666 ( .A1(STATEBS16_REG_SCAN_IN), .A2(READY_N), .ZN(n3853) );
  NOR2_X1 U4667 ( .A1(n5387), .A2(n3853), .ZN(n5980) );
  INV_X1 U4668 ( .A(EBX_REG_1__SCAN_IN), .ZN(n6878) );
  NAND2_X1 U4669 ( .A1(n5273), .A2(n6878), .ZN(n3773) );
  INV_X2 U4670 ( .A(n3776), .ZN(n5344) );
  NAND2_X1 U4671 ( .A1(n4140), .A2(n6009), .ZN(n3777) );
  NAND2_X1 U4672 ( .A1(n3778), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3771)
         );
  OAI211_X1 U4673 ( .C1(n5344), .C2(EBX_REG_1__SCAN_IN), .A(n3777), .B(n3771), 
        .ZN(n3772) );
  INV_X1 U4674 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3774) );
  OAI22_X1 U4675 ( .A1(n3777), .A2(n3774), .B1(n3778), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4743) );
  XNOR2_X1 U4676 ( .A(n3775), .B(n4743), .ZN(n4633) );
  INV_X1 U4677 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U4678 ( .A1(n5273), .A2(n5461), .ZN(n3782) );
  NAND2_X1 U4679 ( .A1(n5189), .A2(n5461), .ZN(n3780) );
  NAND2_X1 U4680 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3779)
         );
  NAND3_X1 U4681 ( .A1(n3780), .A2(n3912), .A3(n3779), .ZN(n3781) );
  AND2_X1 U4682 ( .A1(n3782), .A2(n3781), .ZN(n4712) );
  NAND2_X1 U4683 ( .A1(n4713), .A2(n4712), .ZN(n4711) );
  INV_X1 U4684 ( .A(EBX_REG_3__SCAN_IN), .ZN(n3784) );
  NAND2_X1 U4685 ( .A1(n5176), .A2(n3784), .ZN(n3788) );
  INV_X1 U4686 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U4687 ( .A1(n3912), .A2(n6215), .ZN(n3786) );
  NAND2_X1 U4688 ( .A1(n5189), .A2(n3784), .ZN(n3785) );
  NAND3_X1 U4689 ( .A1(n3786), .A2(n3778), .A3(n3785), .ZN(n3787) );
  INV_X1 U4690 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U4691 ( .A1(n5273), .A2(n4426), .ZN(n3792) );
  NAND2_X1 U4692 ( .A1(n5189), .A2(n4426), .ZN(n3790) );
  NAND2_X1 U4693 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3789)
         );
  NAND3_X1 U4694 ( .A1(n3790), .A2(n3912), .A3(n3789), .ZN(n3791) );
  NAND2_X1 U4695 ( .A1(n3792), .A2(n3791), .ZN(n4423) );
  MUX2_X1 U4696 ( .A(n5273), .B(n5197), .S(EBX_REG_6__SCAN_IN), .Z(n3796) );
  NOR2_X1 U4697 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3795)
         );
  NOR2_X1 U4698 ( .A1(n3796), .A2(n3795), .ZN(n4429) );
  NAND2_X1 U4699 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3797)
         );
  NAND2_X1 U4700 ( .A1(n3912), .A2(n3797), .ZN(n3799) );
  INV_X1 U4701 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4716) );
  NAND2_X1 U4702 ( .A1(n5189), .A2(n4716), .ZN(n3798) );
  MUX2_X1 U4703 ( .A(n5197), .B(n3799), .S(n3798), .Z(n4430) );
  NAND2_X1 U4704 ( .A1(n4429), .A2(n4430), .ZN(n3800) );
  INV_X1 U4705 ( .A(EBX_REG_7__SCAN_IN), .ZN(n6732) );
  NAND2_X1 U4706 ( .A1(n5176), .A2(n6732), .ZN(n3804) );
  INV_X1 U4707 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U4708 ( .A1(n3912), .A2(n4699), .ZN(n3802) );
  NAND2_X1 U4709 ( .A1(n5189), .A2(n6732), .ZN(n3801) );
  NAND3_X1 U4710 ( .A1(n3802), .A2(n3111), .A3(n3801), .ZN(n3803) );
  NAND2_X1 U4711 ( .A1(n3804), .A2(n3803), .ZN(n4551) );
  AND2_X2 U4712 ( .A1(n4552), .A2(n4551), .ZN(n4735) );
  MUX2_X1 U4713 ( .A(n3833), .B(n3111), .S(EBX_REG_8__SCAN_IN), .Z(n3805) );
  INV_X1 U4714 ( .A(n3805), .ZN(n3807) );
  NOR2_X1 U4715 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3806)
         );
  NOR2_X1 U4716 ( .A1(n3807), .A2(n3806), .ZN(n4734) );
  NAND2_X1 U4717 ( .A1(n4735), .A2(n4734), .ZN(n4737) );
  INV_X1 U4718 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U4719 ( .A1(n5176), .A2(n6707), .ZN(n3811) );
  INV_X1 U4720 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U4721 ( .A1(n3912), .A2(n6161), .ZN(n3809) );
  NAND2_X1 U4722 ( .A1(n5189), .A2(n6707), .ZN(n3808) );
  NAND3_X1 U4723 ( .A1(n3809), .A2(n3111), .A3(n3808), .ZN(n3810) );
  MUX2_X1 U4724 ( .A(n3833), .B(n3111), .S(EBX_REG_10__SCAN_IN), .Z(n3814) );
  OAI21_X1 U4725 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5345), .A(n3814), 
        .ZN(n4751) );
  INV_X1 U4726 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6787) );
  NAND2_X1 U4727 ( .A1(n5176), .A2(n6787), .ZN(n3818) );
  INV_X1 U4728 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U4729 ( .A1(n3912), .A2(n6156), .ZN(n3816) );
  NAND2_X1 U4730 ( .A1(n5189), .A2(n6787), .ZN(n3815) );
  NAND3_X1 U4731 ( .A1(n3816), .A2(n3111), .A3(n3815), .ZN(n3817) );
  NAND2_X1 U4732 ( .A1(n3818), .A2(n3817), .ZN(n4848) );
  AND2_X2 U4733 ( .A1(n4849), .A2(n4848), .ZN(n4857) );
  INV_X1 U4734 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3819) );
  NAND2_X1 U4735 ( .A1(n5273), .A2(n3819), .ZN(n3822) );
  NAND2_X1 U4736 ( .A1(n3778), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3820) );
  OAI211_X1 U4737 ( .C1(n5344), .C2(EBX_REG_12__SCAN_IN), .A(n3912), .B(n3820), 
        .ZN(n3821) );
  INV_X1 U4738 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U4739 ( .A1(n5176), .A2(n5899), .ZN(n3826) );
  INV_X1 U4740 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U4741 ( .A1(n3912), .A2(n4894), .ZN(n3824) );
  NAND2_X1 U4742 ( .A1(n5189), .A2(n5899), .ZN(n3823) );
  NAND3_X1 U4743 ( .A1(n3824), .A2(n3111), .A3(n3823), .ZN(n3825) );
  MUX2_X1 U4744 ( .A(n3833), .B(n3111), .S(EBX_REG_14__SCAN_IN), .Z(n3827) );
  NAND2_X1 U4745 ( .A1(n3827), .A2(n3124), .ZN(n4888) );
  NOR2_X2 U4746 ( .A1(n5524), .A2(n4888), .ZN(n5453) );
  NAND2_X1 U4747 ( .A1(n5345), .A2(EBX_REG_15__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4748 ( .A1(n5344), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3828) );
  NAND2_X1 U4749 ( .A1(n3829), .A2(n3828), .ZN(n3830) );
  XNOR2_X1 U4750 ( .A(n3830), .B(n3111), .ZN(n5452) );
  NAND2_X1 U4751 ( .A1(n5453), .A2(n5452), .ZN(n5455) );
  NAND2_X1 U4752 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3831) );
  OAI211_X1 U4753 ( .C1(n5344), .C2(EBX_REG_16__SCAN_IN), .A(n3912), .B(n3831), 
        .ZN(n3832) );
  OAI21_X1 U4754 ( .B1(n3833), .B2(EBX_REG_16__SCAN_IN), .A(n3832), .ZN(n4921)
         );
  INV_X1 U4755 ( .A(n3834), .ZN(n5508) );
  INV_X1 U4756 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U4757 ( .A1(n5176), .A2(n5883), .ZN(n3839) );
  INV_X1 U4758 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5820) );
  NAND2_X1 U4759 ( .A1(n3912), .A2(n5820), .ZN(n3837) );
  NAND2_X1 U4760 ( .A1(n5189), .A2(n5883), .ZN(n3835) );
  NAND3_X1 U4761 ( .A1(n3837), .A2(n3778), .A3(n3835), .ZN(n3838) );
  OR2_X2 U4762 ( .A1(n5508), .A2(n5507), .ZN(n5510) );
  INV_X1 U4763 ( .A(n5510), .ZN(n3843) );
  NAND2_X1 U4764 ( .A1(n5345), .A2(EBX_REG_18__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4765 ( .A1(n5344), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3840) );
  NAND2_X1 U4766 ( .A1(n3841), .A2(n3840), .ZN(n5494) );
  OR2_X1 U4767 ( .A1(n5494), .A2(n5197), .ZN(n3907) );
  NAND2_X1 U4768 ( .A1(n5494), .A2(n5197), .ZN(n3842) );
  AND2_X1 U4769 ( .A1(n3907), .A2(n3842), .ZN(n5430) );
  NAND2_X1 U4770 ( .A1(n3843), .A2(n5430), .ZN(n5433) );
  INV_X1 U4771 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6875) );
  NAND2_X1 U4772 ( .A1(n5273), .A2(n6875), .ZN(n3847) );
  NAND2_X1 U4773 ( .A1(n5189), .A2(n6875), .ZN(n3845) );
  NAND2_X1 U4774 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3844) );
  NAND3_X1 U4775 ( .A1(n3845), .A2(n3912), .A3(n3844), .ZN(n3846) );
  NAND2_X1 U4776 ( .A1(n3847), .A2(n3846), .ZN(n3903) );
  XNOR2_X1 U4777 ( .A(n5433), .B(n3903), .ZN(n5724) );
  OAI22_X1 U4778 ( .A1(n5501), .A2(n5753), .B1(n5929), .B2(n5724), .ZN(n3866)
         );
  OR2_X1 U4779 ( .A1(n3848), .A2(STATE_REG_0__SCAN_IN), .ZN(n6536) );
  INV_X1 U4780 ( .A(n3853), .ZN(n3849) );
  NOR2_X1 U4781 ( .A1(n6536), .A2(n3849), .ZN(n4513) );
  NOR2_X1 U4782 ( .A1(n6618), .A2(n4513), .ZN(n5388) );
  NOR2_X1 U4783 ( .A1(EBX_REG_31__SCAN_IN), .A2(n3853), .ZN(n3850) );
  AND2_X1 U4784 ( .A1(n6009), .A2(n3850), .ZN(n3851) );
  OR2_X1 U4785 ( .A1(n5388), .A2(n3851), .ZN(n3852) );
  NAND2_X1 U4786 ( .A1(n3955), .A2(n5934), .ZN(n5971) );
  NAND3_X1 U4787 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4788 ( .A1(n4121), .A2(n6536), .ZN(n4185) );
  AND3_X1 U4789 ( .A1(n4185), .A2(n3853), .A3(n6009), .ZN(n3854) );
  INV_X1 U4790 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6560) );
  INV_X1 U4791 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6556) );
  INV_X1 U4792 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6728) );
  INV_X1 U4793 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6552) );
  NAND3_X1 U4794 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5966) );
  NOR2_X1 U4795 ( .A1(n6552), .A2(n5966), .ZN(n5959) );
  NAND2_X1 U4796 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5959), .ZN(n5936) );
  NOR2_X1 U4797 ( .A1(n6728), .A2(n5936), .ZN(n5937) );
  NAND2_X1 U4798 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5937), .ZN(n4731) );
  NOR2_X1 U4799 ( .A1(n6556), .A2(n4731), .ZN(n5919) );
  NAND3_X1 U4800 ( .A1(n5919), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .ZN(n5912) );
  NOR2_X1 U4801 ( .A1(n6560), .A2(n5912), .ZN(n5910) );
  NAND3_X1 U4802 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n5910), .ZN(n3858) );
  NAND2_X1 U4803 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5893), .ZN(n5879) );
  NAND2_X1 U4804 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5790) );
  OAI211_X1 U4805 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5435), .B(n5790), .ZN(n3855) );
  OAI211_X1 U4806 ( .C1(n5994), .C2(n6875), .A(n5971), .B(n3855), .ZN(n3856)
         );
  INV_X1 U4807 ( .A(n3856), .ZN(n3864) );
  INV_X1 U4808 ( .A(n3858), .ZN(n3859) );
  OAI221_X1 U4809 ( .B1(n5967), .B2(REIP_REG_14__SCAN_IN), .C1(n5967), .C2(
        n3859), .A(n5934), .ZN(n5892) );
  AOI21_X1 U4810 ( .B1(n5979), .B2(n3860), .A(n5892), .ZN(n5878) );
  INV_X1 U4811 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U4812 ( .A1(n5952), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3861)
         );
  NAND2_X1 U4813 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  OR2_X1 U4814 ( .A1(n3866), .A2(n3865), .ZN(U2808) );
  OR2_X1 U4815 ( .A1(n3867), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3868)
         );
  NAND2_X1 U4816 ( .A1(n3868), .A2(n3900), .ZN(n5817) );
  INV_X1 U4817 ( .A(n5817), .ZN(n3885) );
  AOI22_X1 U4818 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5129), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4819 ( .A1(n5128), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4820 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n5109), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4821 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3311), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3869) );
  NAND4_X1 U4822 ( .A1(n3872), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3878)
         );
  AOI22_X1 U4823 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n5076), .B1(n5135), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4824 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5112), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4825 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5111), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4826 ( .A1(n5028), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4827 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3877)
         );
  OR2_X1 U4828 ( .A1(n3878), .A2(n3877), .ZN(n3883) );
  INV_X1 U4829 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3880) );
  NAND2_X1 U4830 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3879)
         );
  OAI211_X1 U4831 ( .C1(n3881), .C2(n3880), .A(n5155), .B(n3879), .ZN(n3882)
         );
  AOI21_X1 U4832 ( .B1(n5091), .B2(n3883), .A(n3882), .ZN(n3884) );
  AOI22_X1 U4833 ( .A1(n5111), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4834 ( .A1(n5135), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5112), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4835 ( .A1(n5028), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4836 ( .A1(n5076), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4837 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4838 ( .A1(n5129), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4839 ( .A1(n3311), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4840 ( .A1(n5128), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4841 ( .A1(n5109), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4842 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  NOR2_X1 U4843 ( .A1(n3895), .A2(n3894), .ZN(n3899) );
  NAND2_X1 U4844 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3896)
         );
  NAND2_X1 U4845 ( .A1(n5155), .A2(n3896), .ZN(n3897) );
  AOI21_X1 U4846 ( .B1(n3385), .B2(EAX_REG_21__SCAN_IN), .A(n3897), .ZN(n3898)
         );
  OAI21_X1 U4847 ( .B1(n5152), .B2(n3899), .A(n3898), .ZN(n3902) );
  XNOR2_X1 U4848 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3900), .ZN(n5579)
         );
  NAND2_X1 U4849 ( .A1(n5579), .A2(n5148), .ZN(n3901) );
  NAND2_X1 U4850 ( .A1(n3902), .A2(n3901), .ZN(n5482) );
  XNOR2_X1 U4851 ( .A(n5492), .B(n5482), .ZN(n5578) );
  INV_X1 U4852 ( .A(n5578), .ZN(n5300) );
  NOR2_X2 U4853 ( .A1(n5510), .A2(n3903), .ZN(n5495) );
  OR2_X1 U4854 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3906)
         );
  INV_X1 U4855 ( .A(EBX_REG_20__SCAN_IN), .ZN(n3904) );
  NAND2_X1 U4856 ( .A1(n5189), .A2(n3904), .ZN(n3905) );
  NAND2_X1 U4857 ( .A1(n3906), .A2(n3905), .ZN(n5498) );
  OAI22_X1 U4858 ( .A1(n5498), .A2(n5197), .B1(EBX_REG_20__SCAN_IN), .B2(
        EBX_REG_18__SCAN_IN), .ZN(n3909) );
  NAND2_X1 U4859 ( .A1(n5498), .A2(n5344), .ZN(n3908) );
  AND3_X1 U4860 ( .A1(n3909), .A2(n3908), .A3(n3907), .ZN(n3910) );
  NAND2_X1 U4861 ( .A1(n5495), .A2(n3910), .ZN(n3918) );
  INV_X1 U4862 ( .A(EBX_REG_21__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4863 ( .A1(n5273), .A2(n3922), .ZN(n3915) );
  NAND2_X1 U4864 ( .A1(n5189), .A2(n3922), .ZN(n3913) );
  NAND2_X1 U4865 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3911) );
  NAND3_X1 U4866 ( .A1(n3913), .A2(n3912), .A3(n3911), .ZN(n3914) );
  NAND2_X1 U4867 ( .A1(n3915), .A2(n3914), .ZN(n3917) );
  OR2_X2 U4868 ( .A1(n3918), .A2(n3917), .ZN(n5488) );
  INV_X1 U4869 ( .A(n5488), .ZN(n3916) );
  AOI21_X1 U4870 ( .B1(n3918), .B2(n3917), .A(n3916), .ZN(n5693) );
  INV_X1 U4871 ( .A(n5693), .ZN(n3919) );
  OAI22_X1 U4872 ( .A1(n5300), .A2(n5753), .B1(n3919), .B2(n5929), .ZN(n3927)
         );
  NAND4_X1 U4873 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5435), .ZN(n5770) );
  NOR2_X1 U4874 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5770), .ZN(n5784) );
  INV_X1 U4875 ( .A(n5784), .ZN(n3925) );
  AOI22_X1 U4876 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n5952), .B1(n5579), 
        .B2(n5986), .ZN(n3924) );
  INV_X1 U4877 ( .A(n5934), .ZN(n5985) );
  INV_X1 U4878 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6572) );
  OR2_X1 U4879 ( .A1(n6572), .A2(n5790), .ZN(n3920) );
  NAND2_X1 U4880 ( .A1(n5395), .A2(n3920), .ZN(n3921) );
  NAND2_X1 U4881 ( .A1(n5878), .A2(n3921), .ZN(n5791) );
  NAND2_X1 U4882 ( .A1(n5791), .A2(REIP_REG_21__SCAN_IN), .ZN(n3923) );
  NAND2_X1 U4883 ( .A1(n3925), .A2(n3127), .ZN(n3926) );
  OR2_X1 U4884 ( .A1(n4189), .A2(n4806), .ZN(n3930) );
  NAND2_X1 U4885 ( .A1(n3970), .A2(n3966), .ZN(n3928) );
  NAND2_X1 U4886 ( .A1(n3928), .A2(n3948), .ZN(n3929) );
  NAND2_X1 U4887 ( .A1(n3930), .A2(n3929), .ZN(n3937) );
  NOR2_X1 U4888 ( .A1(n3937), .A2(n6520), .ZN(n3932) );
  INV_X1 U4889 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6845) );
  NAND3_X1 U4890 ( .A1(n6606), .A2(STATE2_REG_0__SCAN_IN), .A3(n6442), .ZN(
        n3931) );
  OAI21_X1 U4891 ( .B1(n3932), .B2(n6845), .A(n3931), .ZN(U2790) );
  INV_X1 U4892 ( .A(n3933), .ZN(n3935) );
  INV_X1 U4893 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6897) );
  INV_X1 U4894 ( .A(n3955), .ZN(n3934) );
  OAI211_X1 U4895 ( .C1(n3935), .C2(n6897), .A(n3958), .B(n3934), .ZN(U2788)
         );
  INV_X1 U4896 ( .A(MORE_REG_SCAN_IN), .ZN(n6781) );
  NOR2_X1 U4897 ( .A1(n4806), .A2(n5189), .ZN(n3957) );
  NAND2_X1 U4898 ( .A1(n3957), .A2(n6536), .ZN(n6616) );
  INV_X1 U4899 ( .A(READY_N), .ZN(n6617) );
  AND2_X1 U4900 ( .A1(n6616), .A2(n6617), .ZN(n3936) );
  OR2_X1 U4901 ( .A1(n3937), .A2(n3936), .ZN(n4505) );
  AND2_X1 U4902 ( .A1(n4505), .A2(n4518), .ZN(n5862) );
  INV_X1 U4903 ( .A(n4189), .ZN(n3952) );
  NOR2_X1 U4904 ( .A1(n5159), .A2(n4216), .ZN(n3941) );
  NAND2_X1 U4905 ( .A1(n4169), .A2(n4190), .ZN(n4810) );
  NAND2_X1 U4906 ( .A1(n3938), .A2(n5345), .ZN(n3940) );
  OAI211_X1 U4907 ( .C1(n3941), .C2(n4810), .A(n3940), .B(n3939), .ZN(n3993)
         );
  INV_X1 U4908 ( .A(n4018), .ZN(n4060) );
  NOR2_X1 U4909 ( .A1(n3993), .A2(n4060), .ZN(n3945) );
  INV_X1 U4910 ( .A(n3942), .ZN(n3943) );
  NAND2_X1 U4911 ( .A1(n3943), .A2(n6009), .ZN(n3944) );
  MUX2_X1 U4912 ( .A(n6618), .B(n3944), .S(n4037), .Z(n3994) );
  NAND2_X1 U4913 ( .A1(n3998), .A2(n4190), .ZN(n4184) );
  INV_X1 U4914 ( .A(n4184), .ZN(n3946) );
  INV_X1 U4915 ( .A(n3970), .ZN(n3950) );
  INV_X1 U4916 ( .A(n3998), .ZN(n4004) );
  AND2_X1 U4917 ( .A1(n4004), .A2(n4169), .ZN(n3947) );
  NAND2_X1 U4918 ( .A1(n3971), .A2(n4806), .ZN(n4036) );
  NAND2_X1 U4919 ( .A1(n3971), .A2(n3221), .ZN(n4504) );
  AND2_X1 U4920 ( .A1(n4036), .A2(n4504), .ZN(n4202) );
  AOI21_X1 U4921 ( .B1(n4202), .B2(n3948), .A(n4189), .ZN(n3949) );
  AOI21_X1 U4922 ( .B1(n3966), .B2(n3950), .A(n3949), .ZN(n3951) );
  OAI21_X1 U4923 ( .B1(n3952), .B2(n4249), .A(n3951), .ZN(n4506) );
  NAND2_X1 U4924 ( .A1(n4506), .A2(n5862), .ZN(n3953) );
  OAI21_X1 U4925 ( .B1(n6781), .B2(n5862), .A(n3953), .ZN(U3471) );
  INV_X1 U4926 ( .A(n3954), .ZN(n6625) );
  OAI21_X1 U4927 ( .B1(n3955), .B2(READREQUEST_REG_SCAN_IN), .A(n6625), .ZN(
        n3956) );
  OAI21_X1 U4928 ( .B1(n6625), .B2(n3957), .A(n3956), .ZN(U3474) );
  INV_X1 U4929 ( .A(n6618), .ZN(n4656) );
  INV_X1 U4930 ( .A(n3958), .ZN(n3959) );
  OAI21_X2 U4931 ( .B1(n4656), .B2(n6617), .A(n3959), .ZN(n6106) );
  INV_X1 U4932 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6858) );
  INV_X1 U4933 ( .A(DATAI_11_), .ZN(n3960) );
  NOR2_X1 U4934 ( .A1(n6104), .A2(n3960), .ZN(n6095) );
  AOI21_X1 U4935 ( .B1(n6101), .B2(EAX_REG_27__SCAN_IN), .A(n6095), .ZN(n3961)
         );
  OAI21_X1 U4936 ( .B1(n6057), .B2(n6858), .A(n3961), .ZN(U2935) );
  INV_X1 U4937 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6849) );
  INV_X1 U4938 ( .A(n6104), .ZN(n6092) );
  AOI22_X1 U4939 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6101), .B1(n6092), .B2(
        DATAI_0_), .ZN(n3962) );
  OAI21_X1 U4940 ( .B1(n6057), .B2(n6849), .A(n3962), .ZN(U2924) );
  INV_X1 U4941 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6713) );
  AOI22_X1 U4942 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6101), .B1(n6092), .B2(
        DATAI_10_), .ZN(n3963) );
  OAI21_X1 U4943 ( .B1(n6057), .B2(n6713), .A(n3963), .ZN(U2934) );
  INV_X1 U4944 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n6876) );
  AOI22_X1 U4945 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6101), .B1(n6092), .B2(
        DATAI_1_), .ZN(n3964) );
  OAI21_X1 U4946 ( .B1(n6057), .B2(n6876), .A(n3964), .ZN(U2925) );
  INV_X1 U4947 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6772) );
  INV_X1 U4948 ( .A(DATAI_15_), .ZN(n3965) );
  INV_X1 U4949 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6724) );
  OAI222_X1 U4950 ( .A1(n6108), .A2(n6772), .B1(n6104), .B2(n3965), .C1(n6724), 
        .C2(n6057), .ZN(U2954) );
  NOR2_X1 U4951 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6397), .ZN(n6601) );
  NAND2_X1 U4952 ( .A1(n3966), .A2(n4190), .ZN(n5748) );
  NAND2_X1 U4953 ( .A1(n4201), .A2(n6536), .ZN(n3967) );
  NAND2_X1 U4954 ( .A1(n3967), .A2(n6617), .ZN(n3968) );
  AOI21_X1 U4955 ( .B1(n5748), .B2(n4187), .A(n3968), .ZN(n3976) );
  AND2_X1 U4956 ( .A1(n3970), .A2(n6617), .ZN(n4191) );
  INV_X1 U4957 ( .A(n4191), .ZN(n4029) );
  NAND2_X1 U4958 ( .A1(n3994), .A2(n3971), .ZN(n3973) );
  NAND2_X1 U4959 ( .A1(n3973), .A2(n3972), .ZN(n4195) );
  OR2_X1 U4960 ( .A1(n4810), .A2(n4192), .ZN(n3974) );
  OAI211_X1 U4961 ( .C1(n3969), .C2(n4029), .A(n4195), .B(n3974), .ZN(n3975)
         );
  AOI21_X1 U4962 ( .B1(n4189), .B2(n3976), .A(n3975), .ZN(n3979) );
  INV_X1 U4963 ( .A(n4036), .ZN(n3977) );
  NAND2_X1 U4964 ( .A1(n4189), .A2(n3977), .ZN(n3978) );
  INV_X1 U4965 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6826) );
  NAND2_X1 U4966 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n6527) );
  NOR2_X1 U4967 ( .A1(n6765), .A2(n6527), .ZN(n6600) );
  INV_X1 U4968 ( .A(n6600), .ZN(n3980) );
  OAI22_X1 U4969 ( .A1(n4491), .A2(n6520), .B1(n6826), .B2(n3980), .ZN(n3982)
         );
  INV_X1 U4970 ( .A(n6609), .ZN(n3985) );
  INV_X1 U4971 ( .A(n3969), .ZN(n4076) );
  INV_X1 U4972 ( .A(n6325), .ZN(n6358) );
  OR2_X1 U4973 ( .A1(n3394), .A2(n6358), .ZN(n3981) );
  XNOR2_X1 U4974 ( .A(n3981), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5968)
         );
  NAND4_X1 U4975 ( .A1(n3982), .A2(n6606), .A3(n4076), .A4(n5968), .ZN(n3983)
         );
  OAI21_X1 U4976 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(U3455) );
  INV_X1 U4977 ( .A(n3986), .ZN(n3989) );
  INV_X1 U4978 ( .A(n3987), .ZN(n3988) );
  NAND2_X1 U4979 ( .A1(n3989), .A2(n3988), .ZN(n4001) );
  INV_X1 U4980 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3990) );
  INV_X1 U4981 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6237) );
  AOI22_X1 U4982 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3990), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6237), .ZN(n4022) );
  NAND2_X1 U4983 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4023) );
  INV_X1 U4984 ( .A(n4023), .ZN(n4000) );
  INV_X1 U4985 ( .A(n5983), .ZN(n5740) );
  NAND2_X1 U4986 ( .A1(n4032), .A2(n4187), .ZN(n3992) );
  NOR2_X1 U4987 ( .A1(n3993), .A2(n3992), .ZN(n3995) );
  AND3_X1 U4988 ( .A1(n3996), .A2(n3995), .A3(n3994), .ZN(n3997) );
  AND2_X1 U4989 ( .A1(n3997), .A2(n3969), .ZN(n4012) );
  NOR2_X1 U4990 ( .A1(n5748), .A2(n6699), .ZN(n4064) );
  AOI21_X1 U4991 ( .B1(n3998), .B2(n4001), .A(n4064), .ZN(n3999) );
  OAI21_X1 U4992 ( .B1(n5740), .B2(n4012), .A(n3999), .ZN(n4489) );
  AOI222_X1 U4993 ( .A1(n4001), .A2(n6605), .B1(n4022), .B2(n4000), .C1(n4489), 
        .C2(n6606), .ZN(n4003) );
  NAND2_X1 U4994 ( .A1(n6609), .A2(n6699), .ZN(n4002) );
  OAI21_X1 U4995 ( .B1(n6609), .B2(n4003), .A(n4002), .ZN(U3460) );
  INV_X1 U4996 ( .A(n5748), .ZN(n4488) );
  AOI21_X1 U4997 ( .B1(n4488), .B2(n6606), .A(n6609), .ZN(n4008) );
  OAI22_X1 U4998 ( .A1(n4831), .A2(n4012), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4004), .ZN(n4486) );
  OAI22_X1 U4999 ( .A1(n6708), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4521), .ZN(n4005) );
  AOI21_X1 U5000 ( .B1(n4486), .B2(n6606), .A(n4005), .ZN(n4006) );
  OAI22_X1 U5001 ( .A1(n4008), .A2(n4007), .B1(n6609), .B2(n4006), .ZN(U3461)
         );
  INV_X1 U5002 ( .A(n4020), .ZN(n4051) );
  AOI21_X1 U5003 ( .B1(n4051), .B2(n6605), .A(n6609), .ZN(n4028) );
  INV_X1 U5004 ( .A(n4011), .ZN(n5464) );
  INV_X1 U5005 ( .A(n4012), .ZN(n4048) );
  XNOR2_X1 U5006 ( .A(n4020), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4017)
         );
  NOR2_X1 U5007 ( .A1(n5748), .A2(n3131), .ZN(n4013) );
  MUX2_X1 U5008 ( .A(n4013), .B(n4064), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4014) );
  INV_X1 U5009 ( .A(n4014), .ZN(n4016) );
  NAND2_X1 U5010 ( .A1(n4249), .A2(n4036), .ZN(n4054) );
  NAND2_X1 U5011 ( .A1(n4054), .A2(n4017), .ZN(n4015) );
  OAI211_X1 U5012 ( .C1(n4018), .C2(n4017), .A(n4016), .B(n4015), .ZN(n4019)
         );
  AOI21_X1 U5013 ( .B1(n5464), .B2(n4048), .A(n4019), .ZN(n4044) );
  NOR2_X1 U5014 ( .A1(n4044), .A2(n6521), .ZN(n4025) );
  NAND3_X1 U5015 ( .A1(n4020), .A2(n4027), .A3(n6605), .ZN(n4021) );
  OAI21_X1 U5016 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4024) );
  NOR2_X1 U5017 ( .A1(n4025), .A2(n4024), .ZN(n4026) );
  OAI22_X1 U5018 ( .A1(n4028), .A2(n4027), .B1(n6609), .B2(n4026), .ZN(U3459)
         );
  OR2_X1 U5019 ( .A1(n6520), .A2(n4029), .ZN(n4033) );
  NAND4_X1 U5020 ( .A1(n4349), .A2(n5383), .A3(n4518), .A4(n4031), .ZN(n4418)
         );
  OAI22_X1 U5021 ( .A1(n3969), .A2(n4033), .B1(n4032), .B2(n4418), .ZN(n4034)
         );
  INV_X1 U5022 ( .A(n4034), .ZN(n4035) );
  NAND2_X1 U5023 ( .A1(n4037), .A2(n5161), .ZN(n4040) );
  XNOR2_X1 U5024 ( .A(n4039), .B(n4038), .ZN(n4833) );
  INV_X1 U5025 ( .A(n4040), .ZN(n4041) );
  INV_X1 U5026 ( .A(DATAI_0_), .ZN(n6075) );
  INV_X1 U5027 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6056) );
  OAI222_X1 U5028 ( .A1(n5796), .A2(n4833), .B1(n4336), .B2(n6075), .C1(n5382), 
        .C2(n6056), .ZN(U2891) );
  OAI21_X1 U5029 ( .B1(n4043), .B2(n4042), .A(n3391), .ZN(n5982) );
  INV_X1 U5030 ( .A(DATAI_1_), .ZN(n6077) );
  INV_X1 U5031 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6052) );
  OAI222_X1 U5032 ( .A1(n5982), .A2(n5796), .B1(n4336), .B2(n6077), .C1(n5382), 
        .C2(n6052), .ZN(U2890) );
  OR2_X1 U5033 ( .A1(n4044), .A2(n4491), .ZN(n4046) );
  NAND2_X1 U5034 ( .A1(n4491), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U5035 ( .A1(n4046), .A2(n4045), .ZN(n4496) );
  NAND2_X1 U5036 ( .A1(n4767), .A2(n4048), .ZN(n4068) );
  CLKBUF_X1 U5037 ( .A(n4049), .Z(n4072) );
  AOI21_X1 U5038 ( .B1(n4051), .B2(n4050), .A(n4072), .ZN(n4053) );
  NAND3_X1 U5039 ( .A1(n4054), .A2(n4053), .A3(n3289), .ZN(n4066) );
  AOI21_X1 U5040 ( .B1(n4056), .B2(n6699), .A(n4055), .ZN(n4062) );
  AND2_X1 U5041 ( .A1(n6699), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4059)
         );
  OAI211_X1 U5042 ( .C1(n4059), .C2(n4058), .A(n3310), .B(n4057), .ZN(n6604)
         );
  NAND2_X1 U5043 ( .A1(n4060), .A2(n6604), .ZN(n4061) );
  OAI21_X1 U5044 ( .B1(n5748), .B2(n4062), .A(n4061), .ZN(n4063) );
  AOI21_X1 U5045 ( .B1(n4064), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4063), 
        .ZN(n4065) );
  AND2_X1 U5046 ( .A1(n4066), .A2(n4065), .ZN(n4067) );
  NAND2_X1 U5047 ( .A1(n4068), .A2(n4067), .ZN(n6607) );
  INV_X1 U5048 ( .A(n4491), .ZN(n4069) );
  NAND2_X1 U5049 ( .A1(n6607), .A2(n4069), .ZN(n4071) );
  NAND2_X1 U5050 ( .A1(n4491), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4070) );
  NAND2_X1 U5051 ( .A1(n4071), .A2(n4070), .ZN(n4501) );
  NAND3_X1 U5052 ( .A1(n4496), .A2(n6708), .A3(n4501), .ZN(n4074) );
  NOR2_X1 U5053 ( .A1(FLUSH_REG_SCAN_IN), .A2(n6708), .ZN(n4079) );
  NAND2_X1 U5054 ( .A1(n4072), .A2(n4079), .ZN(n4073) );
  NAND2_X1 U5055 ( .A1(n4074), .A2(n4073), .ZN(n4502) );
  INV_X1 U5056 ( .A(n4075), .ZN(n6638) );
  NAND2_X1 U5057 ( .A1(n4502), .A2(n6638), .ZN(n4082) );
  NAND2_X1 U5058 ( .A1(n5968), .A2(n4076), .ZN(n4078) );
  NAND2_X1 U5059 ( .A1(n4491), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4077) );
  NAND2_X1 U5060 ( .A1(n4078), .A2(n4077), .ZN(n4081) );
  AND2_X1 U5061 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4079), .ZN(n4080)
         );
  AOI21_X1 U5062 ( .B1(n4081), .B2(n6708), .A(n4080), .ZN(n4503) );
  NAND2_X1 U5063 ( .A1(n4082), .A2(n4503), .ZN(n4087) );
  OAI21_X1 U5064 ( .B1(n4087), .B2(FLUSH_REG_SCAN_IN), .A(n6600), .ZN(n4083)
         );
  NAND2_X1 U5065 ( .A1(n4353), .A2(n4083), .ZN(n6252) );
  INV_X1 U5066 ( .A(n4558), .ZN(n5743) );
  NAND2_X1 U5067 ( .A1(n5738), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5742) );
  OR3_X1 U5068 ( .A1(n4558), .A2(n3415), .A3(n5742), .ZN(n6357) );
  OAI211_X1 U5069 ( .C1(n6434), .C2(n5743), .A(n4141), .B(n6357), .ZN(n4084)
         );
  INV_X1 U5070 ( .A(n6439), .ZN(n6433) );
  AND2_X1 U5071 ( .A1(n4084), .A2(n6433), .ZN(n6256) );
  NOR2_X1 U5072 ( .A1(n6439), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6326) );
  INV_X1 U5073 ( .A(n6326), .ZN(n4112) );
  INV_X1 U5074 ( .A(n4767), .ZN(n6258) );
  AND2_X1 U5075 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6397), .ZN(n5744) );
  OAI22_X1 U5076 ( .A1(n6434), .A2(n4112), .B1(n6258), .B2(n5744), .ZN(n4085)
         );
  OAI21_X1 U5077 ( .B1(n6256), .B2(n4085), .A(n6252), .ZN(n4086) );
  OAI21_X1 U5078 ( .B1(n6252), .B2(n6320), .A(n4086), .ZN(U3462) );
  NOR2_X1 U5079 ( .A1(n4087), .A2(n6527), .ZN(n4522) );
  OAI22_X1 U5080 ( .A1(n6318), .A2(n6439), .B1(n4831), .B2(n5744), .ZN(n4088)
         );
  OAI21_X1 U5081 ( .B1(n4522), .B2(n4088), .A(n6252), .ZN(n4089) );
  OAI21_X1 U5082 ( .B1(n6252), .B2(n4487), .A(n4089), .ZN(U3465) );
  NAND2_X1 U5083 ( .A1(n4090), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6529) );
  AND2_X1 U5084 ( .A1(n4169), .A2(n4214), .ZN(n4205) );
  INV_X1 U5085 ( .A(n4205), .ZN(n4091) );
  OAI21_X1 U5086 ( .B1(n6618), .B2(n4211), .A(n4091), .ZN(n4092) );
  INV_X1 U5087 ( .A(n4092), .ZN(n4093) );
  NAND2_X1 U5088 ( .A1(n4094), .A2(n4093), .ZN(n4095) );
  NAND2_X1 U5089 ( .A1(n4095), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4221)
         );
  OAI21_X1 U5090 ( .B1(n4095), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4221), 
        .ZN(n4096) );
  INV_X1 U5091 ( .A(n4096), .ZN(n6241) );
  AND2_X1 U5092 ( .A1(n6229), .A2(REIP_REG_0__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U5093 ( .A1(n4097), .A2(n6439), .ZN(n6623) );
  NAND2_X1 U5094 ( .A1(n6623), .A2(n6765), .ZN(n4098) );
  NAND2_X1 U5095 ( .A1(n6765), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4100) );
  INV_X1 U5096 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5861) );
  NAND2_X1 U5097 ( .A1(n5861), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4099) );
  AND2_X1 U5098 ( .A1(n4100), .A2(n4099), .ZN(n4603) );
  INV_X1 U5099 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4101) );
  AOI21_X1 U5100 ( .B1(n5616), .B2(n4603), .A(n4101), .ZN(n4102) );
  AOI211_X1 U5101 ( .C1(n6241), .C2(n6135), .A(n6239), .B(n4102), .ZN(n4103)
         );
  OAI21_X1 U5102 ( .B1(n4833), .B2(n5617), .A(n4103), .ZN(U2986) );
  INV_X1 U5103 ( .A(n3391), .ZN(n4106) );
  INV_X1 U5104 ( .A(n4104), .ZN(n4105) );
  NOR3_X1 U5105 ( .A1(n4107), .A2(n4106), .A3(n4105), .ZN(n4109) );
  NOR2_X1 U5106 ( .A1(n4109), .A2(n4108), .ZN(n6126) );
  INV_X1 U5107 ( .A(n6126), .ZN(n4715) );
  INV_X1 U5108 ( .A(DATAI_2_), .ZN(n6079) );
  INV_X1 U5109 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6050) );
  OAI222_X1 U5110 ( .A1(n4715), .A2(n5796), .B1(n4336), .B2(n6079), .C1(n5382), 
        .C2(n6050), .ZN(U2889) );
  OAI21_X1 U5111 ( .B1(n4108), .B2(n4111), .A(n4110), .ZN(n4819) );
  INV_X1 U5112 ( .A(DATAI_3_), .ZN(n6894) );
  INV_X1 U5113 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6690) );
  OAI222_X1 U5114 ( .A1(n4819), .A2(n5796), .B1(n4336), .B2(n6894), .C1(n5382), 
        .C2(n6690), .ZN(U2888) );
  INV_X1 U5115 ( .A(n5738), .ZN(n4264) );
  OR2_X1 U5116 ( .A1(n6356), .A2(n6354), .ZN(n4122) );
  NAND2_X1 U5117 ( .A1(n4122), .A2(n6137), .ZN(n4113) );
  NAND2_X1 U5118 ( .A1(n4113), .A2(n4112), .ZN(n4115) );
  OR2_X1 U5119 ( .A1(n4011), .A2(n5740), .ZN(n6324) );
  NOR2_X1 U5120 ( .A1(n6324), .A2(n4831), .ZN(n6359) );
  INV_X1 U5121 ( .A(n4180), .ZN(n6944) );
  AOI21_X1 U5122 ( .B1(n6359), .B2(n4767), .A(n6944), .ZN(n4114) );
  NAND2_X1 U5123 ( .A1(n4115), .A2(n4114), .ZN(n4117) );
  AOI21_X1 U5124 ( .B1(n6439), .B2(n4312), .A(n6438), .ZN(n4116) );
  NAND2_X1 U5125 ( .A1(n4117), .A2(n4116), .ZN(n6956) );
  OR2_X1 U5126 ( .A1(n6354), .A2(n6318), .ZN(n4118) );
  NAND2_X1 U5127 ( .A1(n6137), .A2(DATAI_17_), .ZN(n6451) );
  NOR2_X2 U5128 ( .A1(n4355), .A2(n4121), .ZN(n6490) );
  NAND2_X1 U5129 ( .A1(n6490), .A2(n6944), .ZN(n4124) );
  NAND2_X1 U5130 ( .A1(n6137), .A2(DATAI_25_), .ZN(n6408) );
  INV_X1 U5131 ( .A(n6408), .ZN(n6493) );
  NAND2_X1 U5132 ( .A1(n6947), .A2(n6493), .ZN(n4123) );
  OAI211_X1 U5133 ( .C1(n6950), .C2(n6451), .A(n4124), .B(n4123), .ZN(n4127)
         );
  NOR2_X2 U5134 ( .A1(n6077), .A2(n4353), .ZN(n6491) );
  INV_X1 U5135 ( .A(n6491), .ZN(n4628) );
  NAND2_X1 U5136 ( .A1(n4767), .A2(n6433), .ZN(n6392) );
  INV_X1 U5137 ( .A(n6392), .ZN(n4136) );
  NOR2_X1 U5138 ( .A1(n4628), .A2(n6952), .ZN(n4126) );
  AOI211_X1 U5139 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n6956), .A(n4127), 
        .B(n4126), .ZN(n4128) );
  INV_X1 U5140 ( .A(n4128), .ZN(U3141) );
  NAND2_X1 U5141 ( .A1(n6137), .A2(DATAI_23_), .ZN(n6482) );
  NOR2_X2 U5142 ( .A1(n4355), .A2(n5383), .ZN(n6509) );
  NAND2_X1 U5143 ( .A1(n6509), .A2(n6944), .ZN(n4130) );
  NAND2_X1 U5144 ( .A1(n6137), .A2(DATAI_31_), .ZN(n6430) );
  INV_X1 U5145 ( .A(n6430), .ZN(n6514) );
  NAND2_X1 U5146 ( .A1(n6947), .A2(n6514), .ZN(n4129) );
  OAI211_X1 U5147 ( .C1(n6950), .C2(n6482), .A(n4130), .B(n4129), .ZN(n4132)
         );
  INV_X1 U5148 ( .A(DATAI_7_), .ZN(n6086) );
  NOR2_X2 U5149 ( .A1(n6086), .A2(n4353), .ZN(n6511) );
  INV_X1 U5150 ( .A(n6511), .ZN(n4631) );
  NOR2_X1 U5151 ( .A1(n4631), .A2(n6952), .ZN(n4131) );
  AOI211_X1 U5152 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n6956), .A(n4132), 
        .B(n4131), .ZN(n4133) );
  INV_X1 U5153 ( .A(n4133), .ZN(U3147) );
  OR2_X1 U5154 ( .A1(n6439), .A2(n5861), .ZN(n4134) );
  NAND2_X1 U5155 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4152), .ZN(n4763) );
  OAI21_X1 U5156 ( .B1(n4141), .B2(n4134), .A(n4763), .ZN(n4135) );
  INV_X1 U5157 ( .A(n6438), .ZN(n4382) );
  INV_X1 U5158 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4146) );
  NOR2_X2 U5159 ( .A1(n6894), .A2(n4353), .ZN(n6455) );
  NOR2_X1 U5160 ( .A1(n4487), .A2(n4763), .ZN(n6508) );
  INV_X1 U5161 ( .A(n6508), .ZN(n4139) );
  INV_X1 U5162 ( .A(n4152), .ZN(n4138) );
  NAND2_X1 U5163 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        STATE2_REG_2__SCAN_IN), .ZN(n4137) );
  NOR2_X1 U5164 ( .A1(n4011), .A2(n5983), .ZN(n6286) );
  NAND2_X1 U5165 ( .A1(n4136), .A2(n6286), .ZN(n4762) );
  OAI222_X1 U5166 ( .A1(n4139), .A2(n6439), .B1(n4138), .B2(n4137), .C1(n4831), 
        .C2(n4762), .ZN(n6510) );
  NAND2_X1 U5167 ( .A1(n6455), .A2(n6510), .ZN(n4145) );
  NOR2_X2 U5168 ( .A1(n4355), .A2(n4140), .ZN(n6945) );
  NOR2_X2 U5169 ( .A1(n4141), .A2(n6318), .ZN(n6513) );
  INV_X1 U5170 ( .A(n6513), .ZN(n4368) );
  NAND2_X1 U5171 ( .A1(n6137), .A2(DATAI_19_), .ZN(n6951) );
  NAND2_X1 U5172 ( .A1(n6137), .A2(DATAI_27_), .ZN(n6415) );
  INV_X1 U5173 ( .A(n4141), .ZN(n4142) );
  OAI22_X1 U5174 ( .A1(n4368), .A2(n6951), .B1(n6415), .B2(n6485), .ZN(n4143)
         );
  AOI21_X1 U5175 ( .B1(n6945), .B2(n6508), .A(n4143), .ZN(n4144) );
  OAI211_X1 U5176 ( .C1(n6518), .C2(n4146), .A(n4145), .B(n4144), .ZN(U3127)
         );
  CLKBUF_X1 U5177 ( .A(n4147), .Z(n4283) );
  AND2_X1 U5178 ( .A1(n4110), .A2(n4148), .ZN(n4149) );
  NOR2_X1 U5179 ( .A1(n4283), .A2(n4149), .ZN(n5974) );
  INV_X1 U5180 ( .A(n5974), .ZN(n4427) );
  AOI22_X1 U5181 ( .A1(n5535), .A2(DATAI_4_), .B1(n6005), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4150) );
  OAI21_X1 U5182 ( .B1(n4427), .B2(n5796), .A(n4150), .ZN(U2887) );
  INV_X1 U5183 ( .A(n4156), .ZN(n4151) );
  AOI21_X1 U5184 ( .B1(n4151), .B2(STATEBS16_REG_SCAN_IN), .A(n6439), .ZN(
        n6294) );
  NAND2_X1 U5185 ( .A1(n6286), .A2(n6358), .ZN(n6293) );
  OR2_X1 U5186 ( .A1(n6293), .A2(n4831), .ZN(n4154) );
  NAND2_X1 U5187 ( .A1(n4152), .A2(n6320), .ZN(n6290) );
  NOR2_X1 U5188 ( .A1(n4487), .A2(n6290), .ZN(n4359) );
  INV_X1 U5189 ( .A(n4359), .ZN(n4153) );
  NAND2_X1 U5190 ( .A1(n4154), .A2(n4153), .ZN(n4159) );
  INV_X1 U5191 ( .A(n6290), .ZN(n4155) );
  AOI22_X1 U5192 ( .A1(n6294), .A2(n4159), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4155), .ZN(n4363) );
  INV_X1 U5193 ( .A(n6349), .ZN(n4357) );
  OAI22_X1 U5194 ( .A1(n6451), .A2(n4357), .B1(n4356), .B2(n6408), .ZN(n4157)
         );
  AOI21_X1 U5195 ( .B1(n6490), .B2(n4359), .A(n4157), .ZN(n4162) );
  INV_X1 U5196 ( .A(n6294), .ZN(n4160) );
  AOI21_X1 U5197 ( .B1(n6290), .B2(n6439), .A(n6438), .ZN(n4158) );
  NAND2_X1 U5198 ( .A1(n4360), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4161) );
  OAI211_X1 U5199 ( .C1(n4628), .C2(n4363), .A(n4162), .B(n4161), .ZN(U3061)
         );
  OAI22_X1 U5200 ( .A1(n6482), .A2(n4357), .B1(n4356), .B2(n6430), .ZN(n4163)
         );
  AOI21_X1 U5201 ( .B1(n6509), .B2(n4359), .A(n4163), .ZN(n4165) );
  NAND2_X1 U5202 ( .A1(n4360), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4164) );
  OAI211_X1 U5203 ( .C1(n4631), .C2(n4363), .A(n4165), .B(n4164), .ZN(U3067)
         );
  INV_X1 U5204 ( .A(n6455), .ZN(n6953) );
  OAI22_X1 U5205 ( .A1(n6951), .A2(n4357), .B1(n4356), .B2(n6415), .ZN(n4166)
         );
  AOI21_X1 U5206 ( .B1(n6945), .B2(n4359), .A(n4166), .ZN(n4168) );
  NAND2_X1 U5207 ( .A1(n4360), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4167) );
  OAI211_X1 U5208 ( .C1(n6953), .C2(n4363), .A(n4168), .B(n4167), .ZN(U3063)
         );
  NOR2_X2 U5209 ( .A1(n6075), .A2(n4353), .ZN(n6484) );
  INV_X1 U5210 ( .A(n6484), .ZN(n4667) );
  NOR2_X2 U5211 ( .A1(n4355), .A2(n4169), .ZN(n6483) );
  INV_X1 U5212 ( .A(DATAI_16_), .ZN(n4170) );
  NOR2_X1 U5213 ( .A1(n5617), .A2(n4170), .ZN(n6486) );
  INV_X1 U5214 ( .A(n6486), .ZN(n6448) );
  INV_X1 U5215 ( .A(DATAI_24_), .ZN(n4171) );
  NOR2_X1 U5216 ( .A1(n5617), .A2(n4171), .ZN(n6487) );
  INV_X1 U5217 ( .A(n6487), .ZN(n6405) );
  OAI22_X1 U5218 ( .A1(n6448), .A2(n4357), .B1(n4356), .B2(n6405), .ZN(n4172)
         );
  AOI21_X1 U5219 ( .B1(n6483), .B2(n4359), .A(n4172), .ZN(n4174) );
  NAND2_X1 U5220 ( .A1(n4360), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4173) );
  OAI211_X1 U5221 ( .C1(n4667), .C2(n4363), .A(n4174), .B(n4173), .ZN(U3060)
         );
  NOR2_X2 U5222 ( .A1(n6079), .A2(n4353), .ZN(n6496) );
  INV_X1 U5223 ( .A(n6496), .ZN(n4679) );
  NOR2_X2 U5224 ( .A1(n4355), .A2(n4216), .ZN(n6497) );
  INV_X1 U5225 ( .A(DATAI_18_), .ZN(n4175) );
  NOR2_X1 U5226 ( .A1(n5617), .A2(n4175), .ZN(n6498) );
  INV_X1 U5227 ( .A(n6498), .ZN(n6454) );
  INV_X1 U5228 ( .A(DATAI_26_), .ZN(n4176) );
  NOR2_X1 U5229 ( .A1(n5617), .A2(n4176), .ZN(n6499) );
  INV_X1 U5230 ( .A(n6499), .ZN(n6411) );
  OAI22_X1 U5231 ( .A1(n6454), .A2(n4357), .B1(n4356), .B2(n6411), .ZN(n4177)
         );
  AOI21_X1 U5232 ( .B1(n6497), .B2(n4359), .A(n4177), .ZN(n4179) );
  NAND2_X1 U5233 ( .A1(n4360), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5234 ( .C1(n4679), .C2(n4363), .A(n4179), .B(n4178), .ZN(U3062)
         );
  NOR2_X1 U5235 ( .A1(n4477), .A2(n6405), .ZN(n4182) );
  INV_X1 U5236 ( .A(n6483), .ZN(n4302) );
  OAI22_X1 U5237 ( .A1(n4302), .A2(n4180), .B1(n6448), .B2(n6950), .ZN(n4181)
         );
  AOI211_X1 U5238 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n6956), .A(n4182), 
        .B(n4181), .ZN(n4183) );
  OAI21_X1 U5239 ( .B1(n6952), .B2(n4667), .A(n4183), .ZN(U3140) );
  OR2_X1 U5240 ( .A1(n4189), .A2(n4184), .ZN(n4197) );
  NAND2_X1 U5241 ( .A1(n4185), .A2(n6617), .ZN(n4186) );
  OAI211_X1 U5242 ( .C1(n4187), .C2(n4186), .A(n6009), .B(n5159), .ZN(n4188)
         );
  NAND3_X1 U5243 ( .A1(n4189), .A2(n4216), .A3(n4188), .ZN(n4196) );
  NAND2_X1 U5244 ( .A1(n4190), .A2(n6536), .ZN(n4193) );
  NAND3_X1 U5245 ( .A1(n4193), .A2(n4192), .A3(n4191), .ZN(n4194) );
  NAND4_X1 U5246 ( .A1(n4197), .A2(n4196), .A3(n4195), .A4(n4194), .ZN(n4198)
         );
  OR2_X1 U5247 ( .A1(n4199), .A2(n4349), .ZN(n4200) );
  AND4_X1 U5248 ( .A1(n4202), .A2(n3969), .A3(n4201), .A4(n4200), .ZN(n4203)
         );
  NAND2_X1 U5249 ( .A1(n4211), .A2(n4212), .ZN(n4210) );
  NAND2_X1 U5250 ( .A1(n4210), .A2(n4204), .ZN(n4228) );
  OAI21_X1 U5251 ( .B1(n4204), .B2(n4210), .A(n4228), .ZN(n4206) );
  AOI21_X1 U5252 ( .B1(n4206), .B2(n4656), .A(n4205), .ZN(n4207) );
  OAI21_X1 U5253 ( .B1(n4208), .B2(n4650), .A(n4207), .ZN(n4224) );
  NAND2_X1 U5254 ( .A1(n4224), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6122)
         );
  INV_X1 U5255 ( .A(n4650), .ZN(n4538) );
  NAND2_X1 U5256 ( .A1(n4209), .A2(n4538), .ZN(n4220) );
  OAI21_X1 U5257 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4213) );
  INV_X1 U5258 ( .A(n4213), .ZN(n4218) );
  NAND3_X1 U5259 ( .A1(n4216), .A2(n3220), .A3(n4214), .ZN(n4217) );
  AOI21_X1 U5260 ( .B1(n4656), .B2(n4218), .A(n4217), .ZN(n4219) );
  NAND2_X1 U5261 ( .A1(n4220), .A2(n4219), .ZN(n6133) );
  XNOR2_X1 U5262 ( .A(n4221), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6132)
         );
  NAND2_X1 U5263 ( .A1(n6133), .A2(n6132), .ZN(n6131) );
  INV_X1 U5264 ( .A(n4221), .ZN(n4222) );
  NAND2_X1 U5265 ( .A1(n4222), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4223)
         );
  AND2_X1 U5266 ( .A1(n6131), .A2(n4223), .ZN(n6125) );
  NAND2_X1 U5267 ( .A1(n6122), .A2(n6125), .ZN(n4227) );
  INV_X1 U5268 ( .A(n4224), .ZN(n4226) );
  AND2_X1 U5269 ( .A1(n4227), .A2(n6123), .ZN(n4607) );
  NAND2_X1 U5270 ( .A1(n4228), .A2(n4229), .ZN(n4244) );
  OAI211_X1 U5271 ( .C1(n4229), .C2(n4228), .A(n4244), .B(n4656), .ZN(n4230)
         );
  OAI21_X2 U5272 ( .B1(n4231), .B2(n4650), .A(n4230), .ZN(n4232) );
  XNOR2_X1 U5273 ( .A(n4232), .B(n6215), .ZN(n4609) );
  NAND2_X1 U5274 ( .A1(n4607), .A2(n4609), .ZN(n4234) );
  NAND2_X1 U5275 ( .A1(n4232), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4233)
         );
  NAND2_X1 U5276 ( .A1(n4234), .A2(n4233), .ZN(n4601) );
  NAND2_X1 U5277 ( .A1(n4235), .A2(n4538), .ZN(n4238) );
  XNOR2_X1 U5278 ( .A(n4244), .B(n4242), .ZN(n4236) );
  NAND2_X1 U5279 ( .A1(n4236), .A2(n4656), .ZN(n4237) );
  NAND2_X1 U5280 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  INV_X1 U5281 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6203) );
  XNOR2_X1 U5282 ( .A(n4239), .B(n6203), .ZN(n4602) );
  NAND2_X1 U5283 ( .A1(n4601), .A2(n4602), .ZN(n4241) );
  NAND2_X1 U5284 ( .A1(n4239), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4240)
         );
  NAND2_X1 U5285 ( .A1(n4241), .A2(n4240), .ZN(n4533) );
  INV_X1 U5286 ( .A(n4242), .ZN(n4243) );
  NOR2_X1 U5287 ( .A1(n4244), .A2(n4243), .ZN(n4246) );
  NAND2_X1 U5288 ( .A1(n4246), .A2(n4245), .ZN(n4542) );
  OAI211_X1 U5289 ( .C1(n4246), .C2(n4245), .A(n4542), .B(n4656), .ZN(n4247)
         );
  OAI21_X1 U5290 ( .B1(n4248), .B2(n4650), .A(n4247), .ZN(n4534) );
  INV_X1 U5291 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4259) );
  XNOR2_X1 U5292 ( .A(n4534), .B(n4259), .ZN(n4532) );
  XNOR2_X1 U5293 ( .A(n4533), .B(n4532), .ZN(n4722) );
  INV_X1 U5294 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U5295 ( .B1(n6243), .B2(n6237), .A(n4225), .ZN(n6217) );
  NAND3_X1 U5296 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n6217), .ZN(n4252) );
  NOR2_X1 U5297 ( .A1(n5711), .A2(n4252), .ZN(n4550) );
  OR2_X1 U5298 ( .A1(n4258), .A2(n4250), .ZN(n4892) );
  NAND2_X1 U5299 ( .A1(n5711), .A2(n4892), .ZN(n4898) );
  INV_X1 U5300 ( .A(n6245), .ZN(n4251) );
  INV_X1 U5301 ( .A(n6232), .ZN(n5356) );
  NOR2_X1 U5302 ( .A1(n4259), .A2(n4252), .ZN(n4554) );
  INV_X1 U5303 ( .A(n6229), .ZN(n6205) );
  NAND2_X1 U5304 ( .A1(n6205), .A2(n4258), .ZN(n6244) );
  NAND2_X1 U5305 ( .A1(n6243), .A2(n4898), .ZN(n6249) );
  NAND2_X1 U5306 ( .A1(n4549), .A2(n5711), .ZN(n4254) );
  NAND2_X1 U5307 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U5308 ( .A1(n5708), .A2(n6218), .ZN(n4253) );
  NAND2_X1 U5309 ( .A1(n4254), .A2(n4253), .ZN(n6223) );
  INV_X1 U5310 ( .A(n6223), .ZN(n4255) );
  OAI21_X1 U5311 ( .B1(n5356), .B2(n4554), .A(n4255), .ZN(n6181) );
  OAI21_X1 U5312 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4550), .A(n6181), 
        .ZN(n4263) );
  OR2_X1 U5313 ( .A1(n4199), .A2(n3225), .ZN(n4256) );
  AND2_X1 U5314 ( .A1(n5747), .A2(n4256), .ZN(n4257) );
  XNOR2_X1 U5315 ( .A(n4428), .B(n4430), .ZN(n5954) );
  INV_X1 U5316 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6553) );
  NOR2_X1 U5317 ( .A1(n6205), .A2(n6553), .ZN(n4261) );
  NAND2_X1 U5318 ( .A1(n6245), .A2(n6243), .ZN(n6231) );
  INV_X1 U5319 ( .A(n5326), .ZN(n6224) );
  NAND2_X1 U5320 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6193) );
  NOR2_X1 U5321 ( .A1(n6218), .A2(n6193), .ZN(n4548) );
  AND3_X1 U5322 ( .A1(n6224), .A2(n4548), .A3(n4259), .ZN(n4260) );
  AOI211_X1 U5323 ( .C1(n6247), .C2(n5954), .A(n4261), .B(n4260), .ZN(n4262)
         );
  OAI211_X1 U5324 ( .C1(n6196), .C2(n4722), .A(n4263), .B(n4262), .ZN(U3013)
         );
  NAND2_X1 U5325 ( .A1(n4558), .A2(n4264), .ZN(n4377) );
  INV_X1 U5326 ( .A(n4377), .ZN(n4265) );
  NAND2_X1 U5327 ( .A1(n4011), .A2(n5740), .ZN(n6391) );
  NOR2_X1 U5328 ( .A1(n6391), .A2(n4831), .ZN(n4379) );
  NAND3_X1 U5329 ( .A1(n6320), .A2(n4495), .A3(n4378), .ZN(n4284) );
  NOR2_X1 U5330 ( .A1(n4487), .A2(n4284), .ZN(n4415) );
  AOI21_X1 U5331 ( .B1(n4379), .B2(n6258), .A(n4415), .ZN(n4269) );
  AOI21_X1 U5332 ( .B1(n4270), .B2(STATEBS16_REG_SCAN_IN), .A(n6439), .ZN(
        n4267) );
  AOI22_X1 U5333 ( .A1(n4269), .A2(n4267), .B1(n6439), .B2(n4284), .ZN(n4266)
         );
  NAND2_X1 U5334 ( .A1(n4382), .A2(n4266), .ZN(n4414) );
  INV_X1 U5335 ( .A(n4267), .ZN(n4268) );
  OAI22_X1 U5336 ( .A1(n4269), .A2(n4268), .B1(n6442), .B2(n4284), .ZN(n4413)
         );
  AOI22_X1 U5337 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4414), .B1(n6455), 
        .B2(n4413), .ZN(n4272) );
  INV_X1 U5338 ( .A(n6415), .ZN(n6946) );
  AOI22_X1 U5339 ( .A1(n6946), .A2(n4447), .B1(n6945), .B2(n4415), .ZN(n4271)
         );
  OAI211_X1 U5340 ( .C1(n6951), .C2(n4595), .A(n4272), .B(n4271), .ZN(U3031)
         );
  AOI22_X1 U5341 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4414), .B1(n6511), 
        .B2(n4413), .ZN(n4274) );
  AOI22_X1 U5342 ( .A1(n6514), .A2(n4447), .B1(n6509), .B2(n4415), .ZN(n4273)
         );
  OAI211_X1 U5343 ( .C1(n6482), .C2(n4595), .A(n4274), .B(n4273), .ZN(U3035)
         );
  AOI22_X1 U5344 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4414), .B1(n6491), 
        .B2(n4413), .ZN(n4276) );
  AOI22_X1 U5345 ( .A1(n6493), .A2(n4447), .B1(n6490), .B2(n4415), .ZN(n4275)
         );
  OAI211_X1 U5346 ( .C1(n6451), .C2(n4595), .A(n4276), .B(n4275), .ZN(U3029)
         );
  AOI22_X1 U5347 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4414), .B1(n6484), 
        .B2(n4413), .ZN(n4278) );
  AOI22_X1 U5348 ( .A1(n6483), .A2(n4415), .B1(n4447), .B2(n6487), .ZN(n4277)
         );
  OAI211_X1 U5349 ( .C1(n6448), .C2(n4595), .A(n4278), .B(n4277), .ZN(U3028)
         );
  AOI22_X1 U5350 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4414), .B1(n6496), 
        .B2(n4413), .ZN(n4280) );
  AOI22_X1 U5351 ( .A1(n6497), .A2(n4415), .B1(n4447), .B2(n6499), .ZN(n4279)
         );
  OAI211_X1 U5352 ( .C1(n6454), .C2(n4595), .A(n4280), .B(n4279), .ZN(U3030)
         );
  INV_X1 U5353 ( .A(n4335), .ZN(n4281) );
  OAI21_X1 U5354 ( .B1(n4283), .B2(n4282), .A(n4281), .ZN(n5955) );
  INV_X1 U5355 ( .A(DATAI_5_), .ZN(n6693) );
  INV_X1 U5356 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6044) );
  OAI222_X1 U5357 ( .A1(n5955), .A2(n5796), .B1(n4336), .B2(n6693), .C1(n5382), 
        .C2(n6044), .ZN(U2886) );
  NAND2_X1 U5358 ( .A1(n6391), .A2(n6433), .ZN(n6399) );
  INV_X1 U5359 ( .A(n6950), .ZN(n4342) );
  AOI211_X1 U5360 ( .C1(n6392), .C2(n6399), .A(n4342), .B(n4447), .ZN(n4288)
         );
  OR2_X1 U5361 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4284), .ZN(n4444)
         );
  INV_X1 U5362 ( .A(n4761), .ZN(n4285) );
  NOR2_X1 U5363 ( .A1(n4285), .A2(n6321), .ZN(n4293) );
  OAI21_X1 U5364 ( .B1(n4293), .B2(n6442), .A(n4764), .ZN(n6291) );
  AOI21_X1 U5365 ( .B1(n4444), .B2(STATE2_REG_3__SCAN_IN), .A(n6291), .ZN(
        n4286) );
  NAND2_X1 U5366 ( .A1(n4291), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6288) );
  INV_X1 U5367 ( .A(n6288), .ZN(n6322) );
  AOI21_X1 U5368 ( .B1(n6391), .B2(n6326), .A(n6322), .ZN(n6396) );
  NAND2_X1 U5369 ( .A1(n4286), .A2(n6396), .ZN(n4287) );
  INV_X1 U5370 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4296) );
  INV_X1 U5371 ( .A(n6951), .ZN(n6412) );
  INV_X1 U5372 ( .A(n6945), .ZN(n4289) );
  OAI22_X1 U5373 ( .A1(n4289), .A2(n4444), .B1(n6415), .B2(n6950), .ZN(n4290)
         );
  AOI21_X1 U5374 ( .B1(n6412), .B2(n4447), .A(n4290), .ZN(n4295) );
  INV_X1 U5375 ( .A(n4291), .ZN(n4292) );
  NAND2_X1 U5376 ( .A1(n4292), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6390) );
  INV_X1 U5377 ( .A(n4293), .ZN(n6287) );
  OAI22_X1 U5378 ( .A1(n6400), .A2(n6391), .B1(n6390), .B2(n6287), .ZN(n4448)
         );
  NAND2_X1 U5379 ( .A1(n6455), .A2(n4448), .ZN(n4294) );
  OAI211_X1 U5380 ( .C1(n4451), .C2(n4296), .A(n4295), .B(n4294), .ZN(U3023)
         );
  INV_X1 U5381 ( .A(n6451), .ZN(n6492) );
  INV_X1 U5382 ( .A(n6490), .ZN(n4297) );
  OAI22_X1 U5383 ( .A1(n4297), .A2(n4444), .B1(n6408), .B2(n6950), .ZN(n4298)
         );
  AOI21_X1 U5384 ( .B1(n6492), .B2(n4447), .A(n4298), .ZN(n4300) );
  NAND2_X1 U5385 ( .A1(n6491), .A2(n4448), .ZN(n4299) );
  OAI211_X1 U5386 ( .C1(n4451), .C2(n4301), .A(n4300), .B(n4299), .ZN(U3021)
         );
  OAI22_X1 U5387 ( .A1(n4302), .A2(n4444), .B1(n6405), .B2(n6950), .ZN(n4303)
         );
  AOI21_X1 U5388 ( .B1(n6486), .B2(n4447), .A(n4303), .ZN(n4305) );
  NAND2_X1 U5389 ( .A1(n6484), .A2(n4448), .ZN(n4304) );
  OAI211_X1 U5390 ( .C1(n4451), .C2(n6747), .A(n4305), .B(n4304), .ZN(U3020)
         );
  INV_X1 U5391 ( .A(n6482), .ZN(n6512) );
  INV_X1 U5392 ( .A(n6509), .ZN(n4306) );
  OAI22_X1 U5393 ( .A1(n4306), .A2(n4444), .B1(n6430), .B2(n6950), .ZN(n4307)
         );
  AOI21_X1 U5394 ( .B1(n6512), .B2(n4447), .A(n4307), .ZN(n4309) );
  NAND2_X1 U5395 ( .A1(n6511), .A2(n4448), .ZN(n4308) );
  OAI211_X1 U5396 ( .C1(n4451), .C2(n4310), .A(n4309), .B(n4308), .ZN(U3027)
         );
  NOR3_X1 U5397 ( .A1(n6947), .A2(n6513), .A3(n6439), .ZN(n4311) );
  OAI22_X1 U5398 ( .A1(n4311), .A2(n6326), .B1(n6358), .B2(n6324), .ZN(n4315)
         );
  OAI21_X1 U5399 ( .B1(n6321), .B2(n6442), .A(n4764), .ZN(n4562) );
  AOI21_X1 U5400 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6320), .A(n4562), .ZN(
        n4624) );
  NOR2_X1 U5401 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4312), .ZN(n4475)
         );
  INV_X1 U5402 ( .A(n4475), .ZN(n4313) );
  INV_X1 U5403 ( .A(n6390), .ZN(n6328) );
  AOI21_X1 U5404 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n4313), .A(n6328), .ZN(
        n4314) );
  INV_X1 U5405 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4320) );
  NAND3_X1 U5406 ( .A1(n6322), .A2(n6321), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4316) );
  OAI21_X1 U5407 ( .B1(n6392), .B2(n6324), .A(n4316), .ZN(n4479) );
  AOI22_X1 U5408 ( .A1(n6483), .A2(n4475), .B1(n6487), .B2(n6513), .ZN(n4317)
         );
  OAI21_X1 U5409 ( .B1(n6448), .B2(n4477), .A(n4317), .ZN(n4318) );
  AOI21_X1 U5410 ( .B1(n6484), .B2(n4479), .A(n4318), .ZN(n4319) );
  OAI21_X1 U5411 ( .B1(n4482), .B2(n4320), .A(n4319), .ZN(U3132) );
  INV_X1 U5412 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5413 ( .A1(n6945), .A2(n4475), .B1(n6946), .B2(n6513), .ZN(n4321)
         );
  OAI21_X1 U5414 ( .B1(n6951), .B2(n4477), .A(n4321), .ZN(n4322) );
  AOI21_X1 U5415 ( .B1(n6455), .B2(n4479), .A(n4322), .ZN(n4323) );
  OAI21_X1 U5416 ( .B1(n4482), .B2(n4324), .A(n4323), .ZN(U3135) );
  INV_X1 U5417 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4328) );
  AOI22_X1 U5418 ( .A1(n6490), .A2(n4475), .B1(n6493), .B2(n6513), .ZN(n4325)
         );
  OAI21_X1 U5419 ( .B1(n6451), .B2(n4477), .A(n4325), .ZN(n4326) );
  AOI21_X1 U5420 ( .B1(n6491), .B2(n4479), .A(n4326), .ZN(n4327) );
  OAI21_X1 U5421 ( .B1(n4482), .B2(n4328), .A(n4327), .ZN(U3133) );
  INV_X1 U5422 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4332) );
  AOI22_X1 U5423 ( .A1(n6509), .A2(n4475), .B1(n6514), .B2(n6513), .ZN(n4329)
         );
  OAI21_X1 U5424 ( .B1(n6482), .B2(n4477), .A(n4329), .ZN(n4330) );
  AOI21_X1 U5425 ( .B1(n6511), .B2(n4479), .A(n4330), .ZN(n4331) );
  OAI21_X1 U5426 ( .B1(n4482), .B2(n4332), .A(n4331), .ZN(U3139) );
  OAI21_X1 U5427 ( .B1(n4335), .B2(n4334), .A(n4333), .ZN(n5944) );
  INV_X1 U5428 ( .A(DATAI_6_), .ZN(n6084) );
  OAI222_X1 U5429 ( .A1(n5944), .A2(n5796), .B1(n4336), .B2(n6084), .C1(n5382), 
        .C2(n3478), .ZN(U2885) );
  INV_X1 U5430 ( .A(n6497), .ZN(n4337) );
  OAI22_X1 U5431 ( .A1(n4337), .A2(n4444), .B1(n6411), .B2(n6950), .ZN(n4338)
         );
  AOI21_X1 U5432 ( .B1(n6498), .B2(n4447), .A(n4338), .ZN(n4340) );
  NAND2_X1 U5433 ( .A1(n6496), .A2(n4448), .ZN(n4339) );
  OAI211_X1 U5434 ( .C1(n4451), .C2(n4341), .A(n4340), .B(n4339), .ZN(U3022)
         );
  AOI22_X1 U5435 ( .A1(n6497), .A2(n6944), .B1(n6498), .B2(n4342), .ZN(n4343)
         );
  OAI21_X1 U5436 ( .B1(n6411), .B2(n4477), .A(n4343), .ZN(n4344) );
  AOI21_X1 U5437 ( .B1(INSTQUEUE_REG_15__2__SCAN_IN), .B2(n6956), .A(n4344), 
        .ZN(n4345) );
  OAI21_X1 U5438 ( .B1(n6952), .B2(n4679), .A(n4345), .ZN(U3142) );
  NOR2_X2 U5439 ( .A1(n6693), .A2(n4353), .ZN(n6503) );
  INV_X1 U5440 ( .A(n6503), .ZN(n4682) );
  NOR2_X2 U5441 ( .A1(n4355), .A2(n5162), .ZN(n6502) );
  NAND2_X1 U5442 ( .A1(n6137), .A2(DATAI_21_), .ZN(n6380) );
  NAND2_X1 U5443 ( .A1(n6137), .A2(DATAI_29_), .ZN(n6468) );
  OAI22_X1 U5444 ( .A1(n6380), .A2(n4357), .B1(n4356), .B2(n6468), .ZN(n4346)
         );
  AOI21_X1 U5445 ( .B1(n6502), .B2(n4359), .A(n4346), .ZN(n4348) );
  NAND2_X1 U5446 ( .A1(n4360), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4347) );
  OAI211_X1 U5447 ( .C1(n4682), .C2(n4363), .A(n4348), .B(n4347), .ZN(U3065)
         );
  INV_X1 U5448 ( .A(DATAI_4_), .ZN(n6808) );
  NOR2_X2 U5449 ( .A1(n6808), .A2(n4353), .ZN(n6460) );
  INV_X1 U5450 ( .A(n6460), .ZN(n4691) );
  NOR2_X2 U5451 ( .A1(n4355), .A2(n4349), .ZN(n6459) );
  NAND2_X1 U5452 ( .A1(n6137), .A2(DATAI_20_), .ZN(n6377) );
  NAND2_X1 U5453 ( .A1(n6137), .A2(DATAI_28_), .ZN(n6463) );
  OAI22_X1 U5454 ( .A1(n6377), .A2(n4357), .B1(n4356), .B2(n6463), .ZN(n4350)
         );
  AOI21_X1 U5455 ( .B1(n6459), .B2(n4359), .A(n4350), .ZN(n4352) );
  NAND2_X1 U5456 ( .A1(n4360), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4351) );
  OAI211_X1 U5457 ( .C1(n4691), .C2(n4363), .A(n4352), .B(n4351), .ZN(U3064)
         );
  NOR2_X2 U5458 ( .A1(n6084), .A2(n4353), .ZN(n6471) );
  INV_X1 U5459 ( .A(n6471), .ZN(n4685) );
  NOR2_X2 U5460 ( .A1(n4355), .A2(n4354), .ZN(n6470) );
  NAND2_X1 U5461 ( .A1(n6137), .A2(DATAI_22_), .ZN(n6474) );
  NAND2_X1 U5462 ( .A1(n6137), .A2(DATAI_30_), .ZN(n6423) );
  OAI22_X1 U5463 ( .A1(n6474), .A2(n4357), .B1(n4356), .B2(n6423), .ZN(n4358)
         );
  AOI21_X1 U5464 ( .B1(n6470), .B2(n4359), .A(n4358), .ZN(n4362) );
  NAND2_X1 U5465 ( .A1(n4360), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4361) );
  OAI211_X1 U5466 ( .C1(n4685), .C2(n4363), .A(n4362), .B(n4361), .ZN(U3066)
         );
  INV_X1 U5467 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U5468 ( .A1(n6460), .A2(n6510), .ZN(n4366) );
  OAI22_X1 U5469 ( .A1(n4368), .A2(n6377), .B1(n6463), .B2(n6485), .ZN(n4364)
         );
  AOI21_X1 U5470 ( .B1(n6459), .B2(n6508), .A(n4364), .ZN(n4365) );
  OAI211_X1 U5471 ( .C1(n6518), .C2(n4367), .A(n4366), .B(n4365), .ZN(U3128)
         );
  INV_X1 U5472 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5473 ( .A1(n6471), .A2(n6510), .ZN(n4371) );
  OAI22_X1 U5474 ( .A1(n4368), .A2(n6474), .B1(n6423), .B2(n6485), .ZN(n4369)
         );
  AOI21_X1 U5475 ( .B1(n6470), .B2(n6508), .A(n4369), .ZN(n4370) );
  OAI211_X1 U5476 ( .C1(n6518), .C2(n4372), .A(n4371), .B(n4370), .ZN(U3130)
         );
  INV_X1 U5477 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4376) );
  AOI22_X1 U5478 ( .A1(n6497), .A2(n4475), .B1(n6499), .B2(n6513), .ZN(n4373)
         );
  OAI21_X1 U5479 ( .B1(n6454), .B2(n4477), .A(n4373), .ZN(n4374) );
  AOI21_X1 U5480 ( .B1(n6496), .B2(n4479), .A(n4374), .ZN(n4375) );
  OAI21_X1 U5481 ( .B1(n4482), .B2(n4376), .A(n4375), .ZN(U3134) );
  NAND3_X1 U5482 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4495), .A3(n4378), .ZN(n6393) );
  NOR2_X1 U5483 ( .A1(n4487), .A2(n6393), .ZN(n4406) );
  AOI21_X1 U5484 ( .B1(n4379), .B2(n4767), .A(n4406), .ZN(n4385) );
  AOI21_X1 U5485 ( .B1(n4380), .B2(STATEBS16_REG_SCAN_IN), .A(n6439), .ZN(
        n4383) );
  AOI22_X1 U5486 ( .A1(n4385), .A2(n4383), .B1(n6439), .B2(n6393), .ZN(n4381)
         );
  NAND2_X1 U5487 ( .A1(n4382), .A2(n4381), .ZN(n4405) );
  INV_X1 U5488 ( .A(n4383), .ZN(n4384) );
  OAI22_X1 U5489 ( .A1(n4385), .A2(n4384), .B1(n6442), .B2(n6393), .ZN(n4404)
         );
  AOI22_X1 U5490 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4405), .B1(n6511), 
        .B2(n4404), .ZN(n4388) );
  AOI22_X1 U5491 ( .A1(n4406), .A2(n6509), .B1(n6426), .B2(n6514), .ZN(n4387)
         );
  OAI211_X1 U5492 ( .C1(n4625), .C2(n6482), .A(n4388), .B(n4387), .ZN(U3099)
         );
  AOI22_X1 U5493 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4405), .B1(n6491), 
        .B2(n4404), .ZN(n4390) );
  AOI22_X1 U5494 ( .A1(n4406), .A2(n6490), .B1(n6426), .B2(n6493), .ZN(n4389)
         );
  OAI211_X1 U5495 ( .C1(n4625), .C2(n6451), .A(n4390), .B(n4389), .ZN(U3093)
         );
  AOI22_X1 U5496 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4405), .B1(n6455), 
        .B2(n4404), .ZN(n4392) );
  AOI22_X1 U5497 ( .A1(n4406), .A2(n6945), .B1(n6426), .B2(n6946), .ZN(n4391)
         );
  OAI211_X1 U5498 ( .C1(n4625), .C2(n6951), .A(n4392), .B(n4391), .ZN(U3095)
         );
  AOI22_X1 U5499 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4405), .B1(n6484), 
        .B2(n4404), .ZN(n4394) );
  AOI22_X1 U5500 ( .A1(n6483), .A2(n4406), .B1(n6426), .B2(n6487), .ZN(n4393)
         );
  OAI211_X1 U5501 ( .C1(n6448), .C2(n4625), .A(n4394), .B(n4393), .ZN(U3092)
         );
  AOI22_X1 U5502 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4405), .B1(n6496), 
        .B2(n4404), .ZN(n4396) );
  AOI22_X1 U5503 ( .A1(n6497), .A2(n4406), .B1(n6426), .B2(n6499), .ZN(n4395)
         );
  OAI211_X1 U5504 ( .C1(n4625), .C2(n6454), .A(n4396), .B(n4395), .ZN(U3094)
         );
  NAND2_X1 U5505 ( .A1(n4333), .A2(n4397), .ZN(n4398) );
  AND2_X1 U5506 ( .A1(n4483), .A2(n4398), .ZN(n5933) );
  INV_X1 U5507 ( .A(n5933), .ZN(n4639) );
  AOI22_X1 U5508 ( .A1(n5535), .A2(DATAI_7_), .B1(n6005), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4399) );
  OAI21_X1 U5509 ( .B1(n4639), .B2(n5796), .A(n4399), .ZN(U2884) );
  AOI22_X1 U5510 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4405), .B1(n6503), 
        .B2(n4404), .ZN(n4401) );
  INV_X1 U5511 ( .A(n6468), .ZN(n6505) );
  AOI22_X1 U5512 ( .A1(n4406), .A2(n6502), .B1(n6426), .B2(n6505), .ZN(n4400)
         );
  OAI211_X1 U5513 ( .C1(n4625), .C2(n6380), .A(n4401), .B(n4400), .ZN(U3097)
         );
  AOI22_X1 U5514 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4405), .B1(n6460), 
        .B2(n4404), .ZN(n4403) );
  INV_X1 U5515 ( .A(n6463), .ZN(n6374) );
  AOI22_X1 U5516 ( .A1(n4406), .A2(n6459), .B1(n6426), .B2(n6374), .ZN(n4402)
         );
  OAI211_X1 U5517 ( .C1(n4625), .C2(n6377), .A(n4403), .B(n4402), .ZN(U3096)
         );
  AOI22_X1 U5518 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4405), .B1(n6471), 
        .B2(n4404), .ZN(n4408) );
  INV_X1 U5519 ( .A(n6423), .ZN(n6469) );
  AOI22_X1 U5520 ( .A1(n4406), .A2(n6470), .B1(n6426), .B2(n6469), .ZN(n4407)
         );
  OAI211_X1 U5521 ( .C1(n4625), .C2(n6474), .A(n4408), .B(n4407), .ZN(U3098)
         );
  AOI22_X1 U5522 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4414), .B1(n6503), 
        .B2(n4413), .ZN(n4410) );
  AOI22_X1 U5523 ( .A1(n6505), .A2(n4447), .B1(n6502), .B2(n4415), .ZN(n4409)
         );
  OAI211_X1 U5524 ( .C1(n6380), .C2(n4595), .A(n4410), .B(n4409), .ZN(U3033)
         );
  AOI22_X1 U5525 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4414), .B1(n6460), 
        .B2(n4413), .ZN(n4412) );
  AOI22_X1 U5526 ( .A1(n6374), .A2(n4447), .B1(n6459), .B2(n4415), .ZN(n4411)
         );
  OAI211_X1 U5527 ( .C1(n6377), .C2(n4595), .A(n4412), .B(n4411), .ZN(U3032)
         );
  AOI22_X1 U5528 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4414), .B1(n6471), 
        .B2(n4413), .ZN(n4417) );
  AOI22_X1 U5529 ( .A1(n6469), .A2(n4447), .B1(n6470), .B2(n4415), .ZN(n4416)
         );
  OAI211_X1 U5530 ( .C1(n6474), .C2(n4595), .A(n4417), .B(n4416), .ZN(U3034)
         );
  INV_X1 U5531 ( .A(n4418), .ZN(n4419) );
  NAND3_X1 U5532 ( .A1(n4420), .A2(n5189), .A3(n4419), .ZN(n4421) );
  OAI21_X4 U5533 ( .B1(n4422), .B2(n6520), .A(n4421), .ZN(n5525) );
  NAND2_X2 U5534 ( .A1(n5525), .A2(n5161), .ZN(n5515) );
  OAI21_X1 U5535 ( .B1(n4711), .B2(n4707), .A(n4423), .ZN(n4424) );
  AND2_X1 U5536 ( .A1(n4424), .A2(n4428), .ZN(n6195) );
  INV_X1 U5537 ( .A(n6195), .ZN(n4425) );
  OAI222_X1 U5538 ( .A1(n4427), .A2(n5515), .B1(n5525), .B2(n4426), .C1(n4425), 
        .C2(n5516), .ZN(U2855) );
  INV_X1 U5539 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4433) );
  INV_X1 U5540 ( .A(n4428), .ZN(n4431) );
  AOI21_X1 U5541 ( .B1(n4431), .B2(n4430), .A(n4429), .ZN(n4432) );
  OR2_X1 U5542 ( .A1(n4432), .A2(n4552), .ZN(n5943) );
  OAI222_X1 U5543 ( .A1(n5944), .A2(n5515), .B1(n5525), .B2(n4433), .C1(n5943), 
        .C2(n5516), .ZN(U2853) );
  INV_X1 U5544 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4438) );
  INV_X1 U5545 ( .A(n6474), .ZN(n6420) );
  INV_X1 U5546 ( .A(n6470), .ZN(n4434) );
  OAI22_X1 U5547 ( .A1(n4434), .A2(n4444), .B1(n6423), .B2(n6950), .ZN(n4435)
         );
  AOI21_X1 U5548 ( .B1(n6420), .B2(n4447), .A(n4435), .ZN(n4437) );
  NAND2_X1 U5549 ( .A1(n6471), .A2(n4448), .ZN(n4436) );
  OAI211_X1 U5550 ( .C1(n4451), .C2(n4438), .A(n4437), .B(n4436), .ZN(U3026)
         );
  INV_X1 U5551 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4443) );
  INV_X1 U5552 ( .A(n6380), .ZN(n6504) );
  INV_X1 U5553 ( .A(n6502), .ZN(n4439) );
  OAI22_X1 U5554 ( .A1(n4439), .A2(n4444), .B1(n6468), .B2(n6950), .ZN(n4440)
         );
  AOI21_X1 U5555 ( .B1(n6504), .B2(n4447), .A(n4440), .ZN(n4442) );
  NAND2_X1 U5556 ( .A1(n6503), .A2(n4448), .ZN(n4441) );
  OAI211_X1 U5557 ( .C1(n4451), .C2(n4443), .A(n4442), .B(n4441), .ZN(U3025)
         );
  INV_X1 U5558 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n6830) );
  INV_X1 U5559 ( .A(n6377), .ZN(n6458) );
  INV_X1 U5560 ( .A(n6459), .ZN(n4445) );
  OAI22_X1 U5561 ( .A1(n4445), .A2(n4444), .B1(n6463), .B2(n6950), .ZN(n4446)
         );
  AOI21_X1 U5562 ( .B1(n6458), .B2(n4447), .A(n4446), .ZN(n4450) );
  NAND2_X1 U5563 ( .A1(n6460), .A2(n4448), .ZN(n4449) );
  OAI211_X1 U5564 ( .C1(n4451), .C2(n6830), .A(n4450), .B(n4449), .ZN(U3024)
         );
  NAND2_X1 U5565 ( .A1(n6502), .A2(n6944), .ZN(n4453) );
  NAND2_X1 U5566 ( .A1(n6947), .A2(n6505), .ZN(n4452) );
  OAI211_X1 U5567 ( .C1(n6950), .C2(n6380), .A(n4453), .B(n4452), .ZN(n4455)
         );
  NOR2_X1 U5568 ( .A1(n4682), .A2(n6952), .ZN(n4454) );
  AOI211_X1 U5569 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n6956), .A(n4455), 
        .B(n4454), .ZN(n4456) );
  INV_X1 U5570 ( .A(n4456), .ZN(U3145) );
  NAND2_X1 U5571 ( .A1(n6459), .A2(n6944), .ZN(n4458) );
  NAND2_X1 U5572 ( .A1(n6947), .A2(n6374), .ZN(n4457) );
  OAI211_X1 U5573 ( .C1(n6950), .C2(n6377), .A(n4458), .B(n4457), .ZN(n4460)
         );
  NOR2_X1 U5574 ( .A1(n4691), .A2(n6952), .ZN(n4459) );
  AOI211_X1 U5575 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n6956), .A(n4460), 
        .B(n4459), .ZN(n4461) );
  INV_X1 U5576 ( .A(n4461), .ZN(U3144) );
  NAND2_X1 U5577 ( .A1(n6470), .A2(n6944), .ZN(n4463) );
  NAND2_X1 U5578 ( .A1(n6947), .A2(n6469), .ZN(n4462) );
  OAI211_X1 U5579 ( .C1(n6950), .C2(n6474), .A(n4463), .B(n4462), .ZN(n4465)
         );
  NOR2_X1 U5580 ( .A1(n4685), .A2(n6952), .ZN(n4464) );
  AOI211_X1 U5581 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n6956), .A(n4465), 
        .B(n4464), .ZN(n4466) );
  INV_X1 U5582 ( .A(n4466), .ZN(U3146) );
  INV_X1 U5583 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4470) );
  AOI22_X1 U5584 ( .A1(n6502), .A2(n4475), .B1(n6505), .B2(n6513), .ZN(n4467)
         );
  OAI21_X1 U5585 ( .B1(n6380), .B2(n4477), .A(n4467), .ZN(n4468) );
  AOI21_X1 U5586 ( .B1(n6503), .B2(n4479), .A(n4468), .ZN(n4469) );
  OAI21_X1 U5587 ( .B1(n4482), .B2(n4470), .A(n4469), .ZN(U3137) );
  INV_X1 U5588 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4474) );
  AOI22_X1 U5589 ( .A1(n6459), .A2(n4475), .B1(n6374), .B2(n6513), .ZN(n4471)
         );
  OAI21_X1 U5590 ( .B1(n6377), .B2(n4477), .A(n4471), .ZN(n4472) );
  AOI21_X1 U5591 ( .B1(n6460), .B2(n4479), .A(n4472), .ZN(n4473) );
  OAI21_X1 U5592 ( .B1(n4482), .B2(n4474), .A(n4473), .ZN(U3136) );
  INV_X1 U5593 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U5594 ( .A1(n6470), .A2(n4475), .B1(n6469), .B2(n6513), .ZN(n4476)
         );
  OAI21_X1 U5595 ( .B1(n6474), .B2(n4477), .A(n4476), .ZN(n4478) );
  AOI21_X1 U5596 ( .B1(n6471), .B2(n4479), .A(n4478), .ZN(n4480) );
  OAI21_X1 U5597 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(U3138) );
  XOR2_X1 U5598 ( .A(n4484), .B(n4483), .Z(n4662) );
  AOI22_X1 U5599 ( .A1(n5535), .A2(DATAI_8_), .B1(n6005), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4485) );
  OAI21_X1 U5600 ( .B1(n4745), .B2(n5796), .A(n4485), .ZN(U2883) );
  AOI211_X1 U5601 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n4488), .A(n4487), .B(n4486), .ZN(n4492) );
  INV_X1 U5602 ( .A(n4489), .ZN(n4490) );
  OAI22_X1 U5603 ( .A1(n4492), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n4491), .B2(n4490), .ZN(n4494) );
  NAND2_X1 U5604 ( .A1(n4492), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4493) );
  OAI211_X1 U5605 ( .C1(n4496), .C2(n4495), .A(n4494), .B(n4493), .ZN(n4499)
         );
  NAND2_X1 U5606 ( .A1(n4496), .A2(n4495), .ZN(n4498) );
  INV_X1 U5607 ( .A(n4501), .ZN(n4497) );
  AOI22_X1 U5608 ( .A1(n4499), .A2(n4498), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n4497), .ZN(n4500) );
  AOI21_X1 U5609 ( .B1(n6320), .B2(n4501), .A(n4500), .ZN(n4512) );
  INV_X1 U5610 ( .A(n4502), .ZN(n4511) );
  INV_X1 U5611 ( .A(n4503), .ZN(n4509) );
  INV_X1 U5612 ( .A(n4504), .ZN(n4508) );
  AOI21_X1 U5613 ( .B1(n6781), .B2(n6826), .A(n4505), .ZN(n4507) );
  NOR4_X1 U5614 ( .A1(n4509), .A2(n4508), .A3(n4507), .A4(n4506), .ZN(n4510)
         );
  OAI211_X1 U5615 ( .C1(n4512), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n4511), .B(n4510), .ZN(n4519) );
  INV_X1 U5616 ( .A(n4513), .ZN(n4516) );
  NOR3_X1 U5617 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6442), .A3(n6617), .ZN(
        n4514) );
  OAI22_X1 U5618 ( .A1(n5747), .A2(n4516), .B1(n4515), .B2(n4514), .ZN(n6526)
         );
  AOI221_X1 U5619 ( .B1(n6708), .B2(n6765), .C1(n6708), .C2(n4519), .A(n6526), 
        .ZN(n6602) );
  INV_X1 U5620 ( .A(n6602), .ZN(n4520) );
  AOI221_X1 U5621 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4520), .C1(n6617), .C2(
        n4520), .A(n6765), .ZN(n6524) );
  AOI211_X1 U5622 ( .C1(n4519), .C2(n4518), .A(n4517), .B(n6524), .ZN(n4526)
         );
  OAI21_X1 U5623 ( .B1(n6621), .B2(n4521), .A(n4520), .ZN(n4524) );
  INV_X1 U5624 ( .A(n4522), .ZN(n4523) );
  MUX2_X1 U5625 ( .A(n4524), .B(n4523), .S(STATE2_REG_0__SCAN_IN), .Z(n4525)
         );
  NAND2_X1 U5626 ( .A1(n4526), .A2(n4525), .ZN(U3148) );
  NAND2_X1 U5627 ( .A1(n4527), .A2(n4538), .ZN(n4531) );
  INV_X1 U5628 ( .A(n4542), .ZN(n4528) );
  NAND2_X1 U5629 ( .A1(n4528), .A2(n4541), .ZN(n4654) );
  XNOR2_X1 U5630 ( .A(n4654), .B(n4655), .ZN(n4529) );
  NAND2_X1 U5631 ( .A1(n4529), .A2(n4656), .ZN(n4530) );
  NAND2_X1 U5632 ( .A1(n4531), .A2(n4530), .ZN(n4640) );
  XNOR2_X1 U5633 ( .A(n4640), .B(n4699), .ZN(n4644) );
  NAND2_X1 U5634 ( .A1(n4533), .A2(n4532), .ZN(n4536) );
  NAND2_X1 U5635 ( .A1(n4534), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4535)
         );
  NAND2_X1 U5636 ( .A1(n4536), .A2(n4535), .ZN(n4723) );
  NAND2_X1 U5637 ( .A1(n4653), .A2(n4540), .ZN(n4545) );
  XNOR2_X1 U5638 ( .A(n4542), .B(n4541), .ZN(n4543) );
  NAND2_X1 U5639 ( .A1(n4543), .A2(n4656), .ZN(n4544) );
  NAND2_X1 U5640 ( .A1(n4545), .A2(n4544), .ZN(n4546) );
  INV_X1 U5641 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6189) );
  XNOR2_X1 U5642 ( .A(n4546), .B(n6189), .ZN(n4725) );
  NAND2_X1 U5643 ( .A1(n4723), .A2(n4725), .ZN(n4643) );
  NAND2_X1 U5644 ( .A1(n4546), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4641)
         );
  NAND2_X1 U5645 ( .A1(n4643), .A2(n4641), .ZN(n4547) );
  XNOR2_X1 U5646 ( .A(n4644), .B(n4547), .ZN(n4672) );
  NAND3_X1 U5647 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4548), .ZN(n4891) );
  INV_X1 U5648 ( .A(n5711), .ZN(n6221) );
  NOR2_X1 U5649 ( .A1(n6221), .A2(n4549), .ZN(n5704) );
  INV_X1 U5650 ( .A(n5704), .ZN(n4896) );
  NAND3_X1 U5651 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4550), .ZN(n4889) );
  AOI22_X1 U5652 ( .A1(n5708), .A2(n4891), .B1(n4896), .B2(n4889), .ZN(n4701)
         );
  INV_X1 U5653 ( .A(n4701), .ZN(n6175) );
  NOR2_X1 U5654 ( .A1(n4552), .A2(n4551), .ZN(n4553) );
  OR2_X1 U5655 ( .A1(n4735), .A2(n4553), .ZN(n5928) );
  NAND2_X1 U5656 ( .A1(n6229), .A2(REIP_REG_7__SCAN_IN), .ZN(n4669) );
  OAI21_X1 U5657 ( .B1(n6218), .B2(n5326), .A(n5711), .ZN(n6192) );
  NAND2_X1 U5658 ( .A1(n4554), .A2(n6192), .ZN(n6185) );
  NOR2_X1 U5659 ( .A1(n6189), .A2(n6185), .ZN(n6171) );
  NAND2_X1 U5660 ( .A1(n4699), .A2(n6171), .ZN(n4555) );
  OAI211_X1 U5661 ( .C1(n5928), .C2(n6207), .A(n4669), .B(n4555), .ZN(n4556)
         );
  AOI21_X1 U5662 ( .B1(n6175), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4556), 
        .ZN(n4557) );
  OAI21_X1 U5663 ( .B1(n6196), .B2(n4672), .A(n4557), .ZN(U3011) );
  INV_X1 U5664 ( .A(n4595), .ZN(n4559) );
  NOR2_X1 U5665 ( .A1(n4559), .A2(n6280), .ZN(n4560) );
  NAND2_X1 U5666 ( .A1(n4011), .A2(n5983), .ZN(n4617) );
  OAI22_X1 U5667 ( .A1(n4560), .A2(n6326), .B1(n4767), .B2(n4617), .ZN(n4561)
         );
  NAND2_X1 U5668 ( .A1(n4619), .A2(n6320), .ZN(n6263) );
  NOR2_X1 U5669 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6263), .ZN(n4593)
         );
  AOI21_X1 U5670 ( .B1(n4561), .B2(n6397), .A(n4593), .ZN(n4564) );
  AOI21_X1 U5671 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(
        STATE2_REG_2__SCAN_IN), .A(n4562), .ZN(n6331) );
  INV_X1 U5672 ( .A(n6331), .ZN(n4563) );
  INV_X1 U5673 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4569) );
  NAND3_X1 U5674 ( .A1(n6328), .A2(n6321), .A3(n6320), .ZN(n4565) );
  OAI21_X1 U5675 ( .B1(n6400), .B2(n4617), .A(n4565), .ZN(n4597) );
  AOI22_X1 U5676 ( .A1(n6483), .A2(n4593), .B1(n6486), .B2(n6280), .ZN(n4566)
         );
  OAI21_X1 U5677 ( .B1(n6405), .B2(n4595), .A(n4566), .ZN(n4567) );
  AOI21_X1 U5678 ( .B1(n6484), .B2(n4597), .A(n4567), .ZN(n4568) );
  OAI21_X1 U5679 ( .B1(n4600), .B2(n4569), .A(n4568), .ZN(U3036) );
  INV_X1 U5680 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4573) );
  AOI22_X1 U5681 ( .A1(n6470), .A2(n4593), .B1(n6420), .B2(n6280), .ZN(n4570)
         );
  OAI21_X1 U5682 ( .B1(n6423), .B2(n4595), .A(n4570), .ZN(n4571) );
  AOI21_X1 U5683 ( .B1(n6471), .B2(n4597), .A(n4571), .ZN(n4572) );
  OAI21_X1 U5684 ( .B1(n4600), .B2(n4573), .A(n4572), .ZN(U3042) );
  INV_X1 U5685 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6909) );
  AOI22_X1 U5686 ( .A1(n6509), .A2(n4593), .B1(n6512), .B2(n6280), .ZN(n4574)
         );
  OAI21_X1 U5687 ( .B1(n6430), .B2(n4595), .A(n4574), .ZN(n4575) );
  AOI21_X1 U5688 ( .B1(n6511), .B2(n4597), .A(n4575), .ZN(n4576) );
  OAI21_X1 U5689 ( .B1(n4600), .B2(n6909), .A(n4576), .ZN(U3043) );
  INV_X1 U5690 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5691 ( .A1(n6490), .A2(n4593), .B1(n6492), .B2(n6280), .ZN(n4577)
         );
  OAI21_X1 U5692 ( .B1(n6408), .B2(n4595), .A(n4577), .ZN(n4578) );
  AOI21_X1 U5693 ( .B1(n6491), .B2(n4597), .A(n4578), .ZN(n4579) );
  OAI21_X1 U5694 ( .B1(n4600), .B2(n4580), .A(n4579), .ZN(U3037) );
  INV_X1 U5695 ( .A(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U5696 ( .A1(n6497), .A2(n4593), .B1(n6498), .B2(n6280), .ZN(n4581)
         );
  OAI21_X1 U5697 ( .B1(n6411), .B2(n4595), .A(n4581), .ZN(n4582) );
  AOI21_X1 U5698 ( .B1(n6496), .B2(n4597), .A(n4582), .ZN(n4583) );
  OAI21_X1 U5699 ( .B1(n4600), .B2(n4584), .A(n4583), .ZN(U3038) );
  INV_X1 U5700 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4588) );
  AOI22_X1 U5701 ( .A1(n6459), .A2(n4593), .B1(n6458), .B2(n6280), .ZN(n4585)
         );
  OAI21_X1 U5702 ( .B1(n6463), .B2(n4595), .A(n4585), .ZN(n4586) );
  AOI21_X1 U5703 ( .B1(n6460), .B2(n4597), .A(n4586), .ZN(n4587) );
  OAI21_X1 U5704 ( .B1(n4600), .B2(n4588), .A(n4587), .ZN(U3040) );
  INV_X1 U5705 ( .A(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4592) );
  AOI22_X1 U5706 ( .A1(n6502), .A2(n4593), .B1(n6504), .B2(n6280), .ZN(n4589)
         );
  OAI21_X1 U5707 ( .B1(n6468), .B2(n4595), .A(n4589), .ZN(n4590) );
  AOI21_X1 U5708 ( .B1(n6503), .B2(n4597), .A(n4590), .ZN(n4591) );
  OAI21_X1 U5709 ( .B1(n4600), .B2(n4592), .A(n4591), .ZN(U3041) );
  INV_X1 U5710 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5711 ( .A1(n6945), .A2(n4593), .B1(n6412), .B2(n6280), .ZN(n4594)
         );
  OAI21_X1 U5712 ( .B1(n6415), .B2(n4595), .A(n4594), .ZN(n4596) );
  AOI21_X1 U5713 ( .B1(n6455), .B2(n4597), .A(n4596), .ZN(n4598) );
  OAI21_X1 U5714 ( .B1(n4600), .B2(n4599), .A(n4598), .ZN(U3039) );
  XNOR2_X1 U5715 ( .A(n4601), .B(n4602), .ZN(n6197) );
  AND2_X1 U5716 ( .A1(n6229), .A2(REIP_REG_4__SCAN_IN), .ZN(n6194) );
  AOI21_X1 U5717 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6194), 
        .ZN(n4604) );
  OAI21_X1 U5718 ( .B1(n6140), .B2(n5978), .A(n4604), .ZN(n4605) );
  AOI21_X1 U5719 ( .B1(n5974), .B2(n6137), .A(n4605), .ZN(n4606) );
  OAI21_X1 U5720 ( .B1(n6121), .B2(n6197), .A(n4606), .ZN(U2982) );
  INV_X1 U5721 ( .A(n4607), .ZN(n4608) );
  XNOR2_X1 U5722 ( .A(n4609), .B(n4608), .ZN(n6209) );
  INV_X1 U5723 ( .A(n6209), .ZN(n4614) );
  INV_X1 U5724 ( .A(n4819), .ZN(n4612) );
  AOI22_X1 U5725 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n4610) );
  OAI21_X1 U5726 ( .B1(n6140), .B2(n4812), .A(n4610), .ZN(n4611) );
  AOI21_X1 U5727 ( .B1(n4612), .B2(n6137), .A(n4611), .ZN(n4613) );
  OAI21_X1 U5728 ( .B1(n4614), .B2(n6121), .A(n4613), .ZN(U2983) );
  NOR2_X1 U5729 ( .A1(n6434), .A2(n6353), .ZN(n4615) );
  NAND2_X1 U5730 ( .A1(n4615), .A2(n6254), .ZN(n6467) );
  NAND2_X1 U5731 ( .A1(n4625), .A2(n6467), .ZN(n4616) );
  AOI21_X1 U5732 ( .B1(n4616), .B2(STATEBS16_REG_SCAN_IN), .A(n6439), .ZN(
        n4622) );
  INV_X1 U5733 ( .A(n4617), .ZN(n6257) );
  NOR2_X1 U5734 ( .A1(n6390), .A2(n6320), .ZN(n4618) );
  AOI22_X1 U5735 ( .A1(n4622), .A2(n6437), .B1(n6321), .B2(n4618), .ZN(n4692)
         );
  NAND2_X1 U5736 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4619), .ZN(n6443) );
  NOR2_X1 U5737 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6443), .ZN(n4687)
         );
  INV_X1 U5738 ( .A(n6437), .ZN(n4621) );
  INV_X1 U5739 ( .A(n4687), .ZN(n4620) );
  AOI22_X1 U5740 ( .A1(n4622), .A2(n4621), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n4620), .ZN(n4623) );
  NAND3_X1 U5741 ( .A1(n4624), .A2(n4623), .A3(n6288), .ZN(n4686) );
  AOI22_X1 U5742 ( .A1(n6490), .A2(n4687), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n4686), .ZN(n4627) );
  AOI22_X1 U5743 ( .A1(n4688), .A2(n6493), .B1(n6475), .B2(n6492), .ZN(n4626)
         );
  OAI211_X1 U5744 ( .C1(n4692), .C2(n4628), .A(n4627), .B(n4626), .ZN(U3101)
         );
  AOI22_X1 U5745 ( .A1(n6509), .A2(n4687), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n4686), .ZN(n4630) );
  AOI22_X1 U5746 ( .A1(n4688), .A2(n6514), .B1(n6475), .B2(n6512), .ZN(n4629)
         );
  OAI211_X1 U5747 ( .C1(n4692), .C2(n4631), .A(n4630), .B(n4629), .ZN(U3107)
         );
  INV_X1 U5748 ( .A(n5981), .ZN(n4632) );
  OAI21_X1 U5749 ( .B1(n5189), .B2(n4633), .A(n4632), .ZN(n6230) );
  AOI22_X1 U5750 ( .A1(n5480), .A2(n6230), .B1(n5479), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4634) );
  OAI21_X1 U5751 ( .B1(n5982), .B2(n5515), .A(n4634), .ZN(U2858) );
  AOI22_X1 U5752 ( .A1(n6945), .A2(n4687), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n4686), .ZN(n4636) );
  AOI22_X1 U5753 ( .A1(n4688), .A2(n6946), .B1(n6475), .B2(n6412), .ZN(n4635)
         );
  OAI211_X1 U5754 ( .C1(n4692), .C2(n6953), .A(n4636), .B(n4635), .ZN(U3103)
         );
  INV_X1 U5755 ( .A(n5928), .ZN(n4637) );
  AOI22_X1 U5756 ( .A1(n4637), .A2(n5480), .B1(n5479), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4638) );
  OAI21_X1 U5757 ( .B1(n4639), .B2(n5515), .A(n4638), .ZN(U2852) );
  NAND2_X1 U5758 ( .A1(n4640), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4645)
         );
  AND2_X1 U5759 ( .A1(n4641), .A2(n4645), .ZN(n4642) );
  NAND2_X1 U5760 ( .A1(n4643), .A2(n4642), .ZN(n4648) );
  INV_X1 U5761 ( .A(n4644), .ZN(n4646) );
  NAND2_X1 U5762 ( .A1(n4646), .A2(n4645), .ZN(n4647) );
  AND2_X2 U5763 ( .A1(n4648), .A2(n4647), .ZN(n4694) );
  INV_X1 U5764 ( .A(n4655), .ZN(n4649) );
  NOR3_X1 U5765 ( .A1(n4651), .A2(n4650), .A3(n4649), .ZN(n4652) );
  INV_X1 U5766 ( .A(n4654), .ZN(n4657) );
  NAND3_X1 U5767 ( .A1(n4657), .A2(n4656), .A3(n4655), .ZN(n4658) );
  NAND2_X1 U5768 ( .A1(n5257), .A2(n4658), .ZN(n4695) );
  INV_X1 U5769 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4700) );
  XNOR2_X1 U5770 ( .A(n4695), .B(n4700), .ZN(n4693) );
  INV_X1 U5771 ( .A(n4693), .ZN(n4659) );
  XNOR2_X1 U5772 ( .A(n4694), .B(n4659), .ZN(n6172) );
  INV_X1 U5773 ( .A(n6172), .ZN(n4664) );
  AOI22_X1 U5774 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4660) );
  OAI21_X1 U5775 ( .B1(n6140), .B2(n4733), .A(n4660), .ZN(n4661) );
  AOI21_X1 U5776 ( .B1(n4662), .B2(n6137), .A(n4661), .ZN(n4663) );
  OAI21_X1 U5777 ( .B1(n4664), .B2(n6121), .A(n4663), .ZN(U2978) );
  AOI22_X1 U5778 ( .A1(n6483), .A2(n4687), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n4686), .ZN(n4666) );
  AOI22_X1 U5779 ( .A1(n4688), .A2(n6487), .B1(n6475), .B2(n6486), .ZN(n4665)
         );
  OAI211_X1 U5780 ( .C1(n4692), .C2(n4667), .A(n4666), .B(n4665), .ZN(U3100)
         );
  NAND2_X1 U5781 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4668)
         );
  OAI211_X1 U5782 ( .C1(n6140), .C2(n5931), .A(n4669), .B(n4668), .ZN(n4670)
         );
  AOI21_X1 U5783 ( .B1(n5933), .B2(n6137), .A(n4670), .ZN(n4671) );
  OAI21_X1 U5784 ( .B1(n4672), .B2(n6121), .A(n4671), .ZN(U2979) );
  OAI21_X1 U5785 ( .B1(n4675), .B2(n4674), .A(n4673), .ZN(n5922) );
  AOI22_X1 U5786 ( .A1(n5535), .A2(DATAI_9_), .B1(n6005), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4676) );
  OAI21_X1 U5787 ( .B1(n5922), .B2(n5796), .A(n4676), .ZN(U2882) );
  AOI22_X1 U5788 ( .A1(n6497), .A2(n4687), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n4686), .ZN(n4678) );
  AOI22_X1 U5789 ( .A1(n4688), .A2(n6499), .B1(n6475), .B2(n6498), .ZN(n4677)
         );
  OAI211_X1 U5790 ( .C1(n4692), .C2(n4679), .A(n4678), .B(n4677), .ZN(U3102)
         );
  AOI22_X1 U5791 ( .A1(n6502), .A2(n4687), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n4686), .ZN(n4681) );
  AOI22_X1 U5792 ( .A1(n4688), .A2(n6505), .B1(n6475), .B2(n6504), .ZN(n4680)
         );
  OAI211_X1 U5793 ( .C1(n4692), .C2(n4682), .A(n4681), .B(n4680), .ZN(U3105)
         );
  AOI22_X1 U5794 ( .A1(n6470), .A2(n4687), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n4686), .ZN(n4684) );
  AOI22_X1 U5795 ( .A1(n4688), .A2(n6469), .B1(n6475), .B2(n6420), .ZN(n4683)
         );
  OAI211_X1 U5796 ( .C1(n4692), .C2(n4685), .A(n4684), .B(n4683), .ZN(U3106)
         );
  AOI22_X1 U5797 ( .A1(n6459), .A2(n4687), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n4686), .ZN(n4690) );
  AOI22_X1 U5798 ( .A1(n4688), .A2(n6374), .B1(n6475), .B2(n6458), .ZN(n4689)
         );
  OAI211_X1 U5799 ( .C1(n4692), .C2(n4691), .A(n4690), .B(n4689), .ZN(U3104)
         );
  NAND2_X1 U5800 ( .A1(n4694), .A2(n4693), .ZN(n4697) );
  NAND2_X1 U5801 ( .A1(n4695), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4696)
         );
  XNOR2_X1 U5802 ( .A(n5698), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4698)
         );
  XNOR2_X1 U5803 ( .A(n4867), .B(n4698), .ZN(n4843) );
  NOR2_X1 U5804 ( .A1(n4700), .A2(n4699), .ZN(n6180) );
  OAI21_X1 U5805 ( .B1(n5356), .B2(n6180), .A(n4701), .ZN(n6165) );
  NAND2_X1 U5806 ( .A1(n6180), .A2(n6171), .ZN(n6170) );
  INV_X1 U5807 ( .A(n4752), .ZN(n4702) );
  AOI21_X1 U5808 ( .B1(n4703), .B2(n4737), .A(n4702), .ZN(n5918) );
  NAND2_X1 U5809 ( .A1(n5918), .A2(n6247), .ZN(n4704) );
  NAND2_X1 U5810 ( .A1(n6229), .A2(REIP_REG_9__SCAN_IN), .ZN(n4838) );
  OAI211_X1 U5811 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6170), .A(n4704), 
        .B(n4838), .ZN(n4705) );
  AOI21_X1 U5812 ( .B1(n6165), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n4705), 
        .ZN(n4706) );
  OAI21_X1 U5813 ( .B1(n4843), .B2(n6196), .A(n4706), .ZN(U3009) );
  INV_X1 U5814 ( .A(n4707), .ZN(n4708) );
  XNOR2_X1 U5815 ( .A(n4711), .B(n4708), .ZN(n6204) );
  AOI22_X1 U5816 ( .A1(n5480), .A2(n6204), .B1(n5479), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4709) );
  OAI21_X1 U5817 ( .B1(n4819), .B2(n5515), .A(n4709), .ZN(U2856) );
  AOI22_X1 U5818 ( .A1(n5918), .A2(n5480), .B1(n5479), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n4710) );
  OAI21_X1 U5819 ( .B1(n5922), .B2(n5515), .A(n4710), .ZN(U2850) );
  OAI21_X1 U5820 ( .B1(n4713), .B2(n4712), .A(n4711), .ZN(n5466) );
  INV_X1 U5821 ( .A(n5466), .ZN(n6219) );
  AOI22_X1 U5822 ( .A1(n5480), .A2(n6219), .B1(n5479), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4714) );
  OAI21_X1 U5823 ( .B1(n4715), .B2(n5515), .A(n4714), .ZN(U2857) );
  INV_X1 U5824 ( .A(n5954), .ZN(n4717) );
  OAI222_X1 U5825 ( .A1(n5955), .A2(n5515), .B1(n5516), .B2(n4717), .C1(n4716), 
        .C2(n5525), .ZN(U2854) );
  OAI22_X1 U5826 ( .A1(n5616), .A2(n4718), .B1(n6205), .B2(n6553), .ZN(n4720)
         );
  NOR2_X1 U5827 ( .A1(n5955), .A2(n5617), .ZN(n4719) );
  AOI211_X1 U5828 ( .C1(n6117), .C2(n5956), .A(n4720), .B(n4719), .ZN(n4721)
         );
  OAI21_X1 U5829 ( .B1(n6121), .B2(n4722), .A(n4721), .ZN(U2981) );
  XOR2_X1 U5830 ( .A(n4725), .B(n4724), .Z(n6187) );
  NAND2_X1 U5831 ( .A1(n6187), .A2(n6135), .ZN(n4730) );
  INV_X1 U5832 ( .A(n5951), .ZN(n4728) );
  NAND2_X1 U5833 ( .A1(n6229), .A2(REIP_REG_6__SCAN_IN), .ZN(n6183) );
  OAI21_X1 U5834 ( .B1(n5616), .B2(n4726), .A(n6183), .ZN(n4727) );
  AOI21_X1 U5835 ( .B1(n4728), .B2(n6117), .A(n4727), .ZN(n4729) );
  OAI211_X1 U5836 ( .C1(n5617), .C2(n5944), .A(n4730), .B(n4729), .ZN(U2980)
         );
  OAI21_X1 U5837 ( .B1(n5967), .B2(n4731), .A(n6556), .ZN(n4741) );
  OAI21_X1 U5838 ( .B1(n5919), .B2(n5967), .A(n5934), .ZN(n5917) );
  NAND2_X1 U5839 ( .A1(n5969), .A2(EBX_REG_8__SCAN_IN), .ZN(n4732) );
  OAI211_X1 U5840 ( .C1(n5977), .C2(n4733), .A(n4732), .B(n5971), .ZN(n4740)
         );
  OR2_X1 U5841 ( .A1(n4735), .A2(n4734), .ZN(n4736) );
  NAND2_X1 U5842 ( .A1(n4737), .A2(n4736), .ZN(n6173) );
  OAI22_X1 U5843 ( .A1(n4738), .A2(n5989), .B1(n5929), .B2(n6173), .ZN(n4739)
         );
  AOI211_X1 U5844 ( .C1(n4741), .C2(n5917), .A(n4740), .B(n4739), .ZN(n4742)
         );
  OAI21_X1 U5845 ( .B1(n4745), .B2(n5753), .A(n4742), .ZN(U2819) );
  NOR2_X1 U5846 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4744)
         );
  OR2_X1 U5847 ( .A1(n4744), .A2(n4743), .ZN(n6242) );
  OAI222_X1 U5848 ( .A1(n5516), .A2(n6242), .B1(n5525), .B2(n3774), .C1(n5515), 
        .C2(n4833), .ZN(U2859) );
  INV_X1 U5849 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4746) );
  OAI222_X1 U5850 ( .A1(n6173), .A2(n5516), .B1(n5525), .B2(n4746), .C1(n5515), 
        .C2(n4745), .ZN(U2851) );
  INV_X1 U5851 ( .A(n4673), .ZN(n4749) );
  INV_X1 U5852 ( .A(n4747), .ZN(n4748) );
  OAI21_X1 U5853 ( .B1(n4749), .B2(n4748), .A(n4845), .ZN(n4828) );
  AOI22_X1 U5854 ( .A1(n5535), .A2(DATAI_10_), .B1(n6005), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4750) );
  OAI21_X1 U5855 ( .B1(n4828), .B2(n5796), .A(n4750), .ZN(U2881) );
  AND2_X1 U5856 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  OR2_X1 U5857 ( .A1(n4753), .A2(n4849), .ZN(n6162) );
  OAI22_X1 U5858 ( .A1(n5929), .A2(n6162), .B1(n4824), .B2(n5977), .ZN(n4758)
         );
  INV_X1 U5859 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6843) );
  INV_X1 U5860 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6559) );
  NOR2_X1 U5861 ( .A1(n6843), .A2(n6559), .ZN(n4756) );
  OAI211_X1 U5862 ( .C1(REIP_REG_9__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(
        n5919), .B(n5979), .ZN(n4755) );
  AOI22_X1 U5863 ( .A1(PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n5952), .B1(
        EBX_REG_10__SCAN_IN), .B2(n5969), .ZN(n4754) );
  OAI211_X1 U5864 ( .C1(n4756), .C2(n4755), .A(n4754), .B(n5971), .ZN(n4757)
         );
  AOI211_X1 U5865 ( .C1(n5917), .C2(REIP_REG_10__SCAN_IN), .A(n4758), .B(n4757), .ZN(n4759) );
  OAI21_X1 U5866 ( .B1(n4828), .B2(n5753), .A(n4759), .ZN(U2817) );
  NOR2_X1 U5867 ( .A1(n6434), .A2(n6318), .ZN(n4760) );
  NOR2_X1 U5868 ( .A1(n4761), .A2(n6321), .ZN(n4765) );
  INV_X1 U5869 ( .A(n4765), .ZN(n6389) );
  OAI21_X1 U5870 ( .B1(n6389), .B2(n6288), .A(n4762), .ZN(n4799) );
  NAND2_X1 U5871 ( .A1(n6496), .A2(n4799), .ZN(n4774) );
  NOR2_X1 U5872 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4763), .ZN(n4803)
         );
  INV_X1 U5873 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4771) );
  INV_X1 U5874 ( .A(n4803), .ZN(n4769) );
  OAI21_X1 U5875 ( .B1(n4765), .B2(n6442), .A(n4764), .ZN(n6394) );
  AOI21_X1 U5876 ( .B1(n6485), .B2(n6481), .A(n5861), .ZN(n4766) );
  AOI211_X1 U5877 ( .C1(n6286), .C2(n4767), .A(n4766), .B(n6439), .ZN(n4768)
         );
  AOI211_X1 U5878 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4769), .A(n6394), .B(
        n4768), .ZN(n4770) );
  OAI22_X1 U5879 ( .A1(n6485), .A2(n6454), .B1(n4771), .B2(n4800), .ZN(n4772)
         );
  AOI21_X1 U5880 ( .B1(n6497), .B2(n4803), .A(n4772), .ZN(n4773) );
  OAI211_X1 U5881 ( .C1(n6481), .C2(n6411), .A(n4774), .B(n4773), .ZN(U3118)
         );
  NAND2_X1 U5882 ( .A1(n6491), .A2(n4799), .ZN(n4778) );
  INV_X1 U5883 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4775) );
  OAI22_X1 U5884 ( .A1(n6485), .A2(n6451), .B1(n4775), .B2(n4800), .ZN(n4776)
         );
  AOI21_X1 U5885 ( .B1(n6490), .B2(n4803), .A(n4776), .ZN(n4777) );
  OAI211_X1 U5886 ( .C1(n6481), .C2(n6408), .A(n4778), .B(n4777), .ZN(U3117)
         );
  NAND2_X1 U5887 ( .A1(n6455), .A2(n4799), .ZN(n4782) );
  INV_X1 U5888 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5889 ( .A1(n6485), .A2(n6951), .B1(n4779), .B2(n4800), .ZN(n4780)
         );
  AOI21_X1 U5890 ( .B1(n6945), .B2(n4803), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5891 ( .C1(n6481), .C2(n6415), .A(n4782), .B(n4781), .ZN(U3119)
         );
  NAND2_X1 U5892 ( .A1(n6511), .A2(n4799), .ZN(n4786) );
  INV_X1 U5893 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4783) );
  OAI22_X1 U5894 ( .A1(n6485), .A2(n6482), .B1(n4783), .B2(n4800), .ZN(n4784)
         );
  AOI21_X1 U5895 ( .B1(n6509), .B2(n4803), .A(n4784), .ZN(n4785) );
  OAI211_X1 U5896 ( .C1(n6481), .C2(n6430), .A(n4786), .B(n4785), .ZN(U3123)
         );
  NAND2_X1 U5897 ( .A1(n6484), .A2(n4799), .ZN(n4790) );
  INV_X1 U5898 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4787) );
  OAI22_X1 U5899 ( .A1(n6485), .A2(n6448), .B1(n4787), .B2(n4800), .ZN(n4788)
         );
  AOI21_X1 U5900 ( .B1(n6483), .B2(n4803), .A(n4788), .ZN(n4789) );
  OAI211_X1 U5901 ( .C1(n6405), .C2(n6481), .A(n4790), .B(n4789), .ZN(U3116)
         );
  NAND2_X1 U5902 ( .A1(n6460), .A2(n4799), .ZN(n4794) );
  INV_X1 U5903 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4791) );
  OAI22_X1 U5904 ( .A1(n6485), .A2(n6377), .B1(n4791), .B2(n4800), .ZN(n4792)
         );
  AOI21_X1 U5905 ( .B1(n6459), .B2(n4803), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5906 ( .C1(n6481), .C2(n6463), .A(n4794), .B(n4793), .ZN(U3120)
         );
  NAND2_X1 U5907 ( .A1(n6471), .A2(n4799), .ZN(n4798) );
  INV_X1 U5908 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4795) );
  OAI22_X1 U5909 ( .A1(n6485), .A2(n6474), .B1(n4795), .B2(n4800), .ZN(n4796)
         );
  AOI21_X1 U5910 ( .B1(n6470), .B2(n4803), .A(n4796), .ZN(n4797) );
  OAI211_X1 U5911 ( .C1(n6481), .C2(n6423), .A(n4798), .B(n4797), .ZN(U3122)
         );
  NAND2_X1 U5912 ( .A1(n6503), .A2(n4799), .ZN(n4805) );
  INV_X1 U5913 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4801) );
  OAI22_X1 U5914 ( .A1(n6485), .A2(n6380), .B1(n4801), .B2(n4800), .ZN(n4802)
         );
  AOI21_X1 U5915 ( .B1(n6502), .B2(n4803), .A(n4802), .ZN(n4804) );
  OAI211_X1 U5916 ( .C1(n6481), .C2(n6468), .A(n4805), .B(n4804), .ZN(U3121)
         );
  NAND2_X1 U5917 ( .A1(n4809), .A2(n4806), .ZN(n4807) );
  NAND2_X1 U5918 ( .A1(n4807), .A2(n5753), .ZN(n5991) );
  INV_X1 U5919 ( .A(n5991), .ZN(n4834) );
  INV_X1 U5920 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6745) );
  INV_X1 U5921 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6548) );
  AOI211_X1 U5922 ( .C1(n5979), .C2(n6745), .A(n5985), .B(n6548), .ZN(n5467)
         );
  INV_X1 U5923 ( .A(n5966), .ZN(n4808) );
  OAI21_X1 U5924 ( .B1(n4808), .B2(n5967), .A(n5934), .ZN(n5964) );
  OAI21_X1 U5925 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5467), .A(n5964), .ZN(n4818)
         );
  INV_X1 U5926 ( .A(n4809), .ZN(n4811) );
  NOR2_X1 U5927 ( .A1(n4811), .A2(n4810), .ZN(n5984) );
  INV_X1 U5928 ( .A(n5984), .ZN(n4832) );
  INV_X1 U5929 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4813) );
  OAI22_X1 U5930 ( .A1(n4813), .A2(n5989), .B1(n5977), .B2(n4812), .ZN(n4814)
         );
  AOI21_X1 U5931 ( .B1(n5969), .B2(EBX_REG_3__SCAN_IN), .A(n4814), .ZN(n4815)
         );
  OAI21_X1 U5932 ( .B1(n6258), .B2(n4832), .A(n4815), .ZN(n4816) );
  AOI21_X1 U5933 ( .B1(n5965), .B2(n6204), .A(n4816), .ZN(n4817) );
  OAI211_X1 U5934 ( .C1(n4834), .C2(n4819), .A(n4818), .B(n4817), .ZN(U2824)
         );
  INV_X1 U5935 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4820) );
  OAI222_X1 U5936 ( .A1(n4828), .A2(n5515), .B1(n5525), .B2(n4820), .C1(n5516), 
        .C2(n6162), .ZN(U2849) );
  NOR2_X1 U5937 ( .A1(n5568), .A2(n6161), .ZN(n4869) );
  OR2_X1 U5938 ( .A1(n4867), .A2(n4869), .ZN(n4821) );
  NAND2_X1 U5939 ( .A1(n5698), .A2(n6161), .ZN(n4872) );
  NAND2_X1 U5940 ( .A1(n4821), .A2(n4872), .ZN(n4823) );
  INV_X1 U5941 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6160) );
  NOR2_X1 U5942 ( .A1(n5822), .A2(n6160), .ZN(n4868) );
  AND2_X1 U5943 ( .A1(n5822), .A2(n6160), .ZN(n4871) );
  NOR2_X1 U5944 ( .A1(n4868), .A2(n4871), .ZN(n4822) );
  XNOR2_X1 U5945 ( .A(n4823), .B(n4822), .ZN(n6166) );
  NAND2_X1 U5946 ( .A1(n6166), .A2(n6135), .ZN(n4827) );
  AND2_X1 U5947 ( .A1(n6229), .A2(REIP_REG_10__SCAN_IN), .ZN(n6163) );
  NOR2_X1 U5948 ( .A1(n6140), .A2(n4824), .ZN(n4825) );
  AOI211_X1 U5949 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6163), 
        .B(n4825), .ZN(n4826) );
  OAI211_X1 U5950 ( .C1(n5617), .C2(n4828), .A(n4827), .B(n4826), .ZN(U2976)
         );
  NAND2_X1 U5951 ( .A1(n5989), .A2(n5977), .ZN(n4829) );
  AOI22_X1 U5952 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n4829), .B1(n5969), 
        .B2(EBX_REG_0__SCAN_IN), .ZN(n4830) );
  OAI21_X1 U5953 ( .B1(n4832), .B2(n4831), .A(n4830), .ZN(n4836) );
  OAI22_X1 U5954 ( .A1(n5929), .A2(n6242), .B1(n4834), .B2(n4833), .ZN(n4835)
         );
  AOI211_X1 U5955 ( .C1(REIP_REG_0__SCAN_IN), .C2(n5395), .A(n4836), .B(n4835), 
        .ZN(n4837) );
  INV_X1 U5956 ( .A(n4837), .ZN(U2827) );
  INV_X1 U5957 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n4839) );
  OAI21_X1 U5958 ( .B1(n5616), .B2(n4839), .A(n4838), .ZN(n4841) );
  NOR2_X1 U5959 ( .A1(n5922), .A2(n5617), .ZN(n4840) );
  AOI211_X1 U5960 ( .C1(n6117), .C2(n5923), .A(n4841), .B(n4840), .ZN(n4842)
         );
  OAI21_X1 U5961 ( .B1(n4843), .B2(n6121), .A(n4842), .ZN(U2977) );
  INV_X1 U5962 ( .A(n4844), .ZN(n4855) );
  AOI21_X1 U5963 ( .B1(n4846), .B2(n4845), .A(n4844), .ZN(n6118) );
  INV_X1 U5964 ( .A(n6118), .ZN(n4853) );
  AOI22_X1 U5965 ( .A1(n5535), .A2(DATAI_11_), .B1(n6005), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4847) );
  OAI21_X1 U5966 ( .B1(n4853), .B2(n5796), .A(n4847), .ZN(U2880) );
  INV_X1 U5967 ( .A(n4848), .ZN(n4851) );
  INV_X1 U5968 ( .A(n4849), .ZN(n4850) );
  AOI21_X1 U5969 ( .B1(n4851), .B2(n4850), .A(n4857), .ZN(n6152) );
  AOI22_X1 U5970 ( .A1(n6152), .A2(n5480), .B1(n5479), .B2(EBX_REG_11__SCAN_IN), .ZN(n4852) );
  OAI21_X1 U5971 ( .B1(n4853), .B2(n5515), .A(n4852), .ZN(U2848) );
  XNOR2_X1 U5972 ( .A(n4855), .B(n4854), .ZN(n4883) );
  INV_X1 U5973 ( .A(n4879), .ZN(n4863) );
  OAI21_X1 U5974 ( .B1(n4857), .B2(n4856), .A(n5522), .ZN(n4858) );
  INV_X1 U5975 ( .A(n4858), .ZN(n6142) );
  OAI21_X1 U5976 ( .B1(n5910), .B2(n5967), .A(n5934), .ZN(n5909) );
  AOI22_X1 U5977 ( .A1(n5965), .A2(n6142), .B1(REIP_REG_12__SCAN_IN), .B2(
        n5909), .ZN(n4861) );
  NAND2_X1 U5978 ( .A1(n5979), .A2(n5910), .ZN(n4859) );
  NOR2_X1 U5979 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4859), .ZN(n5904) );
  AOI211_X1 U5980 ( .C1(n5969), .C2(EBX_REG_12__SCAN_IN), .A(n5953), .B(n5904), 
        .ZN(n4860) );
  OAI211_X1 U5981 ( .C1(n6891), .C2(n5989), .A(n4861), .B(n4860), .ZN(n4862)
         );
  AOI21_X1 U5982 ( .B1(n5986), .B2(n4863), .A(n4862), .ZN(n4864) );
  OAI21_X1 U5983 ( .B1(n4883), .B2(n5753), .A(n4864), .ZN(U2815) );
  AOI22_X1 U5984 ( .A1(n6142), .A2(n5480), .B1(n5479), .B2(EBX_REG_12__SCAN_IN), .ZN(n4865) );
  OAI21_X1 U5985 ( .B1(n4883), .B2(n5515), .A(n4865), .ZN(U2847) );
  AOI22_X1 U5986 ( .A1(n5535), .A2(DATAI_12_), .B1(n6005), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n4866) );
  OAI21_X1 U5987 ( .B1(n4883), .B2(n5796), .A(n4866), .ZN(U2879) );
  INV_X1 U5988 ( .A(n4867), .ZN(n4870) );
  NAND2_X1 U5989 ( .A1(n5698), .A2(n6156), .ZN(n6110) );
  INV_X1 U5990 ( .A(n4871), .ZN(n4873) );
  AND2_X1 U5991 ( .A1(n4873), .A2(n4872), .ZN(n6112) );
  AND2_X1 U5992 ( .A1(n6110), .A2(n6112), .ZN(n4874) );
  NAND2_X1 U5993 ( .A1(n6113), .A2(n4874), .ZN(n4875) );
  OR2_X1 U5994 ( .A1(n5822), .A2(n6156), .ZN(n6111) );
  INV_X1 U5995 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U5996 ( .A1(n5568), .A2(n6144), .ZN(n5622) );
  INV_X1 U5997 ( .A(n5622), .ZN(n4876) );
  NAND2_X1 U5998 ( .A1(n5698), .A2(n6144), .ZN(n5624) );
  NAND2_X1 U5999 ( .A1(n4876), .A2(n5624), .ZN(n4877) );
  XNOR2_X1 U6000 ( .A(n5623), .B(n4877), .ZN(n6147) );
  NAND2_X1 U6001 ( .A1(n6147), .A2(n6135), .ZN(n4882) );
  INV_X1 U6002 ( .A(REIP_REG_12__SCAN_IN), .ZN(n4878) );
  NOR2_X1 U6003 ( .A1(n6205), .A2(n4878), .ZN(n6141) );
  NOR2_X1 U6004 ( .A1(n6140), .A2(n4879), .ZN(n4880) );
  AOI211_X1 U6005 ( .C1(n6130), .C2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n6141), 
        .B(n4880), .ZN(n4881) );
  OAI211_X1 U6006 ( .C1(n4883), .C2(n5617), .A(n4882), .B(n4881), .ZN(U2974)
         );
  XNOR2_X1 U6007 ( .A(n5698), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5627)
         );
  INV_X1 U6008 ( .A(n5627), .ZN(n4884) );
  OR2_X1 U6009 ( .A1(n5622), .A2(n4884), .ZN(n4903) );
  OR2_X1 U6010 ( .A1(n5623), .A2(n4903), .ZN(n4885) );
  NAND2_X1 U6011 ( .A1(n5698), .A2(n4894), .ZN(n4905) );
  NAND2_X1 U6012 ( .A1(n5626), .A2(n4905), .ZN(n4887) );
  INV_X1 U6013 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6014 ( .A(n5698), .B(n5315), .ZN(n4886) );
  XNOR2_X1 U6015 ( .A(n4887), .B(n4886), .ZN(n5621) );
  AOI21_X1 U6016 ( .B1(n4888), .B2(n5524), .A(n5453), .ZN(n5888) );
  INV_X1 U6017 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6564) );
  NOR2_X1 U6018 ( .A1(n6205), .A2(n6564), .ZN(n4901) );
  NAND2_X1 U6020 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5850) );
  NAND3_X1 U6021 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6180), .ZN(n4890) );
  INV_X1 U6022 ( .A(n5705), .ZN(n4895) );
  NOR2_X1 U6023 ( .A1(n4891), .A2(n4890), .ZN(n5703) );
  INV_X1 U6024 ( .A(n5703), .ZN(n5851) );
  OR3_X1 U6025 ( .A1(n6243), .A2(n4892), .A3(n5851), .ZN(n4893) );
  AOI211_X1 U6026 ( .C1(n4895), .C2(n4893), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5850), .ZN(n5849) );
  NOR2_X1 U6027 ( .A1(n4894), .A2(n5850), .ZN(n5702) );
  INV_X1 U6028 ( .A(n5702), .ZN(n4917) );
  AOI22_X1 U6029 ( .A1(n5708), .A2(n5851), .B1(n4896), .B2(n4895), .ZN(n6151)
         );
  OAI21_X1 U6030 ( .B1(n5702), .B2(n6245), .A(n6151), .ZN(n4897) );
  AOI211_X1 U6031 ( .C1(n4898), .C2(n5850), .A(n5849), .B(n4897), .ZN(n5857)
         );
  OAI33_X1 U6032 ( .A1(1'b0), .A2(n5857), .A3(n5315), .B1(
        INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5687), .B3(n4917), .ZN(n4900)
         );
  AOI211_X1 U6033 ( .C1(n6247), .C2(n5888), .A(n4901), .B(n4900), .ZN(n4902)
         );
  OAI21_X1 U6034 ( .B1(n5621), .B2(n6196), .A(n4902), .ZN(U3004) );
  NOR2_X1 U6035 ( .A1(n5623), .A2(n4903), .ZN(n4910) );
  NAND2_X1 U6036 ( .A1(n5568), .A2(n5315), .ZN(n4904) );
  AND2_X1 U6037 ( .A1(n4905), .A2(n4904), .ZN(n5603) );
  INV_X1 U6038 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6914) );
  AND2_X1 U6039 ( .A1(n5822), .A2(n6914), .ZN(n5606) );
  INV_X1 U6040 ( .A(n5606), .ZN(n4906) );
  AND2_X1 U6041 ( .A1(n5603), .A2(n4906), .ZN(n4908) );
  NAND2_X1 U6042 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  NOR2_X1 U6043 ( .A1(n4910), .A2(n4909), .ZN(n4911) );
  NOR2_X1 U6044 ( .A1(n4911), .A2(n3112), .ZN(n4912) );
  NAND2_X2 U6045 ( .A1(n4912), .A2(n5605), .ZN(n5819) );
  INV_X1 U6046 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6047 ( .A1(n5568), .A2(n5730), .ZN(n4913) );
  NOR2_X1 U6048 ( .A1(n5568), .A2(n5730), .ZN(n4916) );
  INV_X1 U6049 ( .A(n4913), .ZN(n4914) );
  NOR2_X1 U6050 ( .A1(n4916), .A2(n4914), .ZN(n4915) );
  OAI22_X1 U6051 ( .A1(n5821), .A2(n4916), .B1(n4915), .B2(n5819), .ZN(n5602)
         );
  NAND3_X1 U6052 ( .A1(n5702), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6155), .ZN(n4920) );
  NOR2_X1 U6053 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n4920), .ZN(n5845)
         );
  NOR2_X1 U6054 ( .A1(n5315), .A2(n4917), .ZN(n4918) );
  OAI21_X1 U6055 ( .B1(n5356), .B2(n4918), .A(n6151), .ZN(n5842) );
  OAI21_X1 U6056 ( .B1(n5845), .B2(n5842), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n4919) );
  INV_X1 U6057 ( .A(n4919), .ZN(n4925) );
  NOR3_X1 U6058 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n6914), .A3(n4920), 
        .ZN(n4924) );
  NAND2_X1 U6059 ( .A1(n5455), .A2(n4921), .ZN(n4922) );
  NAND2_X1 U6060 ( .A1(n5508), .A2(n4922), .ZN(n5514) );
  INV_X1 U6061 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6731) );
  OAI22_X1 U6062 ( .A1(n5514), .A2(n6207), .B1(n6731), .B2(n6205), .ZN(n4923)
         );
  NOR3_X1 U6063 ( .A1(n4925), .A2(n4924), .A3(n4923), .ZN(n4926) );
  OAI21_X1 U6064 ( .B1(n5602), .B2(n6196), .A(n4926), .ZN(U3002) );
  OAI21_X1 U6065 ( .B1(n4929), .B2(n4928), .A(n4927), .ZN(n5889) );
  AOI22_X1 U6066 ( .A1(n5888), .A2(n5480), .B1(EBX_REG_14__SCAN_IN), .B2(n5479), .ZN(n4930) );
  OAI21_X1 U6067 ( .B1(n5889), .B2(n5515), .A(n4930), .ZN(U2845) );
  AOI22_X1 U6068 ( .A1(n5535), .A2(DATAI_14_), .B1(n6005), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4931) );
  OAI21_X1 U6069 ( .B1(n5889), .B2(n5796), .A(n4931), .ZN(U2877) );
  INV_X1 U6070 ( .A(n5821), .ZN(n4932) );
  NAND2_X1 U6071 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6072 ( .A1(n4932), .A2(n3115), .ZN(n5260) );
  NAND2_X1 U6073 ( .A1(n5820), .A2(n5730), .ZN(n5818) );
  OAI21_X1 U6074 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5818), .A(n5731), 
        .ZN(n4933) );
  NAND2_X2 U6075 ( .A1(n5260), .A2(n4933), .ZN(n5588) );
  AND2_X1 U6076 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5323) );
  INV_X1 U6077 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6742) );
  INV_X1 U6078 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5713) );
  NOR2_X1 U6079 ( .A1(n6742), .A2(n5713), .ZN(n5712) );
  NAND2_X1 U6080 ( .A1(n5323), .A2(n5712), .ZN(n5316) );
  NAND2_X1 U6081 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5327) );
  NOR2_X1 U6082 ( .A1(n5316), .A2(n5327), .ZN(n4934) );
  NOR2_X1 U6083 ( .A1(n5568), .A2(n6742), .ZN(n5585) );
  AOI21_X1 U6084 ( .B1(n5588), .B2(n4934), .A(n5585), .ZN(n4938) );
  NOR2_X1 U6085 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4935) );
  INV_X1 U6086 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5684) );
  NAND4_X1 U6087 ( .A1(n4935), .A2(n5557), .A3(n5684), .A4(n5713), .ZN(n4936)
         );
  OAI21_X1 U6088 ( .B1(n5588), .B2(n4936), .A(n5731), .ZN(n4937) );
  AND2_X2 U6089 ( .A1(n4938), .A2(n4937), .ZN(n5549) );
  XNOR2_X1 U6090 ( .A(n5698), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5550)
         );
  NAND2_X2 U6091 ( .A1(n5549), .A2(n5550), .ZN(n5548) );
  INV_X1 U6092 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U6093 ( .A1(n5698), .A2(n6774), .ZN(n4939) );
  INV_X1 U6094 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4940) );
  XNOR2_X1 U6095 ( .A(n5698), .B(n4940), .ZN(n4941) );
  XNOR2_X1 U6096 ( .A(n5234), .B(n4941), .ZN(n5657) );
  AOI22_X1 U6097 ( .A1(n5128), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6098 ( .A1(n5129), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4944) );
  AOI22_X1 U6099 ( .A1(n5109), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4943) );
  AOI22_X1 U6100 ( .A1(n5135), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5112), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4942) );
  NAND4_X1 U6101 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n4951)
         );
  AOI22_X1 U6102 ( .A1(n3311), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6103 ( .A1(n5111), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4948) );
  AOI22_X1 U6104 ( .A1(n5075), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4947) );
  AOI22_X1 U6105 ( .A1(n5110), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4946) );
  NAND4_X1 U6106 ( .A1(n4949), .A2(n4948), .A3(n4947), .A4(n4946), .ZN(n4950)
         );
  NOR2_X1 U6107 ( .A1(n4951), .A2(n4950), .ZN(n5019) );
  AOI22_X1 U6108 ( .A1(n5111), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3294), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4955) );
  AOI22_X1 U6109 ( .A1(n5128), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4954) );
  AOI22_X1 U6110 ( .A1(n5129), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6111 ( .A1(n5028), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4952) );
  NAND4_X1 U6112 ( .A1(n4955), .A2(n4954), .A3(n4953), .A4(n4952), .ZN(n4961)
         );
  AOI22_X1 U6113 ( .A1(n5135), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4959) );
  AOI22_X1 U6114 ( .A1(n3311), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4958) );
  AOI22_X1 U6115 ( .A1(n5109), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6116 ( .A1(n5112), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4956) );
  NAND4_X1 U6117 ( .A1(n4959), .A2(n4958), .A3(n4957), .A4(n4956), .ZN(n4960)
         );
  OR2_X1 U6118 ( .A1(n4961), .A2(n4960), .ZN(n4991) );
  AOI22_X1 U6119 ( .A1(n5111), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6120 ( .A1(n5128), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4964) );
  AOI22_X1 U6121 ( .A1(n5129), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4963) );
  AOI22_X1 U6122 ( .A1(n5028), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4962) );
  NAND4_X1 U6123 ( .A1(n4965), .A2(n4964), .A3(n4963), .A4(n4962), .ZN(n4971)
         );
  AOI22_X1 U6124 ( .A1(n5135), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4969) );
  AOI22_X1 U6125 ( .A1(n3311), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U6126 ( .A1(n5109), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4967) );
  INV_X1 U6127 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6879) );
  AOI22_X1 U6128 ( .A1(n5112), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4966) );
  NAND4_X1 U6129 ( .A1(n4969), .A2(n4968), .A3(n4967), .A4(n4966), .ZN(n4970)
         );
  OR2_X1 U6130 ( .A1(n4971), .A2(n4970), .ZN(n4990) );
  NAND2_X1 U6131 ( .A1(n4991), .A2(n4990), .ZN(n5018) );
  OR2_X1 U6132 ( .A1(n5019), .A2(n5018), .ZN(n5039) );
  AOI22_X1 U6133 ( .A1(n5128), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4975) );
  AOI22_X1 U6134 ( .A1(n5111), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4974) );
  AOI22_X1 U6135 ( .A1(n5135), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U6136 ( .A1(n5110), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4972) );
  NAND4_X1 U6137 ( .A1(n4975), .A2(n4974), .A3(n4973), .A4(n4972), .ZN(n4981)
         );
  AOI22_X1 U6138 ( .A1(n5112), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4979) );
  AOI22_X1 U6139 ( .A1(n3294), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4978) );
  AOI22_X1 U6140 ( .A1(n5076), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U6141 ( .A1(n5129), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4976) );
  NAND4_X1 U6142 ( .A1(n4979), .A2(n4978), .A3(n4977), .A4(n4976), .ZN(n4980)
         );
  NOR2_X1 U6143 ( .A1(n4981), .A2(n4980), .ZN(n5040) );
  XOR2_X1 U6144 ( .A(n5039), .B(n5040), .Z(n4982) );
  NAND2_X1 U6145 ( .A1(n4982), .A2(n5091), .ZN(n4984) );
  AOI22_X1 U6146 ( .A1(n3385), .A2(EAX_REG_25__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6442), .ZN(n4983) );
  NAND2_X1 U6147 ( .A1(n4984), .A2(n4983), .ZN(n4988) );
  INV_X1 U6148 ( .A(n4985), .ZN(n4986) );
  XNOR2_X1 U6149 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .B(n4986), .ZN(n5762)
         );
  NOR2_X1 U6150 ( .A1(n5762), .A2(n5155), .ZN(n4987) );
  AOI21_X1 U6151 ( .B1(n4988), .B2(n5155), .A(n4987), .ZN(n4989) );
  INV_X1 U6152 ( .A(n4989), .ZN(n5254) );
  XNOR2_X1 U6153 ( .A(n4991), .B(n4990), .ZN(n4995) );
  NAND2_X1 U6154 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4992)
         );
  NAND2_X1 U6155 ( .A1(n5155), .A2(n4992), .ZN(n4993) );
  AOI21_X1 U6156 ( .B1(n5149), .B2(EAX_REG_23__SCAN_IN), .A(n4993), .ZN(n4994)
         );
  OAI21_X1 U6157 ( .B1(n5152), .B2(n4995), .A(n4994), .ZN(n4998) );
  INV_X1 U6158 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4996) );
  XNOR2_X1 U6159 ( .A(n5015), .B(n4996), .ZN(n5775) );
  NAND2_X1 U6160 ( .A1(n5775), .A2(n5148), .ZN(n4997) );
  AOI22_X1 U6161 ( .A1(n5128), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n5002) );
  AOI22_X1 U6162 ( .A1(n3301), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n5135), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5001) );
  AOI22_X1 U6163 ( .A1(n5112), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5000) );
  AOI22_X1 U6164 ( .A1(n5028), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4999) );
  NAND4_X1 U6165 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5008)
         );
  AOI22_X1 U6166 ( .A1(n5111), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5006) );
  AOI22_X1 U6167 ( .A1(n5110), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5005) );
  AOI22_X1 U6168 ( .A1(n5076), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5004) );
  AOI22_X1 U6169 ( .A1(n5136), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5003) );
  NAND4_X1 U6170 ( .A1(n5006), .A2(n5005), .A3(n5004), .A4(n5003), .ZN(n5007)
         );
  NOR2_X1 U6171 ( .A1(n5008), .A2(n5007), .ZN(n5012) );
  NAND2_X1 U6172 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5009)
         );
  NAND2_X1 U6173 ( .A1(n5155), .A2(n5009), .ZN(n5010) );
  AOI21_X1 U6174 ( .B1(n5149), .B2(EAX_REG_22__SCAN_IN), .A(n5010), .ZN(n5011)
         );
  OAI21_X1 U6175 ( .B1(n5152), .B2(n5012), .A(n5011), .ZN(n5017) );
  NOR2_X1 U6176 ( .A1(n5013), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5014)
         );
  NOR2_X1 U6177 ( .A1(n5015), .A2(n5014), .ZN(n5571) );
  NAND2_X1 U6178 ( .A1(n5571), .A2(n5148), .ZN(n5016) );
  NAND2_X1 U6179 ( .A1(n5017), .A2(n5016), .ZN(n5486) );
  NOR2_X1 U6180 ( .A1(n5482), .A2(n5486), .ZN(n5262) );
  AND2_X1 U6181 ( .A1(n5263), .A2(n5262), .ZN(n5414) );
  INV_X1 U6182 ( .A(n5018), .ZN(n5020) );
  XNOR2_X1 U6183 ( .A(n5020), .B(n5019), .ZN(n5026) );
  NAND2_X1 U6184 ( .A1(n5149), .A2(EAX_REG_24__SCAN_IN), .ZN(n5023) );
  XNOR2_X1 U6185 ( .A(n5021), .B(n5422), .ZN(n5563) );
  NAND2_X1 U6186 ( .A1(n5563), .A2(n5148), .ZN(n5022) );
  OAI211_X1 U6187 ( .C1(n5422), .C2(n5024), .A(n5023), .B(n5022), .ZN(n5025)
         );
  AOI21_X1 U6188 ( .B1(n5091), .B2(n5026), .A(n5025), .ZN(n5418) );
  INV_X1 U6189 ( .A(n5418), .ZN(n5027) );
  AND2_X1 U6190 ( .A1(n5414), .A2(n5027), .ZN(n5253) );
  AND2_X1 U6191 ( .A1(n5254), .A2(n5253), .ZN(n5051) );
  AOI22_X1 U6192 ( .A1(n5128), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5032) );
  AOI22_X1 U6193 ( .A1(n5129), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n5031) );
  AOI22_X1 U6194 ( .A1(n5112), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5030) );
  AOI22_X1 U6195 ( .A1(n5075), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5029) );
  NAND4_X1 U6196 ( .A1(n5032), .A2(n5031), .A3(n5030), .A4(n5029), .ZN(n5038)
         );
  AOI22_X1 U6197 ( .A1(n5111), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5036) );
  AOI22_X1 U6198 ( .A1(n5109), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5035) );
  AOI22_X1 U6199 ( .A1(n5135), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5034) );
  AOI22_X1 U6200 ( .A1(n5104), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5033) );
  NAND4_X1 U6201 ( .A1(n5036), .A2(n5035), .A3(n5034), .A4(n5033), .ZN(n5037)
         );
  NOR2_X1 U6202 ( .A1(n5038), .A2(n5037), .ZN(n5084) );
  OR2_X1 U6203 ( .A1(n5040), .A2(n5039), .ZN(n5083) );
  XNOR2_X1 U6204 ( .A(n5084), .B(n5083), .ZN(n5044) );
  NAND2_X1 U6205 ( .A1(n6442), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5041)
         );
  NAND2_X1 U6206 ( .A1(n5155), .A2(n5041), .ZN(n5042) );
  AOI21_X1 U6207 ( .B1(n3385), .B2(EAX_REG_26__SCAN_IN), .A(n5042), .ZN(n5043)
         );
  OAI21_X1 U6208 ( .B1(n5044), .B2(n5152), .A(n5043), .ZN(n5050) );
  INV_X1 U6209 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5047) );
  INV_X1 U6210 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6211 ( .A1(n5047), .A2(n5046), .ZN(n5048) );
  NAND2_X1 U6212 ( .A1(n5094), .A2(n5048), .ZN(n5751) );
  OR2_X1 U6213 ( .A1(n5751), .A2(n5155), .ZN(n5049) );
  AND2_X2 U6214 ( .A1(n5492), .A2(n5099), .ZN(n5402) );
  AND2_X1 U6215 ( .A1(n5491), .A2(n5051), .ZN(n5052) );
  NOR2_X1 U6216 ( .A1(n5054), .A2(n5053), .ZN(n5055) );
  OR2_X2 U6217 ( .A1(n5402), .A2(n5055), .ZN(n5478) );
  INV_X1 U6218 ( .A(n5478), .ZN(n5797) );
  AND2_X1 U6219 ( .A1(n6229), .A2(REIP_REG_26__SCAN_IN), .ZN(n5652) );
  AOI21_X1 U6220 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5652), 
        .ZN(n5056) );
  OAI21_X1 U6221 ( .B1(n6140), .B2(n5751), .A(n5056), .ZN(n5057) );
  AOI21_X1 U6222 ( .B1(n5797), .B2(n6137), .A(n5057), .ZN(n5058) );
  OAI21_X1 U6223 ( .B1(n6121), .B2(n5657), .A(n5058), .ZN(U2960) );
  INV_X1 U6224 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6225 ( .A1(n5096), .A2(n5225), .ZN(n5060) );
  NAND2_X1 U6226 ( .A1(n5102), .A2(n5060), .ZN(n5336) );
  AOI22_X1 U6227 ( .A1(n5135), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5064) );
  AOI22_X1 U6228 ( .A1(n3311), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5063) );
  AOI22_X1 U6229 ( .A1(n5129), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5062) );
  AOI22_X1 U6230 ( .A1(n3301), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5061) );
  NAND4_X1 U6231 ( .A1(n5064), .A2(n5063), .A3(n5062), .A4(n5061), .ZN(n5070)
         );
  AOI22_X1 U6232 ( .A1(n5128), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5028), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5068) );
  AOI22_X1 U6233 ( .A1(n5111), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5109), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5067) );
  AOI22_X1 U6234 ( .A1(n5110), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5066) );
  AOI22_X1 U6235 ( .A1(n5112), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5065) );
  NAND4_X1 U6236 ( .A1(n5068), .A2(n5067), .A3(n5066), .A4(n5065), .ZN(n5069)
         );
  NOR2_X1 U6237 ( .A1(n5070), .A2(n5069), .ZN(n5120) );
  AOI22_X1 U6238 ( .A1(n5128), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5111), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5074) );
  AOI22_X1 U6239 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5109), .B1(n5135), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U6240 ( .A1(n5028), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5072) );
  AOI22_X1 U6241 ( .A1(n5112), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5071) );
  NAND4_X1 U6242 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5082)
         );
  AOI22_X1 U6243 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5129), .B1(n5110), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n5080) );
  AOI22_X1 U6244 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3311), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U6245 ( .A1(n3301), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5078) );
  AOI22_X1 U6246 ( .A1(n5076), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5077) );
  NAND4_X1 U6247 ( .A1(n5080), .A2(n5079), .A3(n5078), .A4(n5077), .ZN(n5081)
         );
  NOR2_X1 U6248 ( .A1(n5082), .A2(n5081), .ZN(n5089) );
  OR2_X1 U6249 ( .A1(n5084), .A2(n5083), .ZN(n5090) );
  OR2_X1 U6250 ( .A1(n5089), .A2(n5090), .ZN(n5119) );
  XNOR2_X1 U6251 ( .A(n5120), .B(n5119), .ZN(n5087) );
  AOI21_X1 U6252 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6442), .A(n5148), 
        .ZN(n5086) );
  NAND2_X1 U6253 ( .A1(n5149), .A2(EAX_REG_28__SCAN_IN), .ZN(n5085) );
  OAI211_X1 U6254 ( .C1(n5087), .C2(n5152), .A(n5086), .B(n5085), .ZN(n5088)
         );
  OAI21_X1 U6255 ( .B1(n5155), .B2(n5336), .A(n5088), .ZN(n5220) );
  XOR2_X1 U6256 ( .A(n5090), .B(n5089), .Z(n5092) );
  NAND2_X1 U6257 ( .A1(n5092), .A2(n5091), .ZN(n5098) );
  INV_X1 U6258 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n6788) );
  NOR2_X1 U6259 ( .A1(n6788), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5093) );
  AOI211_X1 U6260 ( .C1(n3385), .C2(EAX_REG_27__SCAN_IN), .A(n5148), .B(n5093), 
        .ZN(n5097) );
  NAND2_X1 U6261 ( .A1(n5094), .A2(n6788), .ZN(n5095) );
  AND2_X1 U6262 ( .A1(n5096), .A2(n5095), .ZN(n5408) );
  AOI22_X1 U6263 ( .A1(n5098), .A2(n5097), .B1(n5148), .B2(n5408), .ZN(n5401)
         );
  INV_X1 U6264 ( .A(n5218), .ZN(n5100) );
  NOR2_X1 U6265 ( .A1(n5220), .A2(n5100), .ZN(n5101) );
  NAND2_X1 U6266 ( .A1(n5491), .A2(n5101), .ZN(n5219) );
  NAND2_X1 U6267 ( .A1(n5102), .A2(n5284), .ZN(n5103) );
  AND2_X1 U6268 ( .A1(n5127), .A2(n5103), .ZN(n5243) );
  OAI21_X1 U6269 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5284), .A(n5155), .ZN(
        n5123) );
  AOI22_X1 U6270 ( .A1(n5128), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5108) );
  AOI22_X1 U6271 ( .A1(n3311), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5107) );
  AOI22_X1 U6272 ( .A1(n3294), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5106) );
  AOI22_X1 U6273 ( .A1(n5076), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5105) );
  NAND4_X1 U6274 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n5118)
         );
  AOI22_X1 U6275 ( .A1(n5109), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5135), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U6276 ( .A1(n5111), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n5115) );
  AOI22_X1 U6277 ( .A1(n5028), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5114) );
  AOI22_X1 U6278 ( .A1(n5112), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5113) );
  NAND4_X1 U6279 ( .A1(n5116), .A2(n5115), .A3(n5114), .A4(n5113), .ZN(n5117)
         );
  NOR2_X1 U6280 ( .A1(n5118), .A2(n5117), .ZN(n5144) );
  OR2_X1 U6281 ( .A1(n5120), .A2(n5119), .ZN(n5145) );
  XNOR2_X1 U6282 ( .A(n5144), .B(n5145), .ZN(n5121) );
  NOR2_X1 U6283 ( .A1(n5121), .A2(n5152), .ZN(n5122) );
  AOI211_X1 U6284 ( .C1(n3385), .C2(EAX_REG_29__SCAN_IN), .A(n5123), .B(n5122), 
        .ZN(n5124) );
  AOI21_X1 U6285 ( .B1(n5148), .B2(n5243), .A(n5124), .ZN(n5241) );
  INV_X1 U6286 ( .A(n5241), .ZN(n5125) );
  OR2_X2 U6287 ( .A1(n3699), .A2(n5156), .ZN(n5240) );
  INV_X1 U6288 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5126) );
  XNOR2_X1 U6289 ( .A(n5127), .B(n5126), .ZN(n5368) );
  AOI22_X1 U6290 ( .A1(n5111), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3301), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5134) );
  AOI22_X1 U6291 ( .A1(n5128), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5110), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U6292 ( .A1(n5129), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5104), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U6293 ( .A1(n5028), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5130), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5131) );
  NAND4_X1 U6294 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n5143)
         );
  AOI22_X1 U6295 ( .A1(n5135), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5076), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5141) );
  AOI22_X1 U6296 ( .A1(n3351), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5140) );
  AOI22_X1 U6297 ( .A1(n5109), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5075), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U6298 ( .A1(n5112), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5138) );
  NAND4_X1 U6299 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n5142)
         );
  NOR2_X1 U6300 ( .A1(n5143), .A2(n5142), .ZN(n5147) );
  NOR2_X1 U6301 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  XOR2_X1 U6302 ( .A(n5147), .B(n5146), .Z(n5153) );
  AOI21_X1 U6303 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6442), .A(n5148), 
        .ZN(n5151) );
  NAND2_X1 U6304 ( .A1(n5149), .A2(EAX_REG_30__SCAN_IN), .ZN(n5150) );
  OAI211_X1 U6305 ( .C1(n5153), .C2(n5152), .A(n5151), .B(n5150), .ZN(n5154)
         );
  OAI21_X1 U6306 ( .B1(n5155), .B2(n5368), .A(n5154), .ZN(n5158) );
  OR2_X1 U6307 ( .A1(n5156), .A2(n5158), .ZN(n5157) );
  AOI21_X1 U6308 ( .B1(n5240), .B2(n5158), .A(n5308), .ZN(n5370) );
  INV_X1 U6309 ( .A(n5370), .ZN(n5249) );
  INV_X1 U6310 ( .A(n5159), .ZN(n5160) );
  AOI22_X1 U6311 ( .A1(n6002), .A2(DATAI_30_), .B1(n6005), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5165) );
  AND2_X1 U6312 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  NAND2_X1 U6313 ( .A1(n6006), .A2(DATAI_14_), .ZN(n5164) );
  OAI211_X1 U6314 ( .C1(n5249), .C2(n5796), .A(n5165), .B(n5164), .ZN(U2861)
         );
  NAND3_X1 U6315 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5206) );
  NOR2_X1 U6316 ( .A1(n5770), .A2(n5206), .ZN(n5754) );
  AND3_X1 U6317 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5208) );
  AND2_X1 U6318 ( .A1(n5754), .A2(n5208), .ZN(n5407) );
  AND2_X1 U6319 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5211) );
  INV_X1 U6320 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6593) );
  AND2_X1 U6321 ( .A1(n6593), .A2(REIP_REG_29__SCAN_IN), .ZN(n5216) );
  MUX2_X1 U6322 ( .A(n5273), .B(n5197), .S(EBX_REG_23__SCAN_IN), .Z(n5167) );
  NOR2_X1 U6323 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5166)
         );
  NOR2_X1 U6324 ( .A1(n5167), .A2(n5166), .ZN(n5292) );
  INV_X1 U6325 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U6326 ( .A1(n5176), .A2(n6717), .ZN(n5172) );
  INV_X1 U6327 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6328 ( .A1(n3912), .A2(n5168), .ZN(n5170) );
  NAND2_X1 U6329 ( .A1(n5189), .A2(n6717), .ZN(n5169) );
  NAND3_X1 U6330 ( .A1(n5170), .A2(n5169), .A3(n3111), .ZN(n5171) );
  NAND2_X1 U6331 ( .A1(n5172), .A2(n5171), .ZN(n5291) );
  NAND2_X1 U6332 ( .A1(n5292), .A2(n5291), .ZN(n5173) );
  MUX2_X1 U6333 ( .A(n5273), .B(n5197), .S(EBX_REG_25__SCAN_IN), .Z(n5175) );
  NOR2_X1 U6334 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5174)
         );
  NOR2_X1 U6335 ( .A1(n5175), .A2(n5174), .ZN(n5250) );
  INV_X1 U6336 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6337 ( .A1(n5176), .A2(n5421), .ZN(n5181) );
  INV_X1 U6338 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6339 ( .A1(n3912), .A2(n5177), .ZN(n5179) );
  NAND2_X1 U6340 ( .A1(n5189), .A2(n5421), .ZN(n5178) );
  NAND3_X1 U6341 ( .A1(n5179), .A2(n3111), .A3(n5178), .ZN(n5180) );
  NAND2_X1 U6342 ( .A1(n5181), .A2(n5180), .ZN(n5419) );
  NAND2_X1 U6343 ( .A1(n5250), .A2(n5419), .ZN(n5182) );
  NAND2_X1 U6344 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5183) );
  NAND2_X1 U6345 ( .A1(n3912), .A2(n5183), .ZN(n5185) );
  INV_X1 U6346 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6347 ( .A1(n5189), .A2(n5477), .ZN(n5184) );
  MUX2_X1 U6348 ( .A(n5197), .B(n5185), .S(n5184), .Z(n5474) );
  AND2_X2 U6349 ( .A1(n5475), .A2(n5474), .ZN(n5403) );
  MUX2_X1 U6350 ( .A(n5273), .B(n5197), .S(EBX_REG_27__SCAN_IN), .Z(n5187) );
  NOR2_X1 U6351 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5186)
         );
  NOR2_X1 U6352 ( .A1(n5187), .A2(n5186), .ZN(n5404) );
  AND2_X2 U6353 ( .A1(n5403), .A2(n5404), .ZN(n5406) );
  NAND2_X1 U6354 ( .A1(n3111), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5188) );
  NAND2_X1 U6355 ( .A1(n3912), .A2(n5188), .ZN(n5191) );
  INV_X1 U6356 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6357 ( .A1(n5189), .A2(n5298), .ZN(n5190) );
  MUX2_X1 U6358 ( .A(n5197), .B(n5191), .S(n5190), .Z(n5223) );
  NAND2_X1 U6359 ( .A1(n5406), .A2(n5223), .ZN(n5195) );
  OR2_X1 U6360 ( .A1(n5345), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5271)
         );
  OAI21_X1 U6361 ( .B1(EBX_REG_29__SCAN_IN), .B2(n5344), .A(n5271), .ZN(n5192)
         );
  NAND2_X1 U6362 ( .A1(n5345), .A2(EBX_REG_30__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6363 ( .A1(n5344), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6364 ( .A1(n5194), .A2(n5193), .ZN(n5342) );
  INV_X1 U6365 ( .A(n5279), .ZN(n5276) );
  NAND2_X1 U6366 ( .A1(n5200), .A2(n5276), .ZN(n5196) );
  NAND3_X1 U6367 ( .A1(n5341), .A2(n5342), .A3(n5196), .ZN(n5202) );
  INV_X1 U6368 ( .A(n5342), .ZN(n5199) );
  NAND2_X1 U6369 ( .A1(n5279), .A2(n5197), .ZN(n5198) );
  NAND3_X1 U6370 ( .A1(n5200), .A2(n5199), .A3(n5198), .ZN(n5201) );
  INV_X1 U6371 ( .A(n5368), .ZN(n5203) );
  AOI22_X1 U6372 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5952), .B1(n5986), 
        .B2(n5203), .ZN(n5205) );
  NAND2_X1 U6373 ( .A1(n5969), .A2(EBX_REG_30__SCAN_IN), .ZN(n5204) );
  OAI211_X1 U6374 ( .C1(n5376), .C2(n5929), .A(n5205), .B(n5204), .ZN(n5215)
         );
  AND2_X1 U6375 ( .A1(n5395), .A2(n5206), .ZN(n5207) );
  NOR2_X1 U6376 ( .A1(n5791), .A2(n5207), .ZN(n5773) );
  INV_X1 U6377 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6378 ( .A1(n5395), .A2(n5209), .ZN(n5210) );
  NAND2_X1 U6379 ( .A1(n5773), .A2(n5210), .ZN(n5755) );
  INV_X1 U6380 ( .A(n5211), .ZN(n5212) );
  AND2_X1 U6381 ( .A1(n5979), .A2(n5212), .ZN(n5213) );
  INV_X1 U6382 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6587) );
  OR2_X1 U6383 ( .A1(n5289), .A2(n6587), .ZN(n5396) );
  AND3_X1 U6384 ( .A1(n5396), .A2(REIP_REG_30__SCAN_IN), .A3(n5395), .ZN(n5214) );
  OAI21_X1 U6385 ( .B1(n5249), .B2(n5753), .A(n5217), .ZN(U2797) );
  NAND2_X1 U6386 ( .A1(n5492), .A2(n5218), .ZN(n5400) );
  NOR2_X1 U6387 ( .A1(n3699), .A2(n5219), .ZN(n5242) );
  AOI21_X2 U6388 ( .B1(n5220), .B2(n5400), .A(n5242), .ZN(n5338) );
  INV_X1 U6389 ( .A(n5338), .ZN(n5297) );
  AOI22_X1 U6390 ( .A1(n6002), .A2(DATAI_28_), .B1(n6005), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U6391 ( .A1(n6006), .A2(DATAI_12_), .ZN(n5221) );
  OAI211_X1 U6392 ( .C1(n5297), .C2(n5796), .A(n5222), .B(n5221), .ZN(U2863)
         );
  OR2_X1 U6393 ( .A1(n5406), .A2(n5223), .ZN(n5224) );
  NAND2_X1 U6394 ( .A1(n5279), .A2(n5224), .ZN(n5318) );
  NAND3_X1 U6395 ( .A1(n5407), .A2(REIP_REG_27__SCAN_IN), .A3(n6586), .ZN(
        n5228) );
  OAI22_X1 U6396 ( .A1(n5225), .A2(n5989), .B1(n5977), .B2(n5336), .ZN(n5226)
         );
  AOI21_X1 U6397 ( .B1(n5969), .B2(EBX_REG_28__SCAN_IN), .A(n5226), .ZN(n5227)
         );
  OAI211_X1 U6398 ( .C1(n5929), .C2(n5318), .A(n5228), .B(n5227), .ZN(n5229)
         );
  AOI21_X1 U6399 ( .B1(n5289), .B2(REIP_REG_28__SCAN_IN), .A(n5229), .ZN(n5230) );
  OAI21_X1 U6400 ( .B1(n5297), .B2(n5753), .A(n5230), .ZN(U2799) );
  AOI22_X1 U6401 ( .A1(n6006), .A2(DATAI_3_), .B1(n6005), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6402 ( .A1(n6002), .A2(DATAI_19_), .ZN(n5231) );
  OAI211_X1 U6403 ( .C1(n5501), .C2(n5796), .A(n5232), .B(n5231), .ZN(U2872)
         );
  NAND2_X1 U6404 ( .A1(n5822), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5233) );
  NOR2_X2 U6405 ( .A1(n5234), .A2(n5233), .ZN(n5538) );
  INV_X1 U6406 ( .A(n5548), .ZN(n5236) );
  NOR2_X1 U6407 ( .A1(n5568), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5235)
         );
  NOR2_X1 U6408 ( .A1(n5539), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5237)
         );
  AOI21_X1 U6409 ( .B1(n5538), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5237), 
        .ZN(n5314) );
  AND2_X1 U6410 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5351) );
  NOR2_X1 U6411 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5238) );
  NOR2_X1 U6412 ( .A1(n5351), .A2(n5238), .ZN(n5320) );
  NOR2_X1 U6413 ( .A1(n5314), .A2(n5320), .ZN(n5239) );
  XNOR2_X1 U6414 ( .A(n5239), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5641)
         );
  OAI21_X1 U6415 ( .B1(n5242), .B2(n5241), .A(n5240), .ZN(n5281) );
  INV_X1 U6416 ( .A(n5281), .ZN(n5246) );
  INV_X1 U6417 ( .A(n5243), .ZN(n5283) );
  AND2_X1 U6418 ( .A1(n6229), .A2(REIP_REG_29__SCAN_IN), .ZN(n5634) );
  AOI21_X1 U6419 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5634), 
        .ZN(n5244) );
  OAI21_X1 U6420 ( .B1(n6140), .B2(n5283), .A(n5244), .ZN(n5245) );
  AOI21_X1 U6421 ( .B1(n5246), .B2(n6137), .A(n5245), .ZN(n5247) );
  OAI21_X1 U6422 ( .B1(n5641), .B2(n6121), .A(n5247), .ZN(U2957) );
  INV_X1 U6423 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5248) );
  OAI222_X1 U6424 ( .A1(n5515), .A2(n5249), .B1(n5525), .B2(n5248), .C1(n5376), 
        .C2(n5516), .ZN(U2829) );
  INV_X1 U6425 ( .A(n5420), .ZN(n5251) );
  AOI21_X1 U6426 ( .B1(n5251), .B2(n5419), .A(n5250), .ZN(n5252) );
  NOR2_X1 U6427 ( .A1(n5252), .A2(n5475), .ZN(n5763) );
  INV_X1 U6428 ( .A(n5763), .ZN(n5658) );
  NAND2_X1 U6429 ( .A1(n5492), .A2(n5253), .ZN(n5415) );
  XNOR2_X2 U6430 ( .A(n5415), .B(n5254), .ZN(n5800) );
  INV_X1 U6431 ( .A(n5800), .ZN(n5255) );
  INV_X1 U6432 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6748) );
  OAI222_X1 U6433 ( .A1(n5516), .A2(n5658), .B1(n5515), .B2(n5255), .C1(n5525), 
        .C2(n6748), .ZN(U2834) );
  INV_X1 U6434 ( .A(n5316), .ZN(n5256) );
  NAND2_X1 U6435 ( .A1(n5257), .A2(n5256), .ZN(n5259) );
  NAND2_X1 U6436 ( .A1(n5698), .A2(n6742), .ZN(n5586) );
  NOR2_X1 U6437 ( .A1(n5731), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5258)
         );
  OAI22_X1 U6438 ( .A1(n5700), .A2(n5258), .B1(n5822), .B2(n5713), .ZN(n5576)
         );
  XNOR2_X1 U6439 ( .A(n5698), .B(n5684), .ZN(n5577) );
  NOR2_X1 U6440 ( .A1(n5576), .A2(n5577), .ZN(n5575) );
  NOR2_X1 U6441 ( .A1(n5568), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5567)
         );
  NAND2_X1 U6442 ( .A1(n5575), .A2(n5567), .ZN(n5556) );
  OAI21_X1 U6443 ( .B1(n3108), .B2(n5259), .A(n5556), .ZN(n5261) );
  XNOR2_X1 U6444 ( .A(n5261), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5679)
         );
  AND2_X2 U6445 ( .A1(n5492), .A2(n5262), .ZN(n5484) );
  XNOR2_X2 U6446 ( .A(n5484), .B(n5264), .ZN(n5803) );
  INV_X1 U6447 ( .A(n5775), .ZN(n5266) );
  NAND2_X1 U6448 ( .A1(n6229), .A2(REIP_REG_23__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U6449 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5265)
         );
  OAI211_X1 U6450 ( .C1(n6140), .C2(n5266), .A(n5673), .B(n5265), .ZN(n5267)
         );
  AOI21_X1 U6451 ( .B1(n5803), .B2(n6137), .A(n5267), .ZN(n5268) );
  OAI21_X1 U6452 ( .B1(n5679), .B2(n6121), .A(n5268), .ZN(U2963) );
  AOI22_X1 U6453 ( .A1(n6002), .A2(DATAI_29_), .B1(n6005), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6454 ( .A1(n6006), .A2(DATAI_13_), .ZN(n5269) );
  OAI211_X1 U6455 ( .C1(n5281), .C2(n5796), .A(n5270), .B(n5269), .ZN(U2862)
         );
  INV_X1 U6456 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5282) );
  INV_X1 U6457 ( .A(n5271), .ZN(n5272) );
  MUX2_X1 U6458 ( .A(EBX_REG_29__SCAN_IN), .B(n5272), .S(n3111), .Z(n5275) );
  AND2_X1 U6459 ( .A1(n5273), .A2(n5282), .ZN(n5274) );
  NOR2_X1 U6460 ( .A1(n5275), .A2(n5274), .ZN(n5277) );
  NAND2_X1 U6461 ( .A1(n5276), .A2(n5277), .ZN(n5343) );
  INV_X1 U6462 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6463 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6464 ( .A1(n5343), .A2(n5280), .ZN(n5633) );
  OAI222_X1 U6465 ( .A1(n5282), .A2(n5525), .B1(n5516), .B2(n5633), .C1(n5281), 
        .C2(n5515), .ZN(U2830) );
  NAND2_X1 U6466 ( .A1(n5391), .A2(n6587), .ZN(n5287) );
  OAI22_X1 U6467 ( .A1(n5284), .A2(n5989), .B1(n5977), .B2(n5283), .ZN(n5285)
         );
  AOI21_X1 U6468 ( .B1(n5969), .B2(EBX_REG_29__SCAN_IN), .A(n5285), .ZN(n5286)
         );
  OAI211_X1 U6469 ( .C1(n5929), .C2(n5633), .A(n5287), .B(n5286), .ZN(n5288)
         );
  AOI21_X1 U6470 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5289), .A(n5288), .ZN(n5290) );
  OAI21_X1 U6471 ( .B1(n5281), .B2(n5753), .A(n5290), .ZN(U2798) );
  INV_X1 U6472 ( .A(n5803), .ZN(n5296) );
  INV_X1 U6473 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5295) );
  INV_X1 U6474 ( .A(n5291), .ZN(n5487) );
  INV_X1 U6475 ( .A(n5292), .ZN(n5293) );
  OAI21_X1 U6476 ( .B1(n5488), .B2(n5487), .A(n5293), .ZN(n5294) );
  NAND2_X1 U6477 ( .A1(n5294), .A2(n5420), .ZN(n5771) );
  OAI222_X1 U6478 ( .A1(n5296), .A2(n5515), .B1(n5525), .B2(n5295), .C1(n5771), 
        .C2(n5516), .ZN(U2836) );
  OAI222_X1 U6479 ( .A1(n5298), .A2(n5525), .B1(n5516), .B2(n5318), .C1(n5297), 
        .C2(n5515), .ZN(U2831) );
  AOI22_X1 U6480 ( .A1(n5693), .A2(n5480), .B1(n5479), .B2(EBX_REG_21__SCAN_IN), .ZN(n5299) );
  OAI21_X1 U6481 ( .B1(n5300), .B2(n5515), .A(n5299), .ZN(U2838) );
  INV_X1 U6482 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5301) );
  NAND3_X1 U6483 ( .A1(n5301), .A2(n5313), .A3(n5645), .ZN(n5302) );
  NOR2_X2 U6484 ( .A1(n5539), .A2(n5302), .ZN(n5361) );
  INV_X1 U6485 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U6486 ( .A1(n5361), .A2(n6924), .ZN(n5364) );
  NAND2_X1 U6487 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5355) );
  INV_X1 U6488 ( .A(n5355), .ZN(n5303) );
  AOI22_X1 U6489 ( .A1(n3385), .A2(EAX_REG_31__SCAN_IN), .B1(n5306), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6490 ( .A(n5308), .B(n5307), .ZN(n5386) );
  AND2_X1 U6491 ( .A1(n6229), .A2(REIP_REG_31__SCAN_IN), .ZN(n5349) );
  AOI21_X1 U6492 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5349), 
        .ZN(n5309) );
  OAI21_X1 U6493 ( .B1(n6140), .B2(n5310), .A(n5309), .ZN(n5311) );
  AOI21_X1 U6494 ( .B1(n5386), .B2(n6137), .A(n5311), .ZN(n5312) );
  OAI21_X1 U6495 ( .B1(n5360), .B2(n6121), .A(n5312), .ZN(U2955) );
  XNOR2_X1 U6496 ( .A(n5314), .B(n5313), .ZN(n5340) );
  NOR3_X1 U6497 ( .A1(n5730), .A2(n6914), .A3(n5315), .ZN(n5701) );
  NAND2_X1 U6498 ( .A1(n5702), .A2(n5701), .ZN(n5729) );
  NOR2_X1 U6499 ( .A1(n5709), .A2(n5729), .ZN(n5321) );
  NAND2_X1 U6500 ( .A1(n5321), .A2(n6155), .ZN(n5720) );
  NOR2_X1 U6501 ( .A1(n5720), .A2(n5316), .ZN(n5677) );
  INV_X1 U6502 ( .A(n5327), .ZN(n5317) );
  AND2_X1 U6503 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5330) );
  AND2_X1 U6504 ( .A1(n6229), .A2(REIP_REG_28__SCAN_IN), .ZN(n5334) );
  NOR2_X1 U6505 ( .A1(n5318), .A2(n6207), .ZN(n5319) );
  AOI211_X1 U6506 ( .C1(n5646), .C2(n5320), .A(n5334), .B(n5319), .ZN(n5333)
         );
  NAND2_X1 U6507 ( .A1(n5712), .A2(n5321), .ZN(n5683) );
  NAND2_X1 U6508 ( .A1(n5683), .A2(n6232), .ZN(n5322) );
  NAND2_X1 U6509 ( .A1(n6151), .A2(n5322), .ZN(n5694) );
  INV_X1 U6510 ( .A(n5323), .ZN(n5324) );
  AND2_X1 U6511 ( .A1(n6232), .A2(n5324), .ZN(n5325) );
  NOR2_X1 U6512 ( .A1(n5694), .A2(n5325), .ZN(n5674) );
  NAND2_X1 U6513 ( .A1(n5326), .A2(n5711), .ZN(n5328) );
  NAND2_X1 U6514 ( .A1(n5328), .A2(n5327), .ZN(n5329) );
  NAND2_X1 U6515 ( .A1(n5674), .A2(n5329), .ZN(n5662) );
  INV_X1 U6516 ( .A(n5662), .ZN(n5667) );
  INV_X1 U6517 ( .A(n5330), .ZN(n5651) );
  NAND2_X1 U6518 ( .A1(n6232), .A2(n5651), .ZN(n5331) );
  INV_X1 U6519 ( .A(n5353), .ZN(n5647) );
  NAND2_X1 U6520 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5332) );
  OAI211_X1 U6521 ( .C1(n5340), .C2(n6196), .A(n5333), .B(n5332), .ZN(U2990)
         );
  AOI21_X1 U6522 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5334), 
        .ZN(n5335) );
  OAI21_X1 U6523 ( .B1(n6140), .B2(n5336), .A(n5335), .ZN(n5337) );
  AOI21_X1 U6524 ( .B1(n5338), .B2(n6137), .A(n5337), .ZN(n5339) );
  OAI21_X1 U6525 ( .B1(n5340), .B2(n6121), .A(n5339), .ZN(U2958) );
  AOI22_X1 U6526 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5345), .B1(n5344), .B2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5346) );
  XNOR2_X1 U6527 ( .A(n5347), .B(n5346), .ZN(n5472) );
  INV_X1 U6528 ( .A(n5472), .ZN(n5350) );
  NAND2_X1 U6529 ( .A1(n5646), .A2(n5351), .ZN(n5637) );
  NOR3_X1 U6530 ( .A1(n5637), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5355), 
        .ZN(n5348) );
  OR2_X1 U6531 ( .A1(n5662), .A2(n6232), .ZN(n5378) );
  INV_X1 U6532 ( .A(n5351), .ZN(n5352) );
  NAND2_X1 U6533 ( .A1(n5378), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U6534 ( .A1(n5354), .A2(n5353), .ZN(n5639) );
  NOR2_X1 U6535 ( .A1(n5356), .A2(n5303), .ZN(n5357) );
  OAI21_X1 U6536 ( .B1(n5639), .B2(n5357), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n5358) );
  OAI211_X1 U6537 ( .C1(n5360), .C2(n6196), .A(n5359), .B(n5358), .ZN(U2987)
         );
  NAND2_X1 U6538 ( .A1(n3114), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5365) );
  INV_X1 U6539 ( .A(n5361), .ZN(n5362) );
  NAND3_X1 U6540 ( .A1(n5365), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5362), .ZN(n5363) );
  OAI211_X1 U6541 ( .C1(n5365), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5364), .B(n5363), .ZN(n5366) );
  INV_X1 U6542 ( .A(n5366), .ZN(n5381) );
  AND2_X1 U6543 ( .A1(n6229), .A2(REIP_REG_30__SCAN_IN), .ZN(n5372) );
  AOI21_X1 U6544 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5372), 
        .ZN(n5367) );
  OAI21_X1 U6545 ( .B1(n6140), .B2(n5368), .A(n5367), .ZN(n5369) );
  AOI21_X1 U6546 ( .B1(n5370), .B2(n6137), .A(n5369), .ZN(n5371) );
  OAI21_X1 U6547 ( .B1(n5381), .B2(n6121), .A(n5371), .ZN(U2956) );
  INV_X1 U6548 ( .A(n5372), .ZN(n5375) );
  NAND2_X1 U6549 ( .A1(n6924), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5373) );
  OR2_X1 U6550 ( .A1(n5637), .A2(n5373), .ZN(n5374) );
  OAI211_X1 U6551 ( .C1(n5376), .C2(n6207), .A(n5375), .B(n5374), .ZN(n5377)
         );
  INV_X1 U6552 ( .A(n5377), .ZN(n5380) );
  OAI211_X1 U6553 ( .C1(n5639), .C2(n5301), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5378), .ZN(n5379) );
  OAI211_X1 U6554 ( .C1(n5381), .C2(n6196), .A(n5380), .B(n5379), .ZN(U2988)
         );
  NAND3_X1 U6555 ( .A1(n5386), .A2(n5383), .A3(n5382), .ZN(n5385) );
  AOI22_X1 U6556 ( .A1(n6002), .A2(DATAI_31_), .B1(n6005), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6557 ( .A1(n5385), .A2(n5384), .ZN(U2860) );
  INV_X1 U6558 ( .A(n5386), .ZN(n5399) );
  INV_X1 U6559 ( .A(n5387), .ZN(n5389) );
  AOI22_X1 U6560 ( .A1(n5389), .A2(n5388), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), 
        .B2(n5952), .ZN(n5393) );
  INV_X1 U6561 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5390) );
  NAND4_X1 U6562 ( .A1(n5391), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n5390), .ZN(n5392) );
  OAI211_X1 U6563 ( .C1(n5472), .C2(n5929), .A(n5393), .B(n5392), .ZN(n5394)
         );
  INV_X1 U6564 ( .A(n5394), .ZN(n5398) );
  OAI211_X1 U6565 ( .C1(n5396), .C2(n6593), .A(REIP_REG_31__SCAN_IN), .B(n5395), .ZN(n5397) );
  OAI211_X1 U6566 ( .C1(n5399), .C2(n5753), .A(n5398), .B(n5397), .ZN(U2796)
         );
  NOR2_X1 U6567 ( .A1(n5403), .A2(n5404), .ZN(n5405) );
  OR2_X1 U6568 ( .A1(n5406), .A2(n5405), .ZN(n5642) );
  INV_X1 U6569 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U6570 ( .A1(n5407), .A2(n6583), .ZN(n5411) );
  INV_X1 U6571 ( .A(n5408), .ZN(n5544) );
  OAI22_X1 U6572 ( .A1(n6788), .A2(n5989), .B1(n5977), .B2(n5544), .ZN(n5409)
         );
  AOI21_X1 U6573 ( .B1(n5969), .B2(EBX_REG_27__SCAN_IN), .A(n5409), .ZN(n5410)
         );
  OAI211_X1 U6574 ( .C1(n5929), .C2(n5642), .A(n5411), .B(n5410), .ZN(n5412)
         );
  AOI21_X1 U6575 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5755), .A(n5412), .ZN(n5413) );
  OAI21_X1 U6576 ( .B1(n5542), .B2(n5753), .A(n5413), .ZN(U2800) );
  NAND2_X1 U6577 ( .A1(n5492), .A2(n5414), .ZN(n5417) );
  INV_X1 U6578 ( .A(n5415), .ZN(n5416) );
  XNOR2_X1 U6579 ( .A(n5420), .B(n5419), .ZN(n5670) );
  INV_X1 U6580 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6578) );
  OAI22_X1 U6581 ( .A1(n5773), .A2(n6578), .B1(n5563), .B2(n5977), .ZN(n5424)
         );
  OAI22_X1 U6582 ( .A1(n5422), .A2(n5989), .B1(n5421), .B2(n5994), .ZN(n5423)
         );
  AOI211_X1 U6583 ( .C1(n5670), .C2(n5965), .A(n5424), .B(n5423), .ZN(n5425)
         );
  NAND2_X1 U6584 ( .A1(n5754), .A2(n6578), .ZN(n5764) );
  OAI211_X1 U6585 ( .C1(n5533), .C2(n5753), .A(n5425), .B(n5764), .ZN(U2803)
         );
  NAND2_X1 U6586 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  INV_X1 U6587 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U6588 ( .A1(n5510), .A2(n5431), .ZN(n5432) );
  INV_X1 U6589 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6569) );
  AOI22_X1 U6590 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n5952), .B1(
        EBX_REG_18__SCAN_IN), .B2(n5969), .ZN(n5434) );
  OAI211_X1 U6591 ( .C1(n5878), .C2(n6569), .A(n5434), .B(n5971), .ZN(n5437)
         );
  INV_X1 U6592 ( .A(n5435), .ZN(n5789) );
  OAI22_X1 U6593 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5789), .B1(n5828), .B2(
        n5977), .ZN(n5436) );
  AOI211_X1 U6594 ( .C1(n5965), .C2(n5832), .A(n5437), .B(n5436), .ZN(n5438)
         );
  OAI21_X1 U6595 ( .B1(n5504), .B2(n5753), .A(n5438), .ZN(U2809) );
  OAI21_X1 U6596 ( .B1(n5439), .B2(n5441), .A(n5440), .ZN(n6001) );
  INV_X1 U6597 ( .A(n5514), .ZN(n5447) );
  INV_X1 U6598 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5513) );
  INV_X1 U6599 ( .A(n5600), .ZN(n5442) );
  OAI22_X1 U6600 ( .A1(n5994), .A2(n5513), .B1(n5977), .B2(n5442), .ZN(n5446)
         );
  INV_X1 U6601 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6566) );
  AOI21_X1 U6602 ( .B1(n6731), .B2(n6566), .A(n5879), .ZN(n5443) );
  NAND2_X1 U6603 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5880) );
  AOI22_X1 U6604 ( .A1(n5443), .A2(n5880), .B1(REIP_REG_16__SCAN_IN), .B2(
        n5892), .ZN(n5444) );
  OAI211_X1 U6605 ( .C1(n5989), .C2(n5597), .A(n5444), .B(n5971), .ZN(n5445)
         );
  AOI211_X1 U6606 ( .C1(n5447), .C2(n5965), .A(n5446), .B(n5445), .ZN(n5448)
         );
  OAI21_X1 U6607 ( .B1(n6001), .B2(n5753), .A(n5448), .ZN(U2811) );
  AND2_X1 U6608 ( .A1(n4927), .A2(n5449), .ZN(n5450) );
  OR2_X1 U6609 ( .A1(n5450), .A2(n5439), .ZN(n5614) );
  INV_X1 U6610 ( .A(n5451), .ZN(n5611) );
  OR2_X1 U6611 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  NAND2_X1 U6612 ( .A1(n5455), .A2(n5454), .ZN(n5843) );
  OAI22_X1 U6613 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5879), .B1(n5929), .B2(
        n5843), .ZN(n5458) );
  AOI22_X1 U6614 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5969), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5892), .ZN(n5456) );
  OAI211_X1 U6615 ( .C1(n5989), .C2(n6758), .A(n5456), .B(n5971), .ZN(n5457)
         );
  AOI211_X1 U6616 ( .C1(n5986), .C2(n5611), .A(n5458), .B(n5457), .ZN(n5459)
         );
  OAI21_X1 U6617 ( .B1(n5614), .B2(n5753), .A(n5459), .ZN(U2812) );
  OAI22_X1 U6618 ( .A1(n6129), .A2(n5977), .B1(n5989), .B2(n5460), .ZN(n5463)
         );
  NOR2_X1 U6619 ( .A1(n5994), .A2(n5461), .ZN(n5462) );
  AOI211_X1 U6620 ( .C1(n5984), .C2(n5464), .A(n5463), .B(n5462), .ZN(n5465)
         );
  OAI21_X1 U6621 ( .B1(n5929), .B2(n5466), .A(n5465), .ZN(n5469) );
  AOI221_X1 U6622 ( .B1(n6745), .B2(n6548), .C1(n5967), .C2(n6548), .A(n5467), 
        .ZN(n5468) );
  AOI211_X1 U6623 ( .C1(n6126), .C2(n5991), .A(n5469), .B(n5468), .ZN(n5470)
         );
  INV_X1 U6624 ( .A(n5470), .ZN(U2825) );
  INV_X1 U6625 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5471) );
  OAI22_X1 U6626 ( .A1(n5472), .A2(n5516), .B1(n5471), .B2(n5525), .ZN(U2828)
         );
  INV_X1 U6627 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5473) );
  OAI222_X1 U6628 ( .A1(n5473), .A2(n5525), .B1(n5516), .B2(n5642), .C1(n5542), 
        .C2(n5515), .ZN(U2832) );
  NOR2_X1 U6629 ( .A1(n5475), .A2(n5474), .ZN(n5476) );
  OR2_X1 U6630 ( .A1(n5403), .A2(n5476), .ZN(n5759) );
  OAI222_X1 U6631 ( .A1(n5515), .A2(n5478), .B1(n5525), .B2(n5477), .C1(n5759), 
        .C2(n5516), .ZN(U2833) );
  AOI22_X1 U6632 ( .A1(n5670), .A2(n5480), .B1(n5479), .B2(EBX_REG_24__SCAN_IN), .ZN(n5481) );
  OAI21_X1 U6633 ( .B1(n5533), .B2(n5515), .A(n5481), .ZN(U2835) );
  INV_X1 U6634 ( .A(n5482), .ZN(n5483) );
  NAND2_X1 U6635 ( .A1(n5492), .A2(n5483), .ZN(n5485) );
  AOI21_X2 U6636 ( .B1(n5486), .B2(n5485), .A(n5484), .ZN(n5806) );
  INV_X1 U6637 ( .A(n5515), .ZN(n5527) );
  XNOR2_X1 U6638 ( .A(n5488), .B(n5487), .ZN(n5787) );
  OAI22_X1 U6639 ( .A1(n5787), .A2(n5516), .B1(n6717), .B2(n5525), .ZN(n5489)
         );
  AOI21_X1 U6640 ( .B1(n5806), .B2(n5527), .A(n5489), .ZN(n5490) );
  INV_X1 U6641 ( .A(n5490), .ZN(U2837) );
  INV_X1 U6642 ( .A(n5491), .ZN(n5493) );
  AOI21_X1 U6643 ( .B1(n5493), .B2(n3699), .A(n5492), .ZN(n5813) );
  INV_X1 U6644 ( .A(n5813), .ZN(n5500) );
  INV_X1 U6645 ( .A(n5494), .ZN(n5496) );
  MUX2_X1 U6646 ( .A(n3111), .B(n5496), .S(n5495), .Z(n5499) );
  XNOR2_X1 U6647 ( .A(n5499), .B(n5498), .ZN(n5795) );
  OAI222_X1 U6648 ( .A1(n5500), .A2(n5515), .B1(n5516), .B2(n5795), .C1(n5525), 
        .C2(n3904), .ZN(U2839) );
  OAI22_X1 U6649 ( .A1(n5724), .A2(n5516), .B1(n6875), .B2(n5525), .ZN(n5502)
         );
  AOI21_X1 U6650 ( .B1(n5595), .B2(n5527), .A(n5502), .ZN(n5503) );
  INV_X1 U6651 ( .A(n5503), .ZN(U2840) );
  INV_X1 U6652 ( .A(n5832), .ZN(n5505) );
  INV_X1 U6653 ( .A(EBX_REG_18__SCAN_IN), .ZN(n6816) );
  OAI222_X1 U6654 ( .A1(n5516), .A2(n5505), .B1(n5525), .B2(n6816), .C1(n5515), 
        .C2(n5504), .ZN(U2841) );
  XOR2_X1 U6655 ( .A(n5506), .B(n5440), .Z(n5998) );
  NAND2_X1 U6656 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  NAND2_X1 U6657 ( .A1(n5510), .A2(n5509), .ZN(n5887) );
  OAI22_X1 U6658 ( .A1(n5887), .A2(n5516), .B1(n5883), .B2(n5525), .ZN(n5511)
         );
  AOI21_X1 U6659 ( .B1(n5998), .B2(n5527), .A(n5511), .ZN(n5512) );
  INV_X1 U6660 ( .A(n5512), .ZN(U2842) );
  OAI222_X1 U6661 ( .A1(n5514), .A2(n5516), .B1(n5513), .B2(n5525), .C1(n6001), 
        .C2(n5515), .ZN(U2843) );
  INV_X1 U6662 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6684) );
  OAI222_X1 U6663 ( .A1(n5843), .A2(n5516), .B1(n5525), .B2(n6684), .C1(n5515), 
        .C2(n5614), .ZN(U2844) );
  INV_X1 U6664 ( .A(n5517), .ZN(n5518) );
  AOI21_X1 U6665 ( .B1(n5520), .B2(n5519), .A(n5518), .ZN(n5903) );
  NAND2_X1 U6666 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  NAND2_X1 U6667 ( .A1(n5524), .A2(n5523), .ZN(n5898) );
  OAI22_X1 U6668 ( .A1(n5898), .A2(n5516), .B1(n5899), .B2(n5525), .ZN(n5526)
         );
  AOI21_X1 U6669 ( .B1(n5903), .B2(n5527), .A(n5526), .ZN(n5528) );
  INV_X1 U6670 ( .A(n5528), .ZN(U2846) );
  AOI22_X1 U6671 ( .A1(n6002), .A2(DATAI_27_), .B1(n6005), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U6672 ( .A1(n6006), .A2(DATAI_11_), .ZN(n5529) );
  OAI211_X1 U6673 ( .C1(n5542), .C2(n5796), .A(n5530), .B(n5529), .ZN(U2864)
         );
  AOI22_X1 U6674 ( .A1(n6002), .A2(DATAI_24_), .B1(n6005), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6675 ( .A1(n6006), .A2(DATAI_8_), .ZN(n5531) );
  OAI211_X1 U6676 ( .C1(n5533), .C2(n5796), .A(n5532), .B(n5531), .ZN(U2867)
         );
  AOI22_X1 U6677 ( .A1(n5535), .A2(DATAI_15_), .B1(n6005), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5534) );
  OAI21_X1 U6678 ( .B1(n5614), .B2(n5796), .A(n5534), .ZN(U2876) );
  INV_X1 U6679 ( .A(n5903), .ZN(n5537) );
  AOI22_X1 U6680 ( .A1(n5535), .A2(DATAI_13_), .B1(n6005), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5536) );
  OAI21_X1 U6681 ( .B1(n5537), .B2(n5796), .A(n5536), .ZN(U2878) );
  INV_X1 U6682 ( .A(n5538), .ZN(n5540) );
  NAND2_X1 U6683 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  XNOR2_X1 U6684 ( .A(n5541), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5650)
         );
  INV_X1 U6685 ( .A(n5542), .ZN(n5546) );
  AND2_X1 U6686 ( .A1(n6229), .A2(REIP_REG_27__SCAN_IN), .ZN(n5644) );
  AOI21_X1 U6687 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5644), 
        .ZN(n5543) );
  OAI21_X1 U6688 ( .B1(n6140), .B2(n5544), .A(n5543), .ZN(n5545) );
  AOI21_X1 U6689 ( .B1(n5546), .B2(n6137), .A(n5545), .ZN(n5547) );
  OAI21_X1 U6690 ( .B1(n5650), .B2(n6121), .A(n5547), .ZN(U2959) );
  OAI21_X1 U6691 ( .B1(n5550), .B2(n5549), .A(n5548), .ZN(n5551) );
  INV_X1 U6692 ( .A(n5551), .ZN(n5665) );
  INV_X1 U6693 ( .A(n5762), .ZN(n5553) );
  AND2_X1 U6694 ( .A1(n6229), .A2(REIP_REG_25__SCAN_IN), .ZN(n5660) );
  AOI21_X1 U6695 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n5660), 
        .ZN(n5552) );
  OAI21_X1 U6696 ( .B1(n6140), .B2(n5553), .A(n5552), .ZN(n5554) );
  AOI21_X1 U6697 ( .B1(n5800), .B2(n6137), .A(n5554), .ZN(n5555) );
  OAI21_X1 U6698 ( .B1(n5665), .B2(n6121), .A(n5555), .ZN(U2961) );
  NAND2_X1 U6699 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  NAND2_X1 U6700 ( .A1(n5560), .A2(n5559), .ZN(n5561) );
  XNOR2_X1 U6701 ( .A(n5561), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5672)
         );
  AND2_X1 U6702 ( .A1(n6229), .A2(REIP_REG_24__SCAN_IN), .ZN(n5669) );
  AOI21_X1 U6703 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5669), 
        .ZN(n5562) );
  OAI21_X1 U6704 ( .B1(n6140), .B2(n5563), .A(n5562), .ZN(n5564) );
  AOI21_X1 U6705 ( .B1(n5565), .B2(n6137), .A(n5564), .ZN(n5566) );
  OAI21_X1 U6706 ( .B1(n5672), .B2(n6121), .A(n5566), .ZN(U2962) );
  AOI21_X1 U6707 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5568), .A(n5567), 
        .ZN(n5570) );
  XOR2_X1 U6708 ( .A(n5570), .B(n5569), .Z(n5690) );
  INV_X1 U6709 ( .A(n5571), .ZN(n5779) );
  AND2_X1 U6710 ( .A1(n6229), .A2(REIP_REG_22__SCAN_IN), .ZN(n5681) );
  AOI21_X1 U6711 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5681), 
        .ZN(n5572) );
  OAI21_X1 U6712 ( .B1(n6140), .B2(n5779), .A(n5572), .ZN(n5573) );
  AOI21_X1 U6713 ( .B1(n5806), .B2(n6137), .A(n5573), .ZN(n5574) );
  OAI21_X1 U6714 ( .B1(n5690), .B2(n6121), .A(n5574), .ZN(U2964) );
  AOI21_X1 U6715 ( .B1(n5577), .B2(n5576), .A(n5575), .ZN(n5697) );
  INV_X1 U6716 ( .A(n5579), .ZN(n5582) );
  INV_X1 U6717 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5580) );
  NOR2_X1 U6718 ( .A1(n6205), .A2(n5580), .ZN(n5692) );
  AOI21_X1 U6719 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5692), 
        .ZN(n5581) );
  OAI21_X1 U6720 ( .B1(n6140), .B2(n5582), .A(n5581), .ZN(n5583) );
  AOI21_X1 U6721 ( .B1(n5578), .B2(n6137), .A(n5583), .ZN(n5584) );
  OAI21_X1 U6722 ( .B1(n5697), .B2(n6121), .A(n5584), .ZN(U2965) );
  INV_X1 U6723 ( .A(n5585), .ZN(n5587) );
  NAND2_X1 U6724 ( .A1(n5587), .A2(n5586), .ZN(n5590) );
  XOR2_X1 U6725 ( .A(n5590), .B(n5589), .Z(n5728) );
  INV_X1 U6726 ( .A(n5591), .ZN(n5593) );
  AND2_X1 U6727 ( .A1(n6229), .A2(REIP_REG_19__SCAN_IN), .ZN(n5721) );
  AOI21_X1 U6728 ( .B1(n6130), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5721), 
        .ZN(n5592) );
  OAI21_X1 U6729 ( .B1(n6140), .B2(n5593), .A(n5592), .ZN(n5594) );
  AOI21_X1 U6730 ( .B1(n5595), .B2(n6137), .A(n5594), .ZN(n5596) );
  OAI21_X1 U6731 ( .B1(n5728), .B2(n6121), .A(n5596), .ZN(U2967) );
  INV_X1 U6732 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5597) );
  OAI22_X1 U6733 ( .A1(n5616), .A2(n5597), .B1(n6205), .B2(n6731), .ZN(n5599)
         );
  NOR2_X1 U6734 ( .A1(n6001), .A2(n5617), .ZN(n5598) );
  AOI211_X1 U6735 ( .C1(n6117), .C2(n5600), .A(n5599), .B(n5598), .ZN(n5601)
         );
  OAI21_X1 U6736 ( .B1(n6121), .B2(n5602), .A(n5601), .ZN(U2970) );
  AND2_X1 U6737 ( .A1(n5626), .A2(n5603), .ZN(n5604) );
  NOR2_X1 U6738 ( .A1(n5604), .A2(n3112), .ZN(n5609) );
  INV_X1 U6739 ( .A(n5605), .ZN(n5607) );
  NOR2_X1 U6740 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  XNOR2_X1 U6741 ( .A(n5609), .B(n5608), .ZN(n5846) );
  NAND2_X1 U6742 ( .A1(n5846), .A2(n6135), .ZN(n5613) );
  OAI22_X1 U6743 ( .A1(n5616), .A2(n6758), .B1(n6205), .B2(n6566), .ZN(n5610)
         );
  AOI21_X1 U6744 ( .B1(n5611), .B2(n6117), .A(n5610), .ZN(n5612) );
  OAI211_X1 U6745 ( .C1(n5617), .C2(n5614), .A(n5613), .B(n5612), .ZN(U2971)
         );
  INV_X1 U6746 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5615) );
  OAI22_X1 U6747 ( .A1(n5616), .A2(n5615), .B1(n6205), .B2(n6564), .ZN(n5619)
         );
  NOR2_X1 U6748 ( .A1(n5889), .A2(n5617), .ZN(n5618) );
  AOI211_X1 U6749 ( .C1(n6117), .C2(n5890), .A(n5619), .B(n5618), .ZN(n5620)
         );
  OAI21_X1 U6750 ( .B1(n6121), .B2(n5621), .A(n5620), .ZN(U2972) );
  OR2_X1 U6751 ( .A1(n5623), .A2(n5622), .ZN(n5625) );
  NAND2_X1 U6752 ( .A1(n5625), .A2(n5624), .ZN(n5628) );
  OAI21_X1 U6753 ( .B1(n5628), .B2(n5627), .A(n5626), .ZN(n5629) );
  INV_X1 U6754 ( .A(n5629), .ZN(n5852) );
  AOI22_X1 U6755 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5630) );
  OAI21_X1 U6756 ( .B1(n6140), .B2(n5901), .A(n5630), .ZN(n5631) );
  AOI21_X1 U6757 ( .B1(n5903), .B2(n6137), .A(n5631), .ZN(n5632) );
  OAI21_X1 U6758 ( .B1(n5852), .B2(n6121), .A(n5632), .ZN(U2973) );
  INV_X1 U6759 ( .A(n5633), .ZN(n5635) );
  AOI21_X1 U6760 ( .B1(n5635), .B2(n6247), .A(n5634), .ZN(n5636) );
  OAI21_X1 U6761 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5637), .A(n5636), 
        .ZN(n5638) );
  AOI21_X1 U6762 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5639), .A(n5638), 
        .ZN(n5640) );
  OAI21_X1 U6763 ( .B1(n5641), .B2(n6196), .A(n5640), .ZN(U2989) );
  INV_X1 U6764 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5645) );
  NOR2_X1 U6765 ( .A1(n5642), .A2(n6207), .ZN(n5643) );
  AOI211_X1 U6766 ( .C1(n5646), .C2(n5645), .A(n5644), .B(n5643), .ZN(n5649)
         );
  NAND2_X1 U6767 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U6768 ( .C1(n5650), .C2(n6196), .A(n5649), .B(n5648), .ZN(U2991)
         );
  OAI211_X1 U6769 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5661), .B(n5651), .ZN(n5654) );
  INV_X1 U6770 ( .A(n5652), .ZN(n5653) );
  OAI211_X1 U6771 ( .C1(n6207), .C2(n5759), .A(n5654), .B(n5653), .ZN(n5655)
         );
  AOI21_X1 U6772 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5662), .A(n5655), 
        .ZN(n5656) );
  OAI21_X1 U6773 ( .B1(n5657), .B2(n6196), .A(n5656), .ZN(U2992) );
  NOR2_X1 U6774 ( .A1(n5658), .A2(n6207), .ZN(n5659) );
  AOI211_X1 U6775 ( .C1(n5661), .C2(n6774), .A(n5660), .B(n5659), .ZN(n5664)
         );
  NAND2_X1 U6776 ( .A1(n5662), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5663) );
  OAI211_X1 U6777 ( .C1(n5665), .C2(n6196), .A(n5664), .B(n5663), .ZN(U2993)
         );
  AOI21_X1 U6778 ( .B1(n5677), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5666) );
  NOR2_X1 U6779 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  AOI211_X1 U6780 ( .C1(n6247), .C2(n5670), .A(n5669), .B(n5668), .ZN(n5671)
         );
  OAI21_X1 U6781 ( .B1(n5672), .B2(n6196), .A(n5671), .ZN(U2994) );
  OAI21_X1 U6782 ( .B1(n5771), .B2(n6207), .A(n5673), .ZN(n5676) );
  NOR2_X1 U6783 ( .A1(n5674), .A2(n5557), .ZN(n5675) );
  AOI211_X1 U6784 ( .C1(n5677), .C2(n5557), .A(n5676), .B(n5675), .ZN(n5678)
         );
  OAI21_X1 U6785 ( .B1(n5679), .B2(n6196), .A(n5678), .ZN(U2995) );
  INV_X1 U6786 ( .A(n5787), .ZN(n5682) );
  NOR4_X1 U6787 ( .A1(n5687), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n5683), 
        .A4(n5684), .ZN(n5680) );
  AOI211_X1 U6788 ( .C1(n6247), .C2(n5682), .A(n5681), .B(n5680), .ZN(n5689)
         );
  INV_X1 U6789 ( .A(n5683), .ZN(n5685) );
  NAND2_X1 U6790 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NOR2_X1 U6791 ( .A1(n5687), .A2(n5686), .ZN(n5691) );
  OAI21_X1 U6792 ( .B1(n5694), .B2(n5691), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5688) );
  OAI211_X1 U6793 ( .C1(n5690), .C2(n6196), .A(n5689), .B(n5688), .ZN(U2996)
         );
  AOI211_X1 U6794 ( .C1(n6247), .C2(n5693), .A(n5692), .B(n5691), .ZN(n5696)
         );
  NAND2_X1 U6795 ( .A1(n5694), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5695) );
  OAI211_X1 U6796 ( .C1(n5697), .C2(n6196), .A(n5696), .B(n5695), .ZN(U2997)
         );
  XNOR2_X1 U6797 ( .A(n5698), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5699)
         );
  XNOR2_X1 U6798 ( .A(n5700), .B(n5699), .ZN(n5814) );
  INV_X1 U6799 ( .A(n5814), .ZN(n5719) );
  NAND3_X1 U6800 ( .A1(n5703), .A2(n5702), .A3(n5701), .ZN(n5707) );
  NOR2_X1 U6801 ( .A1(n5820), .A2(n5729), .ZN(n5837) );
  AOI21_X1 U6802 ( .B1(n5705), .B2(n5837), .A(n5704), .ZN(n5706) );
  AOI21_X1 U6803 ( .B1(n5708), .B2(n5707), .A(n5706), .ZN(n5834) );
  NAND2_X1 U6804 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  OAI211_X1 U6805 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5711), .A(n5834), .B(n5710), .ZN(n5726) );
  NOR2_X1 U6806 ( .A1(n5712), .A2(n5720), .ZN(n5715) );
  NAND2_X1 U6807 ( .A1(n5713), .A2(n6742), .ZN(n5714) );
  AOI22_X1 U6808 ( .A1(n6229), .A2(REIP_REG_20__SCAN_IN), .B1(n5715), .B2(
        n5714), .ZN(n5716) );
  OAI21_X1 U6809 ( .B1(n5795), .B2(n6207), .A(n5716), .ZN(n5717) );
  AOI21_X1 U6810 ( .B1(n5726), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5717), 
        .ZN(n5718) );
  OAI21_X1 U6811 ( .B1(n5719), .B2(n6196), .A(n5718), .ZN(U2998) );
  INV_X1 U6812 ( .A(n5720), .ZN(n5722) );
  AOI21_X1 U6813 ( .B1(n5722), .B2(n6742), .A(n5721), .ZN(n5723) );
  OAI21_X1 U6814 ( .B1(n5724), .B2(n6207), .A(n5723), .ZN(n5725) );
  AOI21_X1 U6815 ( .B1(n5726), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5725), 
        .ZN(n5727) );
  OAI21_X1 U6816 ( .B1(n5728), .B2(n6196), .A(n5727), .ZN(U2999) );
  NOR2_X1 U6817 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5729), .ZN(n5835)
         );
  INV_X1 U6818 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6567) );
  NOR2_X1 U6819 ( .A1(n6205), .A2(n6567), .ZN(n5736) );
  NAND2_X1 U6820 ( .A1(n5731), .A2(n5730), .ZN(n5733) );
  NAND3_X1 U6821 ( .A1(n5819), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5822), .ZN(n5732) );
  OAI21_X1 U6822 ( .B1(n5819), .B2(n5733), .A(n5732), .ZN(n5734) );
  XNOR2_X1 U6823 ( .A(n5734), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5831)
         );
  OAI22_X1 U6824 ( .A1(n5834), .A2(n5820), .B1(n5831), .B2(n6196), .ZN(n5735)
         );
  AOI211_X1 U6825 ( .C1(n5835), .C2(n6155), .A(n5736), .B(n5735), .ZN(n5737)
         );
  OAI21_X1 U6826 ( .B1(n6207), .B2(n5887), .A(n5737), .ZN(U3001) );
  OAI211_X1 U6827 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5738), .A(n5742), .B(
        n6433), .ZN(n5739) );
  OAI21_X1 U6828 ( .B1(n5740), .B2(n5744), .A(n5739), .ZN(n5741) );
  MUX2_X1 U6829 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5741), .S(n6252), 
        .Z(U3464) );
  NOR2_X1 U6830 ( .A1(n5743), .A2(n5742), .ZN(n6255) );
  AOI21_X1 U6831 ( .B1(n5743), .B2(n5742), .A(n6255), .ZN(n5745) );
  OAI22_X1 U6832 ( .A1(n5745), .A2(n6439), .B1(n4011), .B2(n5744), .ZN(n5746)
         );
  MUX2_X1 U6833 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5746), .S(n6252), 
        .Z(U3463) );
  AND2_X1 U6834 ( .A1(n5748), .A2(n5747), .ZN(n5749) );
  INV_X2 U6835 ( .A(n6626), .ZN(n6053) );
  NOR2_X4 U6836 ( .A1(n6045), .A2(n6053), .ZN(n6047) );
  AND2_X1 U6837 ( .A1(n6047), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  OAI22_X1 U6838 ( .A1(n5047), .A2(n5989), .B1(n5751), .B2(n5977), .ZN(n5752)
         );
  AOI21_X1 U6839 ( .B1(EBX_REG_26__SCAN_IN), .B2(n5969), .A(n5752), .ZN(n5758)
         );
  INV_X1 U6840 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U6841 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5754), .ZN(n5760) );
  INV_X1 U6842 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6582) );
  OAI21_X1 U6843 ( .B1(n6580), .B2(n5760), .A(n6582), .ZN(n5756) );
  AOI22_X1 U6844 ( .A1(n5797), .A2(n5945), .B1(n5756), .B2(n5755), .ZN(n5757)
         );
  OAI211_X1 U6845 ( .C1(n5759), .C2(n5929), .A(n5758), .B(n5757), .ZN(U2801)
         );
  AOI22_X1 U6846 ( .A1(PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n5952), .B1(
        EBX_REG_25__SCAN_IN), .B2(n5969), .ZN(n5769) );
  INV_X1 U6847 ( .A(n5760), .ZN(n5761) );
  AOI22_X1 U6848 ( .A1(n5762), .A2(n5986), .B1(n5761), .B2(n6580), .ZN(n5768)
         );
  AOI22_X1 U6849 ( .A1(n5800), .A2(n5945), .B1(n5965), .B2(n5763), .ZN(n5767)
         );
  AOI21_X1 U6850 ( .B1(n5764), .B2(n5773), .A(n6580), .ZN(n5765) );
  INV_X1 U6851 ( .A(n5765), .ZN(n5766) );
  NAND4_X1 U6852 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(U2802)
         );
  NOR2_X1 U6853 ( .A1(n5580), .A2(n5770), .ZN(n5778) );
  AOI21_X1 U6854 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5778), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5772) );
  OAI22_X1 U6855 ( .A1(n5773), .A2(n5772), .B1(n5771), .B2(n5929), .ZN(n5774)
         );
  AOI22_X1 U6856 ( .A1(n5775), .A2(n5986), .B1(EBX_REG_23__SCAN_IN), .B2(n5969), .ZN(n5776) );
  OAI211_X1 U6857 ( .C1(n4996), .C2(n5989), .A(n5777), .B(n5776), .ZN(U2804)
         );
  INV_X1 U6858 ( .A(n5778), .ZN(n5782) );
  INV_X1 U6859 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6795) );
  OAI22_X1 U6860 ( .A1(n6795), .A2(n5989), .B1(n5977), .B2(n5779), .ZN(n5780)
         );
  AOI21_X1 U6861 ( .B1(n5969), .B2(EBX_REG_22__SCAN_IN), .A(n5780), .ZN(n5781)
         );
  OAI21_X1 U6862 ( .B1(n5782), .B2(REIP_REG_22__SCAN_IN), .A(n5781), .ZN(n5783) );
  AOI21_X1 U6863 ( .B1(n5806), .B2(n5945), .A(n5783), .ZN(n5786) );
  OAI21_X1 U6864 ( .B1(n5784), .B2(n5791), .A(REIP_REG_22__SCAN_IN), .ZN(n5785) );
  OAI211_X1 U6865 ( .C1(n5929), .C2(n5787), .A(n5786), .B(n5785), .ZN(U2805)
         );
  OAI22_X1 U6866 ( .A1(n5817), .A2(n5977), .B1(n3904), .B2(n5994), .ZN(n5788)
         );
  AOI21_X1 U6867 ( .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n5952), .A(n5788), 
        .ZN(n5794) );
  OAI21_X1 U6868 ( .B1(n5790), .B2(n5789), .A(n6572), .ZN(n5792) );
  AOI22_X1 U6869 ( .A1(n5813), .A2(n5945), .B1(n5792), .B2(n5791), .ZN(n5793)
         );
  OAI211_X1 U6870 ( .C1(n5795), .C2(n5929), .A(n5794), .B(n5793), .ZN(U2807)
         );
  AOI22_X1 U6871 ( .A1(n5797), .A2(n6003), .B1(n6002), .B2(DATAI_26_), .ZN(
        n5799) );
  AOI22_X1 U6872 ( .A1(n6006), .A2(DATAI_10_), .B1(n6005), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U6873 ( .A1(n5799), .A2(n5798), .ZN(U2865) );
  AOI22_X1 U6874 ( .A1(n5800), .A2(n6003), .B1(n6002), .B2(DATAI_25_), .ZN(
        n5802) );
  AOI22_X1 U6875 ( .A1(n6006), .A2(DATAI_9_), .B1(n6005), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U6876 ( .A1(n5802), .A2(n5801), .ZN(U2866) );
  AOI22_X1 U6877 ( .A1(n5803), .A2(n6003), .B1(n6002), .B2(DATAI_23_), .ZN(
        n5805) );
  AOI22_X1 U6878 ( .A1(n6006), .A2(DATAI_7_), .B1(n6005), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U6879 ( .A1(n5805), .A2(n5804), .ZN(U2868) );
  AOI22_X1 U6880 ( .A1(n5806), .A2(n6003), .B1(n6002), .B2(DATAI_22_), .ZN(
        n5808) );
  AOI22_X1 U6881 ( .A1(n6006), .A2(DATAI_6_), .B1(n6005), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U6882 ( .A1(n5808), .A2(n5807), .ZN(U2869) );
  AOI22_X1 U6883 ( .A1(n5578), .A2(n6003), .B1(n6002), .B2(DATAI_21_), .ZN(
        n5810) );
  AOI22_X1 U6884 ( .A1(n6006), .A2(DATAI_5_), .B1(n6005), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6885 ( .A1(n5810), .A2(n5809), .ZN(U2870) );
  AOI22_X1 U6886 ( .A1(n5813), .A2(n6003), .B1(n6002), .B2(DATAI_20_), .ZN(
        n5812) );
  AOI22_X1 U6887 ( .A1(n6006), .A2(DATAI_4_), .B1(n6005), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U6888 ( .A1(n5812), .A2(n5811), .ZN(U2871) );
  AOI22_X1 U6889 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_20__SCAN_IN), .ZN(n5816) );
  AOI22_X1 U6890 ( .A1(n5814), .A2(n6135), .B1(n5813), .B2(n6137), .ZN(n5815)
         );
  OAI211_X1 U6891 ( .C1(n6140), .C2(n5817), .A(n5816), .B(n5815), .ZN(U2966)
         );
  AOI22_X1 U6892 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_18__SCAN_IN), .ZN(n5827) );
  NOR2_X1 U6893 ( .A1(n5819), .A2(n5818), .ZN(n5824) );
  NOR2_X1 U6894 ( .A1(n5821), .A2(n5820), .ZN(n5823) );
  MUX2_X1 U6895 ( .A(n5824), .B(n5823), .S(n5822), .Z(n5825) );
  XOR2_X1 U6896 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5825), .Z(n5833) );
  AOI22_X1 U6897 ( .A1(n5833), .A2(n6135), .B1(n6137), .B2(n5995), .ZN(n5826)
         );
  OAI211_X1 U6898 ( .C1(n6140), .C2(n5828), .A(n5827), .B(n5826), .ZN(U2968)
         );
  AOI22_X1 U6899 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n5830) );
  AOI22_X1 U6900 ( .A1(n5998), .A2(n6137), .B1(n5881), .B2(n6117), .ZN(n5829)
         );
  OAI211_X1 U6901 ( .C1(n5831), .C2(n6121), .A(n5830), .B(n5829), .ZN(U2969)
         );
  AOI22_X1 U6902 ( .A1(n5833), .A2(n6240), .B1(n6247), .B2(n5832), .ZN(n5841)
         );
  NAND2_X1 U6903 ( .A1(n6229), .A2(REIP_REG_18__SCAN_IN), .ZN(n5840) );
  INV_X1 U6904 ( .A(n5834), .ZN(n5836) );
  OAI221_X1 U6905 ( .B1(n5836), .B2(n6143), .C1(n5836), .C2(n5835), .A(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5839) );
  INV_X1 U6906 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6790) );
  NAND3_X1 U6907 ( .A1(n5837), .A2(n6790), .A3(n6155), .ZN(n5838) );
  NAND4_X1 U6908 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(U3000)
         );
  INV_X1 U6909 ( .A(n5842), .ZN(n5848) );
  OAI22_X1 U6910 ( .A1(n5843), .A2(n6207), .B1(n6566), .B2(n6205), .ZN(n5844)
         );
  AOI211_X1 U6911 ( .C1(n5846), .C2(n6240), .A(n5845), .B(n5844), .ZN(n5847)
         );
  OAI21_X1 U6912 ( .B1(n5848), .B2(n6914), .A(n5847), .ZN(U3003) );
  NOR2_X1 U6913 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5849), .ZN(n5856)
         );
  NOR4_X1 U6914 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6245), .A3(n5851), 
        .A4(n5850), .ZN(n5854) );
  OAI22_X1 U6915 ( .A1(n5852), .A2(n6196), .B1(n6207), .B2(n5898), .ZN(n5853)
         );
  AOI211_X1 U6916 ( .C1(REIP_REG_13__SCAN_IN), .C2(n6229), .A(n5854), .B(n5853), .ZN(n5855) );
  OAI21_X1 U6917 ( .B1(n5857), .B2(n5856), .A(n5855), .ZN(U3005) );
  INV_X1 U6918 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6534) );
  AOI21_X1 U6919 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6534), .A(n6538), .ZN(n5859) );
  INV_X1 U6920 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6681) );
  AOI21_X1 U6921 ( .B1(n5859), .B2(n6681), .A(n6629), .ZN(U2789) );
  NOR2_X1 U6922 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5860) );
  OAI21_X1 U6923 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5860), .A(n6589), .ZN(n5858)
         );
  OAI21_X1 U6924 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6589), .A(n5858), .ZN(
        U2791) );
  OAI21_X1 U6925 ( .B1(BS16_N), .B2(n5860), .A(n6599), .ZN(n6597) );
  OAI21_X1 U6926 ( .B1(n6599), .B2(n5861), .A(n6597), .ZN(U2792) );
  OAI21_X1 U6927 ( .B1(n5862), .B2(n6826), .A(n6121), .ZN(U2793) );
  NOR4_X1 U6928 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n5866) );
  NOR4_X1 U6929 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(
        DATAWIDTH_REG_13__SCAN_IN), .A3(DATAWIDTH_REG_14__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n5865) );
  NOR4_X1 U6930 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5864) );
  NOR4_X1 U6931 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5863) );
  NAND4_X1 U6932 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n5872)
         );
  NOR4_X1 U6933 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5870)
         );
  AOI211_X1 U6934 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_5__SCAN_IN), .B(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n5869) );
  NOR4_X1 U6935 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n5868) );
  NOR4_X1 U6936 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(n5867) );
  NAND4_X1 U6937 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(n5871)
         );
  NOR2_X1 U6938 ( .A1(n5872), .A2(n5871), .ZN(n6615) );
  INV_X1 U6939 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5874) );
  NOR3_X1 U6940 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5875) );
  OAI21_X1 U6941 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5875), .A(n6615), .ZN(n5873)
         );
  OAI21_X1 U6942 ( .B1(n6615), .B2(n5874), .A(n5873), .ZN(U2794) );
  INV_X1 U6943 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6598) );
  AOI21_X1 U6944 ( .B1(n6745), .B2(n6598), .A(n5875), .ZN(n5877) );
  INV_X1 U6945 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5876) );
  INV_X1 U6946 ( .A(n6615), .ZN(n6612) );
  AOI22_X1 U6947 ( .A1(n6615), .A2(n5877), .B1(n5876), .B2(n6612), .ZN(U2795)
         );
  AOI221_X1 U6948 ( .B1(n5880), .B2(n6567), .C1(n5879), .C2(n6567), .A(n5878), 
        .ZN(n5885) );
  AOI22_X1 U6949 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n5952), .B1(n5881), 
        .B2(n5986), .ZN(n5882) );
  OAI211_X1 U6950 ( .C1(n5994), .C2(n5883), .A(n5971), .B(n5882), .ZN(n5884)
         );
  AOI211_X1 U6951 ( .C1(n5998), .C2(n5945), .A(n5885), .B(n5884), .ZN(n5886)
         );
  OAI21_X1 U6952 ( .B1(n5929), .B2(n5887), .A(n5886), .ZN(U2810) );
  AOI22_X1 U6953 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n5952), .B1(
        EBX_REG_14__SCAN_IN), .B2(n5969), .ZN(n5897) );
  AOI21_X1 U6954 ( .B1(n5888), .B2(n5965), .A(n5953), .ZN(n5896) );
  INV_X1 U6955 ( .A(n5889), .ZN(n5891) );
  AOI22_X1 U6956 ( .A1(n5891), .A2(n5945), .B1(n5986), .B2(n5890), .ZN(n5895)
         );
  OAI21_X1 U6957 ( .B1(REIP_REG_14__SCAN_IN), .B2(n5893), .A(n5892), .ZN(n5894) );
  NAND4_X1 U6958 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(U2813)
         );
  OAI22_X1 U6959 ( .A1(n5899), .A2(n5994), .B1(n5929), .B2(n5898), .ZN(n5900)
         );
  AOI211_X1 U6960 ( .C1(n5952), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5953), 
        .B(n5900), .ZN(n5908) );
  INV_X1 U6961 ( .A(n5901), .ZN(n5902) );
  AOI22_X1 U6962 ( .A1(n5903), .A2(n5945), .B1(n5902), .B2(n5986), .ZN(n5907)
         );
  OAI21_X1 U6963 ( .B1(n5904), .B2(n5909), .A(REIP_REG_13__SCAN_IN), .ZN(n5906) );
  INV_X1 U6964 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6562) );
  NAND4_X1 U6965 ( .A1(n5979), .A2(REIP_REG_12__SCAN_IN), .A3(n5910), .A4(
        n6562), .ZN(n5905) );
  NAND4_X1 U6966 ( .A1(n5908), .A2(n5907), .A3(n5906), .A4(n5905), .ZN(U2814)
         );
  AOI22_X1 U6967 ( .A1(n5965), .A2(n6152), .B1(REIP_REG_11__SCAN_IN), .B2(
        n5909), .ZN(n5916) );
  OR2_X1 U6968 ( .A1(n5967), .A2(n5910), .ZN(n5911) );
  OAI22_X1 U6969 ( .A1(n6787), .A2(n5994), .B1(n5912), .B2(n5911), .ZN(n5913)
         );
  AOI211_X1 U6970 ( .C1(n5952), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5953), 
        .B(n5913), .ZN(n5915) );
  AOI22_X1 U6971 ( .A1(n6118), .A2(n5945), .B1(n5986), .B2(n6116), .ZN(n5914)
         );
  NAND3_X1 U6972 ( .A1(n5916), .A2(n5915), .A3(n5914), .ZN(U2816) );
  AOI22_X1 U6973 ( .A1(n5965), .A2(n5918), .B1(REIP_REG_9__SCAN_IN), .B2(n5917), .ZN(n5927) );
  NAND2_X1 U6974 ( .A1(n5979), .A2(n5919), .ZN(n5920) );
  OAI22_X1 U6975 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5920), .B1(n6707), .B2(n5994), .ZN(n5921) );
  AOI211_X1 U6976 ( .C1(n5952), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5953), 
        .B(n5921), .ZN(n5926) );
  INV_X1 U6977 ( .A(n5922), .ZN(n5924) );
  AOI22_X1 U6978 ( .A1(n5924), .A2(n5945), .B1(n5986), .B2(n5923), .ZN(n5925)
         );
  NAND3_X1 U6979 ( .A1(n5927), .A2(n5926), .A3(n5925), .ZN(U2818) );
  OAI22_X1 U6980 ( .A1(n6732), .A2(n5994), .B1(n5929), .B2(n5928), .ZN(n5930)
         );
  AOI211_X1 U6981 ( .C1(n5952), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5953), 
        .B(n5930), .ZN(n5941) );
  INV_X1 U6982 ( .A(n5931), .ZN(n5932) );
  AOI22_X1 U6983 ( .A1(n5933), .A2(n5945), .B1(n5932), .B2(n5986), .ZN(n5940)
         );
  INV_X1 U6984 ( .A(n5936), .ZN(n5935) );
  OAI21_X1 U6985 ( .B1(n5935), .B2(n5967), .A(n5934), .ZN(n5958) );
  NOR3_X1 U6986 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5967), .A3(n5936), .ZN(n5942)
         );
  OAI21_X1 U6987 ( .B1(n5958), .B2(n5942), .A(REIP_REG_7__SCAN_IN), .ZN(n5939)
         );
  INV_X1 U6988 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6555) );
  NAND3_X1 U6989 ( .A1(n5979), .A2(n5937), .A3(n6555), .ZN(n5938) );
  NAND4_X1 U6990 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(U2820)
         );
  AOI211_X1 U6991 ( .C1(n5969), .C2(EBX_REG_6__SCAN_IN), .A(n5953), .B(n5942), 
        .ZN(n5949) );
  INV_X1 U6992 ( .A(n5943), .ZN(n6182) );
  AOI22_X1 U6993 ( .A1(n5965), .A2(n6182), .B1(REIP_REG_6__SCAN_IN), .B2(n5958), .ZN(n5948) );
  INV_X1 U6994 ( .A(n5944), .ZN(n5946) );
  AOI22_X1 U6995 ( .A1(n5946), .A2(n5945), .B1(PHYADDRPOINTER_REG_6__SCAN_IN), 
        .B2(n5952), .ZN(n5947) );
  AND3_X1 U6996 ( .A1(n5949), .A2(n5948), .A3(n5947), .ZN(n5950) );
  OAI21_X1 U6997 ( .B1(n5951), .B2(n5977), .A(n5950), .ZN(U2821) );
  AOI22_X1 U6998 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n5952), .B1(
        EBX_REG_5__SCAN_IN), .B2(n5969), .ZN(n5963) );
  AOI21_X1 U6999 ( .B1(n5965), .B2(n5954), .A(n5953), .ZN(n5962) );
  INV_X1 U7000 ( .A(n5955), .ZN(n5957) );
  AOI22_X1 U7001 ( .A1(n5957), .A2(n5991), .B1(n5956), .B2(n5986), .ZN(n5961)
         );
  OAI221_X1 U7002 ( .B1(REIP_REG_5__SCAN_IN), .B2(n5979), .C1(
        REIP_REG_5__SCAN_IN), .C2(n5959), .A(n5958), .ZN(n5960) );
  NAND4_X1 U7003 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(U2822)
         );
  AOI22_X1 U7004 ( .A1(n5965), .A2(n6195), .B1(REIP_REG_4__SCAN_IN), .B2(n5964), .ZN(n5976) );
  NOR3_X1 U7005 ( .A1(n5967), .A2(REIP_REG_4__SCAN_IN), .A3(n5966), .ZN(n5973)
         );
  AOI22_X1 U7006 ( .A1(EBX_REG_4__SCAN_IN), .A2(n5969), .B1(n5968), .B2(n5984), 
        .ZN(n5970) );
  OAI211_X1 U7007 ( .C1(n5989), .C2(n6794), .A(n5971), .B(n5970), .ZN(n5972)
         );
  AOI211_X1 U7008 ( .C1(n5974), .C2(n5991), .A(n5973), .B(n5972), .ZN(n5975)
         );
  OAI211_X1 U7009 ( .C1(n5978), .C2(n5977), .A(n5976), .B(n5975), .ZN(U2823)
         );
  AOI22_X1 U7010 ( .A1(n5981), .A2(n5980), .B1(n5979), .B2(n6745), .ZN(n5993)
         );
  INV_X1 U7011 ( .A(n5982), .ZN(n6136) );
  INV_X1 U7012 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6677) );
  NAND2_X1 U7013 ( .A1(n5984), .A2(n5983), .ZN(n5988) );
  AOI22_X1 U7014 ( .A1(n5986), .A2(n6677), .B1(n5985), .B2(REIP_REG_1__SCAN_IN), .ZN(n5987) );
  OAI211_X1 U7015 ( .C1(n6677), .C2(n5989), .A(n5988), .B(n5987), .ZN(n5990)
         );
  AOI21_X1 U7016 ( .B1(n6136), .B2(n5991), .A(n5990), .ZN(n5992) );
  OAI211_X1 U7017 ( .C1(n6878), .C2(n5994), .A(n5993), .B(n5992), .ZN(U2826)
         );
  AOI22_X1 U7018 ( .A1(n5995), .A2(n6003), .B1(n6002), .B2(DATAI_18_), .ZN(
        n5997) );
  AOI22_X1 U7019 ( .A1(n6006), .A2(DATAI_2_), .B1(n6005), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5996) );
  NAND2_X1 U7020 ( .A1(n5997), .A2(n5996), .ZN(U2873) );
  AOI22_X1 U7021 ( .A1(n5998), .A2(n6003), .B1(n6002), .B2(DATAI_17_), .ZN(
        n6000) );
  AOI22_X1 U7022 ( .A1(n6006), .A2(DATAI_1_), .B1(n6005), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7023 ( .A1(n6000), .A2(n5999), .ZN(U2874) );
  INV_X1 U7024 ( .A(n6001), .ZN(n6004) );
  AOI22_X1 U7025 ( .A1(n6004), .A2(n6003), .B1(n6002), .B2(DATAI_16_), .ZN(
        n6008) );
  AOI22_X1 U7026 ( .A1(n6006), .A2(DATAI_0_), .B1(n6005), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7027 ( .A1(n6008), .A2(n6007), .ZN(U2875) );
  INV_X1 U7028 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6907) );
  NAND2_X1 U7029 ( .A1(n6045), .A2(n6009), .ZN(n6025) );
  AOI22_X1 U7030 ( .A1(DATAO_REG_30__SCAN_IN), .A2(n6047), .B1(n6053), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6010) );
  OAI21_X1 U7031 ( .B1(n6907), .B2(n6025), .A(n6010), .ZN(U2893) );
  INV_X1 U7032 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6012) );
  AOI22_X1 U7033 ( .A1(n6053), .A2(UWORD_REG_13__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n6011) );
  OAI21_X1 U7034 ( .B1(n6012), .B2(n6025), .A(n6011), .ZN(U2894) );
  INV_X1 U7035 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6070) );
  AOI22_X1 U7036 ( .A1(n6053), .A2(UWORD_REG_12__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n6013) );
  OAI21_X1 U7037 ( .B1(n6070), .B2(n6025), .A(n6013), .ZN(U2895) );
  AOI22_X1 U7038 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6029), .B1(n6047), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n6014) );
  OAI21_X1 U7039 ( .B1(n6858), .B2(n6626), .A(n6014), .ZN(U2896) );
  AOI22_X1 U7040 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6029), .B1(n6047), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n6015) );
  OAI21_X1 U7041 ( .B1(n6713), .B2(n6626), .A(n6015), .ZN(U2897) );
  INV_X1 U7042 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6921) );
  AOI22_X1 U7043 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6029), .B1(n6053), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6016) );
  OAI21_X1 U7044 ( .B1(n6921), .B2(n6039), .A(n6016), .ZN(U2898) );
  INV_X1 U7045 ( .A(EAX_REG_24__SCAN_IN), .ZN(n6066) );
  AOI22_X1 U7046 ( .A1(n6053), .A2(UWORD_REG_8__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n6017) );
  OAI21_X1 U7047 ( .B1(n6066), .B2(n6025), .A(n6017), .ZN(U2899) );
  INV_X1 U7048 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6019) );
  AOI22_X1 U7049 ( .A1(n6053), .A2(UWORD_REG_7__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n6018) );
  OAI21_X1 U7050 ( .B1(n6019), .B2(n6025), .A(n6018), .ZN(U2900) );
  INV_X1 U7051 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6813) );
  INV_X1 U7052 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6726) );
  INV_X1 U7053 ( .A(UWORD_REG_6__SCAN_IN), .ZN(n6020) );
  OAI222_X1 U7054 ( .A1(n6039), .A2(n6813), .B1(n6025), .B2(n6726), .C1(n6626), 
        .C2(n6020), .ZN(U2901) );
  INV_X1 U7055 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6022) );
  AOI22_X1 U7056 ( .A1(n6053), .A2(UWORD_REG_5__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n6021) );
  OAI21_X1 U7057 ( .B1(n6022), .B2(n6025), .A(n6021), .ZN(U2902) );
  INV_X1 U7058 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n6710) );
  AOI22_X1 U7059 ( .A1(EAX_REG_20__SCAN_IN), .A2(n6029), .B1(n6047), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n6023) );
  OAI21_X1 U7060 ( .B1(n6710), .B2(n6626), .A(n6023), .ZN(U2903) );
  INV_X1 U7061 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6026) );
  AOI22_X1 U7062 ( .A1(n6053), .A2(UWORD_REG_3__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n6024) );
  OAI21_X1 U7063 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(U2904) );
  INV_X1 U7064 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U7065 ( .A1(EAX_REG_18__SCAN_IN), .A2(n6029), .B1(n6053), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n6027) );
  OAI21_X1 U7066 ( .B1(n6824), .B2(n6039), .A(n6027), .ZN(U2905) );
  AOI22_X1 U7067 ( .A1(EAX_REG_17__SCAN_IN), .A2(n6029), .B1(n6047), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7068 ( .B1(n6876), .B2(n6626), .A(n6028), .ZN(U2906) );
  AOI22_X1 U7069 ( .A1(EAX_REG_16__SCAN_IN), .A2(n6029), .B1(n6047), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n6030) );
  OAI21_X1 U7070 ( .B1(n6849), .B2(n6626), .A(n6030), .ZN(U2907) );
  AOI22_X1 U7071 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6045), .B1(n6047), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6031) );
  OAI21_X1 U7072 ( .B1(n6724), .B2(n6626), .A(n6031), .ZN(U2908) );
  INV_X1 U7073 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6109) );
  AOI22_X1 U7074 ( .A1(n6053), .A2(LWORD_REG_14__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6032) );
  OAI21_X1 U7075 ( .B1(n6109), .B2(n6055), .A(n6032), .ZN(U2909) );
  INV_X1 U7076 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6034) );
  AOI22_X1 U7077 ( .A1(n6053), .A2(LWORD_REG_13__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U7078 ( .B1(n6034), .B2(n6055), .A(n6033), .ZN(U2910) );
  INV_X1 U7079 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6100) );
  AOI22_X1 U7080 ( .A1(n6053), .A2(LWORD_REG_12__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6035) );
  OAI21_X1 U7081 ( .B1(n6100), .B2(n6055), .A(n6035), .ZN(U2911) );
  INV_X1 U7082 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6097) );
  AOI22_X1 U7083 ( .A1(n6053), .A2(LWORD_REG_11__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6036) );
  OAI21_X1 U7084 ( .B1(n6097), .B2(n6055), .A(n6036), .ZN(U2912) );
  INV_X1 U7085 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7086 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6045), .B1(n6053), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6037) );
  OAI21_X1 U7087 ( .B1(n6683), .B2(n6039), .A(n6037), .ZN(U2913) );
  INV_X1 U7088 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7089 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6045), .B1(n6053), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6038) );
  OAI21_X1 U7090 ( .B1(n6751), .B2(n6039), .A(n6038), .ZN(U2914) );
  INV_X1 U7091 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6089) );
  AOI22_X1 U7092 ( .A1(n6053), .A2(LWORD_REG_8__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6040) );
  OAI21_X1 U7093 ( .B1(n6089), .B2(n6055), .A(n6040), .ZN(U2915) );
  AOI22_X1 U7094 ( .A1(n6053), .A2(LWORD_REG_7__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6041) );
  OAI21_X1 U7095 ( .B1(n3495), .B2(n6055), .A(n6041), .ZN(U2916) );
  AOI22_X1 U7096 ( .A1(n6053), .A2(LWORD_REG_6__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6042) );
  OAI21_X1 U7097 ( .B1(n3478), .B2(n6055), .A(n6042), .ZN(U2917) );
  AOI22_X1 U7098 ( .A1(n6053), .A2(LWORD_REG_5__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6043) );
  OAI21_X1 U7099 ( .B1(n6044), .B2(n6055), .A(n6043), .ZN(U2918) );
  INV_X1 U7100 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7101 ( .A1(EAX_REG_4__SCAN_IN), .A2(n6045), .B1(n6047), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6046) );
  OAI21_X1 U7102 ( .B1(n6743), .B2(n6626), .A(n6046), .ZN(U2919) );
  AOI22_X1 U7103 ( .A1(n6053), .A2(LWORD_REG_3__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6048) );
  OAI21_X1 U7104 ( .B1(n6690), .B2(n6055), .A(n6048), .ZN(U2920) );
  AOI22_X1 U7105 ( .A1(n6053), .A2(LWORD_REG_2__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7106 ( .B1(n6050), .B2(n6055), .A(n6049), .ZN(U2921) );
  AOI22_X1 U7107 ( .A1(n6053), .A2(LWORD_REG_1__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6051) );
  OAI21_X1 U7108 ( .B1(n6052), .B2(n6055), .A(n6051), .ZN(U2922) );
  AOI22_X1 U7109 ( .A1(n6053), .A2(LWORD_REG_0__SCAN_IN), .B1(n6047), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U7110 ( .B1(n6056), .B2(n6055), .A(n6054), .ZN(U2923) );
  AOI22_X1 U7111 ( .A1(n6102), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6101), .ZN(n6058) );
  OAI21_X1 U7112 ( .B1(n6104), .B2(n6079), .A(n6058), .ZN(U2926) );
  AOI22_X1 U7113 ( .A1(n6106), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6101), .ZN(n6059) );
  OAI21_X1 U7114 ( .B1(n6104), .B2(n6894), .A(n6059), .ZN(U2927) );
  AOI22_X1 U7115 ( .A1(n6102), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6101), .ZN(n6060) );
  OAI21_X1 U7116 ( .B1(n6104), .B2(n6808), .A(n6060), .ZN(U2928) );
  AOI22_X1 U7117 ( .A1(n6102), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6101), .ZN(n6061) );
  OAI21_X1 U7118 ( .B1(n6104), .B2(n6693), .A(n6061), .ZN(U2929) );
  AOI22_X1 U7119 ( .A1(n6102), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6101), .ZN(n6062) );
  OAI21_X1 U7120 ( .B1(n6104), .B2(n6084), .A(n6062), .ZN(U2930) );
  AOI22_X1 U7121 ( .A1(n6102), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6101), .ZN(n6063) );
  OAI21_X1 U7122 ( .B1(n6104), .B2(n6086), .A(n6063), .ZN(U2931) );
  INV_X1 U7123 ( .A(DATAI_8_), .ZN(n6064) );
  NOR2_X1 U7124 ( .A1(n6104), .A2(n6064), .ZN(n6087) );
  AOI21_X1 U7125 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n6106), .A(n6087), .ZN(n6065) );
  OAI21_X1 U7126 ( .B1(n6066), .B2(n6108), .A(n6065), .ZN(U2932) );
  AOI22_X1 U7127 ( .A1(n6102), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n6101), .ZN(n6067) );
  NAND2_X1 U7128 ( .A1(n6092), .A2(DATAI_9_), .ZN(n6090) );
  NAND2_X1 U7129 ( .A1(n6067), .A2(n6090), .ZN(U2933) );
  INV_X1 U7130 ( .A(DATAI_12_), .ZN(n6068) );
  NOR2_X1 U7131 ( .A1(n6104), .A2(n6068), .ZN(n6098) );
  AOI21_X1 U7132 ( .B1(UWORD_REG_12__SCAN_IN), .B2(n6106), .A(n6098), .ZN(
        n6069) );
  OAI21_X1 U7133 ( .B1(n6070), .B2(n6108), .A(n6069), .ZN(U2936) );
  INV_X1 U7134 ( .A(DATAI_13_), .ZN(n6832) );
  AOI22_X1 U7135 ( .A1(n6102), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n6101), .ZN(n6071) );
  OAI21_X1 U7136 ( .B1(n6104), .B2(n6832), .A(n6071), .ZN(U2937) );
  INV_X1 U7137 ( .A(DATAI_14_), .ZN(n6072) );
  NOR2_X1 U7138 ( .A1(n6104), .A2(n6072), .ZN(n6105) );
  AOI21_X1 U7139 ( .B1(UWORD_REG_14__SCAN_IN), .B2(n6106), .A(n6105), .ZN(
        n6073) );
  OAI21_X1 U7140 ( .B1(n6907), .B2(n6108), .A(n6073), .ZN(U2938) );
  AOI22_X1 U7141 ( .A1(n6102), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6101), .ZN(n6074) );
  OAI21_X1 U7142 ( .B1(n6104), .B2(n6075), .A(n6074), .ZN(U2939) );
  AOI22_X1 U7143 ( .A1(n6106), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6101), .ZN(n6076) );
  OAI21_X1 U7144 ( .B1(n6104), .B2(n6077), .A(n6076), .ZN(U2940) );
  AOI22_X1 U7145 ( .A1(n6106), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6101), .ZN(n6078) );
  OAI21_X1 U7146 ( .B1(n6104), .B2(n6079), .A(n6078), .ZN(U2941) );
  AOI22_X1 U7147 ( .A1(n6106), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6101), .ZN(n6080) );
  OAI21_X1 U7148 ( .B1(n6104), .B2(n6894), .A(n6080), .ZN(U2942) );
  AOI22_X1 U7149 ( .A1(n6102), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6101), .ZN(n6081) );
  OAI21_X1 U7150 ( .B1(n6104), .B2(n6808), .A(n6081), .ZN(U2943) );
  AOI22_X1 U7151 ( .A1(n6102), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6101), .ZN(n6082) );
  OAI21_X1 U7152 ( .B1(n6104), .B2(n6693), .A(n6082), .ZN(U2944) );
  AOI22_X1 U7153 ( .A1(n6102), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6101), .ZN(n6083) );
  OAI21_X1 U7154 ( .B1(n6104), .B2(n6084), .A(n6083), .ZN(U2945) );
  AOI22_X1 U7155 ( .A1(n6102), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6101), .ZN(n6085) );
  OAI21_X1 U7156 ( .B1(n6104), .B2(n6086), .A(n6085), .ZN(U2946) );
  AOI21_X1 U7157 ( .B1(LWORD_REG_8__SCAN_IN), .B2(n6106), .A(n6087), .ZN(n6088) );
  OAI21_X1 U7158 ( .B1(n6089), .B2(n6108), .A(n6088), .ZN(U2947) );
  AOI22_X1 U7159 ( .A1(n6102), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n6101), .ZN(n6091) );
  NAND2_X1 U7160 ( .A1(n6091), .A2(n6090), .ZN(U2948) );
  AOI22_X1 U7161 ( .A1(n6106), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n6101), .ZN(n6094) );
  NAND2_X1 U7162 ( .A1(n6092), .A2(DATAI_10_), .ZN(n6093) );
  NAND2_X1 U7163 ( .A1(n6094), .A2(n6093), .ZN(U2949) );
  AOI21_X1 U7164 ( .B1(LWORD_REG_11__SCAN_IN), .B2(n6106), .A(n6095), .ZN(
        n6096) );
  OAI21_X1 U7165 ( .B1(n6097), .B2(n6108), .A(n6096), .ZN(U2950) );
  AOI21_X1 U7166 ( .B1(LWORD_REG_12__SCAN_IN), .B2(n6106), .A(n6098), .ZN(
        n6099) );
  OAI21_X1 U7167 ( .B1(n6100), .B2(n6108), .A(n6099), .ZN(U2951) );
  AOI22_X1 U7168 ( .A1(n6102), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n6101), .ZN(n6103) );
  OAI21_X1 U7169 ( .B1(n6104), .B2(n6832), .A(n6103), .ZN(U2952) );
  AOI21_X1 U7170 ( .B1(LWORD_REG_14__SCAN_IN), .B2(n6106), .A(n6105), .ZN(
        n6107) );
  OAI21_X1 U7171 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(U2953) );
  NAND2_X1 U7172 ( .A1(n6111), .A2(n6110), .ZN(n6115) );
  AND2_X1 U7173 ( .A1(n6113), .A2(n6112), .ZN(n6114) );
  XOR2_X1 U7174 ( .A(n6115), .B(n6114), .Z(n6159) );
  AOI22_X1 U7175 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_11__SCAN_IN), .ZN(n6120) );
  AOI22_X1 U7176 ( .A1(n6118), .A2(n6137), .B1(n6117), .B2(n6116), .ZN(n6119)
         );
  OAI211_X1 U7177 ( .C1(n6159), .C2(n6121), .A(n6120), .B(n6119), .ZN(U2975)
         );
  AOI22_X1 U7178 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7179 ( .A1(n6123), .A2(n6122), .ZN(n6124) );
  XOR2_X1 U7180 ( .A(n6125), .B(n6124), .Z(n6222) );
  AOI22_X1 U7181 ( .A1(n6222), .A2(n6135), .B1(n6137), .B2(n6126), .ZN(n6127)
         );
  OAI211_X1 U7182 ( .C1(n6140), .C2(n6129), .A(n6128), .B(n6127), .ZN(U2984)
         );
  AOI22_X1 U7183 ( .A1(n6130), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6229), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n6139) );
  OAI21_X1 U7184 ( .B1(n6133), .B2(n6132), .A(n6131), .ZN(n6134) );
  INV_X1 U7185 ( .A(n6134), .ZN(n6234) );
  AOI22_X1 U7186 ( .A1(n6137), .A2(n6136), .B1(n6234), .B2(n6135), .ZN(n6138)
         );
  OAI211_X1 U7187 ( .C1(PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n6140), .A(n6139), 
        .B(n6138), .ZN(U2985) );
  AOI21_X1 U7188 ( .B1(n6142), .B2(n6247), .A(n6141), .ZN(n6150) );
  OAI21_X1 U7189 ( .B1(n6143), .B2(n6221), .A(n6156), .ZN(n6145) );
  AOI21_X1 U7190 ( .B1(n6151), .B2(n6145), .A(n6144), .ZN(n6146) );
  AOI21_X1 U7191 ( .B1(n6147), .B2(n6240), .A(n6146), .ZN(n6149) );
  NAND3_X1 U7192 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6144), .A3(n6155), .ZN(n6148) );
  NAND3_X1 U7193 ( .A1(n6150), .A2(n6149), .A3(n6148), .ZN(U3006) );
  INV_X1 U7194 ( .A(n6151), .ZN(n6157) );
  INV_X1 U7195 ( .A(n6152), .ZN(n6153) );
  OAI22_X1 U7196 ( .A1(n6153), .A2(n6207), .B1(n6560), .B2(n6205), .ZN(n6154)
         );
  AOI221_X1 U7197 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6157), .C1(
        n6156), .C2(n6155), .A(n6154), .ZN(n6158) );
  OAI21_X1 U7198 ( .B1(n6159), .B2(n6196), .A(n6158), .ZN(U3007) );
  AOI22_X1 U7199 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6161), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n6160), .ZN(n6169) );
  INV_X1 U7200 ( .A(n6162), .ZN(n6164) );
  AOI21_X1 U7201 ( .B1(n6164), .B2(n6247), .A(n6163), .ZN(n6168) );
  AOI22_X1 U7202 ( .A1(n6166), .A2(n6240), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6165), .ZN(n6167) );
  OAI211_X1 U7203 ( .C1(n6170), .C2(n6169), .A(n6168), .B(n6167), .ZN(U3008)
         );
  OAI21_X1 U7204 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6171), .ZN(n6179) );
  NAND2_X1 U7205 ( .A1(n6172), .A2(n6240), .ZN(n6177) );
  OAI22_X1 U7206 ( .A1(n6173), .A2(n6207), .B1(n6556), .B2(n6205), .ZN(n6174)
         );
  AOI21_X1 U7207 ( .B1(n6175), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6174), 
        .ZN(n6176) );
  AND2_X1 U7208 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  OAI21_X1 U7209 ( .B1(n6180), .B2(n6179), .A(n6178), .ZN(U3010) );
  INV_X1 U7210 ( .A(n6181), .ZN(n6190) );
  NAND2_X1 U7211 ( .A1(n6247), .A2(n6182), .ZN(n6184) );
  OAI211_X1 U7212 ( .C1(n6185), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n6184), 
        .B(n6183), .ZN(n6186) );
  AOI21_X1 U7213 ( .B1(n6187), .B2(n6240), .A(n6186), .ZN(n6188) );
  OAI21_X1 U7214 ( .B1(n6190), .B2(n6189), .A(n6188), .ZN(U3012) );
  INV_X1 U7215 ( .A(n6217), .ZN(n6191) );
  AOI21_X1 U7216 ( .B1(n6221), .B2(n6191), .A(n6223), .ZN(n6216) );
  NAND2_X1 U7217 ( .A1(n6217), .A2(n6192), .ZN(n6212) );
  OAI21_X1 U7218 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6193), .ZN(n6200) );
  AOI21_X1 U7219 ( .B1(n6247), .B2(n6195), .A(n6194), .ZN(n6199) );
  OR2_X1 U7220 ( .A1(n6197), .A2(n6196), .ZN(n6198) );
  OAI211_X1 U7221 ( .C1(n6212), .C2(n6200), .A(n6199), .B(n6198), .ZN(n6201)
         );
  INV_X1 U7222 ( .A(n6201), .ZN(n6202) );
  OAI21_X1 U7223 ( .B1(n6216), .B2(n6203), .A(n6202), .ZN(U3014) );
  INV_X1 U7224 ( .A(n6204), .ZN(n6206) );
  INV_X1 U7225 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6550) );
  OAI22_X1 U7226 ( .A1(n6207), .A2(n6206), .B1(n6550), .B2(n6205), .ZN(n6208)
         );
  INV_X1 U7227 ( .A(n6208), .ZN(n6211) );
  NAND2_X1 U7228 ( .A1(n6209), .A2(n6240), .ZN(n6210) );
  OAI211_X1 U7229 ( .C1(n6212), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6211), 
        .B(n6210), .ZN(n6213) );
  INV_X1 U7230 ( .A(n6213), .ZN(n6214) );
  OAI21_X1 U7231 ( .B1(n6216), .B2(n6215), .A(n6214), .ZN(U3015) );
  OAI21_X1 U7232 ( .B1(n6218), .B2(n6243), .A(n6217), .ZN(n6220) );
  AOI22_X1 U7233 ( .A1(n6221), .A2(n6220), .B1(n6247), .B2(n6219), .ZN(n6228)
         );
  AOI22_X1 U7234 ( .A1(n6223), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6240), 
        .B2(n6222), .ZN(n6227) );
  NAND2_X1 U7235 ( .A1(n6229), .A2(REIP_REG_2__SCAN_IN), .ZN(n6226) );
  NAND3_X1 U7236 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6224), .A3(n4225), 
        .ZN(n6225) );
  NAND4_X1 U7237 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(U3016)
         );
  AOI22_X1 U7238 ( .A1(n6247), .A2(n6230), .B1(n6229), .B2(REIP_REG_1__SCAN_IN), .ZN(n6236) );
  AND2_X1 U7239 ( .A1(n6231), .A2(n6237), .ZN(n6233) );
  AOI22_X1 U7240 ( .A1(n6234), .A2(n6240), .B1(n6233), .B2(n6232), .ZN(n6235)
         );
  OAI211_X1 U7241 ( .C1(n6238), .C2(n6237), .A(n6236), .B(n6235), .ZN(U3017)
         );
  AOI21_X1 U7242 ( .B1(n6241), .B2(n6240), .A(n6239), .ZN(n6251) );
  INV_X1 U7243 ( .A(n6242), .ZN(n6248) );
  AOI21_X1 U7244 ( .B1(n6245), .B2(n6244), .A(n6243), .ZN(n6246) );
  AOI21_X1 U7245 ( .B1(n6248), .B2(n6247), .A(n6246), .ZN(n6250) );
  NAND3_X1 U7246 ( .A1(n6251), .A2(n6250), .A3(n6249), .ZN(U3018) );
  NOR2_X1 U7247 ( .A1(n6253), .A2(n6252), .ZN(U3019) );
  NOR2_X1 U7248 ( .A1(n6431), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6281)
         );
  AOI22_X1 U7249 ( .A1(n6483), .A2(n6281), .B1(n6487), .B2(n6280), .ZN(n6267)
         );
  INV_X1 U7250 ( .A(n6255), .ZN(n6435) );
  AOI21_X1 U7251 ( .B1(n6433), .B2(n6435), .A(n6256), .ZN(n6265) );
  NAND3_X1 U7252 ( .A1(n6258), .A2(n6257), .A3(n6436), .ZN(n6260) );
  INV_X1 U7253 ( .A(n6281), .ZN(n6259) );
  AND2_X1 U7254 ( .A1(n6260), .A2(n6259), .ZN(n6264) );
  INV_X1 U7255 ( .A(n6264), .ZN(n6262) );
  AOI21_X1 U7256 ( .B1(n6439), .B2(n6263), .A(n6438), .ZN(n6261) );
  OAI21_X1 U7257 ( .B1(n6265), .B2(n6262), .A(n6261), .ZN(n6283) );
  OAI22_X1 U7258 ( .A1(n6265), .A2(n6264), .B1(n6263), .B2(n6442), .ZN(n6282)
         );
  AOI22_X1 U7259 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6283), .B1(n6484), 
        .B2(n6282), .ZN(n6266) );
  OAI211_X1 U7260 ( .C1(n6448), .C2(n6317), .A(n6267), .B(n6266), .ZN(U3044)
         );
  AOI22_X1 U7261 ( .A1(n6490), .A2(n6281), .B1(n6493), .B2(n6280), .ZN(n6269)
         );
  AOI22_X1 U7262 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6283), .B1(n6491), 
        .B2(n6282), .ZN(n6268) );
  OAI211_X1 U7263 ( .C1(n6451), .C2(n6317), .A(n6269), .B(n6268), .ZN(U3045)
         );
  AOI22_X1 U7264 ( .A1(n6497), .A2(n6281), .B1(n6499), .B2(n6280), .ZN(n6271)
         );
  AOI22_X1 U7265 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6283), .B1(n6496), 
        .B2(n6282), .ZN(n6270) );
  OAI211_X1 U7266 ( .C1(n6454), .C2(n6317), .A(n6271), .B(n6270), .ZN(U3046)
         );
  AOI22_X1 U7267 ( .A1(n6945), .A2(n6281), .B1(n6946), .B2(n6280), .ZN(n6273)
         );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6283), .B1(n6455), 
        .B2(n6282), .ZN(n6272) );
  OAI211_X1 U7269 ( .C1(n6951), .C2(n6317), .A(n6273), .B(n6272), .ZN(U3047)
         );
  AOI22_X1 U7270 ( .A1(n6459), .A2(n6281), .B1(n6374), .B2(n6280), .ZN(n6275)
         );
  AOI22_X1 U7271 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6283), .B1(n6460), 
        .B2(n6282), .ZN(n6274) );
  OAI211_X1 U7272 ( .C1(n6377), .C2(n6317), .A(n6275), .B(n6274), .ZN(U3048)
         );
  AOI22_X1 U7273 ( .A1(n6502), .A2(n6281), .B1(n6505), .B2(n6280), .ZN(n6277)
         );
  AOI22_X1 U7274 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6283), .B1(n6503), 
        .B2(n6282), .ZN(n6276) );
  OAI211_X1 U7275 ( .C1(n6380), .C2(n6317), .A(n6277), .B(n6276), .ZN(U3049)
         );
  AOI22_X1 U7276 ( .A1(n6470), .A2(n6281), .B1(n6469), .B2(n6280), .ZN(n6279)
         );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6283), .B1(n6471), 
        .B2(n6282), .ZN(n6278) );
  OAI211_X1 U7278 ( .C1(n6474), .C2(n6317), .A(n6279), .B(n6278), .ZN(U3050)
         );
  AOI22_X1 U7279 ( .A1(n6509), .A2(n6281), .B1(n6514), .B2(n6280), .ZN(n6285)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6283), .B1(n6511), 
        .B2(n6282), .ZN(n6284) );
  OAI211_X1 U7281 ( .C1(n6482), .C2(n6317), .A(n6285), .B(n6284), .ZN(U3051)
         );
  INV_X1 U7282 ( .A(n6286), .ZN(n6289) );
  OAI22_X1 U7283 ( .A1(n6289), .A2(n6400), .B1(n6288), .B2(n6287), .ZN(n6312)
         );
  NOR2_X1 U7284 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6290), .ZN(n6311)
         );
  AOI22_X1 U7285 ( .A1(n6484), .A2(n6312), .B1(n6483), .B2(n6311), .ZN(n6298)
         );
  INV_X1 U7286 ( .A(n6311), .ZN(n6292) );
  AOI211_X1 U7287 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6292), .A(n6328), .B(
        n6291), .ZN(n6296) );
  OAI211_X1 U7288 ( .C1(n6317), .C2(n6326), .A(n6294), .B(n6293), .ZN(n6295)
         );
  NAND2_X1 U7289 ( .A1(n6296), .A2(n6295), .ZN(n6314) );
  AOI22_X1 U7290 ( .A1(n6314), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6486), 
        .B2(n6313), .ZN(n6297) );
  OAI211_X1 U7291 ( .C1(n6405), .C2(n6317), .A(n6298), .B(n6297), .ZN(U3052)
         );
  AOI22_X1 U7292 ( .A1(n6491), .A2(n6312), .B1(n6490), .B2(n6311), .ZN(n6300)
         );
  AOI22_X1 U7293 ( .A1(n6314), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n6492), 
        .B2(n6313), .ZN(n6299) );
  OAI211_X1 U7294 ( .C1(n6408), .C2(n6317), .A(n6300), .B(n6299), .ZN(U3053)
         );
  AOI22_X1 U7295 ( .A1(n6497), .A2(n6311), .B1(n6496), .B2(n6312), .ZN(n6302)
         );
  AOI22_X1 U7296 ( .A1(n6314), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n6498), 
        .B2(n6313), .ZN(n6301) );
  OAI211_X1 U7297 ( .C1(n6411), .C2(n6317), .A(n6302), .B(n6301), .ZN(U3054)
         );
  AOI22_X1 U7298 ( .A1(n6455), .A2(n6312), .B1(n6945), .B2(n6311), .ZN(n6304)
         );
  AOI22_X1 U7299 ( .A1(n6314), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n6412), 
        .B2(n6313), .ZN(n6303) );
  OAI211_X1 U7300 ( .C1(n6415), .C2(n6317), .A(n6304), .B(n6303), .ZN(U3055)
         );
  AOI22_X1 U7301 ( .A1(n6460), .A2(n6312), .B1(n6459), .B2(n6311), .ZN(n6306)
         );
  AOI22_X1 U7302 ( .A1(n6314), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6458), 
        .B2(n6313), .ZN(n6305) );
  OAI211_X1 U7303 ( .C1(n6463), .C2(n6317), .A(n6306), .B(n6305), .ZN(U3056)
         );
  AOI22_X1 U7304 ( .A1(n6503), .A2(n6312), .B1(n6502), .B2(n6311), .ZN(n6308)
         );
  AOI22_X1 U7305 ( .A1(n6314), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6504), 
        .B2(n6313), .ZN(n6307) );
  OAI211_X1 U7306 ( .C1(n6468), .C2(n6317), .A(n6308), .B(n6307), .ZN(U3057)
         );
  AOI22_X1 U7307 ( .A1(n6471), .A2(n6312), .B1(n6470), .B2(n6311), .ZN(n6310)
         );
  AOI22_X1 U7308 ( .A1(n6314), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n6420), 
        .B2(n6313), .ZN(n6309) );
  OAI211_X1 U7309 ( .C1(n6423), .C2(n6317), .A(n6310), .B(n6309), .ZN(U3058)
         );
  AOI22_X1 U7310 ( .A1(n6511), .A2(n6312), .B1(n6509), .B2(n6311), .ZN(n6316)
         );
  AOI22_X1 U7311 ( .A1(n6314), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n6512), 
        .B2(n6313), .ZN(n6315) );
  OAI211_X1 U7312 ( .C1(n6430), .C2(n6317), .A(n6316), .B(n6315), .ZN(U3059)
         );
  INV_X1 U7313 ( .A(n6356), .ZN(n6319) );
  NAND3_X1 U7314 ( .A1(n6319), .A2(n6354), .A3(n6318), .ZN(n6371) );
  NAND3_X1 U7315 ( .A1(n6322), .A2(n6321), .A3(n6320), .ZN(n6323) );
  OAI21_X1 U7316 ( .B1(n6400), .B2(n6324), .A(n6323), .ZN(n6348) );
  NOR2_X1 U7317 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6362), .ZN(n6347)
         );
  AOI22_X1 U7318 ( .A1(n6484), .A2(n6348), .B1(n6483), .B2(n6347), .ZN(n6334)
         );
  INV_X1 U7319 ( .A(n6371), .ZN(n6384) );
  NOR3_X1 U7320 ( .A1(n6384), .A2(n6349), .A3(n6439), .ZN(n6327) );
  OAI22_X1 U7321 ( .A1(n6327), .A2(n6326), .B1(n6325), .B2(n6324), .ZN(n6332)
         );
  INV_X1 U7322 ( .A(n6347), .ZN(n6329) );
  AOI21_X1 U7323 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6329), .A(n6328), .ZN(
        n6330) );
  NAND3_X1 U7324 ( .A1(n6332), .A2(n6331), .A3(n6330), .ZN(n6350) );
  AOI22_X1 U7325 ( .A1(n6350), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6487), 
        .B2(n6349), .ZN(n6333) );
  OAI211_X1 U7326 ( .C1(n6448), .C2(n6371), .A(n6334), .B(n6333), .ZN(U3068)
         );
  AOI22_X1 U7327 ( .A1(n6491), .A2(n6348), .B1(n6490), .B2(n6347), .ZN(n6336)
         );
  AOI22_X1 U7328 ( .A1(n6350), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6493), 
        .B2(n6349), .ZN(n6335) );
  OAI211_X1 U7329 ( .C1(n6451), .C2(n6371), .A(n6336), .B(n6335), .ZN(U3069)
         );
  AOI22_X1 U7330 ( .A1(n6497), .A2(n6347), .B1(n6496), .B2(n6348), .ZN(n6338)
         );
  AOI22_X1 U7331 ( .A1(n6350), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6499), 
        .B2(n6349), .ZN(n6337) );
  OAI211_X1 U7332 ( .C1(n6454), .C2(n6371), .A(n6338), .B(n6337), .ZN(U3070)
         );
  AOI22_X1 U7333 ( .A1(n6455), .A2(n6348), .B1(n6945), .B2(n6347), .ZN(n6340)
         );
  AOI22_X1 U7334 ( .A1(n6350), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6946), 
        .B2(n6349), .ZN(n6339) );
  OAI211_X1 U7335 ( .C1(n6951), .C2(n6371), .A(n6340), .B(n6339), .ZN(U3071)
         );
  AOI22_X1 U7336 ( .A1(n6460), .A2(n6348), .B1(n6459), .B2(n6347), .ZN(n6342)
         );
  AOI22_X1 U7337 ( .A1(n6350), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6374), 
        .B2(n6349), .ZN(n6341) );
  OAI211_X1 U7338 ( .C1(n6377), .C2(n6371), .A(n6342), .B(n6341), .ZN(U3072)
         );
  AOI22_X1 U7339 ( .A1(n6503), .A2(n6348), .B1(n6502), .B2(n6347), .ZN(n6344)
         );
  AOI22_X1 U7340 ( .A1(n6350), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6505), 
        .B2(n6349), .ZN(n6343) );
  OAI211_X1 U7341 ( .C1(n6380), .C2(n6371), .A(n6344), .B(n6343), .ZN(U3073)
         );
  AOI22_X1 U7342 ( .A1(n6471), .A2(n6348), .B1(n6470), .B2(n6347), .ZN(n6346)
         );
  AOI22_X1 U7343 ( .A1(n6350), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6469), 
        .B2(n6349), .ZN(n6345) );
  OAI211_X1 U7344 ( .C1(n6474), .C2(n6371), .A(n6346), .B(n6345), .ZN(U3074)
         );
  AOI22_X1 U7345 ( .A1(n6511), .A2(n6348), .B1(n6509), .B2(n6347), .ZN(n6352)
         );
  AOI22_X1 U7346 ( .A1(n6350), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6514), 
        .B2(n6349), .ZN(n6351) );
  OAI211_X1 U7347 ( .C1(n6482), .C2(n6371), .A(n6352), .B(n6351), .ZN(U3075)
         );
  NAND2_X1 U7348 ( .A1(n6354), .A2(n6353), .ZN(n6355) );
  INV_X1 U7349 ( .A(n6429), .ZN(n6398) );
  AOI22_X1 U7350 ( .A1(n6383), .A2(n6483), .B1(n6486), .B2(n6398), .ZN(n6366)
         );
  NAND2_X1 U7351 ( .A1(n6357), .A2(n6433), .ZN(n6364) );
  AOI21_X1 U7352 ( .B1(n6359), .B2(n6358), .A(n6383), .ZN(n6363) );
  INV_X1 U7353 ( .A(n6363), .ZN(n6361) );
  AOI21_X1 U7354 ( .B1(n6439), .B2(n6362), .A(n6438), .ZN(n6360) );
  OAI21_X1 U7355 ( .B1(n6364), .B2(n6361), .A(n6360), .ZN(n6386) );
  OAI22_X1 U7356 ( .A1(n6364), .A2(n6363), .B1(n6362), .B2(n6442), .ZN(n6385)
         );
  AOI22_X1 U7357 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6386), .B1(n6484), 
        .B2(n6385), .ZN(n6365) );
  OAI211_X1 U7358 ( .C1(n6405), .C2(n6371), .A(n6366), .B(n6365), .ZN(U3076)
         );
  AOI22_X1 U7359 ( .A1(n6490), .A2(n6383), .B1(n6492), .B2(n6398), .ZN(n6368)
         );
  AOI22_X1 U7360 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6386), .B1(n6491), 
        .B2(n6385), .ZN(n6367) );
  OAI211_X1 U7361 ( .C1(n6408), .C2(n6371), .A(n6368), .B(n6367), .ZN(U3077)
         );
  AOI22_X1 U7362 ( .A1(n6383), .A2(n6497), .B1(n6498), .B2(n6398), .ZN(n6370)
         );
  AOI22_X1 U7363 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6386), .B1(n6496), 
        .B2(n6385), .ZN(n6369) );
  OAI211_X1 U7364 ( .C1(n6411), .C2(n6371), .A(n6370), .B(n6369), .ZN(U3078)
         );
  AOI22_X1 U7365 ( .A1(n6946), .A2(n6384), .B1(n6945), .B2(n6383), .ZN(n6373)
         );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6386), .B1(n6455), 
        .B2(n6385), .ZN(n6372) );
  OAI211_X1 U7367 ( .C1(n6951), .C2(n6429), .A(n6373), .B(n6372), .ZN(U3079)
         );
  AOI22_X1 U7368 ( .A1(n6374), .A2(n6384), .B1(n6459), .B2(n6383), .ZN(n6376)
         );
  AOI22_X1 U7369 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6386), .B1(n6460), 
        .B2(n6385), .ZN(n6375) );
  OAI211_X1 U7370 ( .C1(n6377), .C2(n6429), .A(n6376), .B(n6375), .ZN(U3080)
         );
  AOI22_X1 U7371 ( .A1(n6505), .A2(n6384), .B1(n6502), .B2(n6383), .ZN(n6379)
         );
  AOI22_X1 U7372 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6386), .B1(n6503), 
        .B2(n6385), .ZN(n6378) );
  OAI211_X1 U7373 ( .C1(n6380), .C2(n6429), .A(n6379), .B(n6378), .ZN(U3081)
         );
  AOI22_X1 U7374 ( .A1(n6469), .A2(n6384), .B1(n6470), .B2(n6383), .ZN(n6382)
         );
  AOI22_X1 U7375 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6386), .B1(n6471), 
        .B2(n6385), .ZN(n6381) );
  OAI211_X1 U7376 ( .C1(n6474), .C2(n6429), .A(n6382), .B(n6381), .ZN(U3082)
         );
  AOI22_X1 U7377 ( .A1(n6514), .A2(n6384), .B1(n6509), .B2(n6383), .ZN(n6388)
         );
  AOI22_X1 U7378 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6386), .B1(n6511), 
        .B2(n6385), .ZN(n6387) );
  OAI211_X1 U7379 ( .C1(n6482), .C2(n6429), .A(n6388), .B(n6387), .ZN(U3083)
         );
  OAI22_X1 U7380 ( .A1(n6392), .A2(n6391), .B1(n6390), .B2(n6389), .ZN(n6425)
         );
  NOR2_X1 U7381 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6393), .ZN(n6424)
         );
  AOI22_X1 U7382 ( .A1(n6484), .A2(n6425), .B1(n6483), .B2(n6424), .ZN(n6404)
         );
  INV_X1 U7383 ( .A(n6394), .ZN(n6395) );
  OAI211_X1 U7384 ( .C1(n6424), .C2(n6397), .A(n6396), .B(n6395), .ZN(n6402)
         );
  AOI211_X1 U7385 ( .C1(n6400), .C2(n6399), .A(n6398), .B(n6426), .ZN(n6401)
         );
  AOI22_X1 U7386 ( .A1(n3128), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6486), 
        .B2(n6426), .ZN(n6403) );
  OAI211_X1 U7387 ( .C1(n6405), .C2(n6429), .A(n6404), .B(n6403), .ZN(U3084)
         );
  AOI22_X1 U7388 ( .A1(n6491), .A2(n6425), .B1(n6490), .B2(n6424), .ZN(n6407)
         );
  AOI22_X1 U7389 ( .A1(n3128), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6426), 
        .B2(n6492), .ZN(n6406) );
  OAI211_X1 U7390 ( .C1(n6408), .C2(n6429), .A(n6407), .B(n6406), .ZN(U3085)
         );
  AOI22_X1 U7391 ( .A1(n6497), .A2(n6424), .B1(n6496), .B2(n6425), .ZN(n6410)
         );
  AOI22_X1 U7392 ( .A1(n3128), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6426), 
        .B2(n6498), .ZN(n6409) );
  OAI211_X1 U7393 ( .C1(n6411), .C2(n6429), .A(n6410), .B(n6409), .ZN(U3086)
         );
  AOI22_X1 U7394 ( .A1(n6455), .A2(n6425), .B1(n6945), .B2(n6424), .ZN(n6414)
         );
  AOI22_X1 U7395 ( .A1(n3128), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6426), 
        .B2(n6412), .ZN(n6413) );
  OAI211_X1 U7396 ( .C1(n6415), .C2(n6429), .A(n6414), .B(n6413), .ZN(U3087)
         );
  AOI22_X1 U7397 ( .A1(n6460), .A2(n6425), .B1(n6459), .B2(n6424), .ZN(n6417)
         );
  AOI22_X1 U7398 ( .A1(n3128), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6426), 
        .B2(n6458), .ZN(n6416) );
  OAI211_X1 U7399 ( .C1(n6463), .C2(n6429), .A(n6417), .B(n6416), .ZN(U3088)
         );
  AOI22_X1 U7400 ( .A1(n6503), .A2(n6425), .B1(n6502), .B2(n6424), .ZN(n6419)
         );
  AOI22_X1 U7401 ( .A1(n3128), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6426), 
        .B2(n6504), .ZN(n6418) );
  OAI211_X1 U7402 ( .C1(n6468), .C2(n6429), .A(n6419), .B(n6418), .ZN(U3089)
         );
  AOI22_X1 U7403 ( .A1(n6471), .A2(n6425), .B1(n6470), .B2(n6424), .ZN(n6422)
         );
  AOI22_X1 U7404 ( .A1(n3128), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6426), 
        .B2(n6420), .ZN(n6421) );
  OAI211_X1 U7405 ( .C1(n6423), .C2(n6429), .A(n6422), .B(n6421), .ZN(U3090)
         );
  AOI22_X1 U7406 ( .A1(n6511), .A2(n6425), .B1(n6509), .B2(n6424), .ZN(n6428)
         );
  AOI22_X1 U7407 ( .A1(n3128), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6426), 
        .B2(n6512), .ZN(n6427) );
  OAI211_X1 U7408 ( .C1(n6430), .C2(n6429), .A(n6428), .B(n6427), .ZN(U3091)
         );
  INV_X1 U7409 ( .A(n6431), .ZN(n6432) );
  AND2_X1 U7410 ( .A1(n6432), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6476)
         );
  AOI22_X1 U7411 ( .A1(n6487), .A2(n6475), .B1(n6483), .B2(n6476), .ZN(n6447)
         );
  OAI21_X1 U7412 ( .B1(n6435), .B2(n6434), .A(n6433), .ZN(n6445) );
  AOI21_X1 U7413 ( .B1(n6437), .B2(n6436), .A(n6476), .ZN(n6444) );
  INV_X1 U7414 ( .A(n6444), .ZN(n6441) );
  AOI21_X1 U7415 ( .B1(n6439), .B2(n6443), .A(n6438), .ZN(n6440) );
  OAI21_X1 U7416 ( .B1(n6445), .B2(n6441), .A(n6440), .ZN(n6478) );
  OAI22_X1 U7417 ( .A1(n6445), .A2(n6444), .B1(n6443), .B2(n6442), .ZN(n6477)
         );
  AOI22_X1 U7418 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6478), .B1(n6484), 
        .B2(n6477), .ZN(n6446) );
  OAI211_X1 U7419 ( .C1(n6448), .C2(n6481), .A(n6447), .B(n6446), .ZN(U3108)
         );
  AOI22_X1 U7420 ( .A1(n6490), .A2(n6476), .B1(n6475), .B2(n6493), .ZN(n6450)
         );
  AOI22_X1 U7421 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6478), .B1(n6491), 
        .B2(n6477), .ZN(n6449) );
  OAI211_X1 U7422 ( .C1(n6451), .C2(n6481), .A(n6450), .B(n6449), .ZN(U3109)
         );
  AOI22_X1 U7423 ( .A1(n6499), .A2(n6475), .B1(n6497), .B2(n6476), .ZN(n6453)
         );
  AOI22_X1 U7424 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6478), .B1(n6496), 
        .B2(n6477), .ZN(n6452) );
  OAI211_X1 U7425 ( .C1(n6454), .C2(n6481), .A(n6453), .B(n6452), .ZN(U3110)
         );
  AOI22_X1 U7426 ( .A1(n6945), .A2(n6476), .B1(n6475), .B2(n6946), .ZN(n6457)
         );
  AOI22_X1 U7427 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6478), .B1(n6455), 
        .B2(n6477), .ZN(n6456) );
  OAI211_X1 U7428 ( .C1(n6951), .C2(n6481), .A(n6457), .B(n6456), .ZN(U3111)
         );
  INV_X1 U7429 ( .A(n6481), .ZN(n6464) );
  AOI22_X1 U7430 ( .A1(n6459), .A2(n6476), .B1(n6464), .B2(n6458), .ZN(n6462)
         );
  AOI22_X1 U7431 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6478), .B1(n6460), 
        .B2(n6477), .ZN(n6461) );
  OAI211_X1 U7432 ( .C1(n6463), .C2(n6467), .A(n6462), .B(n6461), .ZN(U3112)
         );
  AOI22_X1 U7433 ( .A1(n6502), .A2(n6476), .B1(n6464), .B2(n6504), .ZN(n6466)
         );
  AOI22_X1 U7434 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6478), .B1(n6503), 
        .B2(n6477), .ZN(n6465) );
  OAI211_X1 U7435 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n6465), .ZN(U3113)
         );
  AOI22_X1 U7436 ( .A1(n6470), .A2(n6476), .B1(n6475), .B2(n6469), .ZN(n6473)
         );
  AOI22_X1 U7437 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6478), .B1(n6471), 
        .B2(n6477), .ZN(n6472) );
  OAI211_X1 U7438 ( .C1(n6474), .C2(n6481), .A(n6473), .B(n6472), .ZN(U3114)
         );
  AOI22_X1 U7439 ( .A1(n6509), .A2(n6476), .B1(n6475), .B2(n6514), .ZN(n6480)
         );
  AOI22_X1 U7440 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6478), .B1(n6511), 
        .B2(n6477), .ZN(n6479) );
  OAI211_X1 U7441 ( .C1(n6482), .C2(n6481), .A(n6480), .B(n6479), .ZN(U3115)
         );
  INV_X1 U7442 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6827) );
  AOI22_X1 U7443 ( .A1(n6484), .A2(n6510), .B1(n6483), .B2(n6508), .ZN(n6489)
         );
  INV_X1 U7444 ( .A(n6485), .ZN(n6515) );
  AOI22_X1 U7445 ( .A1(n6515), .A2(n6487), .B1(n6513), .B2(n6486), .ZN(n6488)
         );
  OAI211_X1 U7446 ( .C1(n6518), .C2(n6827), .A(n6489), .B(n6488), .ZN(U3124)
         );
  INV_X1 U7447 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6859) );
  AOI22_X1 U7448 ( .A1(n6491), .A2(n6510), .B1(n6490), .B2(n6508), .ZN(n6495)
         );
  AOI22_X1 U7449 ( .A1(n6515), .A2(n6493), .B1(n6513), .B2(n6492), .ZN(n6494)
         );
  OAI211_X1 U7450 ( .C1(n6518), .C2(n6859), .A(n6495), .B(n6494), .ZN(U3125)
         );
  INV_X1 U7451 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6729) );
  AOI22_X1 U7452 ( .A1(n6497), .A2(n6508), .B1(n6496), .B2(n6510), .ZN(n6501)
         );
  AOI22_X1 U7453 ( .A1(n6515), .A2(n6499), .B1(n6513), .B2(n6498), .ZN(n6500)
         );
  OAI211_X1 U7454 ( .C1(n6518), .C2(n6729), .A(n6501), .B(n6500), .ZN(U3126)
         );
  INV_X1 U7455 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U7456 ( .A1(n6503), .A2(n6510), .B1(n6502), .B2(n6508), .ZN(n6507)
         );
  AOI22_X1 U7457 ( .A1(n6515), .A2(n6505), .B1(n6513), .B2(n6504), .ZN(n6506)
         );
  OAI211_X1 U7458 ( .C1(n6518), .C2(n6716), .A(n6507), .B(n6506), .ZN(U3129)
         );
  INV_X1 U7459 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6861) );
  AOI22_X1 U7460 ( .A1(n6511), .A2(n6510), .B1(n6509), .B2(n6508), .ZN(n6517)
         );
  AOI22_X1 U7461 ( .A1(n6515), .A2(n6514), .B1(n6513), .B2(n6512), .ZN(n6516)
         );
  OAI211_X1 U7462 ( .C1(n6518), .C2(n6861), .A(n6517), .B(n6516), .ZN(U3131)
         );
  NOR2_X1 U7463 ( .A1(n6765), .A2(READY_N), .ZN(n6528) );
  INV_X1 U7464 ( .A(n6528), .ZN(n6519) );
  AOI221_X1 U7465 ( .B1(n6521), .B2(n6520), .C1(n6519), .C2(n6520), .A(n6602), 
        .ZN(n6523) );
  AOI211_X1 U7466 ( .C1(STATE2_REG_1__SCAN_IN), .C2(n6524), .A(n6523), .B(
        n6522), .ZN(n6525) );
  OAI21_X1 U7467 ( .B1(n6527), .B2(n6526), .A(n6525), .ZN(U3149) );
  AOI21_X1 U7468 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6528), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6530) );
  OAI21_X1 U7469 ( .B1(n6600), .B2(n6530), .A(n6529), .ZN(U3150) );
  INV_X1 U7470 ( .A(n6599), .ZN(n6595) );
  AND2_X1 U7471 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6595), .ZN(U3151) );
  AND2_X1 U7472 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6595), .ZN(U3152) );
  AND2_X1 U7473 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6595), .ZN(U3153) );
  AND2_X1 U7474 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6595), .ZN(U3154) );
  AND2_X1 U7475 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6595), .ZN(U3155) );
  INV_X1 U7476 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6778) );
  NOR2_X1 U7477 ( .A1(n6599), .A2(n6778), .ZN(U3156) );
  AND2_X1 U7478 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6595), .ZN(U3157) );
  AND2_X1 U7479 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6595), .ZN(U3158) );
  INV_X1 U7480 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6761) );
  NOR2_X1 U7481 ( .A1(n6599), .A2(n6761), .ZN(U3159) );
  INV_X1 U7482 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6763) );
  NOR2_X1 U7483 ( .A1(n6599), .A2(n6763), .ZN(U3160) );
  AND2_X1 U7484 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6595), .ZN(U3161) );
  AND2_X1 U7485 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6595), .ZN(U3162) );
  AND2_X1 U7486 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6595), .ZN(U3163) );
  AND2_X1 U7487 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6595), .ZN(U3164) );
  AND2_X1 U7488 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6595), .ZN(U3165) );
  AND2_X1 U7489 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6595), .ZN(U3166) );
  AND2_X1 U7490 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6595), .ZN(U3167) );
  AND2_X1 U7491 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6595), .ZN(U3168) );
  AND2_X1 U7492 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6595), .ZN(U3169) );
  INV_X1 U7493 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6723) );
  NOR2_X1 U7494 ( .A1(n6599), .A2(n6723), .ZN(U3170) );
  AND2_X1 U7495 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6595), .ZN(U3171) );
  AND2_X1 U7496 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6595), .ZN(U3172) );
  INV_X1 U7497 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6811) );
  NOR2_X1 U7498 ( .A1(n6599), .A2(n6811), .ZN(U3173) );
  AND2_X1 U7499 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6595), .ZN(U3174) );
  AND2_X1 U7500 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6595), .ZN(U3175) );
  AND2_X1 U7501 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6595), .ZN(U3176) );
  INV_X1 U7502 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6777) );
  NOR2_X1 U7503 ( .A1(n6599), .A2(n6777), .ZN(U3177) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6595), .ZN(U3178) );
  INV_X1 U7505 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6775) );
  NOR2_X1 U7506 ( .A1(n6599), .A2(n6775), .ZN(U3179) );
  AND2_X1 U7507 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6595), .ZN(U3180) );
  NAND2_X1 U7508 ( .A1(STATE_REG_1__SCAN_IN), .A2(READY_N), .ZN(n6542) );
  NOR2_X1 U7509 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6531) );
  INV_X1 U7510 ( .A(HOLD), .ZN(n6810) );
  OAI21_X1 U7511 ( .B1(n6531), .B2(n6810), .A(REQUESTPENDING_REG_SCAN_IN), 
        .ZN(n6532) );
  INV_X1 U7512 ( .A(NA_N), .ZN(n6540) );
  AOI221_X1 U7513 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6540), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6545) );
  AOI21_X1 U7514 ( .B1(n6589), .B2(n6532), .A(n6545), .ZN(n6533) );
  OAI21_X1 U7515 ( .B1(STATE_REG_2__SCAN_IN), .B2(n6542), .A(n6533), .ZN(U3181) );
  AND2_X1 U7516 ( .A1(HOLD), .A2(STATE_REG_1__SCAN_IN), .ZN(n6535) );
  INV_X1 U7517 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6865) );
  NOR2_X1 U7518 ( .A1(n6538), .A2(n6865), .ZN(n6541) );
  OAI22_X1 U7519 ( .A1(n6535), .A2(n6541), .B1(n6810), .B2(n6534), .ZN(n6537)
         );
  NAND3_X1 U7520 ( .A1(n6537), .A2(n6536), .A3(n6542), .ZN(U3182) );
  AOI221_X1 U7521 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6617), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6539) );
  AOI221_X1 U7522 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6539), .C2(HOLD), .A(n6538), .ZN(n6544) );
  AOI21_X1 U7523 ( .B1(n6541), .B2(n6540), .A(STATE_REG_2__SCAN_IN), .ZN(n6543) );
  OAI22_X1 U7524 ( .A1(n6545), .A2(n6544), .B1(n6543), .B2(n6542), .ZN(U3183)
         );
  NAND2_X1 U7525 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6629), .ZN(n6585) );
  NOR2_X2 U7526 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6589), .ZN(n6590) );
  AOI22_X1 U7527 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6589), .ZN(n6546) );
  OAI21_X1 U7528 ( .B1(n6745), .B2(n6585), .A(n6546), .ZN(U3184) );
  AOI22_X1 U7529 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6589), .ZN(n6547) );
  OAI21_X1 U7530 ( .B1(n6548), .B2(n6592), .A(n6547), .ZN(U3185) );
  AOI22_X1 U7531 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6589), .ZN(n6549) );
  OAI21_X1 U7532 ( .B1(n6550), .B2(n6592), .A(n6549), .ZN(U3186) );
  AOI22_X1 U7533 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6589), .ZN(n6551) );
  OAI21_X1 U7534 ( .B1(n6552), .B2(n6592), .A(n6551), .ZN(U3187) );
  INV_X1 U7535 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6862) );
  INV_X1 U7536 ( .A(n6590), .ZN(n6588) );
  OAI222_X1 U7537 ( .A1(n6585), .A2(n6553), .B1(n6862), .B2(n6629), .C1(n6728), 
        .C2(n6588), .ZN(U3188) );
  AOI22_X1 U7538 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6589), .ZN(n6554) );
  OAI21_X1 U7539 ( .B1(n6728), .B2(n6592), .A(n6554), .ZN(U3189) );
  INV_X1 U7540 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6680) );
  OAI222_X1 U7541 ( .A1(n6585), .A2(n6555), .B1(n6680), .B2(n6629), .C1(n6556), 
        .C2(n6588), .ZN(U3190) );
  INV_X1 U7542 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U7543 ( .A1(n6588), .A2(n6843), .B1(n6678), .B2(n6629), .C1(n6556), 
        .C2(n6592), .ZN(U3191) );
  AOI22_X1 U7544 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6589), .ZN(n6557) );
  OAI21_X1 U7545 ( .B1(n6843), .B2(n6592), .A(n6557), .ZN(U3192) );
  AOI22_X1 U7546 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6589), .ZN(n6558) );
  OAI21_X1 U7547 ( .B1(n6559), .B2(n6592), .A(n6558), .ZN(U3193) );
  INV_X1 U7548 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6840) );
  OAI222_X1 U7549 ( .A1(n6585), .A2(n6560), .B1(n6840), .B2(n6629), .C1(n4878), 
        .C2(n6588), .ZN(U3194) );
  AOI22_X1 U7550 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6589), .ZN(n6561) );
  OAI21_X1 U7551 ( .B1(n4878), .B2(n6592), .A(n6561), .ZN(U3195) );
  INV_X1 U7552 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6923) );
  OAI222_X1 U7553 ( .A1(n6592), .A2(n6562), .B1(n6923), .B2(n6629), .C1(n6564), 
        .C2(n6588), .ZN(U3196) );
  AOI22_X1 U7554 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6589), .ZN(n6563) );
  OAI21_X1 U7555 ( .B1(n6564), .B2(n6592), .A(n6563), .ZN(U3197) );
  AOI22_X1 U7556 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6589), .ZN(n6565) );
  OAI21_X1 U7557 ( .B1(n6566), .B2(n6592), .A(n6565), .ZN(U3198) );
  INV_X1 U7558 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6829) );
  OAI222_X1 U7559 ( .A1(n6592), .A2(n6731), .B1(n6829), .B2(n6629), .C1(n6567), 
        .C2(n6588), .ZN(U3199) );
  INV_X1 U7560 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6807) );
  OAI222_X1 U7561 ( .A1(n6588), .A2(n6569), .B1(n6807), .B2(n6629), .C1(n6567), 
        .C2(n6592), .ZN(U3200) );
  AOI22_X1 U7562 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6589), .ZN(n6568) );
  OAI21_X1 U7563 ( .B1(n6569), .B2(n6592), .A(n6568), .ZN(U3201) );
  AOI22_X1 U7564 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6589), .ZN(n6570) );
  OAI21_X1 U7565 ( .B1(n6571), .B2(n6592), .A(n6570), .ZN(U3202) );
  INV_X1 U7566 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6842) );
  OAI222_X1 U7567 ( .A1(n6585), .A2(n6572), .B1(n6842), .B2(n6629), .C1(n5580), 
        .C2(n6588), .ZN(U3203) );
  AOI22_X1 U7568 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6589), .ZN(n6573) );
  OAI21_X1 U7569 ( .B1(n5580), .B2(n6592), .A(n6573), .ZN(U3204) );
  INV_X1 U7570 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6574) );
  INV_X1 U7571 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6920) );
  INV_X1 U7572 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6576) );
  OAI222_X1 U7573 ( .A1(n6585), .A2(n6574), .B1(n6920), .B2(n6629), .C1(n6576), 
        .C2(n6588), .ZN(U3205) );
  AOI22_X1 U7574 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6589), .ZN(n6575) );
  OAI21_X1 U7575 ( .B1(n6576), .B2(n6592), .A(n6575), .ZN(U3206) );
  AOI22_X1 U7576 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6589), .ZN(n6577) );
  OAI21_X1 U7577 ( .B1(n6578), .B2(n6592), .A(n6577), .ZN(U3207) );
  AOI22_X1 U7578 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6589), .ZN(n6579) );
  OAI21_X1 U7579 ( .B1(n6580), .B2(n6592), .A(n6579), .ZN(U3208) );
  AOI22_X1 U7580 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6589), .ZN(n6581) );
  OAI21_X1 U7581 ( .B1(n6582), .B2(n6585), .A(n6581), .ZN(U3209) );
  INV_X1 U7582 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6848) );
  INV_X1 U7583 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6586) );
  OAI222_X1 U7584 ( .A1(n6585), .A2(n6583), .B1(n6848), .B2(n6629), .C1(n6586), 
        .C2(n6588), .ZN(U3210) );
  AOI22_X1 U7585 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6589), .ZN(n6584) );
  OAI21_X1 U7586 ( .B1(n6586), .B2(n6585), .A(n6584), .ZN(U3211) );
  INV_X1 U7587 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U7588 ( .A1(n6588), .A2(n6593), .B1(n6766), .B2(n6629), .C1(n6587), 
        .C2(n6592), .ZN(U3212) );
  AOI22_X1 U7589 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6590), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6589), .ZN(n6591) );
  OAI21_X1 U7590 ( .B1(n6593), .B2(n6592), .A(n6591), .ZN(U3213) );
  MUX2_X1 U7591 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6629), .Z(U3445) );
  MUX2_X1 U7592 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6629), .Z(U3446) );
  MUX2_X1 U7593 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6629), .Z(U3447) );
  MUX2_X1 U7594 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6629), .Z(U3448) );
  INV_X1 U7595 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6596) );
  INV_X1 U7596 ( .A(n6597), .ZN(n6594) );
  AOI21_X1 U7597 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(U3451) );
  OAI21_X1 U7598 ( .B1(n6599), .B2(n6598), .A(n6597), .ZN(U3452) );
  AOI211_X1 U7599 ( .C1(n6602), .C2(STATE2_REG_3__SCAN_IN), .A(n6601), .B(
        n6600), .ZN(n6603) );
  INV_X1 U7600 ( .A(n6603), .ZN(U3453) );
  AOI22_X1 U7601 ( .A1(n6607), .A2(n6606), .B1(n6605), .B2(n6604), .ZN(n6608)
         );
  INV_X1 U7602 ( .A(n6608), .ZN(n6610) );
  MUX2_X1 U7603 ( .A(n6610), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6609), 
        .Z(U3456) );
  AOI21_X1 U7604 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6611) );
  AOI22_X1 U7605 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6611), .B2(n6745), .ZN(n6613) );
  INV_X1 U7606 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6906) );
  AOI22_X1 U7607 ( .A1(n6615), .A2(n6613), .B1(n6906), .B2(n6612), .ZN(U3468)
         );
  INV_X1 U7608 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6912) );
  OAI21_X1 U7609 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6615), .ZN(n6614) );
  OAI21_X1 U7610 ( .B1(n6615), .B2(n6912), .A(n6614), .ZN(U3469) );
  INV_X1 U7611 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6760) );
  MUX2_X1 U7612 ( .A(W_R_N_REG_SCAN_IN), .B(n6760), .S(n6629), .Z(U3470) );
  INV_X1 U7613 ( .A(n6616), .ZN(n6620) );
  OAI211_X1 U7614 ( .C1(n6618), .C2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .B(n6617), .ZN(n6619) );
  OAI21_X1 U7615 ( .B1(n6620), .B2(n6619), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6622) );
  NAND2_X1 U7616 ( .A1(n6622), .A2(n6621), .ZN(n6628) );
  INV_X1 U7617 ( .A(n6623), .ZN(n6624) );
  OAI211_X1 U7618 ( .C1(READY_N), .C2(n6626), .A(n6625), .B(n6624), .ZN(n6627)
         );
  MUX2_X1 U7619 ( .A(REQUESTPENDING_REG_SCAN_IN), .B(n6628), .S(n6627), .Z(
        U3472) );
  MUX2_X1 U7620 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6629), .Z(U3473) );
  INV_X1 U7621 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6675) );
  NAND4_X1 U7622 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4588), .A3(n6830), 
        .A4(n6675), .ZN(n6633) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n6697) );
  NAND4_X1 U7624 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(
        INSTQUEUE_REG_2__7__SCAN_IN), .A3(n6697), .A4(n6879), .ZN(n6632) );
  NAND4_X1 U7625 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(
        INSTQUEUE_REG_11__2__SCAN_IN), .A3(INSTQUEUE_REG_10__2__SCAN_IN), .A4(
        n4376), .ZN(n6631) );
  INV_X1 U7626 ( .A(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n6899) );
  NAND4_X1 U7627 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        INSTQUEUE_REG_3__0__SCAN_IN), .A3(INSTQUEUE_REG_10__0__SCAN_IN), .A4(
        n6899), .ZN(n6630) );
  NOR4_X1 U7628 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6640)
         );
  AND4_X1 U7629 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        STATE2_REG_0__SCAN_IN), .A3(INSTQUEUE_REG_7__7__SCAN_IN), .A4(
        INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6636) );
  INV_X1 U7630 ( .A(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n6864) );
  NOR4_X1 U7631 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(
        INSTQUEUE_REG_10__6__SCAN_IN), .A3(n6864), .A4(n6911), .ZN(n6635) );
  INV_X1 U7632 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6883) );
  NOR4_X1 U7633 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        INSTQUEUE_REG_1__0__SCAN_IN), .A3(n6747), .A4(n6883), .ZN(n6634) );
  NAND3_X1 U7634 ( .A1(n6636), .A2(n6635), .A3(n6634), .ZN(n6637) );
  NOR4_X1 U7635 ( .A1(n6638), .A2(DATAWIDTH_REG_5__SCAN_IN), .A3(
        DATAWIDTH_REG_9__SCAN_IN), .A4(n6637), .ZN(n6639) );
  NAND2_X1 U7636 ( .A1(n6640), .A2(n6639), .ZN(n6672) );
  NOR4_X1 U7637 ( .A1(DATAO_REG_30__SCAN_IN), .A2(UWORD_REG_4__SCAN_IN), .A3(
        DATAO_REG_18__SCAN_IN), .A4(ADDRESS_REG_28__SCAN_IN), .ZN(n6644) );
  NOR4_X1 U7638 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(DATAI_27_), .A3(
        ADS_N_REG_SCAN_IN), .A4(n6894), .ZN(n6643) );
  NOR4_X1 U7639 ( .A1(ADDRESS_REG_7__SCAN_IN), .A2(ADDRESS_REG_6__SCAN_IN), 
        .A3(ADDRESS_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6642)
         );
  NOR4_X1 U7640 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(ADDRESS_REG_16__SCAN_IN), 
        .A3(ADDRESS_REG_15__SCAN_IN), .A4(ADDRESS_REG_12__SCAN_IN), .ZN(n6641)
         );
  NAND4_X1 U7641 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6671)
         );
  NOR4_X1 U7642 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(
        INSTQUEUE_REG_10__3__SCAN_IN), .A3(n6716), .A4(n4324), .ZN(n6648) );
  NOR4_X1 U7643 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(
        INSTQUEUE_REG_12__2__SCAN_IN), .A3(INSTQUEUE_REG_9__3__SCAN_IN), .A4(
        INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6647) );
  INV_X1 U7644 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6881) );
  NOR4_X1 U7645 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6881), .A3(n6859), 
        .A4(n6708), .ZN(n6646) );
  NOR4_X1 U7646 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        INSTQUEUE_REG_3__5__SCAN_IN), .A3(INSTQUEUE_REG_5__1__SCAN_IN), .A4(
        INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6645) );
  NAND4_X1 U7647 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6670)
         );
  NAND4_X1 U7648 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6788), .A3(n5580), .A4(
        n6808), .ZN(n6652) );
  NAND4_X1 U7649 ( .A1(n6742), .A2(n6745), .A3(n6731), .A4(n6845), .ZN(n6651)
         );
  NAND4_X1 U7650 ( .A1(DATAO_REG_22__SCAN_IN), .A2(UWORD_REG_11__SCAN_IN), 
        .A3(READREQUEST_REG_SCAN_IN), .A4(DATAO_REG_25__SCAN_IN), .ZN(n6650)
         );
  NAND4_X1 U7651 ( .A1(DATAO_REG_9__SCAN_IN), .A2(ADDRESS_REG_19__SCAN_IN), 
        .A3(ADDRESS_REG_10__SCAN_IN), .A4(n4225), .ZN(n6649) );
  NOR4_X1 U7652 ( .A1(n6652), .A2(n6651), .A3(n6650), .A4(n6649), .ZN(n6668)
         );
  NOR4_X1 U7653 ( .A1(BYTEENABLE_REG_0__SCAN_IN), .A2(ADDRESS_REG_21__SCAN_IN), 
        .A3(REQUESTPENDING_REG_SCAN_IN), .A4(HOLD), .ZN(n6656) );
  NOR4_X1 U7654 ( .A1(MORE_REG_SCAN_IN), .A2(DATAO_REG_10__SCAN_IN), .A3(
        MEMORYFETCH_REG_SCAN_IN), .A4(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6655)
         );
  NOR4_X1 U7655 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(EBX_REG_25__SCAN_IN), .A3(LWORD_REG_4__SCAN_IN), .A4(UWORD_REG_1__SCAN_IN), .ZN(n6654) );
  NOR4_X1 U7656 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(EAX_REG_3__SCAN_IN), 
        .A3(EAX_REG_6__SCAN_IN), .A4(EBX_REG_9__SCAN_IN), .ZN(n6653) );
  AND4_X1 U7657 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6667)
         );
  NAND4_X1 U7658 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(PHYADDRPOINTER_REG_22__SCAN_IN), 
        .A4(DATAI_21_), .ZN(n6660) );
  NAND4_X1 U7659 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(EBX_REG_18__SCAN_IN), .A4(
        EBX_REG_15__SCAN_IN), .ZN(n6659) );
  NAND4_X1 U7660 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A3(EBX_REG_19__SCAN_IN), .A4(
        DATAI_13_), .ZN(n6658) );
  NAND4_X1 U7661 ( .A1(EAX_REG_22__SCAN_IN), .A2(EAX_REG_30__SCAN_IN), .A3(
        DATAI_5_), .A4(DATAI_20_), .ZN(n6657) );
  NOR4_X1 U7662 ( .A1(n6660), .A2(n6659), .A3(n6658), .A4(n6657), .ZN(n6666)
         );
  NAND4_X1 U7663 ( .A1(EBX_REG_11__SCAN_IN), .A2(BYTEENABLE_REG_2__SCAN_IN), 
        .A3(BS16_N), .A4(UWORD_REG_0__SCAN_IN), .ZN(n6664) );
  NAND4_X1 U7664 ( .A1(FLUSH_REG_SCAN_IN), .A2(DATAWIDTH_REG_22__SCAN_IN), 
        .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_26__SCAN_IN), .ZN(
        n6663) );
  NAND4_X1 U7665 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(EBX_REG_7__SCAN_IN), 
        .A3(REIP_REG_6__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n6662) );
  NAND4_X1 U7666 ( .A1(EAX_REG_15__SCAN_IN), .A2(EBX_REG_22__SCAN_IN), .A3(
        EBX_REG_1__SCAN_IN), .A4(UWORD_REG_10__SCAN_IN), .ZN(n6661) );
  NOR4_X1 U7667 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6665)
         );
  NAND4_X1 U7668 ( .A1(n6668), .A2(n6667), .A3(n6666), .A4(n6665), .ZN(n6669)
         );
  NOR4_X1 U7669 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6943)
         );
  INV_X1 U7670 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6674) );
  AOI22_X1 U7671 ( .A1(n6675), .A2(keyinput2), .B1(keyinput38), .B2(n6674), 
        .ZN(n6673) );
  OAI221_X1 U7672 ( .B1(n6675), .B2(keyinput2), .C1(n6674), .C2(keyinput38), 
        .A(n6673), .ZN(n6688) );
  AOI22_X1 U7673 ( .A1(n6678), .A2(keyinput76), .B1(n6677), .B2(keyinput56), 
        .ZN(n6676) );
  OAI221_X1 U7674 ( .B1(n6678), .B2(keyinput76), .C1(n6677), .C2(keyinput56), 
        .A(n6676), .ZN(n6687) );
  AOI22_X1 U7675 ( .A1(n6681), .A2(keyinput55), .B1(keyinput40), .B2(n6680), 
        .ZN(n6679) );
  OAI221_X1 U7676 ( .B1(n6681), .B2(keyinput55), .C1(n6680), .C2(keyinput40), 
        .A(n6679), .ZN(n6686) );
  AOI22_X1 U7677 ( .A1(n6684), .A2(keyinput3), .B1(keyinput94), .B2(n6683), 
        .ZN(n6682) );
  OAI221_X1 U7678 ( .B1(n6684), .B2(keyinput3), .C1(n6683), .C2(keyinput94), 
        .A(n6682), .ZN(n6685) );
  NOR4_X1 U7679 ( .A1(n6688), .A2(n6687), .A3(n6686), .A4(n6685), .ZN(n6740)
         );
  AOI22_X1 U7680 ( .A1(n6691), .A2(keyinput113), .B1(keyinput9), .B2(n6690), 
        .ZN(n6689) );
  OAI221_X1 U7681 ( .B1(n6691), .B2(keyinput113), .C1(n6690), .C2(keyinput9), 
        .A(n6689), .ZN(n6705) );
  INV_X1 U7682 ( .A(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U7683 ( .A1(n6694), .A2(keyinput83), .B1(keyinput25), .B2(n6693), 
        .ZN(n6692) );
  OAI221_X1 U7684 ( .B1(n6694), .B2(keyinput83), .C1(n6693), .C2(keyinput25), 
        .A(n6692), .ZN(n6704) );
  INV_X1 U7685 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6696) );
  AOI22_X1 U7686 ( .A1(n6697), .A2(keyinput61), .B1(keyinput127), .B2(n6696), 
        .ZN(n6695) );
  OAI221_X1 U7687 ( .B1(n6697), .B2(keyinput61), .C1(n6696), .C2(keyinput127), 
        .A(n6695), .ZN(n6703) );
  INV_X1 U7688 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6698) );
  XOR2_X1 U7689 ( .A(n6698), .B(keyinput26), .Z(n6701) );
  XNOR2_X1 U7690 ( .A(n6699), .B(keyinput89), .ZN(n6700) );
  NAND2_X1 U7691 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  NOR4_X1 U7692 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6739)
         );
  AOI22_X1 U7693 ( .A1(n6708), .A2(keyinput30), .B1(keyinput14), .B2(n6707), 
        .ZN(n6706) );
  OAI221_X1 U7694 ( .B1(n6708), .B2(keyinput30), .C1(n6707), .C2(keyinput14), 
        .A(n6706), .ZN(n6721) );
  INV_X1 U7695 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U7696 ( .A1(n6711), .A2(keyinput123), .B1(keyinput115), .B2(n6710), 
        .ZN(n6709) );
  OAI221_X1 U7697 ( .B1(n6711), .B2(keyinput123), .C1(n6710), .C2(keyinput115), 
        .A(n6709), .ZN(n6720) );
  INV_X1 U7698 ( .A(DATAI_20_), .ZN(n6714) );
  AOI22_X1 U7699 ( .A1(n6714), .A2(keyinput112), .B1(keyinput66), .B2(n6713), 
        .ZN(n6712) );
  OAI221_X1 U7700 ( .B1(n6714), .B2(keyinput112), .C1(n6713), .C2(keyinput66), 
        .A(n6712), .ZN(n6719) );
  AOI22_X1 U7701 ( .A1(n6717), .A2(keyinput6), .B1(n6716), .B2(keyinput51), 
        .ZN(n6715) );
  OAI221_X1 U7702 ( .B1(n6717), .B2(keyinput6), .C1(n6716), .C2(keyinput51), 
        .A(n6715), .ZN(n6718) );
  NOR4_X1 U7703 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6738)
         );
  AOI22_X1 U7704 ( .A1(n6724), .A2(keyinput91), .B1(keyinput54), .B2(n6723), 
        .ZN(n6722) );
  OAI221_X1 U7705 ( .B1(n6724), .B2(keyinput91), .C1(n6723), .C2(keyinput54), 
        .A(n6722), .ZN(n6736) );
  AOI22_X1 U7706 ( .A1(n6726), .A2(keyinput122), .B1(keyinput7), .B2(n5580), 
        .ZN(n6725) );
  OAI221_X1 U7707 ( .B1(n6726), .B2(keyinput122), .C1(n5580), .C2(keyinput7), 
        .A(n6725), .ZN(n6735) );
  AOI22_X1 U7708 ( .A1(n6729), .A2(keyinput19), .B1(keyinput68), .B2(n6728), 
        .ZN(n6727) );
  OAI221_X1 U7709 ( .B1(n6729), .B2(keyinput19), .C1(n6728), .C2(keyinput68), 
        .A(n6727), .ZN(n6734) );
  AOI22_X1 U7710 ( .A1(n6732), .A2(keyinput34), .B1(keyinput74), .B2(n6731), 
        .ZN(n6730) );
  OAI221_X1 U7711 ( .B1(n6732), .B2(keyinput34), .C1(n6731), .C2(keyinput74), 
        .A(n6730), .ZN(n6733) );
  NOR4_X1 U7712 ( .A1(n6736), .A2(n6735), .A3(n6734), .A4(n6733), .ZN(n6737)
         );
  NAND4_X1 U7713 ( .A1(n6740), .A2(n6739), .A3(n6738), .A4(n6737), .ZN(n6941)
         );
  AOI22_X1 U7714 ( .A1(n6743), .A2(keyinput64), .B1(n6742), .B2(keyinput22), 
        .ZN(n6741) );
  OAI221_X1 U7715 ( .B1(n6743), .B2(keyinput64), .C1(n6742), .C2(keyinput22), 
        .A(n6741), .ZN(n6755) );
  AOI22_X1 U7716 ( .A1(n4324), .A2(keyinput21), .B1(keyinput90), .B2(n6745), 
        .ZN(n6744) );
  OAI221_X1 U7717 ( .B1(n4324), .B2(keyinput21), .C1(n6745), .C2(keyinput90), 
        .A(n6744), .ZN(n6754) );
  AOI22_X1 U7718 ( .A1(n6748), .A2(keyinput31), .B1(n6747), .B2(keyinput119), 
        .ZN(n6746) );
  OAI221_X1 U7719 ( .B1(n6748), .B2(keyinput31), .C1(n6747), .C2(keyinput119), 
        .A(n6746), .ZN(n6753) );
  INV_X1 U7720 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7721 ( .A1(n6751), .A2(keyinput121), .B1(n6750), .B2(keyinput42), 
        .ZN(n6749) );
  OAI221_X1 U7722 ( .B1(n6751), .B2(keyinput121), .C1(n6750), .C2(keyinput42), 
        .A(n6749), .ZN(n6752) );
  NOR4_X1 U7723 ( .A1(n6755), .A2(n6754), .A3(n6753), .A4(n6752), .ZN(n6805)
         );
  INV_X1 U7724 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6757) );
  AOI22_X1 U7725 ( .A1(n6758), .A2(keyinput67), .B1(n6757), .B2(keyinput100), 
        .ZN(n6756) );
  OAI221_X1 U7726 ( .B1(n6758), .B2(keyinput67), .C1(n6757), .C2(keyinput100), 
        .A(n6756), .ZN(n6770) );
  AOI22_X1 U7727 ( .A1(n6761), .A2(keyinput11), .B1(keyinput0), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7728 ( .B1(n6761), .B2(keyinput11), .C1(n6760), .C2(keyinput0), 
        .A(n6759), .ZN(n6769) );
  AOI22_X1 U7729 ( .A1(n4588), .A2(keyinput78), .B1(keyinput18), .B2(n6763), 
        .ZN(n6762) );
  OAI221_X1 U7730 ( .B1(n4588), .B2(keyinput78), .C1(n6763), .C2(keyinput18), 
        .A(n6762), .ZN(n6768) );
  AOI22_X1 U7731 ( .A1(n6766), .A2(keyinput24), .B1(n6765), .B2(keyinput20), 
        .ZN(n6764) );
  OAI221_X1 U7732 ( .B1(n6766), .B2(keyinput24), .C1(n6765), .C2(keyinput20), 
        .A(n6764), .ZN(n6767) );
  NOR4_X1 U7733 ( .A1(n6770), .A2(n6769), .A3(n6768), .A4(n6767), .ZN(n6804)
         );
  AOI22_X1 U7734 ( .A1(n5313), .A2(keyinput73), .B1(keyinput13), .B2(n6772), 
        .ZN(n6771) );
  OAI221_X1 U7735 ( .B1(n5313), .B2(keyinput73), .C1(n6772), .C2(keyinput13), 
        .A(n6771), .ZN(n6785) );
  AOI22_X1 U7736 ( .A1(n6775), .A2(keyinput28), .B1(n6774), .B2(keyinput111), 
        .ZN(n6773) );
  OAI221_X1 U7737 ( .B1(n6775), .B2(keyinput28), .C1(n6774), .C2(keyinput111), 
        .A(n6773), .ZN(n6784) );
  AOI22_X1 U7738 ( .A1(n6778), .A2(keyinput12), .B1(n6777), .B2(keyinput62), 
        .ZN(n6776) );
  OAI221_X1 U7739 ( .B1(n6778), .B2(keyinput12), .C1(n6777), .C2(keyinput62), 
        .A(n6776), .ZN(n6783) );
  INV_X1 U7740 ( .A(BS16_N), .ZN(n6780) );
  AOI22_X1 U7741 ( .A1(n6781), .A2(keyinput49), .B1(keyinput5), .B2(n6780), 
        .ZN(n6779) );
  OAI221_X1 U7742 ( .B1(n6781), .B2(keyinput49), .C1(n6780), .C2(keyinput5), 
        .A(n6779), .ZN(n6782) );
  NOR4_X1 U7743 ( .A1(n6785), .A2(n6784), .A3(n6783), .A4(n6782), .ZN(n6803)
         );
  AOI22_X1 U7744 ( .A1(n6788), .A2(keyinput109), .B1(keyinput106), .B2(n6787), 
        .ZN(n6786) );
  OAI221_X1 U7745 ( .B1(n6788), .B2(keyinput109), .C1(n6787), .C2(keyinput106), 
        .A(n6786), .ZN(n6801) );
  INV_X1 U7746 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6791) );
  AOI22_X1 U7747 ( .A1(n6791), .A2(keyinput81), .B1(n6790), .B2(keyinput60), 
        .ZN(n6789) );
  OAI221_X1 U7748 ( .B1(n6791), .B2(keyinput81), .C1(n6790), .C2(keyinput60), 
        .A(n6789), .ZN(n6800) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7750 ( .A1(n6794), .A2(keyinput4), .B1(n6793), .B2(keyinput120), 
        .ZN(n6792) );
  OAI221_X1 U7751 ( .B1(n6794), .B2(keyinput4), .C1(n6793), .C2(keyinput120), 
        .A(n6792), .ZN(n6799) );
  XOR2_X1 U7752 ( .A(n6795), .B(keyinput59), .Z(n6797) );
  XNOR2_X1 U7753 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput45), .ZN(
        n6796) );
  NAND2_X1 U7754 ( .A1(n6797), .A2(n6796), .ZN(n6798) );
  NOR4_X1 U7755 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(n6802)
         );
  NAND4_X1 U7756 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6940)
         );
  AOI22_X1 U7757 ( .A1(n6808), .A2(keyinput96), .B1(keyinput80), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7758 ( .B1(n6808), .B2(keyinput96), .C1(n6807), .C2(keyinput80), 
        .A(n6806), .ZN(n6821) );
  AOI22_X1 U7759 ( .A1(n6811), .A2(keyinput71), .B1(keyinput103), .B2(n6810), 
        .ZN(n6809) );
  OAI221_X1 U7760 ( .B1(n6811), .B2(keyinput71), .C1(n6810), .C2(keyinput103), 
        .A(n6809), .ZN(n6820) );
  INV_X1 U7761 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6814) );
  AOI22_X1 U7762 ( .A1(n6814), .A2(keyinput32), .B1(keyinput107), .B2(n6813), 
        .ZN(n6812) );
  OAI221_X1 U7763 ( .B1(n6814), .B2(keyinput32), .C1(n6813), .C2(keyinput107), 
        .A(n6812), .ZN(n6819) );
  INV_X1 U7764 ( .A(DATAI_27_), .ZN(n6817) );
  AOI22_X1 U7765 ( .A1(n6817), .A2(keyinput48), .B1(n6816), .B2(keyinput50), 
        .ZN(n6815) );
  OAI221_X1 U7766 ( .B1(n6817), .B2(keyinput48), .C1(n6816), .C2(keyinput50), 
        .A(n6815), .ZN(n6818) );
  NOR4_X1 U7767 ( .A1(n6821), .A2(n6820), .A3(n6819), .A4(n6818), .ZN(n6873)
         );
  INV_X1 U7768 ( .A(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n6823) );
  AOI22_X1 U7769 ( .A1(n6824), .A2(keyinput82), .B1(n6823), .B2(keyinput95), 
        .ZN(n6822) );
  OAI221_X1 U7770 ( .B1(n6824), .B2(keyinput82), .C1(n6823), .C2(keyinput95), 
        .A(n6822), .ZN(n6837) );
  AOI22_X1 U7771 ( .A1(n6827), .A2(keyinput36), .B1(keyinput85), .B2(n6826), 
        .ZN(n6825) );
  OAI221_X1 U7772 ( .B1(n6827), .B2(keyinput36), .C1(n6826), .C2(keyinput85), 
        .A(n6825), .ZN(n6836) );
  AOI22_X1 U7773 ( .A1(n6830), .A2(keyinput37), .B1(keyinput8), .B2(n6829), 
        .ZN(n6828) );
  OAI221_X1 U7774 ( .B1(n6830), .B2(keyinput37), .C1(n6829), .C2(keyinput8), 
        .A(n6828), .ZN(n6835) );
  INV_X1 U7775 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6833) );
  AOI22_X1 U7776 ( .A1(n6833), .A2(keyinput110), .B1(keyinput52), .B2(n6832), 
        .ZN(n6831) );
  OAI221_X1 U7777 ( .B1(n6833), .B2(keyinput110), .C1(n6832), .C2(keyinput52), 
        .A(n6831), .ZN(n6834) );
  NOR4_X1 U7778 ( .A1(n6837), .A2(n6836), .A3(n6835), .A4(n6834), .ZN(n6872)
         );
  INV_X1 U7779 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6839) );
  AOI22_X1 U7780 ( .A1(n6840), .A2(keyinput33), .B1(n6839), .B2(keyinput43), 
        .ZN(n6838) );
  OAI221_X1 U7781 ( .B1(n6840), .B2(keyinput33), .C1(n6839), .C2(keyinput43), 
        .A(n6838), .ZN(n6853) );
  AOI22_X1 U7782 ( .A1(n6843), .A2(keyinput35), .B1(keyinput29), .B2(n6842), 
        .ZN(n6841) );
  OAI221_X1 U7783 ( .B1(n6843), .B2(keyinput35), .C1(n6842), .C2(keyinput29), 
        .A(n6841), .ZN(n6852) );
  INV_X1 U7784 ( .A(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n6846) );
  AOI22_X1 U7785 ( .A1(n6846), .A2(keyinput99), .B1(keyinput102), .B2(n6845), 
        .ZN(n6844) );
  OAI221_X1 U7786 ( .B1(n6846), .B2(keyinput99), .C1(n6845), .C2(keyinput102), 
        .A(n6844), .ZN(n6851) );
  AOI22_X1 U7787 ( .A1(n6849), .A2(keyinput77), .B1(n6848), .B2(keyinput117), 
        .ZN(n6847) );
  OAI221_X1 U7788 ( .B1(n6849), .B2(keyinput77), .C1(n6848), .C2(keyinput117), 
        .A(n6847), .ZN(n6850) );
  NOR4_X1 U7789 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n6871)
         );
  INV_X1 U7790 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7791 ( .A1(n6856), .A2(keyinput93), .B1(n6855), .B2(keyinput47), 
        .ZN(n6854) );
  OAI221_X1 U7792 ( .B1(n6856), .B2(keyinput93), .C1(n6855), .C2(keyinput47), 
        .A(n6854), .ZN(n6869) );
  AOI22_X1 U7793 ( .A1(n6859), .A2(keyinput79), .B1(keyinput116), .B2(n6858), 
        .ZN(n6857) );
  OAI221_X1 U7794 ( .B1(n6859), .B2(keyinput79), .C1(n6858), .C2(keyinput116), 
        .A(n6857), .ZN(n6868) );
  AOI22_X1 U7795 ( .A1(n6862), .A2(keyinput10), .B1(n6861), .B2(keyinput69), 
        .ZN(n6860) );
  OAI221_X1 U7796 ( .B1(n6862), .B2(keyinput10), .C1(n6861), .C2(keyinput69), 
        .A(n6860), .ZN(n6867) );
  AOI22_X1 U7797 ( .A1(n6865), .A2(keyinput124), .B1(n6864), .B2(keyinput88), 
        .ZN(n6863) );
  OAI221_X1 U7798 ( .B1(n6865), .B2(keyinput124), .C1(n6864), .C2(keyinput88), 
        .A(n6863), .ZN(n6866) );
  NOR4_X1 U7799 ( .A1(n6869), .A2(n6868), .A3(n6867), .A4(n6866), .ZN(n6870)
         );
  NAND4_X1 U7800 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6939)
         );
  AOI22_X1 U7801 ( .A1(n6876), .A2(keyinput46), .B1(n6875), .B2(keyinput97), 
        .ZN(n6874) );
  OAI221_X1 U7802 ( .B1(n6876), .B2(keyinput46), .C1(n6875), .C2(keyinput97), 
        .A(n6874), .ZN(n6889) );
  AOI22_X1 U7803 ( .A1(n6879), .A2(keyinput86), .B1(keyinput92), .B2(n6878), 
        .ZN(n6877) );
  OAI221_X1 U7804 ( .B1(n6879), .B2(keyinput86), .C1(n6878), .C2(keyinput92), 
        .A(n6877), .ZN(n6888) );
  INV_X1 U7805 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U7806 ( .A1(n6882), .A2(keyinput105), .B1(n6881), .B2(keyinput53), 
        .ZN(n6880) );
  OAI221_X1 U7807 ( .B1(n6882), .B2(keyinput105), .C1(n6881), .C2(keyinput53), 
        .A(n6880), .ZN(n6887) );
  XOR2_X1 U7808 ( .A(n6883), .B(keyinput126), .Z(n6885) );
  XNOR2_X1 U7809 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(keyinput27), .ZN(
        n6884) );
  NAND2_X1 U7810 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  NOR4_X1 U7811 ( .A1(n6889), .A2(n6888), .A3(n6887), .A4(n6886), .ZN(n6937)
         );
  INV_X1 U7812 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6892) );
  AOI22_X1 U7813 ( .A1(n6892), .A2(keyinput39), .B1(keyinput15), .B2(n6891), 
        .ZN(n6890) );
  OAI221_X1 U7814 ( .B1(n6892), .B2(keyinput39), .C1(n6891), .C2(keyinput15), 
        .A(n6890), .ZN(n6904) );
  INV_X1 U7815 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6895) );
  AOI22_X1 U7816 ( .A1(n6895), .A2(keyinput16), .B1(keyinput114), .B2(n6894), 
        .ZN(n6893) );
  OAI221_X1 U7817 ( .B1(n6895), .B2(keyinput16), .C1(n6894), .C2(keyinput114), 
        .A(n6893), .ZN(n6903) );
  AOI22_X1 U7818 ( .A1(n4376), .A2(keyinput63), .B1(keyinput101), .B2(n6897), 
        .ZN(n6896) );
  OAI221_X1 U7819 ( .B1(n4376), .B2(keyinput63), .C1(n6897), .C2(keyinput101), 
        .A(n6896), .ZN(n6902) );
  INV_X1 U7820 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6900) );
  AOI22_X1 U7821 ( .A1(n6900), .A2(keyinput87), .B1(n6899), .B2(keyinput65), 
        .ZN(n6898) );
  OAI221_X1 U7822 ( .B1(n6900), .B2(keyinput87), .C1(n6899), .C2(keyinput65), 
        .A(n6898), .ZN(n6901) );
  NOR4_X1 U7823 ( .A1(n6904), .A2(n6903), .A3(n6902), .A4(n6901), .ZN(n6936)
         );
  AOI22_X1 U7824 ( .A1(n6907), .A2(keyinput75), .B1(keyinput98), .B2(n6906), 
        .ZN(n6905) );
  OAI221_X1 U7825 ( .B1(n6907), .B2(keyinput75), .C1(n6906), .C2(keyinput98), 
        .A(n6905), .ZN(n6918) );
  AOI22_X1 U7826 ( .A1(n6909), .A2(keyinput125), .B1(keyinput84), .B2(n4771), 
        .ZN(n6908) );
  OAI221_X1 U7827 ( .B1(n6909), .B2(keyinput125), .C1(n4771), .C2(keyinput84), 
        .A(n6908), .ZN(n6917) );
  AOI22_X1 U7828 ( .A1(n6912), .A2(keyinput72), .B1(n6911), .B2(keyinput108), 
        .ZN(n6910) );
  OAI221_X1 U7829 ( .B1(n6912), .B2(keyinput72), .C1(n6911), .C2(keyinput108), 
        .A(n6910), .ZN(n6916) );
  AOI22_X1 U7830 ( .A1(n3478), .A2(keyinput23), .B1(n6914), .B2(keyinput58), 
        .ZN(n6913) );
  OAI221_X1 U7831 ( .B1(n3478), .B2(keyinput23), .C1(n6914), .C2(keyinput58), 
        .A(n6913), .ZN(n6915) );
  NOR4_X1 U7832 ( .A1(n6918), .A2(n6917), .A3(n6916), .A4(n6915), .ZN(n6935)
         );
  AOI22_X1 U7833 ( .A1(n6921), .A2(keyinput104), .B1(n6920), .B2(keyinput1), 
        .ZN(n6919) );
  OAI221_X1 U7834 ( .B1(n6921), .B2(keyinput104), .C1(n6920), .C2(keyinput1), 
        .A(n6919), .ZN(n6933) );
  AOI22_X1 U7835 ( .A1(n6924), .A2(keyinput44), .B1(keyinput41), .B2(n6923), 
        .ZN(n6922) );
  OAI221_X1 U7836 ( .B1(n6924), .B2(keyinput44), .C1(n6923), .C2(keyinput41), 
        .A(n6922), .ZN(n6932) );
  INV_X1 U7837 ( .A(DATAI_21_), .ZN(n6927) );
  INV_X1 U7838 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U7839 ( .A1(n6927), .A2(keyinput57), .B1(n6926), .B2(keyinput118), 
        .ZN(n6925) );
  OAI221_X1 U7840 ( .B1(n6927), .B2(keyinput57), .C1(n6926), .C2(keyinput118), 
        .A(n6925), .ZN(n6931) );
  INV_X1 U7841 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6929) );
  AOI22_X1 U7842 ( .A1(n6929), .A2(keyinput70), .B1(keyinput17), .B2(n4225), 
        .ZN(n6928) );
  OAI221_X1 U7843 ( .B1(n6929), .B2(keyinput70), .C1(n4225), .C2(keyinput17), 
        .A(n6928), .ZN(n6930) );
  NOR4_X1 U7844 ( .A1(n6933), .A2(n6932), .A3(n6931), .A4(n6930), .ZN(n6934)
         );
  NAND4_X1 U7845 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6938)
         );
  NOR4_X1 U7846 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n6942)
         );
  XNOR2_X1 U7847 ( .A(n6943), .B(n6942), .ZN(n6959) );
  NAND2_X1 U7848 ( .A1(n6945), .A2(n6944), .ZN(n6949) );
  NAND2_X1 U7849 ( .A1(n6947), .A2(n6946), .ZN(n6948) );
  OAI211_X1 U7850 ( .C1(n6951), .C2(n6950), .A(n6949), .B(n6948), .ZN(n6955)
         );
  NOR2_X1 U7851 ( .A1(n6953), .A2(n6952), .ZN(n6954) );
  AOI211_X1 U7852 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n6956), .A(n6955), 
        .B(n6954), .ZN(n6957) );
  INV_X1 U7853 ( .A(n6957), .ZN(n6958) );
  XNOR2_X1 U7854 ( .A(n6959), .B(n6958), .ZN(U3143) );
  CLKBUF_X1 U3552 ( .A(n3338), .Z(n3395) );
  CLKBUF_X1 U3556 ( .A(n3238), .Z(n3996) );
  CLKBUF_X1 U3598 ( .A(n3698), .Z(n5427) );
  CLKBUF_X1 U3680 ( .A(n3991), .Z(n5983) );
  CLKBUF_X1 U3770 ( .A(n4208), .Z(n4558) );
  CLKBUF_X1 U3825 ( .A(n4231), .Z(n6434) );
  CLKBUF_X1 U3830 ( .A(n3703), .Z(n4027) );
  INV_X2 U3887 ( .A(n5382), .ZN(n6005) );
  OAI211_X2 U3896 ( .C1(n5750), .C2(n4036), .A(n4035), .B(n6104), .ZN(n5382)
         );
endmodule

