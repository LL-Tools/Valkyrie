

module b15_C_SARLock_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117,
         n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137,
         n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147,
         n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157,
         n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
         n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
         n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
         n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
         n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207,
         n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217,
         n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
         n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
         n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247,
         n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
         n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267,
         n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277,
         n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287,
         n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297,
         n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307,
         n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317,
         n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327,
         n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347,
         n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357,
         n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367,
         n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
         n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
         n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
         n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
         n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437,
         n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447,
         n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457,
         n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467,
         n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477,
         n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
         n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
         n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527,
         n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537,
         n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547,
         n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557,
         n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567,
         n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577,
         n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587,
         n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
         n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607,
         n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617,
         n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627,
         n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637,
         n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647,
         n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
         n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
         n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
         n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
         n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697,
         n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727,
         n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047;

  NAND2_X1 U3575 ( .A1(n5680), .A2(n4374), .ZN(n4483) );
  NAND2_X2 U3576 ( .A1(n6010), .A2(n5765), .ZN(n6269) );
  NAND2_X1 U3577 ( .A1(n3725), .A2(n3724), .ZN(n4692) );
  NAND2_X1 U3578 ( .A1(n4557), .A2(n4217), .ZN(n4339) );
  NAND2_X1 U3579 ( .A1(n3478), .A2(n3477), .ZN(n3530) );
  INV_X1 U3580 ( .A(n3745), .ZN(n4756) );
  CLKBUF_X2 U3581 ( .A(n3318), .Z(n4166) );
  CLKBUF_X1 U3582 ( .A(n3416), .Z(n4398) );
  CLKBUF_X2 U3583 ( .A(n3345), .Z(n4403) );
  CLKBUF_X2 U3584 ( .A(n3270), .Z(n4014) );
  CLKBUF_X2 U3585 ( .A(n3271), .Z(n4937) );
  CLKBUF_X2 U3586 ( .A(n3411), .Z(n4031) );
  CLKBUF_X2 U3587 ( .A(n3269), .Z(n3133) );
  CLKBUF_X2 U3588 ( .A(n3998), .Z(n4432) );
  CLKBUF_X2 U3589 ( .A(n4122), .Z(n4433) );
  CLKBUF_X2 U3590 ( .A(n3287), .Z(n4431) );
  INV_X1 U3591 ( .A(n3371), .ZN(n3385) );
  AND4_X1 U3592 ( .A1(n3344), .A2(n3343), .A3(n3342), .A4(n3341), .ZN(n3351)
         );
  AND2_X2 U3593 ( .A1(n4934), .A2(n4952), .ZN(n3269) );
  AND2_X2 U3594 ( .A1(n5361), .A2(n4951), .ZN(n3272) );
  AND2_X1 U3595 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4951) );
  AND2_X1 U3596 ( .A1(n3683), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3222)
         );
  CLKBUF_X1 U3597 ( .A(n6151), .Z(n3126) );
  NOR2_X1 U3598 ( .A1(n5152), .A2(n4499), .ZN(n6151) );
  AND2_X1 U3600 ( .A1(n3373), .A2(n3371), .ZN(n5437) );
  OAI22_X1 U3601 ( .A1(n6747), .A2(keyinput51), .B1(n6746), .B2(keyinput120), 
        .ZN(n6745) );
  AND2_X1 U3602 ( .A1(n5508), .A2(n5404), .ZN(n5497) );
  AOI221_X1 U3604 ( .B1(n6747), .B2(keyinput51), .C1(keyinput120), .C2(n6746), 
        .A(n6745), .ZN(n6760) );
  NOR2_X2 U3605 ( .A1(n3371), .A2(n4217), .ZN(n3388) );
  CLKBUF_X2 U3606 ( .A(n4265), .Z(n4672) );
  INV_X1 U3607 ( .A(n3389), .ZN(n4453) );
  NOR2_X2 U3608 ( .A1(n5458), .A2(n5449), .ZN(n5906) );
  NOR2_X1 U3609 ( .A1(n4707), .A2(n5753), .ZN(n6317) );
  INV_X1 U3610 ( .A(n6108), .ZN(n6146) );
  OR2_X1 U3611 ( .A1(n4519), .A2(n4181), .ZN(n5537) );
  OR2_X1 U3612 ( .A1(n5196), .A2(n5195), .ZN(n3127) );
  INV_X1 U3613 ( .A(n3357), .ZN(n3359) );
  AND2_X4 U3614 ( .A1(n4981), .A2(n5119), .ZN(n5118) );
  NAND2_X2 U3615 ( .A1(n3407), .A2(n3406), .ZN(n3484) );
  AND2_X1 U3616 ( .A1(n4952), .A2(n4930), .ZN(n3470) );
  NAND2_X2 U3617 ( .A1(n5953), .A2(n5575), .ZN(n5612) );
  AOI21_X1 U3618 ( .B1(n4697), .B2(n4698), .A(n3540), .ZN(n6225) );
  NAND2_X1 U3619 ( .A1(n3508), .A2(n3509), .ZN(n3545) );
  CLKBUF_X2 U3620 ( .A(n4592), .Z(n4638) );
  AND2_X1 U3621 ( .A1(n3384), .A2(n3383), .ZN(n4195) );
  INV_X1 U3622 ( .A(n3132), .ZN(n3128) );
  NAND2_X2 U3624 ( .A1(n3306), .A2(n3359), .ZN(n4455) );
  INV_X2 U3625 ( .A(n3268), .ZN(n3306) );
  CLKBUF_X2 U3626 ( .A(n3272), .Z(n4424) );
  BUF_X2 U3627 ( .A(n3470), .Z(n4426) );
  INV_X2 U3628 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3217) );
  AOI22_X1 U3629 ( .A1(n3658), .A2(n5558), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5977), .ZN(n3659) );
  AND2_X1 U3630 ( .A1(n5568), .A2(n3188), .ZN(n5549) );
  OR2_X1 U3631 ( .A1(n3656), .A2(n3657), .ZN(n5558) );
  XNOR2_X1 U3632 ( .A(n4524), .B(n4523), .ZN(n5382) );
  NAND2_X1 U3633 ( .A1(n3177), .A2(n3178), .ZN(n5952) );
  XNOR2_X1 U3634 ( .A(n4512), .B(n4452), .ZN(n5556) );
  AND2_X1 U3635 ( .A1(n5493), .A2(n5495), .ZN(n5860) );
  NAND2_X1 U3636 ( .A1(n3198), .A2(n3153), .ZN(n5492) );
  INV_X1 U3637 ( .A(n5395), .ZN(n3198) );
  AOI21_X1 U3638 ( .B1(n3165), .B2(n3167), .A(n3163), .ZN(n3162) );
  AOI21_X1 U3639 ( .B1(n3174), .B2(n3172), .A(n3154), .ZN(n3171) );
  OAI21_X1 U3640 ( .B1(n3634), .B2(n3167), .A(n5179), .ZN(n3166) );
  NAND2_X1 U3641 ( .A1(n3793), .A2(n3792), .ZN(n4827) );
  INV_X2 U3642 ( .A(n3138), .ZN(n5584) );
  XNOR2_X1 U3643 ( .A(n3629), .B(n3617), .ZN(n3783) );
  AOI21_X1 U3644 ( .B1(n3542), .B2(n6225), .A(n3541), .ZN(n6215) );
  NAND2_X1 U3645 ( .A1(n3755), .A2(n3754), .ZN(n4653) );
  INV_X1 U3646 ( .A(n3566), .ZN(n3590) );
  XNOR2_X1 U3647 ( .A(n3566), .B(n3588), .ZN(n3763) );
  AND2_X1 U3648 ( .A1(n3528), .A2(n3539), .ZN(n4697) );
  NAND2_X1 U3649 ( .A1(n3780), .A2(n3779), .ZN(n4718) );
  OAI21_X1 U3650 ( .B1(n4754), .B2(n3904), .A(n4095), .ZN(n3760) );
  NAND2_X1 U3651 ( .A1(n3546), .A2(n4769), .ZN(n3566) );
  INV_X1 U3652 ( .A(n3545), .ZN(n3546) );
  AND2_X1 U3653 ( .A1(n5332), .A2(n5331), .ZN(n5472) );
  NOR2_X1 U3654 ( .A1(n4808), .A2(n4957), .ZN(n6560) );
  NAND2_X1 U3655 ( .A1(n5379), .A2(n4664), .ZN(n5924) );
  NOR2_X1 U3656 ( .A1(n5075), .A2(n3423), .ZN(n6536) );
  NAND2_X2 U3657 ( .A1(n3389), .A2(n6163), .ZN(n5531) );
  NOR2_X1 U3658 ( .A1(n5075), .A2(n4747), .ZN(n6521) );
  NAND2_X2 U3659 ( .A1(n4560), .A2(n3385), .ZN(n4611) );
  OR2_X1 U3660 ( .A1(n4215), .A2(n4214), .ZN(n4385) );
  NAND2_X1 U3661 ( .A1(n3460), .A2(n3627), .ZN(n3531) );
  AOI21_X1 U3662 ( .B1(n3402), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3405), 
        .ZN(n3408) );
  NAND2_X1 U3663 ( .A1(n4279), .A2(n4278), .ZN(n5168) );
  INV_X1 U3664 ( .A(n5166), .ZN(n4279) );
  INV_X1 U3666 ( .A(n5165), .ZN(n4278) );
  AND3_X1 U3667 ( .A1(n4211), .A2(n4217), .A3(n4210), .ZN(n4547) );
  NAND2_X2 U3668 ( .A1(n4195), .A2(n3386), .ZN(n4219) );
  INV_X1 U3669 ( .A(n3382), .ZN(n4211) );
  OR2_X1 U3670 ( .A1(n3687), .A2(n3686), .ZN(n3693) );
  AND2_X1 U3671 ( .A1(n3305), .A2(n3304), .ZN(n3384) );
  AND3_X1 U3672 ( .A1(n3361), .A2(n4223), .A3(n3367), .ZN(n3364) );
  OAI21_X1 U3673 ( .B1(n4269), .B2(n4271), .A(n4270), .ZN(n4641) );
  NAND2_X1 U3674 ( .A1(n3457), .A2(n3456), .ZN(n3518) );
  NOR2_X1 U3675 ( .A1(n3660), .A2(n3140), .ZN(n3378) );
  NAND2_X1 U3676 ( .A1(n4455), .A2(n3423), .ZN(n3355) );
  INV_X1 U3677 ( .A(n4339), .ZN(n4265) );
  OR2_X1 U3678 ( .A1(n4688), .A2(n5367), .ZN(n4383) );
  NAND2_X1 U3679 ( .A1(n3492), .A2(n3491), .ZN(n3722) );
  AND2_X2 U3680 ( .A1(n3385), .A2(n4217), .ZN(n5383) );
  CLKBUF_X1 U3681 ( .A(n3359), .Z(n3360) );
  NAND2_X1 U3682 ( .A1(n3688), .A2(n4382), .ZN(n3703) );
  AND2_X1 U3683 ( .A1(n3423), .A2(n3357), .ZN(n3690) );
  OR2_X1 U3684 ( .A1(n3476), .A2(n3475), .ZN(n3534) );
  OR2_X1 U3685 ( .A1(n3451), .A2(n3450), .ZN(n3533) );
  INV_X1 U3686 ( .A(n3373), .ZN(n4779) );
  OR2_X1 U3687 ( .A1(n3440), .A2(n3439), .ZN(n3621) );
  AND2_X1 U3688 ( .A1(n4217), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3688) );
  CLKBUF_X1 U3689 ( .A(n3362), .Z(n4382) );
  AND2_X1 U3690 ( .A1(n3373), .A2(n4747), .ZN(n4223) );
  INV_X1 U3691 ( .A(n4217), .ZN(n3129) );
  AND4_X2 U3692 ( .A1(n3255), .A2(n3141), .A3(n3254), .A4(n3253), .ZN(n3268)
         );
  AND4_X2 U3693 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n4747)
         );
  NAND2_X1 U3694 ( .A1(n3212), .A2(n3139), .ZN(n3373) );
  NAND4_X2 U3695 ( .A1(n3330), .A2(n3329), .A3(n3328), .A4(n3327), .ZN(n3371)
         );
  AND4_X1 U3696 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3329)
         );
  AND4_X1 U3697 ( .A1(n3231), .A2(n3230), .A3(n3229), .A4(n3228), .ZN(n3213)
         );
  AND4_X1 U3698 ( .A1(n3248), .A2(n3247), .A3(n3246), .A4(n3245), .ZN(n3254)
         );
  AND4_X1 U3699 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3353)
         );
  AND4_X1 U3700 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3281)
         );
  AND4_X1 U3701 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3300)
         );
  AND4_X1 U3702 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3302)
         );
  AND4_X1 U3703 ( .A1(n3240), .A2(n3239), .A3(n3238), .A4(n3237), .ZN(n3255)
         );
  AND4_X1 U3704 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3330)
         );
  AND4_X1 U3705 ( .A1(n3235), .A2(n3234), .A3(n3233), .A4(n3232), .ZN(n3236)
         );
  AND4_X1 U3706 ( .A1(n3322), .A2(n3321), .A3(n3320), .A4(n3319), .ZN(n3328)
         );
  AND4_X1 U3707 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3301)
         );
  AND4_X1 U3708 ( .A1(n3326), .A2(n3325), .A3(n3324), .A4(n3323), .ZN(n3327)
         );
  AND4_X1 U3709 ( .A1(n3252), .A2(n3251), .A3(n3250), .A4(n3249), .ZN(n3253)
         );
  INV_X2 U3710 ( .A(n5955), .ZN(n6226) );
  AND4_X1 U3711 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3352)
         );
  AND4_X1 U3712 ( .A1(n3285), .A2(n3284), .A3(n3283), .A4(n3282), .ZN(n3303)
         );
  AND4_X1 U3713 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3350)
         );
  BUF_X2 U3714 ( .A(n3286), .Z(n4425) );
  BUF_X2 U3715 ( .A(n3335), .Z(n4435) );
  AND2_X2 U3716 ( .A1(n3222), .A2(n3223), .ZN(n3345) );
  AND2_X2 U3717 ( .A1(n4930), .A2(n4917), .ZN(n3271) );
  AND2_X2 U3718 ( .A1(n3223), .A2(n5361), .ZN(n3998) );
  AND2_X2 U3719 ( .A1(n3222), .A2(n4951), .ZN(n3411) );
  AND2_X2 U3720 ( .A1(n4934), .A2(n5361), .ZN(n3286) );
  BUF_X2 U3721 ( .A(n3445), .Z(n4127) );
  AND2_X2 U3722 ( .A1(n4917), .A2(n4951), .ZN(n4122) );
  AND2_X2 U3723 ( .A1(n3217), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4934)
         );
  CLKBUF_X1 U3724 ( .A(n4540), .Z(n6456) );
  AND2_X2 U3725 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4917) );
  OR2_X1 U3726 ( .A1(n3509), .A2(n3508), .ZN(n3510) );
  NAND2_X2 U3727 ( .A1(n3762), .A2(n3761), .ZN(n4651) );
  AND2_X4 U3728 ( .A1(n3782), .A2(n4715), .ZN(n4742) );
  OR2_X2 U3729 ( .A1(n5474), .A2(n5460), .ZN(n5458) );
  NOR2_X2 U3730 ( .A1(n5415), .A2(n3201), .ZN(n5504) );
  AND2_X4 U3731 ( .A1(n3223), .A2(n4952), .ZN(n3336) );
  AND2_X1 U3732 ( .A1(n4952), .A2(n4930), .ZN(n3130) );
  AND2_X1 U3733 ( .A1(n4952), .A2(n4930), .ZN(n3131) );
  NAND2_X2 U3734 ( .A1(n5523), .A2(n5524), .ZN(n5415) );
  NOR2_X4 U3735 ( .A1(n5429), .A2(n5902), .ZN(n5523) );
  AND2_X4 U3736 ( .A1(n4934), .A2(n4917), .ZN(n3318) );
  NOR2_X1 U3737 ( .A1(n5561), .A2(n3136), .ZN(n5925) );
  NOR2_X4 U3738 ( .A1(n5492), .A2(n5562), .ZN(n5561) );
  XNOR2_X2 U3739 ( .A(n3465), .B(n3464), .ZN(n4750) );
  AOI21_X4 U3740 ( .B1(n5299), .B2(n5326), .A(n5327), .ZN(n5325) );
  NAND2_X2 U3741 ( .A1(n5298), .A2(n5300), .ZN(n5299) );
  OR2_X1 U3742 ( .A1(n3459), .A2(n6611), .ZN(n3627) );
  NAND2_X1 U3743 ( .A1(n3423), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3492) );
  NOR2_X1 U3744 ( .A1(n3175), .A2(n5317), .ZN(n3174) );
  INV_X1 U3745 ( .A(n3638), .ZN(n3175) );
  NAND2_X1 U3746 ( .A1(n3357), .A2(n4557), .ZN(n3664) );
  NAND2_X1 U3747 ( .A1(n3129), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3491) );
  OR2_X1 U3748 ( .A1(n6702), .A2(n4476), .ZN(n6096) );
  OR2_X1 U3749 ( .A1(n4559), .A2(n4558), .ZN(n4662) );
  AND2_X1 U3750 ( .A1(n5561), .A2(n3207), .ZN(n4512) );
  AND2_X1 U3751 ( .A1(n4517), .A2(n4180), .ZN(n3207) );
  INV_X1 U3752 ( .A(n5690), .ZN(n3653) );
  INV_X1 U3753 ( .A(n3644), .ZN(n3182) );
  AND2_X1 U3754 ( .A1(n4211), .A2(n4210), .ZN(n4686) );
  INV_X1 U3755 ( .A(n6617), .ZN(n4681) );
  INV_X1 U3756 ( .A(n5556), .ZN(n5378) );
  OAI211_X1 U3757 ( .C1(n3362), .C2(n3363), .A(n3389), .B(n4455), .ZN(n3660)
         );
  AND2_X1 U3758 ( .A1(n3388), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3160) );
  AND2_X1 U3759 ( .A1(n3602), .A2(n3601), .ZN(n3605) );
  NAND2_X1 U3760 ( .A1(n3558), .A2(n3557), .ZN(n3588) );
  NAND2_X1 U3761 ( .A1(n3356), .A2(n3389), .ZN(n3382) );
  AND2_X2 U3762 ( .A1(n4929), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4930)
         );
  NOR2_X1 U3763 ( .A1(n3267), .A2(n4453), .ZN(n3305) );
  AND2_X1 U3764 ( .A1(n3373), .A2(n3363), .ZN(n3267) );
  NAND2_X1 U3765 ( .A1(n3309), .A2(n3308), .ZN(n3383) );
  INV_X1 U3766 ( .A(n3703), .ZN(n3715) );
  NOR2_X1 U3767 ( .A1(n5352), .A2(n6611), .ZN(n4444) );
  INV_X1 U3768 ( .A(n3195), .ZN(n3193) );
  NOR2_X1 U3769 ( .A1(n5194), .A2(n3196), .ZN(n3195) );
  INV_X1 U3770 ( .A(n5128), .ZN(n3196) );
  NOR2_X1 U3771 ( .A1(n4863), .A2(n4983), .ZN(n3206) );
  INV_X1 U3772 ( .A(n3920), .ZN(n3904) );
  INV_X1 U3773 ( .A(n3752), .ZN(n4447) );
  OR2_X1 U3774 ( .A1(n3389), .A2(n6465), .ZN(n3210) );
  AND2_X1 U3775 ( .A1(n3268), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3920) );
  XNOR2_X1 U3776 ( .A(n3530), .B(n3529), .ZN(n3532) );
  NAND2_X1 U3777 ( .A1(n3490), .A2(n3489), .ZN(n4771) );
  NAND2_X1 U3778 ( .A1(n4547), .A2(n4567), .ZN(n4559) );
  INV_X1 U3779 ( .A(n6632), .ZN(n4673) );
  INV_X2 U3780 ( .A(n3210), .ZN(n4521) );
  AND2_X1 U3781 ( .A1(n5022), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4520) );
  OR2_X1 U3782 ( .A1(n4115), .A2(n4114), .ZN(n4155) );
  NAND2_X1 U3783 ( .A1(n3202), .A2(n5589), .ZN(n3201) );
  INV_X1 U3784 ( .A(n3204), .ZN(n3202) );
  INV_X1 U3785 ( .A(n5415), .ZN(n3203) );
  AND2_X1 U3786 ( .A1(n3959), .A2(n3200), .ZN(n3199) );
  NOR2_X1 U3787 ( .A1(n3892), .A2(n5308), .ZN(n3908) );
  AND2_X1 U3788 ( .A1(n4216), .A2(n3690), .ZN(n6593) );
  NAND2_X1 U3789 ( .A1(n3184), .A2(n3135), .ZN(n3183) );
  INV_X1 U3790 ( .A(n3179), .ZN(n3178) );
  OAI21_X1 U3791 ( .B1(n3135), .B2(n3180), .A(n3647), .ZN(n3179) );
  INV_X1 U3792 ( .A(n3174), .ZN(n3173) );
  INV_X1 U3793 ( .A(n3209), .ZN(n3172) );
  NAND2_X1 U3794 ( .A1(n3164), .A2(n3162), .ZN(n5290) );
  INV_X1 U3795 ( .A(n5261), .ZN(n3163) );
  INV_X1 U3796 ( .A(n5178), .ZN(n3167) );
  OR2_X1 U3797 ( .A1(n4865), .A2(n4864), .ZN(n4304) );
  NAND2_X1 U3798 ( .A1(n4920), .A2(n4385), .ZN(n6291) );
  INV_X1 U3799 ( .A(n6411), .ZN(n4957) );
  NOR2_X1 U3800 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4748), .ZN(n6411) );
  NAND2_X1 U3801 ( .A1(n3717), .A2(n4200), .ZN(n3725) );
  AND2_X1 U3802 ( .A1(n4501), .A2(n4500), .ZN(n4502) );
  NOR2_X1 U3803 ( .A1(n4527), .A2(n5351), .ZN(n4479) );
  AND2_X2 U3804 ( .A1(n4461), .A2(n4681), .ZN(n6163) );
  AND2_X1 U3805 ( .A1(n5379), .A2(n5368), .ZN(n6168) );
  AND2_X1 U3806 ( .A1(n5379), .A2(n4665), .ZN(n5547) );
  INV_X1 U3807 ( .A(n4516), .ZN(n4452) );
  OAI211_X1 U3808 ( .C1(n3190), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n3187), .B(n3185), .ZN(n4530) );
  NAND2_X1 U3809 ( .A1(n5568), .A2(n3151), .ZN(n3187) );
  NAND2_X1 U3810 ( .A1(n3190), .A2(n3186), .ZN(n3185) );
  AND2_X1 U3811 ( .A1(n4385), .A2(n4384), .ZN(n6310) );
  NAND2_X2 U3812 ( .A1(n3521), .A2(n3142), .ZN(n3745) );
  INV_X1 U3813 ( .A(n4540), .ZN(n6499) );
  AND2_X1 U3814 ( .A1(n4201), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3686) );
  NOR2_X1 U3815 ( .A1(n3388), .A2(n3678), .ZN(n3702) );
  NAND2_X1 U3816 ( .A1(n3385), .A2(n4199), .ZN(n3156) );
  OR2_X1 U3817 ( .A1(n3600), .A2(n3599), .ZN(n3619) );
  NAND2_X1 U3818 ( .A1(n3604), .A2(n3603), .ZN(n3629) );
  INV_X1 U3819 ( .A(n3605), .ZN(n3603) );
  OR2_X1 U3820 ( .A1(n3556), .A2(n3555), .ZN(n3608) );
  OR2_X1 U3821 ( .A1(n3576), .A2(n3575), .ZN(n3607) );
  NAND2_X1 U3822 ( .A1(n3354), .A2(n3388), .ZN(n3370) );
  NOR2_X1 U3823 ( .A1(n3677), .A2(n3676), .ZN(n3707) );
  NAND2_X1 U3824 ( .A1(n3159), .A2(n3158), .ZN(n3402) );
  NAND2_X1 U3825 ( .A1(n3161), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U3826 ( .A1(n3335), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3260) );
  INV_X1 U3827 ( .A(n5494), .ZN(n4139) );
  INV_X1 U3828 ( .A(n5397), .ZN(n4119) );
  NAND2_X1 U3829 ( .A1(n3205), .A2(n4030), .ZN(n3204) );
  INV_X1 U3830 ( .A(n5512), .ZN(n3205) );
  AND2_X1 U3831 ( .A1(n5457), .A2(n5475), .ZN(n3200) );
  INV_X1 U3832 ( .A(n3784), .ZN(n3791) );
  AND3_X1 U3833 ( .A1(n3661), .A2(n4223), .A3(n3663), .ZN(n4216) );
  AND2_X1 U3834 ( .A1(n5567), .A2(n4249), .ZN(n3188) );
  NAND2_X1 U3835 ( .A1(n3171), .A2(n3173), .ZN(n3170) );
  NAND2_X1 U3836 ( .A1(n4792), .A2(n4196), .ZN(n3157) );
  AND2_X1 U3837 ( .A1(n4223), .A2(n3360), .ZN(n4210) );
  INV_X1 U3838 ( .A(n3503), .ZN(n3504) );
  CLKBUF_X1 U3839 ( .A(n4930), .Z(n4933) );
  NAND2_X1 U3840 ( .A1(n3690), .A2(n5437), .ZN(n4687) );
  AOI21_X1 U3841 ( .B1(n6623), .B2(n4959), .A(n5362), .ZN(n4748) );
  INV_X1 U3842 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U3843 ( .A1(n3703), .A2(n3664), .ZN(n3717) );
  OR2_X1 U3844 ( .A1(n3709), .A2(n3671), .ZN(n3672) );
  AND2_X1 U3845 ( .A1(n6323), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3671)
         );
  AND2_X1 U3846 ( .A1(n4471), .A2(n4545), .ZN(n4543) );
  AND2_X1 U3847 ( .A1(n4235), .A2(n4234), .ZN(n4920) );
  INV_X1 U3848 ( .A(n4642), .ZN(n4375) );
  AND2_X1 U3849 ( .A1(n4325), .A2(n4324), .ZN(n5331) );
  AND2_X1 U3850 ( .A1(n4421), .A2(n4420), .ZN(n4517) );
  OR2_X1 U3851 ( .A1(n4535), .A2(n4447), .ZN(n4420) );
  AND2_X1 U3852 ( .A1(n5552), .A2(n4472), .ZN(n4449) );
  AND2_X1 U3853 ( .A1(n4496), .A2(n4472), .ZN(n4177) );
  NAND2_X1 U3854 ( .A1(n4093), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4115)
         );
  AND2_X1 U3855 ( .A1(n4078), .A2(n4077), .ZN(n5589) );
  AND2_X1 U3856 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4026), .ZN(n4027)
         );
  INV_X1 U3857 ( .A(n4025), .ZN(n4026) );
  AND2_X1 U3858 ( .A1(n4009), .A2(n4008), .ZN(n5524) );
  NOR2_X1 U3859 ( .A1(n3976), .A2(n5436), .ZN(n3977) );
  CLKBUF_X1 U3860 ( .A(n5429), .Z(n5430) );
  NAND2_X1 U3861 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3956), .ZN(n3976)
         );
  NOR2_X1 U3862 ( .A1(n3924), .A2(n3923), .ZN(n3955) );
  NAND2_X1 U3863 ( .A1(n3908), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3924)
         );
  NAND2_X1 U3864 ( .A1(n3137), .A2(n3891), .ZN(n5326) );
  AND3_X1 U3865 ( .A1(n3907), .A2(n3906), .A3(n3905), .ZN(n5327) );
  NAND2_X1 U3866 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3892)
         );
  INV_X1 U3867 ( .A(n3891), .ZN(n3194) );
  NAND2_X1 U3868 ( .A1(n3854), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3855)
         );
  INV_X1 U3869 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U3870 ( .A1(n6950), .A2(n3811), .ZN(n3854) );
  AND2_X1 U3871 ( .A1(n3829), .A2(n3828), .ZN(n4983) );
  CLKBUF_X1 U3872 ( .A(n4981), .Z(n4982) );
  NOR2_X1 U3873 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  INV_X1 U3874 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3785) );
  AND2_X1 U3875 ( .A1(n4740), .A2(n4741), .ZN(n3782) );
  NAND2_X1 U3876 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3767), .ZN(n3786)
         );
  NOR2_X1 U3877 ( .A1(n3773), .A2(n3768), .ZN(n3767) );
  CLKBUF_X1 U3878 ( .A(n4715), .Z(n4716) );
  INV_X1 U3879 ( .A(n3756), .ZN(n3774) );
  NAND2_X1 U3880 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3774), .ZN(n3773)
         );
  NAND2_X1 U3881 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3756) );
  NAND2_X1 U3882 ( .A1(n3744), .A2(n3743), .ZN(n4700) );
  AOI21_X1 U3883 ( .B1(n5568), .B2(n3148), .A(n3189), .ZN(n3186) );
  NOR2_X2 U3884 ( .A1(n5706), .A2(n4356), .ZN(n5508) );
  AND2_X1 U3885 ( .A1(n5906), .A2(n5907), .ZN(n5519) );
  NAND2_X1 U3886 ( .A1(n5472), .A2(n5471), .ZN(n5474) );
  NAND2_X1 U3887 ( .A1(n3642), .A2(n3641), .ZN(n3643) );
  AND2_X1 U3888 ( .A1(n4322), .A2(n4321), .ZN(n5301) );
  INV_X1 U3889 ( .A(n3166), .ZN(n3165) );
  AND2_X1 U3890 ( .A1(n4300), .A2(n4299), .ZN(n4865) );
  INV_X1 U3891 ( .A(n6269), .ZN(n5753) );
  OAI21_X2 U3892 ( .B1(n4754), .B2(n3664), .A(n3515), .ZN(n6223) );
  NAND2_X1 U3893 ( .A1(n4274), .A2(n4273), .ZN(n5166) );
  AND2_X1 U3894 ( .A1(n5765), .A2(n4237), .ZN(n6270) );
  AND2_X1 U3895 ( .A1(n3128), .A2(n4369), .ZN(n4642) );
  OAI21_X1 U3896 ( .B1(n3531), .B2(n3530), .A(n3529), .ZN(n3483) );
  XNOR2_X1 U3897 ( .A(n3427), .B(n3426), .ZN(n3509) );
  AND2_X1 U3898 ( .A1(n4195), .A2(n4194), .ZN(n4471) );
  OR2_X1 U3899 ( .A1(n3363), .A2(n3662), .ZN(n5352) );
  OR2_X1 U3901 ( .A1(n4754), .A2(n4769), .ZN(n6371) );
  OR2_X1 U3902 ( .A1(n6457), .A2(n6372), .ZN(n5015) );
  INV_X1 U3903 ( .A(n3740), .ZN(n6455) );
  NAND2_X1 U3904 ( .A1(n4792), .A2(n4754), .ZN(n6457) );
  OAI21_X1 U3905 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6693), .A(n6411), 
        .ZN(n6462) );
  NOR2_X1 U3906 ( .A1(n5787), .A2(n4751), .ZN(n5207) );
  OR3_X1 U3907 ( .A1(n6693), .A2(STATE2_REG_0__SCAN_IN), .A3(n4748), .ZN(n5075) );
  CLKBUF_X1 U3908 ( .A(n3752), .Z(n4472) );
  INV_X1 U3909 ( .A(n4559), .ZN(n4560) );
  NAND2_X1 U3910 ( .A1(n4541), .A2(n4559), .ZN(n6702) );
  INV_X1 U3911 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6950) );
  INV_X1 U3912 ( .A(n6105), .ZN(n6094) );
  INV_X1 U3913 ( .A(n3126), .ZN(n6140) );
  AND2_X1 U3914 ( .A1(n6096), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6142) );
  INV_X1 U3915 ( .A(n6155), .ZN(n6159) );
  INV_X1 U3916 ( .A(n6163), .ZN(n5529) );
  INV_X1 U3917 ( .A(n5924), .ZN(n6165) );
  NOR2_X2 U3918 ( .A1(n6167), .A2(n5367), .ZN(n6164) );
  NAND2_X1 U3919 ( .A1(n4663), .A2(n4662), .ZN(n5379) );
  NAND2_X1 U3920 ( .A1(n4661), .A2(n4681), .ZN(n4663) );
  OR2_X1 U3921 ( .A1(n4670), .A2(n4660), .ZN(n4661) );
  INV_X1 U3922 ( .A(n5547), .ZN(n5324) );
  AND2_X1 U3923 ( .A1(n4569), .A2(n4568), .ZN(n6185) );
  AND2_X1 U3924 ( .A1(n4567), .A2(n4673), .ZN(n4568) );
  XNOR2_X1 U3925 ( .A(n4478), .B(n5385), .ZN(n4527) );
  OR2_X1 U3926 ( .A1(n4477), .A2(n5554), .ZN(n4478) );
  OR2_X1 U3927 ( .A1(n4417), .A2(n4157), .ZN(n5848) );
  INV_X1 U3928 ( .A(n5969), .ZN(n6222) );
  NAND2_X1 U3929 ( .A1(n5568), .A2(n5567), .ZN(n5559) );
  AND2_X1 U3930 ( .A1(n5716), .A2(n5718), .ZN(n5707) );
  NAND2_X1 U3931 ( .A1(n3183), .A2(n3181), .ZN(n5587) );
  NAND2_X1 U3932 ( .A1(n3169), .A2(n3171), .ZN(n5651) );
  OR2_X1 U3933 ( .A1(n3636), .A2(n3173), .ZN(n3169) );
  NAND2_X1 U3934 ( .A1(n3636), .A2(n3209), .ZN(n3176) );
  NAND2_X1 U3935 ( .A1(n5079), .A2(n3634), .ZN(n5181) );
  INV_X1 U3936 ( .A(n6291), .ZN(n6311) );
  INV_X1 U3937 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6323) );
  OAI21_X1 U3938 ( .B1(n4958), .B2(n6691), .A(n4957), .ZN(n6322) );
  AND2_X2 U3939 ( .A1(n4921), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5361)
         );
  INV_X1 U3940 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5351) );
  INV_X1 U3941 ( .A(n6612), .ZN(n5362) );
  NOR2_X1 U3942 ( .A1(n3484), .A2(n6501), .ZN(n4953) );
  OR2_X1 U3943 ( .A1(n6020), .A2(n4685), .ZN(n6025) );
  INV_X1 U3944 ( .A(n5109), .ZN(n5091) );
  NOR2_X1 U3945 ( .A1(n4799), .A2(n4756), .ZN(n5109) );
  OR2_X1 U3946 ( .A1(n4904), .A2(n4903), .ZN(n6367) );
  INV_X1 U3947 ( .A(n6370), .ZN(n6353) );
  INV_X1 U3948 ( .A(n5100), .ZN(n6449) );
  AND2_X1 U3949 ( .A1(n5048), .A2(n5047), .ZN(n5106) );
  OR3_X1 U3950 ( .A1(n6457), .A2(n4756), .A3(n6455), .ZN(n6497) );
  NOR2_X1 U3951 ( .A1(n5075), .A2(n4779), .ZN(n6529) );
  NOR2_X1 U3952 ( .A1(n5075), .A2(n3268), .ZN(n6544) );
  INV_X1 U3953 ( .A(n6484), .ZN(n6553) );
  NOR2_X1 U3954 ( .A1(n5075), .A2(n4453), .ZN(n7041) );
  NOR2_X1 U3955 ( .A1(n4773), .A2(n4957), .ZN(n6528) );
  NOR2_X1 U3956 ( .A1(n4886), .A2(n4957), .ZN(n6535) );
  NOR2_X1 U3957 ( .A1(n4869), .A2(n4957), .ZN(n6543) );
  NOR2_X1 U3958 ( .A1(n4831), .A2(n4957), .ZN(n6550) );
  INV_X1 U3959 ( .A(n6528), .ZN(n5236) );
  INV_X1 U3960 ( .A(n6550), .ZN(n7044) );
  INV_X1 U3961 ( .A(n6572), .ZN(n5244) );
  NAND2_X1 U3962 ( .A1(n4758), .A2(n4756), .ZN(n6562) );
  AND2_X1 U3963 ( .A1(DATAI_2_), .A2(n6411), .ZN(n6522) );
  INV_X1 U3964 ( .A(n6529), .ZN(n5242) );
  AND2_X1 U3965 ( .A1(DATAI_5_), .A2(n6411), .ZN(n6570) );
  AND2_X1 U3966 ( .A1(n4758), .A2(n3745), .ZN(n6572) );
  INV_X1 U3967 ( .A(n7041), .ZN(n5216) );
  INV_X1 U3968 ( .A(n4822), .ZN(n6577) );
  NAND2_X1 U3969 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4692), .ZN(n6612) );
  INV_X1 U3970 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6693) );
  AOI21_X1 U3971 ( .B1(n4505), .B2(n6143), .A(n4504), .ZN(n4506) );
  NAND2_X1 U3972 ( .A1(n4503), .A2(n4502), .ZN(n4504) );
  INV_X1 U3973 ( .A(n5674), .ZN(n4505) );
  OAI22_X1 U3974 ( .A1(n4467), .A2(n6155), .B1(n5372), .B2(n6163), .ZN(n4468)
         );
  AOI21_X1 U3975 ( .B1(n5966), .B2(n4496), .A(n4188), .ZN(n4189) );
  INV_X1 U3976 ( .A(n4264), .ZN(n4386) );
  AOI21_X1 U3977 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5657), .A(n4396), 
        .ZN(n4397) );
  AND2_X2 U3978 ( .A1(n4952), .A2(n4951), .ZN(n3445) );
  AOI21_X1 U3979 ( .B1(n4749), .B2(n6611), .A(n3504), .ZN(n4755) );
  OR2_X2 U3980 ( .A1(n3266), .A2(n3265), .ZN(n3389) );
  OR2_X1 U3981 ( .A1(n5633), .A2(n5759), .ZN(n3135) );
  NAND2_X1 U3982 ( .A1(n3203), .A2(n4030), .ZN(n5414) );
  NAND2_X1 U3983 ( .A1(n5325), .A2(n3200), .ZN(n5445) );
  AND2_X1 U3984 ( .A1(n5493), .A2(n5562), .ZN(n3136) );
  AND2_X1 U3985 ( .A1(n5118), .A2(n3195), .ZN(n3137) );
  NAND2_X1 U3986 ( .A1(n3484), .A2(n3410), .ZN(n4751) );
  OAI211_X1 U3987 ( .C1(n5118), .C2(n3194), .A(n3152), .B(n3191), .ZN(n5298)
         );
  NAND2_X1 U3988 ( .A1(n3183), .A2(n3644), .ZN(n5616) );
  AND2_X1 U3989 ( .A1(n3629), .A2(n3628), .ZN(n3138) );
  AND2_X2 U3990 ( .A1(n4930), .A2(n3222), .ZN(n3335) );
  NAND2_X1 U3991 ( .A1(n3357), .A2(n3268), .ZN(n3363) );
  NOR2_X1 U3992 ( .A1(n5415), .A2(n3204), .ZN(n5511) );
  AND4_X1 U3993 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n3139)
         );
  AND2_X1 U3994 ( .A1(n3363), .A2(n3362), .ZN(n3140) );
  AND4_X1 U3995 ( .A1(n3244), .A2(n3243), .A3(n3242), .A4(n3241), .ZN(n3141)
         );
  OR2_X1 U3996 ( .A1(n3520), .A2(n3519), .ZN(n3142) );
  NAND2_X1 U3997 ( .A1(n3198), .A2(n4119), .ZN(n5394) );
  OR2_X1 U3998 ( .A1(n5537), .A2(n5955), .ZN(n3143) );
  XNOR2_X1 U3999 ( .A(n3532), .B(n3531), .ZN(n3740) );
  XNOR2_X1 U4000 ( .A(n3579), .B(n3587), .ZN(n3727) );
  AND2_X1 U4001 ( .A1(n5486), .A2(n6310), .ZN(n3144) );
  NAND2_X1 U4002 ( .A1(n3358), .A2(n4687), .ZN(n3145) );
  OR2_X1 U4003 ( .A1(n3511), .A2(n3492), .ZN(n3146) );
  AND2_X1 U4004 ( .A1(n3170), .A2(n5650), .ZN(n3147) );
  NAND2_X1 U4005 ( .A1(n5118), .A2(n5128), .ZN(n5127) );
  AND2_X1 U4006 ( .A1(n3188), .A2(n4259), .ZN(n3148) );
  AND2_X1 U4007 ( .A1(n5325), .A2(n5475), .ZN(n3149) );
  OAI21_X1 U4008 ( .B1(n5079), .B2(n3167), .A(n3165), .ZN(n5262) );
  NAND2_X1 U4009 ( .A1(n3176), .A2(n3638), .ZN(n5316) );
  AND2_X1 U4010 ( .A1(n5584), .A2(n3645), .ZN(n3150) );
  AND2_X1 U4011 ( .A1(n3148), .A2(n3189), .ZN(n3151) );
  OR2_X1 U4012 ( .A1(n3195), .A2(n3194), .ZN(n3152) );
  AND2_X1 U4013 ( .A1(n4139), .A2(n4119), .ZN(n3153) );
  AND3_X1 U4014 ( .A1(n3807), .A2(n3806), .A3(n3805), .ZN(n4863) );
  AND3_X1 U4015 ( .A1(n3875), .A2(n3874), .A3(n3873), .ZN(n5194) );
  NAND2_X1 U4016 ( .A1(n3643), .A2(n5641), .ZN(n5632) );
  INV_X1 U4017 ( .A(n3181), .ZN(n3180) );
  NOR2_X1 U4018 ( .A1(n3150), .A2(n3182), .ZN(n3181) );
  NOR2_X1 U4019 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3752) );
  NAND2_X1 U4020 ( .A1(n4742), .A2(n4827), .ZN(n4860) );
  AND2_X1 U4021 ( .A1(n5584), .A2(n5779), .ZN(n3154) );
  AND2_X1 U4022 ( .A1(n3975), .A2(n3974), .ZN(n3155) );
  INV_X1 U4023 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6611) );
  INV_X1 U4024 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4921) );
  INV_X1 U4025 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n3189) );
  NOR2_X4 U4026 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4952) );
  NOR2_X4 U4027 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4028 ( .A1(n3156), .A2(n3360), .ZN(n3361) );
  NAND2_X1 U4029 ( .A1(n4547), .A2(n3156), .ZN(n3390) );
  NAND2_X1 U4030 ( .A1(n3157), .A2(n3507), .ZN(n3543) );
  XNOR2_X2 U4031 ( .A(n4769), .B(n3545), .ZN(n4792) );
  NAND2_X1 U4032 ( .A1(n3402), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4033 ( .A1(n3160), .A2(n3354), .ZN(n3159) );
  NAND4_X1 U4034 ( .A1(n3358), .A2(n3364), .A3(n4687), .A4(n3378), .ZN(n3161)
         );
  NAND2_X1 U4035 ( .A1(n5079), .A2(n3165), .ZN(n3164) );
  XNOR2_X2 U4036 ( .A(n3484), .B(n4771), .ZN(n4749) );
  NAND2_X1 U4037 ( .A1(n3168), .A2(n3147), .ZN(n3640) );
  NAND2_X1 U4038 ( .A1(n3636), .A2(n3171), .ZN(n3168) );
  INV_X1 U4039 ( .A(n5632), .ZN(n3184) );
  NAND2_X1 U4040 ( .A1(n5632), .A2(n3181), .ZN(n3177) );
  NAND2_X1 U4041 ( .A1(n4193), .A2(n4192), .ZN(n3190) );
  NAND2_X1 U4042 ( .A1(n5118), .A2(n3192), .ZN(n3191) );
  NOR2_X1 U4043 ( .A1(n3193), .A2(n3891), .ZN(n3192) );
  NAND2_X1 U4044 ( .A1(n3197), .A2(n3146), .ZN(n3427) );
  NAND3_X1 U4045 ( .A1(n3484), .A2(n3410), .A3(n6611), .ZN(n3197) );
  NAND2_X1 U4046 ( .A1(n5325), .A2(n3199), .ZN(n5428) );
  AND3_X2 U4047 ( .A1(n4742), .A2(n3206), .A3(n4827), .ZN(n4981) );
  NAND3_X1 U4048 ( .A1(n4742), .A2(n4827), .A3(n3808), .ZN(n4861) );
  AND2_X2 U4049 ( .A1(n5561), .A2(n4180), .ZN(n4519) );
  INV_X1 U4050 ( .A(n5534), .ZN(n4513) );
  NAND2_X1 U4051 ( .A1(n3772), .A2(n3771), .ZN(n4717) );
  NAND2_X1 U4052 ( .A1(n3590), .A2(n3589), .ZN(n3606) );
  AOI21_X1 U4053 ( .B1(n3402), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3398), 
        .ZN(n3399) );
  INV_X1 U4054 ( .A(n3660), .ZN(n3661) );
  AND2_X2 U4055 ( .A1(n3222), .A2(n4934), .ZN(n3270) );
  NOR2_X1 U4056 ( .A1(n4900), .A2(n4792), .ZN(n3208) );
  NAND2_X1 U4057 ( .A1(n6593), .A2(n4567), .ZN(n6034) );
  INV_X1 U4058 ( .A(n6034), .ZN(n4529) );
  NAND2_X1 U4059 ( .A1(n5584), .A2(n6970), .ZN(n3209) );
  INV_X1 U4060 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6024) );
  AND2_X1 U4061 ( .A1(n3216), .A2(n4510), .ZN(n3211) );
  INV_X1 U4062 ( .A(n6143), .ZN(n6115) );
  NOR2_X2 U4063 ( .A1(n5152), .A2(n4486), .ZN(n6143) );
  INV_X1 U4064 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3923) );
  AND4_X1 U4065 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3212)
         );
  INV_X1 U4066 ( .A(n4269), .ZN(n4457) );
  AND3_X1 U4067 ( .A1(n3279), .A2(n3278), .A3(n3277), .ZN(n3214) );
  AND3_X1 U4068 ( .A1(n3262), .A2(n3261), .A3(n3260), .ZN(n3215) );
  INV_X1 U4069 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3768) );
  INV_X1 U4070 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5022) );
  INV_X1 U4071 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6465) );
  OR2_X1 U4072 ( .A1(n6231), .A2(n4535), .ZN(n3216) );
  AND2_X1 U4073 ( .A1(n3693), .A2(n3692), .ZN(n3695) );
  AND2_X1 U4074 ( .A1(n6978), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3682)
         );
  NOR2_X1 U4075 ( .A1(n3377), .A2(n3145), .ZN(n3381) );
  INV_X1 U4076 ( .A(n3534), .ZN(n3479) );
  OR2_X1 U4077 ( .A1(n3502), .A2(n3501), .ZN(n3559) );
  AND2_X1 U4078 ( .A1(n3714), .A2(n3713), .ZN(n4203) );
  AND2_X1 U4079 ( .A1(n3588), .A2(n3587), .ZN(n3589) );
  NOR2_X1 U4080 ( .A1(n3422), .A2(n3421), .ZN(n3511) );
  OR2_X1 U4081 ( .A1(n3703), .A2(n4977), .ZN(n3456) );
  NAND2_X1 U4082 ( .A1(n3530), .A2(n3531), .ZN(n3482) );
  INV_X1 U4083 ( .A(n5446), .ZN(n3959) );
  INV_X1 U4084 ( .A(n4863), .ZN(n3808) );
  NOR2_X1 U4085 ( .A1(n3789), .A2(n4447), .ZN(n3790) );
  AND2_X1 U4086 ( .A1(n4717), .A2(n4718), .ZN(n3781) );
  INV_X1 U4087 ( .A(n4457), .ZN(n4369) );
  INV_X1 U4088 ( .A(n3518), .ZN(n3519) );
  INV_X1 U4089 ( .A(n3453), .ZN(n3454) );
  NAND2_X1 U4090 ( .A1(n3336), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3263) );
  OR2_X1 U4091 ( .A1(n5848), .A2(n4447), .ZN(n4158) );
  NAND2_X1 U4092 ( .A1(n4122), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3341)
         );
  OR2_X1 U4093 ( .A1(n4418), .A2(n4508), .ZN(n4477) );
  OR2_X1 U4094 ( .A1(n5950), .A2(n4447), .ZN(n4117) );
  INV_X1 U4095 ( .A(n5416), .ZN(n4030) );
  INV_X1 U4096 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5308) );
  INV_X1 U4097 ( .A(n3809), .ZN(n3810) );
  NOR2_X1 U4098 ( .A1(n3791), .A2(n3790), .ZN(n3792) );
  AND2_X1 U4099 ( .A1(n3370), .A2(n3369), .ZN(n4232) );
  AND2_X1 U4100 ( .A1(n3672), .A2(n3708), .ZN(n4200) );
  NOR2_X1 U4101 ( .A1(n6659), .A2(n5463), .ZN(n5462) );
  NAND2_X1 U4102 ( .A1(n3129), .A2(n3371), .ZN(n3367) );
  INV_X1 U4103 ( .A(n4444), .ZN(n4415) );
  NOR2_X1 U4104 ( .A1(n4155), .A2(n5571), .ZN(n4156) );
  NOR2_X1 U4105 ( .A1(n4074), .A2(n4073), .ZN(n4093) );
  AND2_X1 U4106 ( .A1(n3955), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3956)
         );
  NAND2_X1 U4107 ( .A1(n3810), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3811)
         );
  AND2_X1 U4108 ( .A1(n5584), .A2(n4323), .ZN(n5642) );
  NOR2_X1 U4109 ( .A1(n6371), .A2(n6372), .ZN(n4780) );
  AND2_X1 U4110 ( .A1(n3404), .A2(n6324), .ZN(n4837) );
  NAND2_X1 U4112 ( .A1(n4027), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4074)
         );
  INV_X1 U4113 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5436) );
  NOR2_X1 U4114 ( .A1(n6746), .A2(n3855), .ZN(n3876) );
  AND2_X1 U4115 ( .A1(n4527), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4491) );
  NAND2_X1 U4116 ( .A1(n6702), .A2(n4489), .ZN(n6098) );
  AND2_X1 U4117 ( .A1(n4293), .A2(n4292), .ZN(n6113) );
  AND2_X1 U4118 ( .A1(n4156), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4417)
         );
  AND2_X1 U4119 ( .A1(n4335), .A2(n4334), .ZN(n5449) );
  INV_X1 U4120 ( .A(n3138), .ZN(n5633) );
  NAND2_X1 U4121 ( .A1(n4385), .A2(n6580), .ZN(n5765) );
  OR2_X1 U4122 ( .A1(n4793), .A2(n4792), .ZN(n4799) );
  AND2_X1 U4123 ( .A1(n4839), .A2(n4838), .ZN(n5041) );
  INV_X1 U4124 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6325) );
  OR2_X1 U4125 ( .A1(n5015), .A2(n3745), .ZN(n5100) );
  INV_X1 U4126 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6584) );
  OR2_X1 U4127 ( .A1(n5489), .A2(n6115), .ZN(n4538) );
  NOR2_X1 U4128 ( .A1(n6798), .A2(n5448), .ZN(n5912) );
  INV_X1 U4129 ( .A(n6098), .ZN(n6121) );
  AND2_X1 U4130 ( .A1(n6096), .A2(n4491), .ZN(n6108) );
  INV_X1 U4131 ( .A(n5531), .ZN(n6160) );
  INV_X1 U4132 ( .A(n5379), .ZN(n6167) );
  OAI21_X1 U4133 ( .B1(n5383), .B2(n6704), .A(n4560), .ZN(n4592) );
  INV_X1 U4134 ( .A(n4662), .ZN(n4637) );
  NAND2_X1 U4135 ( .A1(n3977), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4025)
         );
  NAND2_X1 U4136 ( .A1(n3787), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3809)
         );
  INV_X1 U4137 ( .A(n6231), .ZN(n5966) );
  AND2_X1 U4138 ( .A1(n4692), .A2(n4681), .ZN(n4567) );
  AND2_X1 U4139 ( .A1(n5707), .A2(n4256), .ZN(n5975) );
  AOI21_X2 U4140 ( .B1(n5584), .B2(n6778), .A(n5602), .ZN(n5596) );
  NOR2_X1 U4141 ( .A1(n4323), .A2(n6019), .ZN(n6004) );
  AND2_X1 U4142 ( .A1(n4385), .A2(n4221), .ZN(n6315) );
  AND2_X1 U4143 ( .A1(n4471), .A2(n4557), .ZN(n6580) );
  NOR2_X1 U4144 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6022) );
  OAI21_X1 U4145 ( .B1(n6456), .B2(n4778), .A(n4777), .ZN(n7034) );
  INV_X1 U4146 ( .A(n7036), .ZN(n5043) );
  INV_X1 U4147 ( .A(n6444), .ZN(n6416) );
  INV_X1 U4148 ( .A(n6455), .ZN(n6372) );
  INV_X1 U4149 ( .A(n6415), .ZN(n6447) );
  NOR2_X1 U4150 ( .A1(n4784), .A2(n4957), .ZN(n6514) );
  AND2_X1 U4151 ( .A1(n4997), .A2(n3745), .ZN(n6554) );
  OAI211_X1 U4152 ( .C1(n5205), .C2(n6693), .A(n5204), .B(n5203), .ZN(n5243)
         );
  AND2_X1 U4153 ( .A1(n5351), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3726) );
  INV_X1 U4154 ( .A(n6702), .ZN(n5152) );
  AND2_X1 U4155 ( .A1(n4538), .A2(n4537), .ZN(n4539) );
  INV_X1 U4156 ( .A(n6142), .ZN(n6117) );
  NAND2_X1 U4157 ( .A1(n6096), .A2(n4479), .ZN(n6105) );
  INV_X1 U4158 ( .A(n4468), .ZN(n4469) );
  NAND2_X1 U4159 ( .A1(n6163), .A2(n4453), .ZN(n6155) );
  INV_X1 U4160 ( .A(n6185), .ZN(n6197) );
  NAND2_X1 U4161 ( .A1(n6034), .A2(n4182), .ZN(n5969) );
  OR2_X1 U4162 ( .A1(n6624), .A2(n6499), .ZN(n5955) );
  NAND2_X1 U4163 ( .A1(n5969), .A2(n4185), .ZN(n6231) );
  INV_X1 U4164 ( .A(n6310), .ZN(n6233) );
  INV_X1 U4165 ( .A(n6315), .ZN(n5992) );
  INV_X1 U4166 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6978) );
  NOR2_X1 U4167 ( .A1(n4850), .A2(n4849), .ZN(n5098) );
  INV_X1 U4168 ( .A(n5833), .ZN(n5846) );
  NAND2_X1 U4169 ( .A1(n3208), .A2(n3745), .ZN(n6359) );
  NAND2_X1 U4170 ( .A1(n3208), .A2(n4756), .ZN(n6370) );
  INV_X1 U4171 ( .A(n4772), .ZN(n7045) );
  NAND2_X1 U4172 ( .A1(n4833), .A2(n6372), .ZN(n6406) );
  NAND2_X1 U4173 ( .A1(n6373), .A2(n6372), .ZN(n6444) );
  OR2_X1 U4174 ( .A1(n5015), .A2(n4756), .ZN(n6415) );
  INV_X1 U4175 ( .A(n6514), .ZN(n5222) );
  INV_X1 U4176 ( .A(n6543), .ZN(n5217) );
  OR3_X1 U4177 ( .A1(n6457), .A2(n6455), .A3(n3745), .ZN(n6484) );
  NOR2_X1 U4178 ( .A1(n6507), .A2(n6506), .ZN(n6559) );
  INV_X1 U4179 ( .A(n6515), .ZN(n5226) );
  INV_X1 U4180 ( .A(n6544), .ZN(n5221) );
  INV_X1 U4181 ( .A(n6521), .ZN(n5250) );
  NAND2_X1 U4182 ( .A1(n3726), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6617) );
  INV_X1 U4183 ( .A(n6678), .ZN(n6684) );
  OAI21_X1 U4184 ( .B1(n5537), .B2(n6105), .A(n4506), .ZN(U2799) );
  OAI21_X1 U4185 ( .B1(n5378), .B2(n5531), .A(n4469), .ZN(U2829) );
  OAI211_X1 U4186 ( .C1(n5678), .C2(n6034), .A(n3143), .B(n4189), .ZN(U2958)
         );
  OAI21_X1 U4187 ( .B1(n4515), .B2(n5992), .A(n4397), .ZN(U2989) );
  INV_X1 U4188 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4189 ( .A1(n3270), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3221) );
  INV_X1 U4190 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4929) );
  AND2_X2 U4191 ( .A1(n5361), .A2(n4930), .ZN(n3287) );
  AOI22_X1 U4192 ( .A1(n3286), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3220) );
  AOI22_X1 U4193 ( .A1(n3272), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3219) );
  AOI22_X1 U4194 ( .A1(n3411), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3218) );
  AOI22_X1 U4195 ( .A1(n3335), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4196 ( .A1(n3318), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4197 ( .A1(n3998), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3225) );
  AND2_X4 U4198 ( .A1(n3223), .A2(n4917), .ZN(n3416) );
  AOI22_X1 U4199 ( .A1(n3470), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4200 ( .A1(n3286), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4201 ( .A1(n3272), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4202 ( .A1(n3270), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4203 ( .A1(n3411), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4204 ( .A1(n3998), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3235) );
  AOI22_X1 U4205 ( .A1(n3130), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3234) );
  AOI22_X1 U4206 ( .A1(n3318), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4207 ( .A1(n3335), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3232) );
  NAND2_X2 U4208 ( .A1(n3213), .A2(n3236), .ZN(n3357) );
  NAND2_X1 U4209 ( .A1(n3998), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4210 ( .A1(n3335), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3239) );
  NAND2_X1 U4211 ( .A1(n3131), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4212 ( .A1(n3416), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U4213 ( .A1(n3272), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3244)
         );
  NAND2_X1 U4214 ( .A1(n3318), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3243)
         );
  NAND2_X1 U4215 ( .A1(n3445), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3242)
         );
  NAND2_X1 U4216 ( .A1(n3336), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4217 ( .A1(n3411), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3248)
         );
  NAND2_X1 U4218 ( .A1(n3286), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U4219 ( .A1(n3287), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4220 ( .A1(n4122), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3245)
         );
  NAND2_X1 U4221 ( .A1(n3270), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3252)
         );
  NAND2_X1 U4222 ( .A1(n3269), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3251) );
  NAND2_X1 U4223 ( .A1(n3345), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4224 ( .A1(n3271), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U4225 ( .A1(n3270), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3259) );
  AOI22_X1 U4226 ( .A1(n3286), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3258) );
  AOI22_X1 U4227 ( .A1(n3272), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4228 ( .A1(n3411), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3256) );
  NAND4_X1 U4229 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3266)
         );
  AOI22_X1 U4230 ( .A1(n3998), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3262) );
  AOI22_X1 U4231 ( .A1(n3318), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4232 ( .A1(n3470), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3264) );
  NAND3_X1 U4233 ( .A1(n3215), .A2(n3264), .A3(n3263), .ZN(n3265) );
  AOI22_X1 U4234 ( .A1(n3270), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3269), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4235 ( .A1(n3286), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4236 ( .A1(n3272), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4237 ( .A1(n3411), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4238 ( .A1(n3335), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4239 ( .A1(n3998), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3279) );
  AOI22_X1 U4240 ( .A1(n3470), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4241 ( .A1(n3318), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3445), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3277) );
  NAND3_X1 U4242 ( .A1(n3281), .A2(n3280), .A3(n3214), .ZN(n3362) );
  INV_X2 U4243 ( .A(n3362), .ZN(n3423) );
  NAND2_X1 U4244 ( .A1(n3318), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4245 ( .A1(n3335), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3284) );
  NAND2_X1 U4246 ( .A1(n3445), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3283)
         );
  NAND2_X1 U4247 ( .A1(n3336), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4248 ( .A1(n3286), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4249 ( .A1(n3270), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3290)
         );
  NAND2_X1 U4250 ( .A1(n3287), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4251 ( .A1(n3271), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3288) );
  NAND2_X1 U4252 ( .A1(n3998), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3295) );
  NAND2_X1 U4253 ( .A1(n3345), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3294) );
  NAND2_X1 U4254 ( .A1(n3470), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3293) );
  NAND2_X1 U4255 ( .A1(n3416), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3292) );
  NAND2_X1 U4256 ( .A1(n3269), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3299) );
  NAND2_X1 U4257 ( .A1(n3272), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3298)
         );
  NAND2_X1 U4258 ( .A1(n3411), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3297)
         );
  NAND2_X1 U4259 ( .A1(n4122), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3296)
         );
  INV_X1 U4260 ( .A(n4747), .ZN(n4669) );
  NAND2_X1 U4261 ( .A1(n3355), .A2(n4669), .ZN(n3304) );
  NAND2_X1 U4262 ( .A1(n3355), .A2(n3268), .ZN(n3309) );
  NAND2_X1 U4263 ( .A1(n4455), .A2(n4747), .ZN(n3307) );
  NAND2_X1 U4264 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  NAND2_X1 U4265 ( .A1(n3384), .A2(n3383), .ZN(n3354) );
  NAND2_X1 U4266 ( .A1(n3411), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3313)
         );
  NAND2_X1 U4267 ( .A1(n3269), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3312) );
  NAND2_X1 U4268 ( .A1(n4122), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4269 ( .A1(n3270), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3310)
         );
  NAND2_X1 U4270 ( .A1(n3287), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3317) );
  NAND2_X1 U4271 ( .A1(n3286), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3316) );
  NAND2_X1 U4272 ( .A1(n3272), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3315)
         );
  NAND2_X1 U4273 ( .A1(n3271), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4274 ( .A1(n3998), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4275 ( .A1(n3345), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4276 ( .A1(n3318), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3320)
         );
  NAND2_X1 U4277 ( .A1(n3445), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3319)
         );
  NAND2_X1 U4278 ( .A1(n3335), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U4279 ( .A1(n3470), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U4280 ( .A1(n3336), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4281 ( .A1(n3416), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4282 ( .A1(n3269), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3334) );
  NAND2_X1 U4283 ( .A1(n3270), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3333)
         );
  NAND2_X1 U4284 ( .A1(n3286), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4285 ( .A1(n3411), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3331)
         );
  NAND2_X1 U4286 ( .A1(n3318), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3340)
         );
  NAND2_X1 U4287 ( .A1(n3998), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3339) );
  NAND2_X1 U4288 ( .A1(n3335), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3338) );
  NAND2_X1 U4289 ( .A1(n3336), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4290 ( .A1(n3287), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4291 ( .A1(n3272), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3343)
         );
  NAND2_X1 U4292 ( .A1(n3271), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4293 ( .A1(n3345), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4294 ( .A1(n3131), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3348) );
  NAND2_X1 U4295 ( .A1(n3445), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3347)
         );
  NAND2_X1 U4296 ( .A1(n3416), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3346) );
  NAND4_X4 U4297 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n4217)
         );
  INV_X1 U4298 ( .A(n3355), .ZN(n3356) );
  NAND2_X1 U4299 ( .A1(n3382), .A2(n5383), .ZN(n3358) );
  NAND2_X1 U4300 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6636) );
  OAI21_X1 U4301 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6636), .ZN(n4199) );
  NAND2_X1 U4302 ( .A1(n6022), .A2(n6611), .ZN(n4186) );
  MUX2_X1 U4303 ( .A(n3726), .B(n4186), .S(n6978), .Z(n3365) );
  NAND2_X1 U4304 ( .A1(n3366), .A2(n3365), .ZN(n3430) );
  INV_X1 U4305 ( .A(n3690), .ZN(n3368) );
  INV_X1 U4306 ( .A(n3367), .ZN(n4544) );
  NAND2_X1 U4307 ( .A1(n3368), .A2(n4544), .ZN(n3369) );
  NAND2_X1 U4308 ( .A1(n4223), .A2(n3363), .ZN(n3372) );
  BUF_X4 U4309 ( .A(n3371), .Z(n4557) );
  NAND2_X1 U4310 ( .A1(n4747), .A2(n4557), .ZN(n4456) );
  NAND3_X1 U4311 ( .A1(n3372), .A2(n4217), .A3(n4456), .ZN(n3376) );
  NAND2_X1 U4312 ( .A1(n6022), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6618) );
  INV_X1 U4313 ( .A(n6618), .ZN(n3375) );
  NAND2_X1 U4314 ( .A1(n3362), .A2(n3389), .ZN(n3662) );
  INV_X1 U4315 ( .A(n3662), .ZN(n3374) );
  NAND4_X1 U4316 ( .A1(n3374), .A2(n4747), .A3(n3268), .A4(n4779), .ZN(n4939)
         );
  NAND3_X1 U4317 ( .A1(n3376), .A2(n3375), .A3(n4939), .ZN(n3377) );
  INV_X1 U4318 ( .A(n3378), .ZN(n3379) );
  OAI21_X1 U4319 ( .B1(n3379), .B2(n4779), .A(n4557), .ZN(n3380) );
  NAND3_X1 U4320 ( .A1(n4232), .A2(n3381), .A3(n3380), .ZN(n3428) );
  NAND2_X1 U4321 ( .A1(n3430), .A2(n3428), .ZN(n3461) );
  AND2_X1 U4322 ( .A1(n3690), .A2(n3129), .ZN(n4194) );
  AND2_X1 U4323 ( .A1(n3385), .A2(n4194), .ZN(n3386) );
  NOR2_X1 U4324 ( .A1(n3357), .A2(n3373), .ZN(n3387) );
  NAND3_X1 U4325 ( .A1(n3388), .A2(n4747), .A3(n3387), .ZN(n4688) );
  NAND2_X1 U4326 ( .A1(n3306), .A2(n3389), .ZN(n5367) );
  NAND3_X1 U4327 ( .A1(n3390), .A2(n4219), .A3(n4383), .ZN(n3391) );
  NAND2_X1 U4328 ( .A1(n3391), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3400) );
  INV_X1 U4329 ( .A(n3400), .ZN(n3397) );
  INV_X1 U4330 ( .A(n4186), .ZN(n3392) );
  XNOR2_X1 U4331 ( .A(n6584), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6410)
         );
  NAND2_X1 U4332 ( .A1(n3392), .A2(n6410), .ZN(n3395) );
  INV_X1 U4333 ( .A(n3726), .ZN(n3393) );
  NAND2_X1 U4334 ( .A1(n3393), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4335 ( .A1(n3395), .A2(n3394), .ZN(n3398) );
  OR2_X1 U4336 ( .A1(n3398), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3396)
         );
  NAND2_X1 U4337 ( .A1(n3397), .A2(n3396), .ZN(n3463) );
  NAND2_X1 U4338 ( .A1(n3461), .A2(n3463), .ZN(n3401) );
  NAND2_X1 U4339 ( .A1(n3400), .A2(n3399), .ZN(n3462) );
  NAND2_X1 U4340 ( .A1(n3401), .A2(n3462), .ZN(n3409) );
  INV_X1 U4341 ( .A(n3409), .ZN(n3407) );
  NAND2_X1 U4342 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3403) );
  NAND2_X1 U4343 ( .A1(n3403), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3404) );
  NOR2_X1 U4344 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6584), .ZN(n5800)
         );
  NAND2_X1 U4345 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5800), .ZN(n6324) );
  OAI22_X1 U4346 ( .A1(n4186), .A2(n4837), .B1(n3726), .B2(n6589), .ZN(n3405)
         );
  INV_X1 U4347 ( .A(n3408), .ZN(n3406) );
  NAND2_X1 U4348 ( .A1(n3409), .A2(n3408), .ZN(n3410) );
  AOI22_X1 U4349 ( .A1(n4014), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4350 ( .A1(n4425), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4351 ( .A1(n4424), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4352 ( .A1(n4031), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3412) );
  NAND4_X1 U4353 ( .A1(n3415), .A2(n3414), .A3(n3413), .A4(n3412), .ZN(n3422)
         );
  AOI22_X1 U4354 ( .A1(n4432), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4355 ( .A1(n4166), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4356 ( .A1(n4435), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4357 ( .A1(n3130), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3417) );
  NAND4_X1 U4358 ( .A1(n3420), .A2(n3419), .A3(n3418), .A4(n3417), .ZN(n3421)
         );
  INV_X1 U4359 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n6787) );
  OAI22_X1 U4360 ( .A1(n3703), .A2(n6787), .B1(n3491), .B2(n3511), .ZN(n3425)
         );
  INV_X1 U4361 ( .A(n3425), .ZN(n3426) );
  INV_X1 U4362 ( .A(n3428), .ZN(n3429) );
  XNOR2_X1 U4363 ( .A(n3430), .B(n3429), .ZN(n3746) );
  NAND2_X1 U4364 ( .A1(n3746), .A2(n6611), .ZN(n3516) );
  AOI22_X1 U4365 ( .A1(n4425), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4366 ( .A1(n3272), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3433) );
  AOI22_X1 U4367 ( .A1(n4432), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3432) );
  AOI22_X1 U4368 ( .A1(n3335), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3431) );
  NAND4_X1 U4369 ( .A1(n3434), .A2(n3433), .A3(n3432), .A4(n3431), .ZN(n3440)
         );
  AOI22_X1 U4370 ( .A1(n4031), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4371 ( .A1(n4937), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4372 ( .A1(n3130), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4373 ( .A1(n4014), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3435) );
  NAND4_X1 U4374 ( .A1(n3438), .A2(n3437), .A3(n3436), .A4(n3435), .ZN(n3439)
         );
  NAND2_X1 U4375 ( .A1(n3423), .A2(n3621), .ZN(n3459) );
  INV_X1 U4376 ( .A(n3621), .ZN(n3630) );
  NAND2_X1 U4377 ( .A1(n3630), .A2(n3423), .ZN(n3452) );
  AOI22_X1 U4378 ( .A1(n4014), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4379 ( .A1(n4425), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4432), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4380 ( .A1(n4435), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3130), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4381 ( .A1(n4031), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3441) );
  NAND4_X1 U4382 ( .A1(n3444), .A2(n3443), .A3(n3442), .A4(n3441), .ZN(n3451)
         );
  AOI22_X1 U4383 ( .A1(n3287), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4384 ( .A1(n4403), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4385 ( .A1(n4166), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4386 ( .A1(n3336), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3446) );
  NAND4_X1 U4387 ( .A1(n3449), .A2(n3448), .A3(n3447), .A4(n3446), .ZN(n3450)
         );
  MUX2_X1 U4388 ( .A(n3459), .B(n3452), .S(n3533), .Z(n3453) );
  NAND2_X1 U4389 ( .A1(n3454), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4390 ( .A1(n3516), .A2(n3520), .ZN(n3458) );
  AOI21_X1 U4391 ( .B1(n3129), .B2(n3533), .A(n6611), .ZN(n3455) );
  AND2_X1 U4392 ( .A1(n3455), .A2(n3459), .ZN(n3457) );
  INV_X1 U4393 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U4394 ( .A1(n3458), .A2(n3518), .ZN(n3460) );
  INV_X1 U4395 ( .A(n3461), .ZN(n3465) );
  NAND2_X1 U4396 ( .A1(n3463), .A2(n3462), .ZN(n3464) );
  NAND2_X1 U4397 ( .A1(n4750), .A2(n6611), .ZN(n3478) );
  AOI22_X1 U4398 ( .A1(n4014), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4399 ( .A1(n4425), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4400 ( .A1(n4403), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4401 ( .A1(n4432), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4402 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3476)
         );
  AOI22_X1 U4403 ( .A1(n4424), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4404 ( .A1(n4435), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3470), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4405 ( .A1(n4031), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4406 ( .A1(n4127), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3471) );
  NAND4_X1 U4407 ( .A1(n3474), .A2(n3473), .A3(n3472), .A4(n3471), .ZN(n3475)
         );
  OR2_X1 U4408 ( .A1(n3492), .A2(n3479), .ZN(n3477) );
  INV_X1 U4409 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n6968) );
  OR2_X1 U4410 ( .A1(n3491), .A2(n3479), .ZN(n3481) );
  OR2_X1 U4411 ( .A1(n3492), .A2(n3621), .ZN(n3480) );
  OAI211_X1 U4412 ( .C1(n3703), .C2(n6968), .A(n3481), .B(n3480), .ZN(n3529)
         );
  NAND2_X1 U4413 ( .A1(n3483), .A2(n3482), .ZN(n3508) );
  NAND2_X1 U4414 ( .A1(n3402), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3490) );
  NAND3_X1 U4415 ( .A1(n6325), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6381) );
  INV_X1 U4416 ( .A(n6381), .ZN(n3486) );
  NAND2_X1 U4417 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3486), .ZN(n6377) );
  NAND2_X1 U4418 ( .A1(n6325), .A2(n6377), .ZN(n3487) );
  NAND3_X1 U4419 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5199) );
  INV_X1 U4420 ( .A(n5199), .ZN(n4762) );
  NAND2_X1 U4421 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4762), .ZN(n5146) );
  NAND2_X1 U4422 ( .A1(n3487), .A2(n5146), .ZN(n6409) );
  OAI22_X1 U4423 ( .A1(n4186), .A2(n6409), .B1(n3726), .B2(n6325), .ZN(n3488)
         );
  INV_X1 U4424 ( .A(n3488), .ZN(n3489) );
  AOI22_X1 U4425 ( .A1(n4014), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4426 ( .A1(n4425), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4427 ( .A1(n4424), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4428 ( .A1(n4031), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3493) );
  NAND4_X1 U4429 ( .A1(n3496), .A2(n3495), .A3(n3494), .A4(n3493), .ZN(n3502)
         );
  AOI22_X1 U4430 ( .A1(n4432), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U4431 ( .A1(n4166), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4432 ( .A1(n4435), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4433 ( .A1(n4426), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3497) );
  NAND4_X1 U4434 ( .A1(n3500), .A2(n3499), .A3(n3498), .A4(n3497), .ZN(n3501)
         );
  AOI22_X1 U4435 ( .A1(n3715), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3722), 
        .B2(n3559), .ZN(n3503) );
  INV_X1 U4436 ( .A(n3664), .ZN(n4196) );
  NAND2_X1 U4437 ( .A1(n3534), .A2(n3533), .ZN(n3512) );
  NAND2_X1 U4438 ( .A1(n3512), .A2(n3511), .ZN(n3560) );
  INV_X1 U4439 ( .A(n3559), .ZN(n3505) );
  XNOR2_X1 U4440 ( .A(n3560), .B(n3505), .ZN(n3506) );
  NAND2_X1 U4441 ( .A1(n3506), .A2(n5383), .ZN(n3507) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4280) );
  XNOR2_X1 U4443 ( .A(n3543), .B(n4280), .ZN(n6214) );
  NAND2_X2 U4444 ( .A1(n3545), .A2(n3510), .ZN(n4754) );
  XNOR2_X1 U4445 ( .A(n3512), .B(n3511), .ZN(n3514) );
  NAND2_X1 U4446 ( .A1(n3129), .A2(n3373), .ZN(n3522) );
  INV_X1 U4447 ( .A(n3522), .ZN(n3513) );
  AOI21_X1 U4448 ( .B1(n3514), .B2(n5383), .A(n3513), .ZN(n3515) );
  NAND2_X1 U4449 ( .A1(n6223), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3542)
         );
  NAND2_X1 U4450 ( .A1(n3516), .A2(n3518), .ZN(n3517) );
  NAND2_X1 U4451 ( .A1(n3517), .A2(n3520), .ZN(n3521) );
  NAND2_X1 U4452 ( .A1(n4756), .A2(n4196), .ZN(n3525) );
  INV_X1 U4453 ( .A(n5383), .ZN(n6706) );
  OAI21_X1 U4454 ( .B1(n6706), .B2(n3533), .A(n3522), .ZN(n3523) );
  INV_X1 U4455 ( .A(n3523), .ZN(n3524) );
  NAND2_X1 U4456 ( .A1(n3525), .A2(n3524), .ZN(n4583) );
  NAND2_X1 U4457 ( .A1(n4583), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3526)
         );
  INV_X1 U4458 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U4459 ( .A1(n3526), .A2(n6313), .ZN(n3528) );
  AND2_X1 U4460 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U4461 ( .A1(n4583), .A2(n3527), .ZN(n3539) );
  NAND2_X1 U4462 ( .A1(n3740), .A2(n4196), .ZN(n3538) );
  XNOR2_X1 U4463 ( .A(n3534), .B(n3533), .ZN(n3535) );
  OAI211_X1 U4464 ( .C1(n3535), .C2(n6706), .A(n4223), .B(n3357), .ZN(n3536)
         );
  INV_X1 U4465 ( .A(n3536), .ZN(n3537) );
  NAND2_X1 U4466 ( .A1(n3538), .A2(n3537), .ZN(n4698) );
  INV_X1 U4467 ( .A(n3539), .ZN(n3540) );
  NOR2_X1 U4468 ( .A1(n6223), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3541)
         );
  NAND2_X1 U4469 ( .A1(n6214), .A2(n6215), .ZN(n6216) );
  NAND2_X1 U4470 ( .A1(n3543), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3544)
         );
  NAND2_X1 U4471 ( .A1(n6216), .A2(n3544), .ZN(n4726) );
  INV_X1 U4472 ( .A(n4755), .ZN(n4769) );
  AOI22_X1 U4473 ( .A1(n3133), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4474 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4424), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4475 ( .A1(n4403), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3548) );
  AOI22_X1 U4476 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4426), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3547) );
  NAND4_X1 U4477 ( .A1(n3550), .A2(n3549), .A3(n3548), .A4(n3547), .ZN(n3556)
         );
  AOI22_X1 U4478 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4425), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4479 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4435), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4480 ( .A1(n4432), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3552) );
  AOI22_X1 U4481 ( .A1(n4014), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3551) );
  NAND4_X1 U4482 ( .A1(n3554), .A2(n3553), .A3(n3552), .A4(n3551), .ZN(n3555)
         );
  NAND2_X1 U4483 ( .A1(n3722), .A2(n3608), .ZN(n3558) );
  INV_X1 U4484 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4969) );
  OR2_X1 U4485 ( .A1(n3703), .A2(n4969), .ZN(n3557) );
  NAND2_X1 U4486 ( .A1(n3763), .A2(n4196), .ZN(n3563) );
  NAND2_X1 U4487 ( .A1(n3560), .A2(n3559), .ZN(n3610) );
  XNOR2_X1 U4488 ( .A(n3610), .B(n3608), .ZN(n3561) );
  NAND2_X1 U4489 ( .A1(n3561), .A2(n5383), .ZN(n3562) );
  NAND2_X1 U4490 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  INV_X1 U4491 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4287) );
  XNOR2_X1 U4492 ( .A(n3564), .B(n4287), .ZN(n4724) );
  NAND2_X1 U4493 ( .A1(n4726), .A2(n4724), .ZN(n4725) );
  NAND2_X1 U4494 ( .A1(n3564), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3565)
         );
  NAND2_X1 U4495 ( .A1(n4725), .A2(n3565), .ZN(n6207) );
  NAND2_X1 U4496 ( .A1(n3590), .A2(n3588), .ZN(n3579) );
  AOI22_X1 U4497 ( .A1(n4014), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3570) );
  INV_X1 U4498 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6831) );
  AOI22_X1 U4499 ( .A1(n4425), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4500 ( .A1(n4424), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4501 ( .A1(n4031), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3567) );
  NAND4_X1 U4502 ( .A1(n3570), .A2(n3569), .A3(n3568), .A4(n3567), .ZN(n3576)
         );
  AOI22_X1 U4503 ( .A1(n4432), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4504 ( .A1(n4166), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3573) );
  AOI22_X1 U4505 ( .A1(n4435), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3572) );
  AOI22_X1 U4506 ( .A1(n4426), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3571) );
  NAND4_X1 U4507 ( .A1(n3574), .A2(n3573), .A3(n3572), .A4(n3571), .ZN(n3575)
         );
  NAND2_X1 U4508 ( .A1(n3722), .A2(n3607), .ZN(n3578) );
  INV_X1 U4509 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5097) );
  OR2_X1 U4510 ( .A1(n3703), .A2(n5097), .ZN(n3577) );
  NAND2_X1 U4511 ( .A1(n3578), .A2(n3577), .ZN(n3587) );
  NAND2_X1 U4512 ( .A1(n3727), .A2(n4196), .ZN(n3584) );
  INV_X1 U4513 ( .A(n3608), .ZN(n3580) );
  OR2_X1 U4514 ( .A1(n3610), .A2(n3580), .ZN(n3581) );
  XNOR2_X1 U4515 ( .A(n3581), .B(n3607), .ZN(n3582) );
  NAND2_X1 U4516 ( .A1(n3582), .A2(n5383), .ZN(n3583) );
  NAND2_X1 U4517 ( .A1(n3584), .A2(n3583), .ZN(n3585) );
  INV_X1 U4518 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6283) );
  XNOR2_X1 U4519 ( .A(n3585), .B(n6283), .ZN(n6206) );
  NAND2_X1 U4520 ( .A1(n6207), .A2(n6206), .ZN(n6209) );
  NAND2_X1 U4521 ( .A1(n3585), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3586)
         );
  NAND2_X1 U4522 ( .A1(n6209), .A2(n3586), .ZN(n4813) );
  INV_X1 U4523 ( .A(n3606), .ZN(n3604) );
  NAND2_X1 U4524 ( .A1(n3715), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4525 ( .A1(n4014), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4526 ( .A1(n4425), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4527 ( .A1(n4424), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3592) );
  AOI22_X1 U4528 ( .A1(n4031), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3591) );
  NAND4_X1 U4529 ( .A1(n3594), .A2(n3593), .A3(n3592), .A4(n3591), .ZN(n3600)
         );
  AOI22_X1 U4530 ( .A1(n4432), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4531 ( .A1(n4166), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4532 ( .A1(n4435), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4533 ( .A1(n4426), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3595) );
  NAND4_X1 U4534 ( .A1(n3598), .A2(n3597), .A3(n3596), .A4(n3595), .ZN(n3599)
         );
  NAND2_X1 U4535 ( .A1(n3722), .A2(n3619), .ZN(n3601) );
  NAND2_X1 U4536 ( .A1(n3606), .A2(n3605), .ZN(n3733) );
  NAND3_X1 U4537 ( .A1(n3629), .A2(n3733), .A3(n4196), .ZN(n3613) );
  NAND2_X1 U4538 ( .A1(n3608), .A2(n3607), .ZN(n3609) );
  OR2_X1 U4539 ( .A1(n3610), .A2(n3609), .ZN(n3618) );
  XNOR2_X1 U4540 ( .A(n3618), .B(n3619), .ZN(n3611) );
  NAND2_X1 U4541 ( .A1(n3611), .A2(n5383), .ZN(n3612) );
  NAND2_X1 U4542 ( .A1(n3613), .A2(n3612), .ZN(n3614) );
  INV_X1 U4543 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U4544 ( .A(n3614), .B(n6264), .ZN(n4812) );
  NAND2_X1 U4545 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  NAND2_X1 U4546 ( .A1(n3614), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3615)
         );
  NAND2_X1 U4547 ( .A1(n4811), .A2(n3615), .ZN(n6200) );
  INV_X1 U4548 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4859) );
  NAND2_X1 U4549 ( .A1(n3722), .A2(n3621), .ZN(n3616) );
  OAI21_X1 U4550 ( .B1(n4859), .B2(n3703), .A(n3616), .ZN(n3617) );
  NAND2_X1 U4551 ( .A1(n3783), .A2(n4196), .ZN(n3624) );
  INV_X1 U4552 ( .A(n3618), .ZN(n3620) );
  NAND2_X1 U4553 ( .A1(n3620), .A2(n3619), .ZN(n3631) );
  XNOR2_X1 U4554 ( .A(n3631), .B(n3621), .ZN(n3622) );
  NAND2_X1 U4555 ( .A1(n3622), .A2(n5383), .ZN(n3623) );
  NAND2_X1 U4556 ( .A1(n3624), .A2(n3623), .ZN(n3625) );
  INV_X1 U4557 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6262) );
  XNOR2_X1 U4558 ( .A(n3625), .B(n6262), .ZN(n6199) );
  NAND2_X1 U4559 ( .A1(n6200), .A2(n6199), .ZN(n6198) );
  NAND2_X1 U4560 ( .A1(n3625), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3626)
         );
  NAND2_X1 U4561 ( .A1(n6198), .A2(n3626), .ZN(n5081) );
  NOR2_X1 U4562 ( .A1(n3627), .A2(n3664), .ZN(n3628) );
  OR3_X1 U4563 ( .A1(n3631), .A2(n3630), .A3(n6706), .ZN(n3632) );
  NAND2_X1 U4564 ( .A1(n5584), .A2(n3632), .ZN(n3633) );
  INV_X1 U4565 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6255) );
  XNOR2_X1 U4566 ( .A(n3633), .B(n6255), .ZN(n5080) );
  NAND2_X1 U4567 ( .A1(n5081), .A2(n5080), .ZN(n5079) );
  NAND2_X1 U4568 ( .A1(n3633), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3634)
         );
  INV_X1 U4569 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U4570 ( .A1(n5584), .A2(n5281), .ZN(n5178) );
  NAND2_X1 U4571 ( .A1(n3138), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5179)
         );
  INV_X1 U4572 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3635) );
  NAND2_X1 U4573 ( .A1(n5584), .A2(n3635), .ZN(n5261) );
  INV_X1 U4574 ( .A(n5290), .ZN(n3636) );
  NAND2_X1 U4575 ( .A1(n3138), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U4576 ( .A1(n3138), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3637) );
  AND2_X1 U4577 ( .A1(n5289), .A2(n3637), .ZN(n3638) );
  INV_X1 U4578 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5779) );
  NOR2_X1 U4579 ( .A1(n5584), .A2(n5779), .ZN(n5317) );
  XNOR2_X1 U4580 ( .A(n5633), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5650)
         );
  INV_X1 U4581 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U4582 ( .A1(n5584), .A2(n4318), .ZN(n3639) );
  NAND2_X1 U4583 ( .A1(n3640), .A2(n3639), .ZN(n5640) );
  INV_X1 U4584 ( .A(n5640), .ZN(n3642) );
  INV_X1 U4585 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4323) );
  INV_X1 U4586 ( .A(n5642), .ZN(n3641) );
  NAND2_X1 U4587 ( .A1(n3138), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5641) );
  INV_X1 U4588 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U4589 ( .A1(n5584), .A2(n5759), .ZN(n3644) );
  AND2_X1 U4590 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4254) );
  NAND2_X1 U4591 ( .A1(n4254), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3645) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5743) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5963) );
  INV_X1 U4594 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6947) );
  NAND3_X1 U4595 ( .A1(n5743), .A2(n5963), .A3(n6947), .ZN(n3646) );
  NAND2_X1 U4596 ( .A1(n3138), .A2(n3646), .ZN(n3647) );
  AND2_X1 U4597 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5734) );
  AND2_X1 U4598 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5718) );
  AND2_X1 U4599 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4256) );
  NAND3_X1 U4600 ( .A1(n5734), .A2(n5718), .A3(n4256), .ZN(n3648) );
  NAND2_X1 U4601 ( .A1(n5584), .A2(n3648), .ZN(n3649) );
  NAND2_X1 U4602 ( .A1(n5952), .A2(n3649), .ZN(n3652) );
  NOR2_X1 U4603 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733) );
  NOR2_X1 U4604 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5700) );
  NOR2_X1 U4605 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5717) );
  NAND3_X1 U4606 ( .A1(n5733), .A2(n5700), .A3(n5717), .ZN(n3650) );
  NAND2_X1 U4607 ( .A1(n3138), .A2(n3650), .ZN(n3651) );
  NAND2_X1 U4608 ( .A1(n3652), .A2(n3651), .ZN(n3656) );
  INV_X1 U4609 ( .A(n3656), .ZN(n3654) );
  INV_X1 U4610 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5976) );
  XNOR2_X1 U4611 ( .A(n5633), .B(n5976), .ZN(n5690) );
  NAND2_X1 U4612 ( .A1(n3654), .A2(n3653), .ZN(n4190) );
  NAND2_X1 U4613 ( .A1(n5584), .A2(n5976), .ZN(n3655) );
  AND2_X2 U4614 ( .A1(n4190), .A2(n3655), .ZN(n5568) );
  NAND3_X1 U4615 ( .A1(n5568), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5584), .ZN(n3658) );
  NOR2_X1 U4616 ( .A1(n5633), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5566)
         );
  NAND2_X1 U4617 ( .A1(n5566), .A2(n5976), .ZN(n3657) );
  INV_X1 U4618 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5977) );
  XNOR2_X1 U4619 ( .A(n3659), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5678)
         );
  NAND2_X1 U4620 ( .A1(n5352), .A2(n3129), .ZN(n3663) );
  XNOR2_X1 U4621 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4622 ( .A1(n3682), .A2(n3680), .ZN(n3666) );
  NAND2_X1 U4623 ( .A1(n6584), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4624 ( .A1(n3666), .A2(n3665), .ZN(n3675) );
  XNOR2_X1 U4625 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3673) );
  NAND2_X1 U4626 ( .A1(n3675), .A2(n3673), .ZN(n3668) );
  NAND2_X1 U4627 ( .A1(n6589), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3667) );
  NAND2_X1 U4628 ( .A1(n3668), .A2(n3667), .ZN(n3712) );
  XNOR2_X1 U4629 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3710) );
  NAND2_X1 U4630 ( .A1(n3712), .A2(n3710), .ZN(n3670) );
  NAND2_X1 U4631 ( .A1(n6325), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3669) );
  NAND2_X1 U4632 ( .A1(n3670), .A2(n3669), .ZN(n3709) );
  NAND2_X1 U4633 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6024), .ZN(n3708) );
  INV_X1 U4634 ( .A(n3722), .ZN(n3677) );
  INV_X1 U4635 ( .A(n3673), .ZN(n3674) );
  XNOR2_X1 U4636 ( .A(n3675), .B(n3674), .ZN(n4202) );
  INV_X1 U4637 ( .A(n4202), .ZN(n3676) );
  AND2_X1 U4638 ( .A1(n3385), .A2(n3357), .ZN(n3678) );
  INV_X1 U4639 ( .A(n3702), .ZN(n3706) );
  NAND2_X1 U4640 ( .A1(n3722), .A2(n4557), .ZN(n3679) );
  NAND2_X1 U4641 ( .A1(n3679), .A2(n3357), .ZN(n3687) );
  INV_X1 U4642 ( .A(n3687), .ZN(n3700) );
  INV_X1 U4643 ( .A(n3680), .ZN(n3681) );
  XNOR2_X1 U4644 ( .A(n3681), .B(n3682), .ZN(n4201) );
  INV_X1 U4645 ( .A(n3686), .ZN(n3699) );
  INV_X1 U4646 ( .A(n3682), .ZN(n3685) );
  NAND2_X1 U4647 ( .A1(n3683), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3684) );
  NAND2_X1 U4648 ( .A1(n3685), .A2(n3684), .ZN(n3689) );
  INV_X1 U4649 ( .A(n3689), .ZN(n3694) );
  OAI21_X1 U4650 ( .B1(n3690), .B2(n3689), .A(n3688), .ZN(n3691) );
  NAND2_X1 U4651 ( .A1(n3702), .A2(n3691), .ZN(n3692) );
  NAND3_X1 U4652 ( .A1(n3694), .A2(n3695), .A3(n3722), .ZN(n3698) );
  INV_X1 U4653 ( .A(n4201), .ZN(n3696) );
  OAI21_X1 U4654 ( .B1(n3696), .B2(n3695), .A(n3717), .ZN(n3697) );
  OAI211_X1 U4655 ( .C1(n3700), .C2(n3699), .A(n3698), .B(n3697), .ZN(n3705)
         );
  INV_X1 U4656 ( .A(n3707), .ZN(n3701) );
  OAI211_X1 U4657 ( .C1(n4202), .C2(n3703), .A(n3702), .B(n3701), .ZN(n3704)
         );
  AOI22_X1 U4658 ( .A1(n3707), .A2(n3706), .B1(n3705), .B2(n3704), .ZN(n3720)
         );
  OR2_X1 U4659 ( .A1(n3709), .A2(n3708), .ZN(n3714) );
  INV_X1 U4660 ( .A(n3710), .ZN(n3711) );
  XNOR2_X1 U4661 ( .A(n3712), .B(n3711), .ZN(n3713) );
  NOR2_X1 U4662 ( .A1(n3715), .A2(n4203), .ZN(n3719) );
  INV_X1 U4663 ( .A(n4203), .ZN(n3716) );
  AOI22_X1 U4664 ( .A1(n3717), .A2(n3716), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6611), .ZN(n3718) );
  OAI21_X1 U4665 ( .B1(n3720), .B2(n3719), .A(n3718), .ZN(n3721) );
  AOI21_X1 U4666 ( .B1(n3722), .B2(n4200), .A(n3721), .ZN(n3723) );
  INV_X1 U4667 ( .A(n3723), .ZN(n3724) );
  NAND2_X1 U4668 ( .A1(n3727), .A2(n3920), .ZN(n3732) );
  INV_X1 U4669 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4766) );
  OAI21_X1 U4670 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3767), .A(n3786), 
        .ZN(n6213) );
  NAND2_X1 U4671 ( .A1(n6213), .A2(n4472), .ZN(n3729) );
  NAND2_X1 U4672 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3728)
         );
  OAI211_X1 U4673 ( .C1(n3210), .C2(n4766), .A(n3729), .B(n3728), .ZN(n3730)
         );
  INV_X1 U4674 ( .A(n3730), .ZN(n3731) );
  NAND2_X1 U4675 ( .A1(n3732), .A2(n3731), .ZN(n4740) );
  NAND2_X1 U4676 ( .A1(n3733), .A2(n3920), .ZN(n3739) );
  INV_X1 U4677 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3735) );
  INV_X1 U4678 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6033) );
  OAI21_X1 U4679 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6033), .A(n5022), 
        .ZN(n3734) );
  OAI21_X1 U4680 ( .B1(n3210), .B2(n3735), .A(n3734), .ZN(n3737) );
  XNOR2_X1 U4681 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .B(n3786), .ZN(n6109) );
  NAND2_X1 U4682 ( .A1(n6109), .A2(n4472), .ZN(n3736) );
  NAND2_X1 U4683 ( .A1(n3737), .A2(n3736), .ZN(n3738) );
  NAND2_X1 U4684 ( .A1(n3739), .A2(n3738), .ZN(n4741) );
  NAND2_X1 U4685 ( .A1(n3740), .A2(n3920), .ZN(n3744) );
  OR2_X1 U4686 ( .A1(n5367), .A2(n5022), .ZN(n3766) );
  INV_X1 U4687 ( .A(n3766), .ZN(n3778) );
  INV_X1 U4688 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3741) );
  INV_X1 U4689 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5155) );
  OAI22_X1 U4690 ( .A1(n3210), .A2(n3741), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5155), .ZN(n3742) );
  AOI21_X1 U4691 ( .B1(n3778), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3742), 
        .ZN(n3743) );
  AOI21_X1 U4692 ( .B1(n3745), .B2(n3268), .A(n5022), .ZN(n4586) );
  NAND2_X1 U4693 ( .A1(n3134), .A2(n3920), .ZN(n3751) );
  INV_X1 U4694 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3748) );
  NAND2_X1 U4695 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n5022), .ZN(n3747)
         );
  OAI21_X1 U4696 ( .B1(n3210), .B2(n3748), .A(n3747), .ZN(n3749) );
  AOI21_X1 U4697 ( .B1(n3778), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n3749), 
        .ZN(n3750) );
  NAND2_X1 U4698 ( .A1(n3751), .A2(n3750), .ZN(n4585) );
  NAND2_X1 U4699 ( .A1(n4586), .A2(n4585), .ZN(n4584) );
  OR2_X1 U4700 ( .A1(n4585), .A2(n4447), .ZN(n3753) );
  NAND2_X1 U4701 ( .A1(n4584), .A2(n3753), .ZN(n4699) );
  AND2_X2 U4702 ( .A1(n4700), .A2(n4699), .ZN(n3759) );
  INV_X1 U4703 ( .A(n3759), .ZN(n3755) );
  INV_X1 U4704 ( .A(n4520), .ZN(n4095) );
  INV_X1 U4705 ( .A(n3760), .ZN(n3754) );
  OAI21_X1 U4706 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3756), .ZN(n6230) );
  AOI22_X1 U4707 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4472), 
        .B2(n6230), .ZN(n3758) );
  NAND2_X1 U4708 ( .A1(n4521), .A2(EAX_REG_2__SCAN_IN), .ZN(n3757) );
  OAI211_X1 U4709 ( .C1(n3766), .C2(n3217), .A(n3758), .B(n3757), .ZN(n4652)
         );
  NAND2_X1 U4710 ( .A1(n4653), .A2(n4652), .ZN(n3762) );
  NAND2_X1 U4711 ( .A1(n3759), .A2(n3760), .ZN(n3761) );
  NAND2_X1 U4712 ( .A1(n3763), .A2(n3920), .ZN(n3772) );
  OAI21_X1 U4713 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6033), .A(n5022), 
        .ZN(n3765) );
  NAND2_X1 U4714 ( .A1(n4521), .A2(EAX_REG_4__SCAN_IN), .ZN(n3764) );
  OAI211_X1 U4715 ( .C1(n3766), .C2(n6024), .A(n3765), .B(n3764), .ZN(n3770)
         );
  AOI21_X1 U4716 ( .B1(n3773), .B2(n3768), .A(n3767), .ZN(n6133) );
  NAND2_X1 U4717 ( .A1(n6133), .A2(n4472), .ZN(n3769) );
  NAND2_X1 U4718 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  NAND2_X1 U4719 ( .A1(n4792), .A2(n3920), .ZN(n3780) );
  INV_X1 U4720 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3776) );
  OAI21_X1 U4721 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3774), .A(n3773), 
        .ZN(n6221) );
  AOI22_X1 U4722 ( .A1(n4472), .A2(n6221), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3775) );
  OAI21_X1 U4723 ( .B1(n3210), .B2(n3776), .A(n3775), .ZN(n3777) );
  AOI21_X1 U4724 ( .B1(n3778), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3777), 
        .ZN(n3779) );
  AND2_X2 U4725 ( .A1(n4651), .A2(n3781), .ZN(n4715) );
  NAND2_X1 U4726 ( .A1(n3783), .A2(n3920), .ZN(n3793) );
  AOI22_X1 U4727 ( .A1(n4521), .A2(EAX_REG_7__SCAN_IN), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3784) );
  OR2_X1 U4728 ( .A1(n3787), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3788) );
  NAND2_X1 U4729 ( .A1(n3788), .A2(n3809), .ZN(n6205) );
  INV_X1 U4730 ( .A(n6205), .ZN(n3789) );
  NAND2_X1 U4731 ( .A1(n4521), .A2(EAX_REG_8__SCAN_IN), .ZN(n3807) );
  XNOR2_X1 U4732 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3809), .ZN(n5084) );
  INV_X1 U4733 ( .A(n5084), .ZN(n5269) );
  AOI22_X1 U4734 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4472), 
        .B2(n5269), .ZN(n3806) );
  AOI22_X1 U4735 ( .A1(n4425), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4736 ( .A1(n4432), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4737 ( .A1(n4014), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4738 ( .A1(n4426), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3794) );
  NAND4_X1 U4739 ( .A1(n3797), .A2(n3796), .A3(n3795), .A4(n3794), .ZN(n3803)
         );
  AOI22_X1 U4740 ( .A1(n3133), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4741 ( .A1(n4424), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4742 ( .A1(n4435), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3799) );
  AOI22_X1 U4743 ( .A1(n4403), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3798) );
  NAND4_X1 U4744 ( .A1(n3801), .A2(n3800), .A3(n3799), .A4(n3798), .ZN(n3802)
         );
  NOR2_X1 U4745 ( .A1(n3803), .A2(n3802), .ZN(n3804) );
  OR2_X1 U4746 ( .A1(n3904), .A2(n3804), .ZN(n3805) );
  NAND2_X1 U4747 ( .A1(n3811), .A2(n6950), .ZN(n3813) );
  INV_X1 U4748 ( .A(n3854), .ZN(n3812) );
  NAND2_X1 U4749 ( .A1(n3813), .A2(n3812), .ZN(n5254) );
  NAND2_X1 U4750 ( .A1(n5254), .A2(n3752), .ZN(n3829) );
  AOI22_X1 U4751 ( .A1(n3133), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4752 ( .A1(n4432), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4753 ( .A1(n4425), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4754 ( .A1(n4166), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3814) );
  NAND4_X1 U4755 ( .A1(n3817), .A2(n3816), .A3(n3815), .A4(n3814), .ZN(n3823)
         );
  AOI22_X1 U4756 ( .A1(n4431), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4757 ( .A1(n4426), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4758 ( .A1(n4435), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4759 ( .A1(n4014), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4760 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3822)
         );
  NOR2_X1 U4761 ( .A1(n3823), .A2(n3822), .ZN(n3826) );
  NAND2_X1 U4762 ( .A1(n4521), .A2(EAX_REG_9__SCAN_IN), .ZN(n3825) );
  NAND2_X1 U4763 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3824)
         );
  OAI211_X1 U4764 ( .C1(n3826), .C2(n3904), .A(n3825), .B(n3824), .ZN(n3827)
         );
  INV_X1 U4765 ( .A(n3827), .ZN(n3828) );
  AOI22_X1 U4766 ( .A1(n4425), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4767 ( .A1(n4403), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4768 ( .A1(n4424), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4769 ( .A1(n4127), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4770 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3839)
         );
  AOI22_X1 U4771 ( .A1(n4031), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4772 ( .A1(n4432), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4426), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4773 ( .A1(n4435), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4774 ( .A1(n4014), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4775 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  NOR2_X1 U4776 ( .A1(n3839), .A2(n3838), .ZN(n3843) );
  NAND2_X1 U4777 ( .A1(n4521), .A2(EAX_REG_10__SCAN_IN), .ZN(n3842) );
  XOR2_X1 U4778 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3854), .Z(n6082) );
  INV_X1 U4779 ( .A(n6082), .ZN(n3840) );
  AOI22_X1 U4780 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n3752), 
        .B2(n3840), .ZN(n3841) );
  OAI211_X1 U4781 ( .C1(n3904), .C2(n3843), .A(n3842), .B(n3841), .ZN(n5119)
         );
  AOI22_X1 U4782 ( .A1(n4425), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4783 ( .A1(n4432), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4784 ( .A1(n4424), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4785 ( .A1(n3336), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3844) );
  NAND4_X1 U4786 ( .A1(n3847), .A2(n3846), .A3(n3845), .A4(n3844), .ZN(n3853)
         );
  AOI22_X1 U4787 ( .A1(n4014), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4788 ( .A1(n4435), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4426), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4789 ( .A1(n4031), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4790 ( .A1(n4403), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4791 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3852)
         );
  NOR2_X1 U4792 ( .A1(n3853), .A2(n3852), .ZN(n3860) );
  NAND2_X1 U4793 ( .A1(n4521), .A2(EAX_REG_11__SCAN_IN), .ZN(n3859) );
  INV_X1 U4794 ( .A(n3855), .ZN(n3857) );
  INV_X1 U4795 ( .A(n3876), .ZN(n3856) );
  OAI21_X1 U4796 ( .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n3857), .A(n3856), 
        .ZN(n6067) );
  AOI22_X1 U4797 ( .A1(n4472), .A2(n6067), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3858) );
  OAI211_X1 U4798 ( .C1(n3904), .C2(n3860), .A(n3859), .B(n3858), .ZN(n5128)
         );
  NAND2_X1 U4799 ( .A1(n4521), .A2(EAX_REG_12__SCAN_IN), .ZN(n3875) );
  XOR2_X1 U4800 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3876), .Z(n6060) );
  INV_X1 U4801 ( .A(n6060), .ZN(n3861) );
  AOI22_X1 U4802 ( .A1(n4520), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n3752), 
        .B2(n3861), .ZN(n3874) );
  AOI22_X1 U4803 ( .A1(n4014), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4804 ( .A1(n4425), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4805 ( .A1(n4426), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4806 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4435), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4807 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3871)
         );
  AOI22_X1 U4808 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4424), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4809 ( .A1(n4432), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4810 ( .A1(n3133), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4811 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4166), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3866) );
  NAND4_X1 U4812 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  NOR2_X1 U4813 ( .A1(n3871), .A2(n3870), .ZN(n3872) );
  OR2_X1 U4814 ( .A1(n3904), .A2(n3872), .ZN(n3873) );
  NAND2_X1 U4815 ( .A1(n4521), .A2(EAX_REG_13__SCAN_IN), .ZN(n3879) );
  INV_X1 U4816 ( .A(n3892), .ZN(n3877) );
  XNOR2_X1 U4817 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3877), .ZN(n5652)
         );
  AOI22_X1 U4818 ( .A1(n4472), .A2(n5652), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3878) );
  NAND2_X1 U4819 ( .A1(n3879), .A2(n3878), .ZN(n3891) );
  AOI22_X1 U4820 ( .A1(n3133), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4821 ( .A1(n4425), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4822 ( .A1(n4014), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4823 ( .A1(n3336), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4824 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  AOI22_X1 U4825 ( .A1(n4431), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4432), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4826 ( .A1(n4937), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4426), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4827 ( .A1(n4424), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4828 ( .A1(n4435), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4829 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  NOR2_X1 U4830 ( .A1(n3889), .A2(n3888), .ZN(n3890) );
  NOR2_X1 U4831 ( .A1(n3904), .A2(n3890), .ZN(n5300) );
  NAND2_X1 U4832 ( .A1(n4521), .A2(EAX_REG_14__SCAN_IN), .ZN(n3907) );
  XNOR2_X1 U4833 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3908), .ZN(n5645)
         );
  AOI22_X1 U4834 ( .A1(n4472), .A2(n5645), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4835 ( .A1(n4014), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4836 ( .A1(n4425), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4837 ( .A1(n4432), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4838 ( .A1(n4435), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3893) );
  NAND4_X1 U4839 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3902)
         );
  AOI22_X1 U4840 ( .A1(n4424), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4841 ( .A1(n4426), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4842 ( .A1(n4403), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4843 ( .A1(n3133), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3897) );
  NAND4_X1 U4844 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3901)
         );
  NOR2_X1 U4845 ( .A1(n3902), .A2(n3901), .ZN(n3903) );
  OR2_X1 U4846 ( .A1(n3904), .A2(n3903), .ZN(n3905) );
  XNOR2_X1 U4847 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3924), .ZN(n5636)
         );
  AOI22_X1 U4848 ( .A1(n4014), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4849 ( .A1(n4431), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4850 ( .A1(n4166), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4851 ( .A1(n4435), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3909) );
  NAND4_X1 U4852 ( .A1(n3912), .A2(n3911), .A3(n3910), .A4(n3909), .ZN(n3918)
         );
  AOI22_X1 U4853 ( .A1(n4432), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4854 ( .A1(n4425), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4855 ( .A1(n4426), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4856 ( .A1(n4031), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3913) );
  NAND4_X1 U4857 ( .A1(n3916), .A2(n3915), .A3(n3914), .A4(n3913), .ZN(n3917)
         );
  OR2_X1 U4858 ( .A1(n3918), .A2(n3917), .ZN(n3919) );
  AOI22_X1 U4859 ( .A1(n3920), .A2(n3919), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3922) );
  NAND2_X1 U4860 ( .A1(n4521), .A2(EAX_REG_15__SCAN_IN), .ZN(n3921) );
  OAI211_X1 U4861 ( .C1(n5636), .C2(n4447), .A(n3922), .B(n3921), .ZN(n5475)
         );
  XNOR2_X1 U4862 ( .A(n3955), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5627)
         );
  NAND2_X1 U4863 ( .A1(n5627), .A2(n3752), .ZN(n3940) );
  AOI22_X1 U4864 ( .A1(n4014), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4865 ( .A1(n4424), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4866 ( .A1(n4425), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3926) );
  AOI22_X1 U4867 ( .A1(n4426), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3925) );
  NAND4_X1 U4868 ( .A1(n3928), .A2(n3927), .A3(n3926), .A4(n3925), .ZN(n3934)
         );
  AOI22_X1 U4869 ( .A1(n4031), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4870 ( .A1(n4403), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4871 ( .A1(n4166), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4872 ( .A1(n4435), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3929) );
  NAND4_X1 U4873 ( .A1(n3932), .A2(n3931), .A3(n3930), .A4(n3929), .ZN(n3933)
         );
  OR2_X1 U4874 ( .A1(n3934), .A2(n3933), .ZN(n3938) );
  INV_X1 U4875 ( .A(EAX_REG_16__SCAN_IN), .ZN(n3936) );
  INV_X1 U4876 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3935) );
  OAI22_X1 U4877 ( .A1(n3210), .A2(n3936), .B1(n4095), .B2(n3935), .ZN(n3937)
         );
  AOI21_X1 U4878 ( .B1(n4444), .B2(n3938), .A(n3937), .ZN(n3939) );
  NAND2_X1 U4879 ( .A1(n3940), .A2(n3939), .ZN(n5457) );
  AOI22_X1 U4880 ( .A1(n4014), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4881 ( .A1(n4403), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4882 ( .A1(n4435), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4426), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4883 ( .A1(n4166), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4884 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3950)
         );
  AOI22_X1 U4885 ( .A1(n4425), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4886 ( .A1(n4431), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4887 ( .A1(n3133), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4888 ( .A1(n3336), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4889 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  NOR2_X1 U4890 ( .A1(n3950), .A2(n3949), .ZN(n3954) );
  NAND2_X1 U4891 ( .A1(n6465), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3951)
         );
  NAND2_X1 U4892 ( .A1(n4447), .A2(n3951), .ZN(n3952) );
  AOI21_X1 U4893 ( .B1(n4521), .B2(EAX_REG_17__SCAN_IN), .A(n3952), .ZN(n3953)
         );
  OAI21_X1 U4894 ( .B1(n4415), .B2(n3954), .A(n3953), .ZN(n3958) );
  OAI21_X1 U4895 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3956), .A(n3976), 
        .ZN(n5965) );
  OR2_X1 U4896 ( .A1(n4447), .A2(n5965), .ZN(n3957) );
  NAND2_X1 U4897 ( .A1(n3958), .A2(n3957), .ZN(n5446) );
  AOI22_X1 U4898 ( .A1(n4014), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4899 ( .A1(n4432), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4900 ( .A1(n4431), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4901 ( .A1(n4435), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3960) );
  NAND4_X1 U4902 ( .A1(n3963), .A2(n3962), .A3(n3961), .A4(n3960), .ZN(n3969)
         );
  AOI22_X1 U4903 ( .A1(n4425), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4904 ( .A1(n4166), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4905 ( .A1(n4426), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3336), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4906 ( .A1(n4031), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3964) );
  NAND4_X1 U4907 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3968)
         );
  NOR2_X1 U4908 ( .A1(n3969), .A2(n3968), .ZN(n3973) );
  NAND2_X1 U4909 ( .A1(n5022), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3970)
         );
  NAND2_X1 U4910 ( .A1(n4447), .A2(n3970), .ZN(n3971) );
  AOI21_X1 U4911 ( .B1(n4521), .B2(EAX_REG_18__SCAN_IN), .A(n3971), .ZN(n3972)
         );
  OAI21_X1 U4912 ( .B1(n4415), .B2(n3973), .A(n3972), .ZN(n3975) );
  XNOR2_X1 U4913 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3976), .ZN(n5622)
         );
  NAND2_X1 U4914 ( .A1(n5622), .A2(n3752), .ZN(n3974) );
  NAND2_X1 U4915 ( .A1(n5431), .A2(n3155), .ZN(n5429) );
  OR2_X1 U4916 ( .A1(n3977), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3978)
         );
  NAND2_X1 U4917 ( .A1(n3978), .A2(n4025), .ZN(n5960) );
  AOI22_X1 U4918 ( .A1(n4014), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4919 ( .A1(n4031), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4920 ( .A1(n4432), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4921 ( .A1(n4426), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4922 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3988)
         );
  AOI22_X1 U4923 ( .A1(n4403), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4924 ( .A1(n4431), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4925 ( .A1(n4435), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4926 ( .A1(n4425), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3983) );
  NAND4_X1 U4927 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n3987)
         );
  NOR2_X1 U4928 ( .A1(n3988), .A2(n3987), .ZN(n3989) );
  NOR2_X1 U4929 ( .A1(n4415), .A2(n3989), .ZN(n3993) );
  INV_X1 U4930 ( .A(EAX_REG_19__SCAN_IN), .ZN(n3991) );
  NAND2_X1 U4931 ( .A1(n6465), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3990)
         );
  OAI211_X1 U4932 ( .C1(n3210), .C2(n3991), .A(n4447), .B(n3990), .ZN(n3992)
         );
  OAI22_X1 U4933 ( .A1(n5960), .A2(n4447), .B1(n3993), .B2(n3992), .ZN(n5902)
         );
  AOI22_X1 U4934 ( .A1(n4014), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4935 ( .A1(n4425), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4936 ( .A1(n4424), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3995) );
  AOI22_X1 U4937 ( .A1(n4031), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3994) );
  NAND4_X1 U4938 ( .A1(n3997), .A2(n3996), .A3(n3995), .A4(n3994), .ZN(n4004)
         );
  AOI22_X1 U4939 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4403), .B1(n3998), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4940 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4166), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4941 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4435), .B1(n3336), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4942 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4426), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4943 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4003)
         );
  NOR2_X1 U4944 ( .A1(n4004), .A2(n4003), .ZN(n4007) );
  INV_X1 U4945 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5897) );
  AOI21_X1 U4946 ( .B1(n5897), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4005) );
  AOI21_X1 U4947 ( .B1(n4521), .B2(EAX_REG_20__SCAN_IN), .A(n4005), .ZN(n4006)
         );
  OAI21_X1 U4948 ( .B1(n4415), .B2(n4007), .A(n4006), .ZN(n4009) );
  XNOR2_X1 U4949 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4025), .ZN(n5888)
         );
  NAND2_X1 U4950 ( .A1(n5888), .A2(n4472), .ZN(n4008) );
  AOI22_X1 U4951 ( .A1(n4425), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4952 ( .A1(n4432), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4012) );
  AOI22_X1 U4953 ( .A1(n4403), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4954 ( .A1(n4435), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4010) );
  NAND4_X1 U4955 ( .A1(n4013), .A2(n4012), .A3(n4011), .A4(n4010), .ZN(n4020)
         );
  AOI22_X1 U4956 ( .A1(n4014), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4957 ( .A1(n4431), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4958 ( .A1(n4426), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4959 ( .A1(n4031), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4015) );
  NAND4_X1 U4960 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4019)
         );
  NOR2_X1 U4961 ( .A1(n4020), .A2(n4019), .ZN(n4024) );
  NAND2_X1 U4962 ( .A1(n5022), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4021)
         );
  NAND2_X1 U4963 ( .A1(n4447), .A2(n4021), .ZN(n4022) );
  AOI21_X1 U4964 ( .B1(n4521), .B2(EAX_REG_21__SCAN_IN), .A(n4022), .ZN(n4023)
         );
  OAI21_X1 U4965 ( .B1(n4415), .B2(n4024), .A(n4023), .ZN(n4029) );
  OAI21_X1 U4966 ( .B1(n4027), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4074), 
        .ZN(n5607) );
  OR2_X1 U4967 ( .A1(n5607), .A2(n4447), .ZN(n4028) );
  NAND2_X1 U4968 ( .A1(n4029), .A2(n4028), .ZN(n5416) );
  AOI22_X1 U4969 ( .A1(n4014), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4970 ( .A1(n4425), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4034) );
  INV_X1 U4971 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U4972 ( .A1(n4424), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4973 ( .A1(n4031), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4032) );
  NAND4_X1 U4974 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4041)
         );
  AOI22_X1 U4975 ( .A1(n4432), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4976 ( .A1(n4166), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4977 ( .A1(n4435), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4978 ( .A1(n4426), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U4979 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4040)
         );
  NOR2_X1 U4980 ( .A1(n4041), .A2(n4040), .ZN(n4045) );
  INV_X1 U4981 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4042) );
  AOI21_X1 U4982 ( .B1(n4042), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4043) );
  AOI21_X1 U4983 ( .B1(n4521), .B2(EAX_REG_22__SCAN_IN), .A(n4043), .ZN(n4044)
         );
  OAI21_X1 U4984 ( .B1(n4415), .B2(n4045), .A(n4044), .ZN(n4047) );
  XNOR2_X1 U4985 ( .A(n4074), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5881)
         );
  NAND2_X1 U4986 ( .A1(n5881), .A2(n3752), .ZN(n4046) );
  NAND2_X1 U4987 ( .A1(n4047), .A2(n4046), .ZN(n5512) );
  AOI22_X1 U4988 ( .A1(n4014), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4425), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4989 ( .A1(n4431), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4990 ( .A1(n4435), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4426), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4991 ( .A1(n4127), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U4992 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4057)
         );
  AOI22_X1 U4993 ( .A1(n4031), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4994 ( .A1(n4432), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4995 ( .A1(n3133), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4996 ( .A1(n3318), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U4997 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  NOR2_X1 U4998 ( .A1(n4057), .A2(n4056), .ZN(n4079) );
  AOI22_X1 U4999 ( .A1(n4425), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U5000 ( .A1(n4127), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5001 ( .A1(n4426), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5002 ( .A1(n4014), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4058) );
  NAND4_X1 U5003 ( .A1(n4061), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4067)
         );
  AOI22_X1 U5004 ( .A1(n3133), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4065) );
  AOI22_X1 U5005 ( .A1(n4432), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5006 ( .A1(n3318), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4435), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5007 ( .A1(n4424), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5008 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4066)
         );
  NOR2_X1 U5009 ( .A1(n4067), .A2(n4066), .ZN(n4080) );
  XNOR2_X1 U5010 ( .A(n4079), .B(n4080), .ZN(n4071) );
  NAND2_X1 U5011 ( .A1(n5022), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4068)
         );
  NAND2_X1 U5012 ( .A1(n4447), .A2(n4068), .ZN(n4069) );
  AOI21_X1 U5013 ( .B1(n4521), .B2(EAX_REG_23__SCAN_IN), .A(n4069), .ZN(n4070)
         );
  OAI21_X1 U5014 ( .B1(n4415), .B2(n4071), .A(n4070), .ZN(n4078) );
  INV_X1 U5015 ( .A(n4074), .ZN(n4072) );
  AOI21_X1 U5016 ( .B1(n4072), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4075) );
  NAND2_X1 U5017 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4073) );
  OR2_X1 U5018 ( .A1(n4075), .A2(n4093), .ZN(n5873) );
  INV_X1 U5019 ( .A(n5873), .ZN(n4076) );
  NAND2_X1 U5020 ( .A1(n4076), .A2(n3752), .ZN(n4077) );
  NOR2_X1 U5021 ( .A1(n4080), .A2(n4079), .ZN(n4110) );
  AOI22_X1 U5022 ( .A1(n4014), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5023 ( .A1(n4425), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5024 ( .A1(n4424), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4082) );
  AOI22_X1 U5025 ( .A1(n4031), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4081) );
  NAND4_X1 U5026 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4090)
         );
  AOI22_X1 U5027 ( .A1(n4432), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5028 ( .A1(n4166), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5029 ( .A1(n4435), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5030 ( .A1(n4426), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4085) );
  NAND4_X1 U5031 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4089)
         );
  OR2_X1 U5032 ( .A1(n4090), .A2(n4089), .ZN(n4109) );
  INV_X1 U5033 ( .A(n4109), .ZN(n4091) );
  XNOR2_X1 U5034 ( .A(n4110), .B(n4091), .ZN(n4092) );
  NAND2_X1 U5035 ( .A1(n4092), .A2(n4444), .ZN(n4098) );
  OR2_X1 U5036 ( .A1(n4093), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4094)
         );
  AND2_X1 U5037 ( .A1(n4115), .A2(n4094), .ZN(n5864) );
  INV_X1 U5038 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6808) );
  OAI22_X1 U5039 ( .A1(n5864), .A2(n4447), .B1(n6808), .B2(n4095), .ZN(n4096)
         );
  AOI21_X1 U5040 ( .B1(n4521), .B2(EAX_REG_24__SCAN_IN), .A(n4096), .ZN(n4097)
         );
  NAND2_X1 U5041 ( .A1(n4098), .A2(n4097), .ZN(n5505) );
  NAND2_X1 U5042 ( .A1(n5504), .A2(n5505), .ZN(n5395) );
  AOI22_X1 U5043 ( .A1(n4014), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5044 ( .A1(n4031), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5045 ( .A1(n4432), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4166), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5046 ( .A1(n4426), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4099) );
  NAND4_X1 U5047 ( .A1(n4102), .A2(n4101), .A3(n4100), .A4(n4099), .ZN(n4108)
         );
  AOI22_X1 U5048 ( .A1(n4431), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5049 ( .A1(n4435), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5050 ( .A1(n4403), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5051 ( .A1(n4425), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5052 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4107)
         );
  NOR2_X1 U5053 ( .A1(n4108), .A2(n4107), .ZN(n4121) );
  NAND2_X1 U5054 ( .A1(n4110), .A2(n4109), .ZN(n4120) );
  XNOR2_X1 U5055 ( .A(n4121), .B(n4120), .ZN(n4113) );
  INV_X1 U5056 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4114) );
  OAI21_X1 U5057 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4114), .A(n4447), .ZN(
        n4111) );
  AOI21_X1 U5058 ( .B1(n4521), .B2(EAX_REG_25__SCAN_IN), .A(n4111), .ZN(n4112)
         );
  OAI21_X1 U5059 ( .B1(n4113), .B2(n4415), .A(n4112), .ZN(n4118) );
  NAND2_X1 U5060 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  NAND2_X1 U5061 ( .A1(n4155), .A2(n4116), .ZN(n5950) );
  NAND2_X1 U5062 ( .A1(n4118), .A2(n4117), .ZN(n5397) );
  NOR2_X1 U5063 ( .A1(n4121), .A2(n4120), .ZN(n4141) );
  AOI22_X1 U5064 ( .A1(n4014), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5065 ( .A1(n4425), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5066 ( .A1(n4424), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5067 ( .A1(n4031), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4122), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5068 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4133)
         );
  AOI22_X1 U5069 ( .A1(n4432), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5070 ( .A1(n3318), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5071 ( .A1(n4435), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5072 ( .A1(n4426), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5073 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4132)
         );
  OR2_X1 U5074 ( .A1(n4133), .A2(n4132), .ZN(n4140) );
  XNOR2_X1 U5075 ( .A(n4141), .B(n4140), .ZN(n4136) );
  INV_X1 U5076 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5571) );
  AOI21_X1 U5077 ( .B1(n5571), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4134) );
  AOI21_X1 U5078 ( .B1(n4521), .B2(EAX_REG_26__SCAN_IN), .A(n4134), .ZN(n4135)
         );
  OAI21_X1 U5079 ( .B1(n4136), .B2(n4415), .A(n4135), .ZN(n4138) );
  XNOR2_X1 U5080 ( .A(n4155), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5855)
         );
  NAND2_X1 U5081 ( .A1(n5855), .A2(n4472), .ZN(n4137) );
  NAND2_X1 U5082 ( .A1(n4138), .A2(n4137), .ZN(n5494) );
  NAND2_X1 U5083 ( .A1(n4141), .A2(n4140), .ZN(n4160) );
  AOI22_X1 U5084 ( .A1(n4014), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4145) );
  AOI22_X1 U5085 ( .A1(n4431), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5086 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4166), .B1(n4426), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5087 ( .A1(n4031), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4142) );
  NAND4_X1 U5088 ( .A1(n4145), .A2(n4144), .A3(n4143), .A4(n4142), .ZN(n4151)
         );
  AOI22_X1 U5089 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4432), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5090 ( .A1(n4425), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5091 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n4435), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5092 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3416), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4146) );
  NAND4_X1 U5093 ( .A1(n4149), .A2(n4148), .A3(n4147), .A4(n4146), .ZN(n4150)
         );
  NOR2_X1 U5094 ( .A1(n4151), .A2(n4150), .ZN(n4161) );
  XNOR2_X1 U5095 ( .A(n4160), .B(n4161), .ZN(n4154) );
  INV_X1 U5096 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5849) );
  AOI21_X1 U5097 ( .B1(n5849), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4152) );
  AOI21_X1 U5098 ( .B1(n4521), .B2(EAX_REG_27__SCAN_IN), .A(n4152), .ZN(n4153)
         );
  OAI21_X1 U5099 ( .B1(n4154), .B2(n4415), .A(n4153), .ZN(n4159) );
  NOR2_X1 U5100 ( .A1(n4156), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4157)
         );
  NAND2_X1 U5101 ( .A1(n4159), .A2(n4158), .ZN(n5562) );
  NOR2_X1 U5102 ( .A1(n4161), .A2(n4160), .ZN(n4411) );
  AOI22_X1 U5103 ( .A1(n4014), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4165) );
  AOI22_X1 U5104 ( .A1(n4425), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4431), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5105 ( .A1(n4424), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5106 ( .A1(n4031), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4162) );
  NAND4_X1 U5107 ( .A1(n4165), .A2(n4164), .A3(n4163), .A4(n4162), .ZN(n4172)
         );
  AOI22_X1 U5108 ( .A1(n4432), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5109 ( .A1(n4166), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5110 ( .A1(n4435), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5111 ( .A1(n4426), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U5112 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4171)
         );
  OR2_X1 U5113 ( .A1(n4172), .A2(n4171), .ZN(n4410) );
  INV_X1 U5114 ( .A(n4410), .ZN(n4173) );
  XNOR2_X1 U5115 ( .A(n4411), .B(n4173), .ZN(n4174) );
  NAND2_X1 U5116 ( .A1(n4174), .A2(n4444), .ZN(n4179) );
  NAND2_X1 U5117 ( .A1(n5022), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4175)
         );
  NAND2_X1 U5118 ( .A1(n4447), .A2(n4175), .ZN(n4176) );
  AOI21_X1 U5119 ( .B1(n4521), .B2(EAX_REG_28__SCAN_IN), .A(n4176), .ZN(n4178)
         );
  INV_X1 U5120 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4187) );
  XNOR2_X1 U5121 ( .A(n4417), .B(n4187), .ZN(n4496) );
  AOI21_X1 U5122 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4180) );
  NOR2_X1 U5123 ( .A1(n5561), .A2(n4180), .ZN(n4181) );
  AND2_X1 U5124 ( .A1(n6611), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U5125 ( .A1(n4473), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6624) );
  NOR2_X1 U5126 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n4540) );
  NAND2_X1 U5127 ( .A1(n6499), .A2(n4186), .ZN(n6703) );
  NAND2_X1 U5128 ( .A1(n6703), .A2(n6611), .ZN(n4182) );
  NAND2_X1 U5129 ( .A1(n6611), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4184) );
  NAND2_X1 U5130 ( .A1(n6033), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4183) );
  AND2_X1 U5131 ( .A1(n4184), .A2(n4183), .ZN(n4588) );
  INV_X1 U5132 ( .A(n4588), .ZN(n4185) );
  OR2_X2 U5133 ( .A1(n4186), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6232) );
  INV_X2 U5134 ( .A(n6232), .ZN(n6308) );
  NAND2_X1 U5135 ( .A1(n6308), .A2(REIP_REG_28__SCAN_IN), .ZN(n5673) );
  OAI21_X1 U5136 ( .B1(n5969), .B2(n4187), .A(n5673), .ZN(n4188) );
  NOR2_X1 U5137 ( .A1(n3138), .A2(n5977), .ZN(n5567) );
  NAND2_X1 U5138 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4258) );
  AND2_X1 U5139 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4259) );
  INV_X1 U5140 ( .A(n4190), .ZN(n4193) );
  NOR2_X1 U5141 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4191) );
  NAND2_X1 U5142 ( .A1(n5566), .A2(n4191), .ZN(n4389) );
  NOR3_X1 U5143 ( .A1(n4389), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4192) );
  INV_X1 U5144 ( .A(n4530), .ZN(n4388) );
  INV_X1 U5145 ( .A(n4471), .ZN(n4546) );
  NAND2_X1 U5146 ( .A1(n4211), .A2(n3363), .ZN(n4227) );
  NAND2_X1 U5147 ( .A1(n4196), .A2(n3268), .ZN(n4226) );
  NAND3_X1 U5148 ( .A1(n4227), .A2(n4217), .A3(n4226), .ZN(n4197) );
  NAND2_X1 U5149 ( .A1(n4197), .A2(n4216), .ZN(n4198) );
  NAND2_X1 U5150 ( .A1(n4546), .A2(n4198), .ZN(n4668) );
  NOR2_X1 U5151 ( .A1(n5352), .A2(n4456), .ZN(n4234) );
  INV_X1 U5152 ( .A(n4234), .ZN(n4207) );
  OR2_X1 U5153 ( .A1(n4199), .A2(STATE_REG_0__SCAN_IN), .ZN(n6632) );
  INV_X1 U5154 ( .A(n4200), .ZN(n4205) );
  NAND3_X1 U5155 ( .A1(n4203), .A2(n4202), .A3(n4201), .ZN(n4204) );
  NAND2_X1 U5156 ( .A1(n4205), .A2(n4204), .ZN(n4470) );
  NOR2_X1 U5157 ( .A1(READY_N), .A2(n4470), .ZN(n4655) );
  OAI211_X1 U5158 ( .C1(n3385), .C2(n4673), .A(n4669), .B(n4655), .ZN(n4206)
         );
  OAI21_X1 U5159 ( .B1(n4692), .B2(n4207), .A(n4206), .ZN(n4208) );
  INV_X1 U5160 ( .A(n4208), .ZN(n4209) );
  AOI21_X1 U5161 ( .B1(n4668), .B2(n4209), .A(n6617), .ZN(n4215) );
  OR2_X1 U5162 ( .A1(n4557), .A2(n4673), .ZN(n4488) );
  NAND3_X1 U5163 ( .A1(n4686), .A2(n4488), .A3(n6704), .ZN(n4212) );
  NAND3_X1 U5164 ( .A1(n4212), .A2(n4217), .A3(n5367), .ZN(n4213) );
  AND3_X1 U5165 ( .A1(n4213), .A2(n4567), .A3(n4747), .ZN(n4214) );
  NAND2_X1 U5166 ( .A1(n4216), .A2(n3388), .ZN(n4656) );
  INV_X1 U5167 ( .A(n4656), .ZN(n4919) );
  NOR2_X1 U5168 ( .A1(n4919), .A2(n6593), .ZN(n4549) );
  INV_X1 U5169 ( .A(n4383), .ZN(n4218) );
  AOI22_X1 U5170 ( .A1(n4686), .A2(n4672), .B1(n4218), .B2(n4382), .ZN(n4220)
         );
  NAND3_X1 U5171 ( .A1(n4549), .A2(n4220), .A3(n4219), .ZN(n4221) );
  INV_X1 U5172 ( .A(n5367), .ZN(n4222) );
  OAI22_X1 U5173 ( .A1(n3661), .A2(n3128), .B1(n4747), .B2(n4222), .ZN(n4225)
         );
  NAND2_X1 U5174 ( .A1(n4779), .A2(n4217), .ZN(n4269) );
  AOI21_X1 U5175 ( .B1(n4642), .B2(n4456), .A(n4223), .ZN(n4224) );
  NOR2_X1 U5176 ( .A1(n4225), .A2(n4224), .ZN(n4231) );
  NAND2_X1 U5177 ( .A1(n4227), .A2(n4226), .ZN(n4228) );
  NAND2_X1 U5178 ( .A1(n4228), .A2(n4747), .ZN(n4229) );
  NAND2_X1 U5179 ( .A1(n4229), .A2(n4217), .ZN(n4230) );
  NAND3_X1 U5180 ( .A1(n4232), .A2(n4231), .A3(n4230), .ZN(n4690) );
  OAI21_X1 U5181 ( .B1(n4687), .B2(n4217), .A(n4939), .ZN(n4233) );
  NOR2_X1 U5182 ( .A1(n4690), .A2(n4233), .ZN(n4235) );
  INV_X1 U5183 ( .A(n4235), .ZN(n4236) );
  NAND2_X1 U5184 ( .A1(n4236), .A2(n4385), .ZN(n6010) );
  NAND2_X1 U5185 ( .A1(n6291), .A2(n6010), .ZN(n5768) );
  INV_X1 U5186 ( .A(n5768), .ZN(n4237) );
  INV_X1 U5187 ( .A(n5765), .ZN(n4238) );
  NOR2_X1 U5188 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n4238), .ZN(n4707)
         );
  OR2_X1 U5189 ( .A1(n6317), .A2(n6311), .ZN(n4248) );
  INV_X1 U5190 ( .A(n4256), .ZN(n4247) );
  NOR2_X1 U5191 ( .A1(n6262), .A2(n6255), .ZN(n6250) );
  NAND3_X1 U5192 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6250), .ZN(n4242) );
  NOR2_X1 U5193 ( .A1(n4280), .A2(n4287), .ZN(n6297) );
  INV_X1 U5194 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6320) );
  NOR2_X1 U5195 ( .A1(n6320), .A2(n6313), .ZN(n6284) );
  NAND4_X1 U5196 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n6297), .A4(n6284), .ZN(n5279) );
  NOR2_X1 U5197 ( .A1(n4242), .A2(n5279), .ZN(n5752) );
  NAND2_X1 U5198 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U5199 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5769) );
  NOR2_X1 U5200 ( .A1(n4318), .A2(n5769), .ZN(n5766) );
  NAND2_X1 U5201 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5766), .ZN(n5751) );
  NOR2_X1 U5202 ( .A1(n6003), .A2(n5751), .ZN(n4243) );
  NAND2_X1 U5203 ( .A1(n5752), .A2(n4243), .ZN(n4239) );
  NAND2_X1 U5204 ( .A1(n6269), .A2(n4239), .ZN(n4241) );
  INV_X1 U5205 ( .A(n4385), .ZN(n4240) );
  NAND2_X1 U5206 ( .A1(n4240), .A2(n6232), .ZN(n4640) );
  INV_X1 U5207 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U5208 ( .A1(n6306), .A2(n5768), .ZN(n4646) );
  NAND2_X1 U5209 ( .A1(n4640), .A2(n4646), .ZN(n5755) );
  NAND2_X1 U5210 ( .A1(n6291), .A2(n5755), .ZN(n6267) );
  AND2_X1 U5211 ( .A1(n4241), .A2(n6267), .ZN(n5738) );
  OAI21_X1 U5212 ( .B1(n6313), .B2(n6306), .A(n6320), .ZN(n6305) );
  NAND2_X1 U5213 ( .A1(n6297), .A2(n6305), .ZN(n6279) );
  NOR2_X1 U5214 ( .A1(n6283), .A2(n6279), .ZN(n6271) );
  NAND2_X1 U5215 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6271), .ZN(n5280)
         );
  NOR2_X1 U5216 ( .A1(n5280), .A2(n4242), .ZN(n4252) );
  AND2_X1 U5217 ( .A1(n4252), .A2(n4243), .ZN(n5739) );
  NAND3_X1 U5218 ( .A1(n5739), .A2(n4254), .A3(n5734), .ZN(n4244) );
  OAI21_X1 U5219 ( .B1(n6311), .B2(n6269), .A(n4244), .ZN(n4245) );
  NAND2_X1 U5220 ( .A1(n5738), .A2(n4245), .ZN(n5728) );
  NOR2_X1 U5221 ( .A1(n6270), .A2(n5718), .ZN(n4246) );
  OR2_X1 U5222 ( .A1(n5728), .A2(n4246), .ZN(n5708) );
  AOI21_X1 U5223 ( .B1(n4248), .B2(n4247), .A(n5708), .ZN(n5699) );
  NAND2_X1 U5224 ( .A1(n5699), .A2(n6270), .ZN(n5686) );
  INV_X1 U5225 ( .A(n4258), .ZN(n4249) );
  NAND3_X1 U5226 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5699), .ZN(n5685) );
  INV_X1 U5227 ( .A(n5685), .ZN(n5667) );
  NAND2_X1 U5228 ( .A1(n4249), .A2(n5667), .ZN(n4250) );
  AND2_X1 U5229 ( .A1(n5686), .A2(n4250), .ZN(n5657) );
  INV_X1 U5230 ( .A(n5657), .ZN(n4251) );
  OAI21_X1 U5231 ( .B1(n6270), .B2(n4259), .A(n4251), .ZN(n4263) );
  INV_X1 U5232 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6917) );
  NOR2_X1 U5233 ( .A1(n6232), .A2(n6917), .ZN(n4525) );
  INV_X1 U5234 ( .A(n5734), .ZN(n4255) );
  NAND2_X1 U5235 ( .A1(n6311), .A2(n4252), .ZN(n6011) );
  NAND2_X1 U5236 ( .A1(n6317), .A2(n5752), .ZN(n5778) );
  NAND2_X1 U5237 ( .A1(n6011), .A2(n5778), .ZN(n5764) );
  NAND2_X1 U5238 ( .A1(n5766), .A2(n5764), .ZN(n6019) );
  NAND3_X1 U5239 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n6004), .ZN(n5998) );
  INV_X1 U5240 ( .A(n5998), .ZN(n4253) );
  NAND2_X1 U5241 ( .A1(n4254), .A2(n4253), .ZN(n5988) );
  NOR2_X1 U5242 ( .A1(n4255), .A2(n5988), .ZN(n5716) );
  AND2_X1 U5243 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4257) );
  NAND2_X1 U5244 ( .A1(n5975), .A2(n4257), .ZN(n5669) );
  NOR2_X1 U5245 ( .A1(n5669), .A2(n4258), .ZN(n5659) );
  INV_X1 U5246 ( .A(n5659), .ZN(n4261) );
  INV_X1 U5247 ( .A(n4259), .ZN(n4260) );
  NOR3_X1 U5248 ( .A1(n4261), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n4260), 
        .ZN(n4262) );
  AOI211_X1 U5249 ( .C1(n4263), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n4525), .B(n4262), .ZN(n4264) );
  OAI22_X1 U5250 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4339), .ZN(n4381) );
  NOR2_X2 U5251 ( .A1(n5437), .A2(n4339), .ZN(n4361) );
  INV_X1 U5252 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5153) );
  NAND2_X1 U5253 ( .A1(n4361), .A2(n5153), .ZN(n4268) );
  NAND2_X1 U5254 ( .A1(n4265), .A2(n5153), .ZN(n4266) );
  OAI211_X1 U5255 ( .C1(n5437), .C2(n6313), .A(n4266), .B(n4269), .ZN(n4267)
         );
  NAND2_X1 U5256 ( .A1(n4268), .A2(n4267), .ZN(n4272) );
  INV_X1 U5257 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4271) );
  NAND2_X1 U5258 ( .A1(n5437), .A2(n4271), .ZN(n4270) );
  XNOR2_X1 U5259 ( .A(n4272), .B(n4641), .ZN(n4710) );
  NAND2_X1 U5260 ( .A1(n4710), .A2(n4672), .ZN(n4274) );
  INV_X1 U5261 ( .A(n4272), .ZN(n4273) );
  INV_X1 U5262 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5263 ( .A1(n4361), .A2(n6162), .ZN(n4277) );
  NAND2_X1 U5264 ( .A1(n4672), .A2(n6162), .ZN(n4275) );
  OAI211_X1 U5265 ( .C1(n3132), .C2(n6320), .A(n4275), .B(n4369), .ZN(n4276)
         );
  NAND2_X1 U5266 ( .A1(n4277), .A2(n4276), .ZN(n5165) );
  NAND2_X1 U5267 ( .A1(n4369), .A2(n4280), .ZN(n4282) );
  INV_X1 U5268 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4283) );
  NAND2_X1 U5269 ( .A1(n4672), .A2(n4283), .ZN(n4281) );
  NAND3_X1 U5270 ( .A1(n4282), .A2(n3128), .A3(n4281), .ZN(n4285) );
  NAND2_X1 U5271 ( .A1(n3132), .A2(n4283), .ZN(n4284) );
  AND2_X1 U5272 ( .A1(n4285), .A2(n4284), .ZN(n4705) );
  NOR2_X2 U5273 ( .A1(n5168), .A2(n4705), .ZN(n4721) );
  INV_X1 U5274 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U5275 ( .A1(n4361), .A2(n6827), .ZN(n4289) );
  NAND2_X1 U5276 ( .A1(n4672), .A2(n6827), .ZN(n4286) );
  OAI211_X1 U5277 ( .C1(n3132), .C2(n4287), .A(n4286), .B(n4369), .ZN(n4288)
         );
  AND2_X1 U5278 ( .A1(n4289), .A2(n4288), .ZN(n4720) );
  NAND2_X1 U5279 ( .A1(n4721), .A2(n4720), .ZN(n6114) );
  NAND2_X1 U5280 ( .A1(n4369), .A2(n6283), .ZN(n4291) );
  INV_X1 U5281 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U5282 ( .A1(n4672), .A2(n6158), .ZN(n4290) );
  NAND3_X1 U5283 ( .A1(n4291), .A2(n3128), .A3(n4290), .ZN(n4293) );
  NAND2_X1 U5284 ( .A1(n3132), .A2(n6158), .ZN(n4292) );
  INV_X1 U5285 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U5286 ( .A1(n4361), .A2(n6112), .ZN(n4296) );
  NAND2_X1 U5287 ( .A1(n4672), .A2(n6112), .ZN(n4294) );
  OAI211_X1 U5288 ( .C1(n3132), .C2(n6264), .A(n4294), .B(n4369), .ZN(n4295)
         );
  NAND2_X1 U5289 ( .A1(n4296), .A2(n4295), .ZN(n4744) );
  OR3_X2 U5290 ( .A1(n6114), .A2(n6113), .A3(n4744), .ZN(n4866) );
  OAI21_X1 U5291 ( .B1(n3132), .B2(n6262), .A(n4369), .ZN(n4298) );
  INV_X1 U5292 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4829) );
  NAND2_X1 U5293 ( .A1(n4672), .A2(n4829), .ZN(n4297) );
  NAND2_X1 U5294 ( .A1(n4298), .A2(n4297), .ZN(n4300) );
  NAND2_X1 U5295 ( .A1(n3132), .A2(n4829), .ZN(n4299) );
  INV_X1 U5296 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U5297 ( .A1(n4361), .A2(n6828), .ZN(n4303) );
  NAND2_X1 U5298 ( .A1(n4672), .A2(n6828), .ZN(n4301) );
  OAI211_X1 U5299 ( .C1(n3132), .C2(n6255), .A(n4301), .B(n4369), .ZN(n4302)
         );
  NAND2_X1 U5300 ( .A1(n4303), .A2(n4302), .ZN(n4864) );
  OR2_X2 U5301 ( .A1(n4866), .A2(n4304), .ZN(n5121) );
  INV_X1 U5302 ( .A(n4361), .ZN(n4365) );
  MUX2_X1 U5303 ( .A(n4365), .B(n3128), .S(EBX_REG_10__SCAN_IN), .Z(n4306) );
  NAND2_X1 U5304 ( .A1(n4642), .A2(n3635), .ZN(n4305) );
  AND2_X1 U5305 ( .A1(n4306), .A2(n4305), .ZN(n5122) );
  OAI21_X1 U5306 ( .B1(n3132), .B2(n5281), .A(n4369), .ZN(n4308) );
  INV_X1 U5307 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U5308 ( .A1(n4672), .A2(n4986), .ZN(n4307) );
  NAND2_X1 U5309 ( .A1(n4308), .A2(n4307), .ZN(n4310) );
  NAND2_X1 U5310 ( .A1(n3132), .A2(n4986), .ZN(n4309) );
  NAND2_X1 U5311 ( .A1(n4310), .A2(n4309), .ZN(n5123) );
  NAND2_X1 U5312 ( .A1(n5122), .A2(n5123), .ZN(n4311) );
  NOR2_X2 U5313 ( .A1(n5121), .A2(n4311), .ZN(n5131) );
  NAND2_X1 U5314 ( .A1(n4369), .A2(n6970), .ZN(n4313) );
  INV_X1 U5315 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U5316 ( .A1(n4672), .A2(n6949), .ZN(n4312) );
  NAND3_X1 U5317 ( .A1(n4313), .A2(n3128), .A3(n4312), .ZN(n4315) );
  NAND2_X1 U5318 ( .A1(n3132), .A2(n6949), .ZN(n4314) );
  NAND2_X1 U5319 ( .A1(n4315), .A2(n4314), .ZN(n5130) );
  NAND2_X1 U5320 ( .A1(n5131), .A2(n5130), .ZN(n5196) );
  MUX2_X1 U5321 ( .A(n4365), .B(n3128), .S(EBX_REG_12__SCAN_IN), .Z(n4317) );
  NAND2_X1 U5322 ( .A1(n4642), .A2(n5779), .ZN(n4316) );
  NAND2_X1 U5323 ( .A1(n4317), .A2(n4316), .ZN(n5195) );
  NAND2_X1 U5324 ( .A1(n4369), .A2(n4318), .ZN(n4320) );
  INV_X1 U5325 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U5326 ( .A1(n4672), .A2(n5313), .ZN(n4319) );
  NAND3_X1 U5327 ( .A1(n4320), .A2(n3128), .A3(n4319), .ZN(n4322) );
  NAND2_X1 U5328 ( .A1(n3132), .A2(n5313), .ZN(n4321) );
  NOR2_X2 U5329 ( .A1(n3127), .A2(n5301), .ZN(n5332) );
  MUX2_X1 U5330 ( .A(n4365), .B(n3128), .S(EBX_REG_14__SCAN_IN), .Z(n4325) );
  NAND2_X1 U5331 ( .A1(n4642), .A2(n4323), .ZN(n4324) );
  NAND2_X1 U5332 ( .A1(n4375), .A2(EBX_REG_15__SCAN_IN), .ZN(n4327) );
  NAND2_X1 U5333 ( .A1(n4339), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4326) );
  NAND2_X1 U5334 ( .A1(n4327), .A2(n4326), .ZN(n4328) );
  XNOR2_X1 U5335 ( .A(n4328), .B(n3128), .ZN(n5471) );
  INV_X1 U5336 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U5337 ( .A1(n4361), .A2(n5467), .ZN(n4331) );
  NAND2_X1 U5338 ( .A1(n4672), .A2(n5467), .ZN(n4329) );
  OAI211_X1 U5339 ( .C1(n3132), .C2(n6947), .A(n4329), .B(n4369), .ZN(n4330)
         );
  NAND2_X1 U5340 ( .A1(n4331), .A2(n4330), .ZN(n5460) );
  NAND2_X1 U5341 ( .A1(n4369), .A2(n5963), .ZN(n4333) );
  INV_X1 U5342 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U5343 ( .A1(n4672), .A2(n5526), .ZN(n4332) );
  NAND3_X1 U5344 ( .A1(n4333), .A2(n3128), .A3(n4332), .ZN(n4335) );
  NAND2_X1 U5345 ( .A1(n3132), .A2(n5526), .ZN(n4334) );
  INV_X1 U5346 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U5347 ( .A1(n4361), .A2(n5923), .ZN(n4338) );
  INV_X1 U5348 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6971) );
  NAND2_X1 U5349 ( .A1(n4672), .A2(n5923), .ZN(n4336) );
  OAI211_X1 U5350 ( .C1(n3132), .C2(n6971), .A(n4336), .B(n4369), .ZN(n4337)
         );
  AND2_X1 U5351 ( .A1(n4338), .A2(n4337), .ZN(n5907) );
  INV_X1 U5352 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5576) );
  NOR2_X1 U5353 ( .A1(n4339), .A2(EBX_REG_20__SCAN_IN), .ZN(n4340) );
  AOI21_X1 U5354 ( .B1(n4642), .B2(n5576), .A(n4340), .ZN(n5521) );
  OR2_X1 U5355 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4341)
         );
  INV_X1 U5356 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U5357 ( .A1(n4672), .A2(n5440), .ZN(n5438) );
  NAND2_X1 U5358 ( .A1(n4341), .A2(n5438), .ZN(n5520) );
  NAND2_X1 U5359 ( .A1(n3132), .A2(EBX_REG_20__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U5360 ( .A1(n5520), .A2(n3128), .ZN(n4342) );
  OAI211_X1 U5361 ( .C1(n5521), .C2(n5520), .A(n4343), .B(n4342), .ZN(n4344)
         );
  INV_X1 U5362 ( .A(n4344), .ZN(n4345) );
  NAND2_X1 U5363 ( .A1(n5519), .A2(n4345), .ZN(n5419) );
  INV_X1 U5364 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6778) );
  OAI21_X1 U5365 ( .B1(n3132), .B2(n6778), .A(n4369), .ZN(n4347) );
  INV_X1 U5366 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5518) );
  NAND2_X1 U5367 ( .A1(n4672), .A2(n5518), .ZN(n4346) );
  AOI22_X1 U5368 ( .A1(n4347), .A2(n4346), .B1(n3132), .B2(n5518), .ZN(n5418)
         );
  OR2_X2 U5369 ( .A1(n5419), .A2(n5418), .ZN(n5514) );
  MUX2_X1 U5370 ( .A(n4365), .B(n3128), .S(EBX_REG_22__SCAN_IN), .Z(n4348) );
  OAI21_X1 U5371 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4375), .A(n4348), 
        .ZN(n5515) );
  OR2_X2 U5372 ( .A1(n5514), .A2(n5515), .ZN(n5706) );
  MUX2_X1 U5373 ( .A(n4361), .B(n3132), .S(EBX_REG_24__SCAN_IN), .Z(n4350) );
  NOR2_X1 U5374 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4349)
         );
  NOR2_X1 U5375 ( .A1(n4350), .A2(n4349), .ZN(n5507) );
  INV_X1 U5376 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4351) );
  NAND2_X1 U5377 ( .A1(n4369), .A2(n4351), .ZN(n4353) );
  INV_X1 U5378 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U5379 ( .A1(n4672), .A2(n6717), .ZN(n4352) );
  NAND3_X1 U5380 ( .A1(n4353), .A2(n3128), .A3(n4352), .ZN(n4355) );
  NAND2_X1 U5381 ( .A1(n3132), .A2(n6717), .ZN(n4354) );
  NAND2_X1 U5382 ( .A1(n4355), .A2(n4354), .ZN(n5705) );
  NAND2_X1 U5383 ( .A1(n5507), .A2(n5705), .ZN(n4356) );
  NAND2_X1 U5384 ( .A1(n4369), .A2(n5976), .ZN(n4358) );
  INV_X1 U5385 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5501) );
  NAND2_X1 U5386 ( .A1(n4672), .A2(n5501), .ZN(n4357) );
  NAND3_X1 U5387 ( .A1(n4358), .A2(n3128), .A3(n4357), .ZN(n4360) );
  NAND2_X1 U5388 ( .A1(n3132), .A2(n5501), .ZN(n4359) );
  NAND2_X1 U5389 ( .A1(n4360), .A2(n4359), .ZN(n5404) );
  INV_X1 U5390 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U5391 ( .A1(n4361), .A2(n5863), .ZN(n4364) );
  NAND2_X1 U5392 ( .A1(n4672), .A2(n5863), .ZN(n4362) );
  OAI211_X1 U5393 ( .C1(n3132), .C2(n5977), .A(n4362), .B(n4369), .ZN(n4363)
         );
  AND2_X1 U5394 ( .A1(n4364), .A2(n4363), .ZN(n5496) );
  AND2_X2 U5395 ( .A1(n5497), .A2(n5496), .ZN(n5680) );
  MUX2_X1 U5396 ( .A(n4365), .B(n3128), .S(EBX_REG_28__SCAN_IN), .Z(n4367) );
  OR2_X1 U5397 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4366)
         );
  NAND2_X1 U5398 ( .A1(n4367), .A2(n4366), .ZN(n4481) );
  INV_X1 U5399 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4368) );
  NAND2_X1 U5400 ( .A1(n4369), .A2(n4368), .ZN(n4371) );
  INV_X1 U5401 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U5402 ( .A1(n4672), .A2(n5918), .ZN(n4370) );
  NAND3_X1 U5403 ( .A1(n4371), .A2(n3128), .A3(n4370), .ZN(n4373) );
  NAND2_X1 U5404 ( .A1(n3132), .A2(n5918), .ZN(n4372) );
  AND2_X1 U5405 ( .A1(n4373), .A2(n4372), .ZN(n5679) );
  NOR2_X1 U5406 ( .A1(n4481), .A2(n5679), .ZN(n4374) );
  OR2_X1 U5407 ( .A1(n4375), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4377)
         );
  INV_X1 U5408 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U5409 ( .A1(n4672), .A2(n5490), .ZN(n4376) );
  NAND2_X1 U5410 ( .A1(n4377), .A2(n4376), .ZN(n4462) );
  NAND2_X1 U5411 ( .A1(n4462), .A2(n3128), .ZN(n4379) );
  NAND2_X1 U5412 ( .A1(n3132), .A2(EBX_REG_29__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U5413 ( .A1(n4379), .A2(n4378), .ZN(n4391) );
  OR2_X2 U5414 ( .A1(n4483), .A2(n4391), .ZN(n4393) );
  INV_X1 U5415 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5372) );
  INV_X1 U5416 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5658) );
  OAI22_X1 U5417 ( .A1(n4642), .A2(n5372), .B1(n4672), .B2(n5658), .ZN(n4465)
         );
  NAND2_X1 U5418 ( .A1(n4483), .A2(n3128), .ZN(n4463) );
  OAI211_X2 U5419 ( .C1(n4393), .C2(n4465), .A(n4379), .B(n4463), .ZN(n4380)
         );
  XOR2_X2 U5420 ( .A(n4381), .B(n4380), .Z(n5486) );
  NAND2_X1 U5421 ( .A1(n4686), .A2(n5383), .ZN(n6607) );
  OAI21_X1 U5422 ( .B1(n4383), .B2(n4382), .A(n6607), .ZN(n4384) );
  NOR2_X1 U5423 ( .A1(n4386), .A2(n3144), .ZN(n4387) );
  OAI21_X1 U5424 ( .B1(n4388), .B2(n5992), .A(n4387), .ZN(U2987) );
  NOR2_X1 U5425 ( .A1(n5568), .A2(n4389), .ZN(n5550) );
  NOR2_X1 U5426 ( .A1(n5549), .A2(n5550), .ZN(n4390) );
  INV_X1 U5427 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6830) );
  XNOR2_X1 U5428 ( .A(n4390), .B(n6830), .ZN(n4515) );
  NAND2_X1 U5429 ( .A1(n4483), .A2(n4391), .ZN(n4392) );
  NAND2_X1 U5430 ( .A1(n4393), .A2(n4392), .ZN(n5489) );
  INV_X1 U5431 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6681) );
  OR2_X1 U5432 ( .A1(n6232), .A2(n6681), .ZN(n4507) );
  INV_X1 U5433 ( .A(n4507), .ZN(n4394) );
  AOI21_X1 U5434 ( .B1(n5659), .B2(n6830), .A(n4394), .ZN(n4395) );
  OAI21_X1 U5435 ( .B1(n5489), .B2(n6233), .A(n4395), .ZN(n4396) );
  AOI22_X1 U5436 ( .A1(n4431), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U5437 ( .A1(n4432), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4937), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4401) );
  AOI22_X1 U5438 ( .A1(n3133), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U5439 ( .A1(n3318), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4398), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4399) );
  NAND4_X1 U5440 ( .A1(n4402), .A2(n4401), .A3(n4400), .A4(n4399), .ZN(n4409)
         );
  AOI22_X1 U5441 ( .A1(n4014), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5442 ( .A1(n4425), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4406) );
  AOI22_X1 U5443 ( .A1(n4426), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U5444 ( .A1(n4435), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4404) );
  NAND4_X1 U5445 ( .A1(n4407), .A2(n4406), .A3(n4405), .A4(n4404), .ZN(n4408)
         );
  NOR2_X1 U5446 ( .A1(n4409), .A2(n4408), .ZN(n4423) );
  NAND2_X1 U5447 ( .A1(n4411), .A2(n4410), .ZN(n4422) );
  XNOR2_X1 U5448 ( .A(n4423), .B(n4422), .ZN(n4416) );
  NAND2_X1 U5449 ( .A1(n5022), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4412)
         );
  NAND2_X1 U5450 ( .A1(n4447), .A2(n4412), .ZN(n4413) );
  AOI21_X1 U5451 ( .B1(n4521), .B2(EAX_REG_29__SCAN_IN), .A(n4413), .ZN(n4414)
         );
  OAI21_X1 U5452 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n4421) );
  NAND2_X1 U5453 ( .A1(n4417), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4418)
         );
  INV_X1 U5454 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4508) );
  NAND2_X1 U5455 ( .A1(n4418), .A2(n4508), .ZN(n4419) );
  NAND2_X1 U5456 ( .A1(n4477), .A2(n4419), .ZN(n4535) );
  NOR2_X1 U5457 ( .A1(n4423), .A2(n4422), .ZN(n4443) );
  AOI22_X1 U5458 ( .A1(n3133), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4031), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U5459 ( .A1(n4425), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4424), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4429) );
  AOI22_X1 U5460 ( .A1(n4937), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4127), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4428) );
  AOI22_X1 U5461 ( .A1(n4426), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3416), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4427) );
  NAND4_X1 U5462 ( .A1(n4430), .A2(n4429), .A3(n4428), .A4(n4427), .ZN(n4441)
         );
  AOI22_X1 U5463 ( .A1(n4431), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4403), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U5464 ( .A1(n4432), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3318), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U5465 ( .A1(n4014), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4433), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U5466 ( .A1(n4435), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4436) );
  NAND4_X1 U5467 ( .A1(n4439), .A2(n4438), .A3(n4437), .A4(n4436), .ZN(n4440)
         );
  NOR2_X1 U5468 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  XNOR2_X1 U5469 ( .A(n4443), .B(n4442), .ZN(n4445) );
  NAND2_X1 U5470 ( .A1(n4445), .A2(n4444), .ZN(n4451) );
  NAND2_X1 U5471 ( .A1(n6465), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4446)
         );
  NAND2_X1 U5472 ( .A1(n4447), .A2(n4446), .ZN(n4448) );
  AOI21_X1 U5473 ( .B1(n4521), .B2(EAX_REG_30__SCAN_IN), .A(n4448), .ZN(n4450)
         );
  XNOR2_X1 U5474 ( .A(n4477), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5552)
         );
  AOI21_X1 U5475 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4516) );
  INV_X1 U5476 ( .A(n4692), .ZN(n4657) );
  NAND2_X1 U5477 ( .A1(n4920), .A2(n4657), .ZN(n4680) );
  NAND2_X1 U5478 ( .A1(n3423), .A2(n4453), .ZN(n4454) );
  OR2_X1 U5479 ( .A1(n4455), .A2(n4454), .ZN(n4659) );
  INV_X1 U5480 ( .A(n4659), .ZN(n4459) );
  INV_X1 U5481 ( .A(n4456), .ZN(n4458) );
  NAND3_X1 U5482 ( .A1(n4459), .A2(n4458), .A3(n4457), .ZN(n4460) );
  NAND2_X1 U5483 ( .A1(n4680), .A2(n4460), .ZN(n4461) );
  INV_X1 U5484 ( .A(n4462), .ZN(n4464) );
  OAI21_X1 U5485 ( .B1(n4464), .B2(n4483), .A(n4463), .ZN(n4466) );
  XNOR2_X1 U5486 ( .A(n4466), .B(n4465), .ZN(n5664) );
  INV_X1 U5487 ( .A(n5664), .ZN(n4467) );
  INV_X1 U5488 ( .A(n4470), .ZN(n4545) );
  NAND2_X1 U5489 ( .A1(n4543), .A2(n4681), .ZN(n4541) );
  NAND2_X1 U5490 ( .A1(n5351), .A2(n5022), .ZN(n6623) );
  NOR3_X1 U5491 ( .A1(n6611), .A2(n6693), .A3(n6623), .ZN(n6609) );
  AND2_X1 U5492 ( .A1(n4473), .A2(n4472), .ZN(n6619) );
  INV_X1 U5493 ( .A(n6619), .ZN(n4474) );
  NAND2_X1 U5494 ( .A1(n4474), .A2(n6232), .ZN(n4475) );
  OR2_X1 U5495 ( .A1(n6609), .A2(n4475), .ZN(n4476) );
  INV_X1 U5496 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5554) );
  INV_X1 U5497 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5385) );
  INV_X1 U5498 ( .A(n5679), .ZN(n4480) );
  NAND2_X1 U5499 ( .A1(n5680), .A2(n4480), .ZN(n4482) );
  NAND2_X1 U5500 ( .A1(n4482), .A2(n4481), .ZN(n4484) );
  NAND2_X1 U5501 ( .A1(n4484), .A2(n4483), .ZN(n5674) );
  NOR2_X1 U5502 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4497) );
  INV_X1 U5503 ( .A(n4497), .ZN(n4485) );
  AND2_X1 U5504 ( .A1(n4217), .A2(n4485), .ZN(n4498) );
  NAND3_X1 U5505 ( .A1(n4498), .A2(EBX_REG_31__SCAN_IN), .A3(n4557), .ZN(n4486) );
  INV_X1 U5506 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6676) );
  NAND3_X1 U5507 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n4493) );
  INV_X1 U5508 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6798) );
  INV_X1 U5509 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6659) );
  AND2_X1 U5510 ( .A1(n4217), .A2(n4497), .ZN(n4487) );
  AND2_X1 U5511 ( .A1(n4488), .A2(n4487), .ZN(n4489) );
  INV_X1 U5512 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4490) );
  INV_X1 U5513 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6057) );
  INV_X1 U5514 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6651) );
  INV_X1 U5515 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6934) );
  INV_X1 U5516 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6648) );
  NAND3_X1 U5517 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6130) );
  NOR3_X1 U5518 ( .A1(n6934), .A2(n6648), .A3(n6130), .ZN(n6097) );
  NAND2_X1 U5519 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6097), .ZN(n6089) );
  NOR2_X1 U5520 ( .A1(n6651), .A2(n6089), .ZN(n5268) );
  NAND2_X1 U5521 ( .A1(REIP_REG_8__SCAN_IN), .A2(n5268), .ZN(n5255) );
  NAND2_X1 U5522 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n6076) );
  NOR2_X1 U5523 ( .A1(n5255), .A2(n6076), .ZN(n6065) );
  NAND2_X1 U5524 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6065), .ZN(n6055) );
  NOR2_X1 U5525 ( .A1(n6057), .A2(n6055), .ZN(n5306) );
  NAND2_X1 U5526 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5306), .ZN(n5339) );
  NOR2_X1 U5527 ( .A1(n4490), .A2(n5339), .ZN(n5334) );
  NAND2_X1 U5528 ( .A1(n6121), .A2(n5334), .ZN(n5463) );
  NAND2_X1 U5529 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5462), .ZN(n5448) );
  NAND4_X1 U5530 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5912), .ZN(n5871) );
  NOR2_X1 U5531 ( .A1(n4493), .A2(n5871), .ZN(n5400) );
  NAND2_X1 U5532 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5400), .ZN(n5403) );
  NOR2_X1 U5533 ( .A1(n5409), .A2(n5403), .ZN(n5856) );
  NAND2_X1 U5534 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5856), .ZN(n5854) );
  OR3_X1 U5535 ( .A1(n6676), .A2(n5854), .A3(REIP_REG_28__SCAN_IN), .ZN(n4503)
         );
  NAND2_X1 U5536 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4533) );
  INV_X1 U5537 ( .A(n4533), .ZN(n4495) );
  INV_X1 U5538 ( .A(n6096), .ZN(n6131) );
  INV_X1 U5539 ( .A(n5334), .ZN(n5336) );
  NAND3_X1 U5540 ( .A1(REIP_REG_15__SCAN_IN), .A2(REIP_REG_17__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n4492) );
  NOR3_X1 U5541 ( .A1(n6131), .A2(n5336), .A3(n4492), .ZN(n5434) );
  NAND4_X1 U5542 ( .A1(n5434), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(REIP_REG_18__SCAN_IN), .ZN(n5422) );
  NOR2_X1 U5543 ( .A1(n5422), .A2(n4493), .ZN(n5399) );
  NAND4_X1 U5544 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5399), .ZN(n4494) );
  NAND2_X1 U5545 ( .A1(n6098), .A2(n6096), .ZN(n6129) );
  NAND2_X1 U5546 ( .A1(n4494), .A2(n6129), .ZN(n5857) );
  OAI21_X1 U5547 ( .B1(n6098), .B2(n4495), .A(n5857), .ZN(n5373) );
  AOI22_X1 U5548 ( .A1(n4496), .A2(n6108), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5373), .ZN(n4501) );
  NAND2_X1 U5549 ( .A1(n4673), .A2(n4497), .ZN(n6608) );
  INV_X1 U5550 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5487) );
  AOI22_X1 U5551 ( .A1(n5383), .A2(n6608), .B1(n4498), .B2(n5487), .ZN(n4499)
         );
  AOI22_X1 U5552 ( .A1(EBX_REG_28__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6142), .ZN(n4500) );
  OAI21_X1 U5553 ( .B1(n5969), .B2(n4508), .A(n4507), .ZN(n4509) );
  INV_X1 U5554 ( .A(n4509), .ZN(n4510) );
  NOR2_X1 U5555 ( .A1(n4519), .A2(n4517), .ZN(n4511) );
  OR2_X2 U5556 ( .A1(n4512), .A2(n4511), .ZN(n5534) );
  NAND2_X1 U5557 ( .A1(n4513), .A2(n6226), .ZN(n4514) );
  OAI211_X1 U5558 ( .C1(n4515), .C2(n6034), .A(n3211), .B(n4514), .ZN(U2957)
         );
  AND2_X1 U5559 ( .A1(n4517), .A2(n4516), .ZN(n4518) );
  NAND2_X1 U5560 ( .A1(n4519), .A2(n4518), .ZN(n4524) );
  AOI22_X1 U5561 ( .A1(n4521), .A2(EAX_REG_31__SCAN_IN), .B1(n4520), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4522) );
  INV_X1 U5562 ( .A(n4522), .ZN(n4523) );
  AOI21_X1 U5563 ( .B1(n6222), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4525), 
        .ZN(n4526) );
  OAI21_X1 U5564 ( .B1(n6231), .B2(n4527), .A(n4526), .ZN(n4528) );
  AOI21_X1 U5565 ( .B1(n5382), .B2(n6226), .A(n4528), .ZN(n4532) );
  NAND2_X1 U5566 ( .A1(n4530), .A2(n4529), .ZN(n4531) );
  NAND2_X1 U5567 ( .A1(n4532), .A2(n4531), .ZN(U2955) );
  NOR2_X1 U5568 ( .A1(n5854), .A2(n4533), .ZN(n5386) );
  AOI22_X1 U5569 ( .A1(EBX_REG_29__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6142), .ZN(n4534) );
  OAI21_X1 U5570 ( .B1(n4535), .B2(n6146), .A(n4534), .ZN(n4536) );
  AOI221_X1 U5571 ( .B1(n5386), .B2(n6681), .C1(n5373), .C2(
        REIP_REG_29__SCAN_IN), .A(n4536), .ZN(n4537) );
  OAI21_X1 U5572 ( .B1(n5534), .B2(n6105), .A(n4539), .ZN(U2798) );
  NAND2_X1 U5573 ( .A1(n6456), .A2(n5351), .ZN(n6029) );
  INV_X1 U5574 ( .A(n6029), .ZN(n4554) );
  AOI211_X1 U5575 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4541), .A(n4554), .B(
        n4560), .ZN(n4542) );
  INV_X1 U5576 ( .A(n4542), .ZN(U2788) );
  OAI22_X1 U5577 ( .A1(n4543), .A2(n4547), .B1(n3388), .B2(n4692), .ZN(n6027)
         );
  OR2_X1 U5578 ( .A1(n5383), .A2(n4544), .ZN(n4556) );
  AOI21_X1 U5579 ( .B1(n4556), .B2(n6632), .A(READY_N), .ZN(n6705) );
  NOR2_X1 U5580 ( .A1(n6027), .A2(n6705), .ZN(n6594) );
  NOR2_X1 U5581 ( .A1(n6594), .A2(n6617), .ZN(n6036) );
  INV_X1 U5582 ( .A(MORE_REG_SCAN_IN), .ZN(n6912) );
  NOR2_X1 U5583 ( .A1(n4546), .A2(n4545), .ZN(n4551) );
  INV_X1 U5584 ( .A(n4547), .ZN(n4548) );
  AOI21_X1 U5585 ( .B1(n4549), .B2(n4548), .A(n4692), .ZN(n4550) );
  AOI211_X1 U5586 ( .C1(n4920), .C2(n4692), .A(n4551), .B(n4550), .ZN(n6597)
         );
  INV_X1 U5587 ( .A(n6597), .ZN(n4552) );
  NAND2_X1 U5588 ( .A1(n4552), .A2(n6036), .ZN(n4553) );
  OAI21_X1 U5589 ( .B1(n6036), .B2(n6912), .A(n4553), .ZN(U3471) );
  OAI21_X1 U5590 ( .B1(n4554), .B2(READREQUEST_REG_SCAN_IN), .A(n5152), .ZN(
        n4555) );
  OAI21_X1 U5591 ( .B1(n5152), .B2(n4556), .A(n4555), .ZN(U3474) );
  INV_X1 U5592 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5593 ( .A1(n4557), .A2(n6704), .ZN(n4558) );
  NAND2_X1 U5594 ( .A1(n4637), .A2(DATAI_4_), .ZN(n4606) );
  INV_X1 U5595 ( .A(READY_N), .ZN(n6704) );
  NAND2_X1 U5596 ( .A1(n4592), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4561) );
  OAI211_X1 U5597 ( .C1(n4574), .C2(n4611), .A(n4606), .B(n4561), .ZN(U2928)
         );
  NAND2_X1 U5598 ( .A1(n4637), .A2(DATAI_3_), .ZN(n4608) );
  NAND2_X1 U5599 ( .A1(n4592), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4562) );
  OAI211_X1 U5600 ( .C1(n3991), .C2(n4611), .A(n4608), .B(n4562), .ZN(U2927)
         );
  INV_X1 U5601 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4572) );
  NAND2_X1 U5602 ( .A1(n4637), .A2(DATAI_5_), .ZN(n4604) );
  NAND2_X1 U5603 ( .A1(n4592), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4563) );
  OAI211_X1 U5604 ( .C1(n4572), .C2(n4611), .A(n4604), .B(n4563), .ZN(U2929)
         );
  INV_X1 U5605 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4581) );
  NAND2_X1 U5606 ( .A1(n4637), .A2(DATAI_8_), .ZN(n4594) );
  NAND2_X1 U5607 ( .A1(n4592), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4564) );
  OAI211_X1 U5608 ( .C1(n4581), .C2(n4611), .A(n4594), .B(n4564), .ZN(U2932)
         );
  INV_X1 U5609 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U5610 ( .A1(n4637), .A2(DATAI_7_), .ZN(n4599) );
  NAND2_X1 U5611 ( .A1(n4592), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4565) );
  OAI211_X1 U5612 ( .C1(n6899), .C2(n4611), .A(n4599), .B(n4565), .ZN(U2931)
         );
  INV_X1 U5613 ( .A(EAX_REG_22__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U5614 ( .A1(n4637), .A2(DATAI_6_), .ZN(n4616) );
  NAND2_X1 U5615 ( .A1(n4592), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4566) );
  OAI211_X1 U5616 ( .C1(n6921), .C2(n4611), .A(n4616), .B(n4566), .ZN(U2930)
         );
  INV_X1 U5617 ( .A(n6580), .ZN(n4941) );
  NAND2_X1 U5618 ( .A1(n4941), .A2(n6607), .ZN(n4569) );
  NAND2_X1 U5619 ( .A1(n6185), .A2(n4217), .ZN(n4739) );
  NAND2_X1 U5620 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4959) );
  OR2_X1 U5621 ( .A1(n4959), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6604) );
  INV_X2 U5622 ( .A(n6604), .ZN(n6195) );
  NOR2_X4 U5623 ( .A1(n6195), .A2(n6185), .ZN(n5847) );
  AOI22_X1 U5624 ( .A1(n6195), .A2(UWORD_REG_3__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4570) );
  OAI21_X1 U5625 ( .B1(n3991), .B2(n4739), .A(n4570), .ZN(U2904) );
  AOI22_X1 U5626 ( .A1(n6195), .A2(UWORD_REG_5__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5627 ( .B1(n4572), .B2(n4739), .A(n4571), .ZN(U2902) );
  AOI22_X1 U5628 ( .A1(n6195), .A2(UWORD_REG_4__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5629 ( .B1(n4574), .B2(n4739), .A(n4573), .ZN(U2903) );
  INV_X1 U5630 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4636) );
  AOI22_X1 U5631 ( .A1(n6195), .A2(UWORD_REG_2__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5632 ( .B1(n4636), .B2(n4739), .A(n4575), .ZN(U2905) );
  INV_X1 U5633 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4614) );
  AOI22_X1 U5634 ( .A1(n6195), .A2(UWORD_REG_9__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4576) );
  OAI21_X1 U5635 ( .B1(n4614), .B2(n4739), .A(n4576), .ZN(U2898) );
  INV_X1 U5636 ( .A(EAX_REG_28__SCAN_IN), .ZN(n6813) );
  AOI22_X1 U5637 ( .A1(n6195), .A2(UWORD_REG_12__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5638 ( .B1(n6813), .B2(n4739), .A(n4577), .ZN(U2895) );
  INV_X1 U5639 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4628) );
  AOI22_X1 U5640 ( .A1(n6195), .A2(UWORD_REG_13__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4578) );
  OAI21_X1 U5641 ( .B1(n4628), .B2(n4739), .A(n4578), .ZN(U2894) );
  AOI22_X1 U5642 ( .A1(n6195), .A2(UWORD_REG_6__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5643 ( .B1(n6921), .B2(n4739), .A(n4579), .ZN(U2901) );
  AOI22_X1 U5644 ( .A1(n6195), .A2(UWORD_REG_8__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4580) );
  OAI21_X1 U5645 ( .B1(n4581), .B2(n4739), .A(n4580), .ZN(U2899) );
  INV_X1 U5646 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4623) );
  AOI22_X1 U5647 ( .A1(n6195), .A2(UWORD_REG_14__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4582) );
  OAI21_X1 U5648 ( .B1(n4623), .B2(n4739), .A(n4582), .ZN(U2893) );
  XOR2_X1 U5649 ( .A(n4583), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n4649) );
  OAI21_X1 U5650 ( .B1(n4586), .B2(n4585), .A(n4584), .ZN(n5193) );
  NAND2_X1 U5651 ( .A1(n6308), .A2(REIP_REG_0__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5652 ( .B1(n5193), .B2(n5955), .A(n4645), .ZN(n4590) );
  INV_X1 U5653 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4587) );
  AOI21_X1 U5654 ( .B1(n4588), .B2(n5969), .A(n4587), .ZN(n4589) );
  AOI211_X1 U5655 ( .C1(n4529), .C2(n4649), .A(n4590), .B(n4589), .ZN(n4591)
         );
  INV_X1 U5656 ( .A(n4591), .ZN(U2986) );
  INV_X1 U5657 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U5658 ( .A1(n4638), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4593) );
  OAI211_X1 U5659 ( .C1(n6184), .C2(n4611), .A(n4594), .B(n4593), .ZN(U2947)
         );
  INV_X1 U5660 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U5661 ( .A1(n4637), .A2(DATAI_10_), .ZN(n4620) );
  NAND2_X1 U5662 ( .A1(n4638), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4595) );
  OAI211_X1 U5663 ( .C1(n6977), .C2(n4611), .A(n4620), .B(n4595), .ZN(U2934)
         );
  INV_X1 U5664 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U5665 ( .A1(n4637), .A2(DATAI_9_), .ZN(n4613) );
  NAND2_X1 U5666 ( .A1(n4638), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4596) );
  OAI211_X1 U5667 ( .C1(n6182), .C2(n4611), .A(n4613), .B(n4596), .ZN(U2948)
         );
  NAND2_X1 U5668 ( .A1(n4637), .A2(DATAI_1_), .ZN(n4631) );
  NAND2_X1 U5669 ( .A1(n4638), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4597) );
  OAI211_X1 U5670 ( .C1(n3741), .C2(n4611), .A(n4631), .B(n4597), .ZN(U2940)
         );
  INV_X1 U5671 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U5672 ( .A1(n4638), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4598) );
  OAI211_X1 U5673 ( .C1(n4830), .C2(n4611), .A(n4599), .B(n4598), .ZN(U2946)
         );
  INV_X1 U5674 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6193) );
  NAND2_X1 U5675 ( .A1(n4637), .A2(DATAI_2_), .ZN(n4635) );
  NAND2_X1 U5676 ( .A1(n4638), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4600) );
  OAI211_X1 U5677 ( .C1(n6193), .C2(n4611), .A(n4635), .B(n4600), .ZN(U2941)
         );
  INV_X1 U5678 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U5679 ( .A1(n4637), .A2(DATAI_14_), .ZN(n4622) );
  NAND2_X1 U5680 ( .A1(n4638), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4601) );
  OAI211_X1 U5681 ( .C1(n6795), .C2(n4611), .A(n4622), .B(n4601), .ZN(U2953)
         );
  INV_X1 U5682 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U5683 ( .A1(n4637), .A2(DATAI_13_), .ZN(n4627) );
  NAND2_X1 U5684 ( .A1(n4638), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4602) );
  OAI211_X1 U5685 ( .C1(n4611), .C2(n6716), .A(n4627), .B(n4602), .ZN(U2952)
         );
  NAND2_X1 U5686 ( .A1(n4638), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4603) );
  OAI211_X1 U5687 ( .C1(n4766), .C2(n4611), .A(n4604), .B(n4603), .ZN(U2944)
         );
  INV_X1 U5688 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U5689 ( .A1(n4638), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4605) );
  OAI211_X1 U5690 ( .C1(n6190), .C2(n4611), .A(n4606), .B(n4605), .ZN(U2943)
         );
  NAND2_X1 U5691 ( .A1(n4638), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4607) );
  OAI211_X1 U5692 ( .C1(n3776), .C2(n4611), .A(n4608), .B(n4607), .ZN(U2942)
         );
  NAND2_X1 U5693 ( .A1(n4637), .A2(DATAI_12_), .ZN(n4625) );
  NAND2_X1 U5694 ( .A1(n4638), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4609) );
  OAI211_X1 U5695 ( .C1(n6813), .C2(n4611), .A(n4625), .B(n4609), .ZN(U2936)
         );
  INV_X1 U5696 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4732) );
  NAND2_X1 U5697 ( .A1(n4637), .A2(DATAI_11_), .ZN(n4618) );
  NAND2_X1 U5698 ( .A1(n4638), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4610) );
  OAI211_X1 U5699 ( .C1(n4611), .C2(n4732), .A(n4618), .B(n4610), .ZN(U2935)
         );
  NAND2_X1 U5700 ( .A1(n4638), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4612) );
  OAI211_X1 U5701 ( .C1(n4614), .C2(n4611), .A(n4613), .B(n4612), .ZN(U2933)
         );
  NAND2_X1 U5702 ( .A1(n4638), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4615) );
  OAI211_X1 U5703 ( .C1(n3735), .C2(n4611), .A(n4616), .B(n4615), .ZN(U2945)
         );
  INV_X1 U5704 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U5705 ( .A1(n4638), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4617) );
  OAI211_X1 U5706 ( .C1(n6178), .C2(n4611), .A(n4618), .B(n4617), .ZN(U2950)
         );
  INV_X1 U5707 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U5708 ( .A1(n4638), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4619) );
  OAI211_X1 U5709 ( .C1(n6180), .C2(n4611), .A(n4620), .B(n4619), .ZN(U2949)
         );
  NAND2_X1 U5710 ( .A1(n4638), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4621) );
  OAI211_X1 U5711 ( .C1(n4623), .C2(n4611), .A(n4622), .B(n4621), .ZN(U2938)
         );
  INV_X1 U5712 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U5713 ( .A1(n4638), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4624) );
  OAI211_X1 U5714 ( .C1(n6176), .C2(n4611), .A(n4625), .B(n4624), .ZN(U2951)
         );
  NAND2_X1 U5715 ( .A1(n4638), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4626) );
  OAI211_X1 U5716 ( .C1(n4628), .C2(n4611), .A(n4627), .B(n4626), .ZN(U2937)
         );
  NAND2_X1 U5717 ( .A1(n4637), .A2(DATAI_0_), .ZN(n4633) );
  NAND2_X1 U5718 ( .A1(n4638), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4629) );
  OAI211_X1 U5719 ( .C1(n3748), .C2(n4611), .A(n4633), .B(n4629), .ZN(U2939)
         );
  INV_X1 U5720 ( .A(EAX_REG_17__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U5721 ( .A1(n4638), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4630) );
  OAI211_X1 U5722 ( .C1(n6766), .C2(n4611), .A(n4631), .B(n4630), .ZN(U2925)
         );
  NAND2_X1 U5723 ( .A1(n4638), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4632) );
  OAI211_X1 U5724 ( .C1(n3936), .C2(n4611), .A(n4633), .B(n4632), .ZN(U2924)
         );
  NAND2_X1 U5725 ( .A1(n4638), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4634) );
  OAI211_X1 U5726 ( .C1(n4636), .C2(n4611), .A(n4635), .B(n4634), .ZN(U2926)
         );
  INV_X1 U5727 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6172) );
  AOI22_X1 U5728 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n4638), .B1(n4637), .B2(
        DATAI_15_), .ZN(n4639) );
  OAI21_X1 U5729 ( .B1(n6172), .B2(n4611), .A(n4639), .ZN(U2954) );
  AOI21_X1 U5730 ( .B1(n4640), .B2(n5765), .A(n6306), .ZN(n4648) );
  INV_X1 U5731 ( .A(n4641), .ZN(n4644) );
  NAND2_X1 U5732 ( .A1(n4642), .A2(n6306), .ZN(n4643) );
  NAND2_X1 U5733 ( .A1(n4644), .A2(n4643), .ZN(n5186) );
  OAI211_X1 U5734 ( .C1(n6233), .C2(n5186), .A(n4646), .B(n4645), .ZN(n4647)
         );
  AOI211_X1 U5735 ( .C1(n4649), .C2(n6315), .A(n4648), .B(n4647), .ZN(n4650)
         );
  INV_X1 U5736 ( .A(n4650), .ZN(U3018) );
  NOR2_X1 U5737 ( .A1(n4653), .A2(n4652), .ZN(n4654) );
  NOR2_X1 U5738 ( .A1(n4651), .A2(n4654), .ZN(n6227) );
  INV_X1 U5739 ( .A(n6227), .ZN(n4667) );
  INV_X1 U5740 ( .A(n4655), .ZN(n4658) );
  OAI22_X1 U5741 ( .A1(n4219), .A2(n4658), .B1(n4657), .B2(n4656), .ZN(n4670)
         );
  NOR2_X1 U5742 ( .A1(n4688), .A2(n4659), .ZN(n4660) );
  NAND2_X1 U5743 ( .A1(n3363), .A2(n3389), .ZN(n4664) );
  INV_X1 U5744 ( .A(n4664), .ZN(n4665) );
  AOI22_X1 U5745 ( .A1(n5547), .A2(DATAI_2_), .B1(n6167), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4666) );
  OAI21_X1 U5746 ( .B1(n4667), .B2(n5924), .A(n4666), .ZN(U2889) );
  INV_X1 U5747 ( .A(DATAI_0_), .ZN(n4808) );
  OAI222_X1 U5748 ( .A1(n5193), .A2(n5924), .B1(n5324), .B2(n4808), .C1(n5379), 
        .C2(n3748), .ZN(U2891) );
  OAI21_X1 U5749 ( .B1(n4669), .B2(n3367), .A(n4668), .ZN(n4671) );
  OR2_X1 U5750 ( .A1(n4671), .A2(n4670), .ZN(n4678) );
  NAND2_X1 U5751 ( .A1(n6580), .A2(n4673), .ZN(n4676) );
  OAI21_X1 U5752 ( .B1(n4673), .B2(n4672), .A(n4686), .ZN(n4675) );
  NAND2_X1 U5753 ( .A1(n4692), .A2(n6704), .ZN(n4674) );
  AOI21_X1 U5754 ( .B1(n4676), .B2(n4675), .A(n4674), .ZN(n4677) );
  NOR2_X1 U5755 ( .A1(n4678), .A2(n4677), .ZN(n4679) );
  NAND2_X1 U5756 ( .A1(n4680), .A2(n4679), .ZN(n6581) );
  NAND2_X1 U5757 ( .A1(n6581), .A2(n4681), .ZN(n4684) );
  OR2_X1 U5758 ( .A1(n6611), .A2(n4959), .ZN(n6691) );
  INV_X1 U5759 ( .A(n6691), .ZN(n4682) );
  NAND2_X1 U5760 ( .A1(n4682), .A2(FLUSH_REG_SCAN_IN), .ZN(n4683) );
  NAND2_X1 U5761 ( .A1(n4684), .A2(n4683), .ZN(n6020) );
  AND2_X1 U5762 ( .A1(n6611), .A2(STATE2_REG_3__SCAN_IN), .ZN(n4685) );
  NOR2_X1 U5763 ( .A1(n6025), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4696)
         );
  INV_X1 U5764 ( .A(n3134), .ZN(n6378) );
  INV_X1 U5765 ( .A(n4686), .ZN(n4689) );
  NAND4_X1 U5766 ( .A1(n4219), .A2(n4689), .A3(n4688), .A4(n4687), .ZN(n4691)
         );
  NOR2_X1 U5767 ( .A1(n4691), .A2(n4690), .ZN(n5358) );
  OAI22_X1 U5768 ( .A1(n6378), .A2(n5358), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n5352), .ZN(n6579) );
  OAI21_X1 U5769 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6612), .A(n6025), 
        .ZN(n5363) );
  NOR2_X1 U5770 ( .A1(n5351), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4693)
         );
  AOI211_X1 U5771 ( .C1(n6579), .C2(n6022), .A(n5363), .B(n4693), .ZN(n4695)
         );
  NAND3_X1 U5772 ( .A1(n6580), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n6022), .ZN(n4694) );
  OAI21_X1 U5773 ( .B1(n4696), .B2(n4695), .A(n4694), .ZN(U3461) );
  XNOR2_X1 U5774 ( .A(n4698), .B(n4697), .ZN(n4714) );
  NOR2_X1 U5775 ( .A1(n4700), .A2(n4699), .ZN(n4701) );
  NOR2_X1 U5776 ( .A1(n3759), .A2(n4701), .ZN(n4734) );
  INV_X1 U5777 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6815) );
  NOR2_X1 U5778 ( .A1(n6232), .A2(n6815), .ZN(n4711) );
  AOI21_X1 U5779 ( .B1(n6222), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4711), 
        .ZN(n4702) );
  OAI21_X1 U5780 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6231), .A(n4702), 
        .ZN(n4703) );
  AOI21_X1 U5781 ( .B1(n4734), .B2(n6226), .A(n4703), .ZN(n4704) );
  OAI21_X1 U5782 ( .B1(n4714), .B2(n6034), .A(n4704), .ZN(U2985) );
  XOR2_X1 U5783 ( .A(n4651), .B(n4718), .Z(n6218) );
  INV_X1 U5784 ( .A(n6218), .ZN(n6148) );
  AOI21_X1 U5785 ( .B1(n4705), .B2(n5168), .A(n4721), .ZN(n6299) );
  AOI22_X1 U5786 ( .A1(n6159), .A2(n6299), .B1(EBX_REG_3__SCAN_IN), .B2(n5529), 
        .ZN(n4706) );
  OAI21_X1 U5787 ( .B1(n6148), .B2(n5531), .A(n4706), .ZN(U2856) );
  NOR2_X1 U5788 ( .A1(n4707), .A2(n6270), .ZN(n4708) );
  MUX2_X1 U5789 ( .A(n4708), .B(n5755), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4709) );
  INV_X1 U5790 ( .A(n4709), .ZN(n4713) );
  XNOR2_X1 U5791 ( .A(n4710), .B(n4672), .ZN(n5156) );
  AOI21_X1 U5792 ( .B1(n6310), .B2(n5156), .A(n4711), .ZN(n4712) );
  OAI211_X1 U5793 ( .C1(n4714), .C2(n5992), .A(n4713), .B(n4712), .ZN(U3017)
         );
  AOI21_X1 U5794 ( .B1(n4651), .B2(n4718), .A(n4717), .ZN(n4719) );
  NOR2_X1 U5795 ( .A1(n4716), .A2(n4719), .ZN(n4728) );
  INV_X1 U5796 ( .A(n4728), .ZN(n6135) );
  OAI21_X1 U5797 ( .B1(n4721), .B2(n4720), .A(n6114), .ZN(n4722) );
  INV_X1 U5798 ( .A(n4722), .ZN(n6290) );
  AOI22_X1 U5799 ( .A1(n6159), .A2(n6290), .B1(EBX_REG_4__SCAN_IN), .B2(n5529), 
        .ZN(n4723) );
  OAI21_X1 U5800 ( .B1(n6135), .B2(n5531), .A(n4723), .ZN(U2855) );
  INV_X1 U5801 ( .A(DATAI_4_), .ZN(n4886) );
  OAI222_X1 U5802 ( .A1(n6135), .A2(n5924), .B1(n5324), .B2(n4886), .C1(n5379), 
        .C2(n6190), .ZN(U2887) );
  OAI21_X1 U5803 ( .B1(n4726), .B2(n4724), .A(n4725), .ZN(n6292) );
  NOR2_X1 U5804 ( .A1(n6232), .A2(n6934), .ZN(n6289) );
  NOR2_X1 U5805 ( .A1(n5969), .A2(n3768), .ZN(n4727) );
  AOI211_X1 U5806 ( .C1(n5966), .C2(n6133), .A(n6289), .B(n4727), .ZN(n4730)
         );
  NAND2_X1 U5807 ( .A1(n4728), .A2(n6226), .ZN(n4729) );
  OAI211_X1 U5808 ( .C1(n6292), .C2(n6034), .A(n4730), .B(n4729), .ZN(U2982)
         );
  AOI22_X1 U5809 ( .A1(n6195), .A2(UWORD_REG_11__SCAN_IN), .B1(
        DATAO_REG_27__SCAN_IN), .B2(n5847), .ZN(n4731) );
  OAI21_X1 U5810 ( .B1(n4732), .B2(n4739), .A(n4731), .ZN(U2896) );
  AOI22_X1 U5811 ( .A1(n6195), .A2(UWORD_REG_10__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4733) );
  OAI21_X1 U5812 ( .B1(n6977), .B2(n4739), .A(n4733), .ZN(U2897) );
  INV_X1 U5813 ( .A(n4734), .ZN(n5163) );
  AOI22_X1 U5814 ( .A1(n6159), .A2(n5156), .B1(EBX_REG_1__SCAN_IN), .B2(n5529), 
        .ZN(n4735) );
  OAI21_X1 U5815 ( .B1(n5163), .B2(n5531), .A(n4735), .ZN(U2858) );
  AOI22_X1 U5816 ( .A1(n6195), .A2(UWORD_REG_0__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4736) );
  OAI21_X1 U5817 ( .B1(n3936), .B2(n4739), .A(n4736), .ZN(U2907) );
  AOI22_X1 U5818 ( .A1(n6195), .A2(UWORD_REG_1__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4737) );
  OAI21_X1 U5819 ( .B1(n6766), .B2(n4739), .A(n4737), .ZN(U2906) );
  AOI22_X1 U5820 ( .A1(n6195), .A2(UWORD_REG_7__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4738) );
  OAI21_X1 U5821 ( .B1(n6899), .B2(n4739), .A(n4738), .ZN(U2900) );
  AOI21_X1 U5822 ( .B1(n4716), .B2(n4740), .A(n4741), .ZN(n4743) );
  NOR2_X1 U5823 ( .A1(n4743), .A2(n4742), .ZN(n4816) );
  INV_X1 U5824 ( .A(n4816), .ZN(n6106) );
  OAI21_X1 U5825 ( .B1(n6114), .B2(n6113), .A(n4744), .ZN(n4745) );
  NAND2_X1 U5826 ( .A1(n4745), .A2(n4866), .ZN(n6102) );
  INV_X1 U5827 ( .A(n6102), .ZN(n6266) );
  AOI22_X1 U5828 ( .A1(n6159), .A2(n6266), .B1(EBX_REG_6__SCAN_IN), .B2(n5529), 
        .ZN(n4746) );
  OAI21_X1 U5829 ( .B1(n6106), .B2(n5531), .A(n4746), .ZN(U2853) );
  OAI222_X1 U5830 ( .A1(n5186), .A2(n6155), .B1(n4271), .B2(n6163), .C1(n5193), 
        .C2(n5531), .ZN(U2859) );
  INV_X1 U5831 ( .A(DATAI_6_), .ZN(n4869) );
  OAI222_X1 U5832 ( .A1(n6106), .A2(n5924), .B1(n5324), .B2(n4869), .C1(n5379), 
        .C2(n3735), .ZN(U2885) );
  INV_X1 U5833 ( .A(DATAI_1_), .ZN(n4784) );
  OAI222_X1 U5834 ( .A1(n5163), .A2(n5924), .B1(n5324), .B2(n4784), .C1(n5379), 
        .C2(n3741), .ZN(U2890) );
  INV_X1 U5835 ( .A(DATAI_3_), .ZN(n4773) );
  OAI222_X1 U5836 ( .A1(n6148), .A2(n5924), .B1(n5324), .B2(n4773), .C1(n5379), 
        .C2(n3776), .ZN(U2888) );
  NAND2_X1 U5837 ( .A1(n4749), .A2(n3134), .ZN(n5017) );
  INV_X1 U5838 ( .A(n5017), .ZN(n4990) );
  INV_X1 U5839 ( .A(n4750), .ZN(n5787) );
  INV_X1 U5840 ( .A(n5146), .ZN(n6567) );
  AOI21_X1 U5841 ( .B1(n4990), .B2(n5207), .A(n6567), .ZN(n4759) );
  OR2_X1 U5842 ( .A1(n4759), .A2(n6499), .ZN(n4753) );
  NAND2_X1 U5843 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4762), .ZN(n4752) );
  NAND2_X1 U5844 ( .A1(n4753), .A2(n4752), .ZN(n6569) );
  NOR2_X1 U5845 ( .A1(n4754), .A2(n4755), .ZN(n4989) );
  AND2_X1 U5846 ( .A1(n4989), .A2(n6372), .ZN(n4758) );
  NAND2_X1 U5847 ( .A1(n6226), .A2(DATAI_26_), .ZN(n6477) );
  NAND2_X1 U5848 ( .A1(n6226), .A2(DATAI_18_), .ZN(n6390) );
  OAI22_X1 U5849 ( .A1(n5244), .A2(n6477), .B1(n6390), .B2(n6562), .ZN(n4757)
         );
  AOI21_X1 U5850 ( .B1(n6522), .B2(n6569), .A(n4757), .ZN(n4764) );
  AND2_X1 U5851 ( .A1(n6456), .A2(n6033), .ZN(n6502) );
  INV_X1 U5852 ( .A(n6502), .ZN(n5801) );
  OAI21_X1 U5853 ( .B1(n4758), .B2(n5955), .A(n5801), .ZN(n4760) );
  NAND2_X1 U5854 ( .A1(n4760), .A2(n4759), .ZN(n4761) );
  INV_X1 U5855 ( .A(n6462), .ZN(n6376) );
  OAI211_X1 U5856 ( .C1(n6456), .C2(n4762), .A(n4761), .B(n6376), .ZN(n4822)
         );
  NAND2_X1 U5857 ( .A1(n4822), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4763)
         );
  OAI211_X1 U5858 ( .C1(n5250), .C2(n5146), .A(n4764), .B(n4763), .ZN(U3142)
         );
  INV_X1 U5859 ( .A(DATAI_5_), .ZN(n4768) );
  INV_X1 U5860 ( .A(n4740), .ZN(n4765) );
  XNOR2_X1 U5861 ( .A(n4716), .B(n4765), .ZN(n6210) );
  INV_X1 U5862 ( .A(n6210), .ZN(n4767) );
  OAI222_X1 U5863 ( .A1(n4768), .A2(n5324), .B1(n5924), .B2(n4767), .C1(n4766), 
        .C2(n5379), .ZN(U2886) );
  INV_X1 U5864 ( .A(n4780), .ZN(n4770) );
  AOI21_X1 U5865 ( .B1(n4770), .B2(n6456), .A(n6502), .ZN(n4774) );
  NOR2_X1 U5866 ( .A1(n4751), .A2(n4750), .ZN(n6500) );
  INV_X1 U5867 ( .A(n4771), .ZN(n6501) );
  AND2_X1 U5868 ( .A1(n6500), .A2(n6501), .ZN(n4901) );
  NAND3_X1 U5869 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6325), .A3(n6584), .ZN(n4898) );
  NOR2_X1 U5870 ( .A1(n6978), .A2(n4898), .ZN(n7040) );
  AOI21_X1 U5871 ( .B1(n4901), .B2(n3134), .A(n7040), .ZN(n4776) );
  OAI22_X1 U5872 ( .A1(n4774), .A2(n4776), .B1(n4898), .B2(n6465), .ZN(n4772)
         );
  INV_X1 U5873 ( .A(n4898), .ZN(n4778) );
  INV_X1 U5874 ( .A(n4774), .ZN(n4775) );
  AOI21_X1 U5875 ( .B1(n4776), .B2(n4775), .A(n6462), .ZN(n4777) );
  NAND2_X1 U5876 ( .A1(n7034), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U5877 ( .A1(n6226), .A2(DATAI_27_), .ZN(n6431) );
  NAND2_X1 U5878 ( .A1(n4780), .A2(n3745), .ZN(n7037) );
  NAND2_X1 U5879 ( .A1(n4780), .A2(n4756), .ZN(n7036) );
  NAND2_X1 U5880 ( .A1(n6226), .A2(DATAI_19_), .ZN(n6480) );
  OAI22_X1 U5881 ( .A1(n6431), .A2(n7037), .B1(n7036), .B2(n6480), .ZN(n4781)
         );
  AOI21_X1 U5882 ( .B1(n6529), .B2(n7040), .A(n4781), .ZN(n4782) );
  OAI211_X1 U5883 ( .C1(n7045), .C2(n5236), .A(n4783), .B(n4782), .ZN(U3063)
         );
  NAND2_X1 U5884 ( .A1(n7034), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4787) );
  NOR2_X1 U5885 ( .A1(n5075), .A2(n3385), .ZN(n6515) );
  NAND2_X1 U5886 ( .A1(n6226), .A2(DATAI_25_), .ZN(n6426) );
  NAND2_X1 U5887 ( .A1(n6226), .A2(DATAI_17_), .ZN(n6474) );
  OAI22_X1 U5888 ( .A1(n6426), .A2(n7037), .B1(n7036), .B2(n6474), .ZN(n4785)
         );
  AOI21_X1 U5889 ( .B1(n6515), .B2(n7040), .A(n4785), .ZN(n4786) );
  OAI211_X1 U5890 ( .C1(n7045), .C2(n5222), .A(n4787), .B(n4786), .ZN(U3061)
         );
  INV_X1 U5891 ( .A(n6522), .ZN(n5065) );
  NAND2_X1 U5892 ( .A1(n7034), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4790) );
  OAI22_X1 U5893 ( .A1(n6477), .A2(n7037), .B1(n7036), .B2(n6390), .ZN(n4788)
         );
  AOI21_X1 U5894 ( .B1(n6521), .B2(n7040), .A(n4788), .ZN(n4789) );
  OAI211_X1 U5895 ( .C1(n7045), .C2(n5065), .A(n4790), .B(n4789), .ZN(U3062)
         );
  NAND3_X1 U5896 ( .A1(n6325), .A2(n6589), .A3(n6584), .ZN(n4846) );
  NOR2_X1 U5897 ( .A1(n6978), .A2(n4846), .ZN(n4791) );
  INV_X1 U5898 ( .A(n4791), .ZN(n5112) );
  NAND2_X1 U5899 ( .A1(n5787), .A2(n4751), .ZN(n6417) );
  NOR2_X1 U5900 ( .A1(n4749), .A2(n6417), .ZN(n4852) );
  AOI21_X1 U5901 ( .B1(n4852), .B2(n3134), .A(n4791), .ZN(n4797) );
  NAND2_X1 U5902 ( .A1(n6455), .A2(n4754), .ZN(n4793) );
  INV_X1 U5903 ( .A(n4799), .ZN(n4794) );
  AOI21_X1 U5904 ( .B1(n4794), .B2(STATEBS16_REG_SCAN_IN), .A(n6499), .ZN(
        n4796) );
  AOI22_X1 U5905 ( .A1(n4797), .A2(n4796), .B1(n6499), .B2(n4846), .ZN(n4795)
         );
  NAND2_X1 U5906 ( .A1(n6376), .A2(n4795), .ZN(n5108) );
  INV_X1 U5907 ( .A(n4796), .ZN(n4798) );
  OAI22_X1 U5908 ( .A1(n4798), .A2(n4797), .B1(n5022), .B2(n4846), .ZN(n5107)
         );
  AOI22_X1 U5909 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5108), .B1(n6522), 
        .B2(n5107), .ZN(n4801) );
  INV_X1 U5910 ( .A(n6477), .ZN(n6523) );
  NOR2_X2 U5911 ( .A1(n4799), .A2(n3745), .ZN(n5840) );
  INV_X1 U5912 ( .A(n6390), .ZN(n6524) );
  AOI22_X1 U5913 ( .A1(n6523), .A2(n5109), .B1(n5840), .B2(n6524), .ZN(n4800)
         );
  OAI211_X1 U5914 ( .C1(n5250), .C2(n5112), .A(n4801), .B(n4800), .ZN(U3030)
         );
  AOI22_X1 U5915 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5108), .B1(n6514), 
        .B2(n5107), .ZN(n4803) );
  INV_X1 U5916 ( .A(n6426), .ZN(n6516) );
  INV_X1 U5917 ( .A(n6474), .ZN(n6517) );
  AOI22_X1 U5918 ( .A1(n6516), .A2(n5109), .B1(n5840), .B2(n6517), .ZN(n4802)
         );
  OAI211_X1 U5919 ( .C1(n5226), .C2(n5112), .A(n4803), .B(n4802), .ZN(U3029)
         );
  INV_X1 U5920 ( .A(DATAI_7_), .ZN(n4831) );
  AOI22_X1 U5921 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5108), .B1(n6550), 
        .B2(n5107), .ZN(n4805) );
  NAND2_X1 U5922 ( .A1(n6226), .A2(DATAI_31_), .ZN(n7038) );
  INV_X1 U5923 ( .A(n7038), .ZN(n6552) );
  NAND2_X1 U5924 ( .A1(n6226), .A2(DATAI_23_), .ZN(n7035) );
  INV_X1 U5925 ( .A(n7035), .ZN(n6555) );
  AOI22_X1 U5926 ( .A1(n6552), .A2(n5109), .B1(n5840), .B2(n6555), .ZN(n4804)
         );
  OAI211_X1 U5927 ( .C1(n5216), .C2(n5112), .A(n4805), .B(n4804), .ZN(U3035)
         );
  AOI22_X1 U5928 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5108), .B1(n6528), 
        .B2(n5107), .ZN(n4807) );
  INV_X1 U5929 ( .A(n6431), .ZN(n6530) );
  INV_X1 U5930 ( .A(n6480), .ZN(n6531) );
  AOI22_X1 U5931 ( .A1(n6530), .A2(n5109), .B1(n5840), .B2(n6531), .ZN(n4806)
         );
  OAI211_X1 U5932 ( .C1(n5242), .C2(n5112), .A(n4807), .B(n4806), .ZN(U3031)
         );
  NOR2_X2 U5933 ( .A1(n5075), .A2(n3129), .ZN(n6561) );
  INV_X1 U5934 ( .A(n6561), .ZN(n5212) );
  AOI22_X1 U5935 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5108), .B1(n6560), 
        .B2(n5107), .ZN(n4810) );
  NAND2_X1 U5936 ( .A1(n6226), .A2(DATAI_24_), .ZN(n6471) );
  INV_X1 U5937 ( .A(n6471), .ZN(n6563) );
  NAND2_X1 U5938 ( .A1(n6226), .A2(DATAI_16_), .ZN(n5810) );
  INV_X1 U5939 ( .A(n5810), .ZN(n6564) );
  AOI22_X1 U5940 ( .A1(n6563), .A2(n5109), .B1(n5840), .B2(n6564), .ZN(n4809)
         );
  OAI211_X1 U5941 ( .C1(n5212), .C2(n5112), .A(n4810), .B(n4809), .ZN(U3028)
         );
  OAI21_X1 U5942 ( .B1(n4813), .B2(n4812), .A(n4811), .ZN(n6272) );
  INV_X1 U5943 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4814) );
  NOR2_X1 U5944 ( .A1(n6232), .A2(n4814), .ZN(n6265) );
  AND2_X1 U5945 ( .A1(n6222), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n4815)
         );
  AOI211_X1 U5946 ( .C1(n5966), .C2(n6109), .A(n6265), .B(n4815), .ZN(n4818)
         );
  NAND2_X1 U5947 ( .A1(n4816), .A2(n6226), .ZN(n4817) );
  OAI211_X1 U5948 ( .C1(n6272), .C2(n6034), .A(n4818), .B(n4817), .ZN(U2980)
         );
  INV_X1 U5949 ( .A(n6560), .ZN(n5208) );
  NAND2_X1 U5950 ( .A1(n7034), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U5951 ( .A1(n6471), .A2(n7037), .B1(n7036), .B2(n5810), .ZN(n4819)
         );
  AOI21_X1 U5952 ( .B1(n6561), .B2(n7040), .A(n4819), .ZN(n4820) );
  OAI211_X1 U5953 ( .C1(n7045), .C2(n5208), .A(n4821), .B(n4820), .ZN(U3060)
         );
  INV_X1 U5954 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4826) );
  INV_X1 U5955 ( .A(n6569), .ZN(n5145) );
  OAI22_X1 U5956 ( .A1(n6562), .A2(n7035), .B1(n5145), .B2(n7044), .ZN(n4824)
         );
  NOR2_X1 U5957 ( .A1(n5216), .A2(n5146), .ZN(n4823) );
  AOI211_X1 U5958 ( .C1(n6572), .C2(n6552), .A(n4824), .B(n4823), .ZN(n4825)
         );
  OAI21_X1 U5959 ( .B1(n6577), .B2(n4826), .A(n4825), .ZN(U3147) );
  INV_X1 U5960 ( .A(n4827), .ZN(n4828) );
  XNOR2_X1 U5961 ( .A(n4742), .B(n4828), .ZN(n6202) );
  INV_X1 U5962 ( .A(n6202), .ZN(n4832) );
  XNOR2_X1 U5963 ( .A(n4866), .B(n4865), .ZN(n6256) );
  OAI222_X1 U5964 ( .A1(n5531), .A2(n4832), .B1(n4829), .B2(n6163), .C1(n6155), 
        .C2(n6256), .ZN(U2852) );
  OAI222_X1 U5965 ( .A1(n5924), .A2(n4832), .B1(n5324), .B2(n4831), .C1(n5379), 
        .C2(n4830), .ZN(U2884) );
  OR2_X1 U5966 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6381), .ZN(n5140)
         );
  NOR2_X1 U5967 ( .A1(n6371), .A2(n4756), .ZN(n4833) );
  AOI21_X1 U5968 ( .B1(n7036), .B2(n6406), .A(n6033), .ZN(n4836) );
  NAND2_X1 U5969 ( .A1(n5207), .A2(n6501), .ZN(n6379) );
  NAND2_X1 U5970 ( .A1(n6379), .A2(n6456), .ZN(n4835) );
  AND2_X1 U5971 ( .A1(n4837), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5806) );
  OAI21_X1 U5972 ( .B1(n6410), .B2(n5022), .A(n6411), .ZN(n5200) );
  AOI211_X1 U5973 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5140), .A(n5806), .B(
        n5200), .ZN(n4834) );
  OAI211_X1 U5974 ( .C1(n4836), .C2(n4835), .A(n4834), .B(n6325), .ZN(n5135)
         );
  NAND2_X1 U5975 ( .A1(n5135), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4842) );
  INV_X1 U5976 ( .A(n4749), .ZN(n6418) );
  NAND3_X1 U5977 ( .A1(n6418), .A2(n5207), .A3(n6456), .ZN(n4839) );
  NOR2_X1 U5978 ( .A1(n4837), .A2(n6465), .ZN(n6413) );
  NAND3_X1 U5979 ( .A1(n6413), .A2(n6410), .A3(n6325), .ZN(n4838) );
  OAI22_X1 U5980 ( .A1(n6406), .A2(n7035), .B1(n5041), .B2(n7044), .ZN(n4840)
         );
  AOI21_X1 U5981 ( .B1(n6552), .B2(n5043), .A(n4840), .ZN(n4841) );
  OAI211_X1 U5982 ( .C1(n5140), .C2(n5216), .A(n4842), .B(n4841), .ZN(U3075)
         );
  NAND2_X1 U5983 ( .A1(n5135), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4845) );
  INV_X1 U5984 ( .A(n5041), .ZN(n5137) );
  OAI22_X1 U5985 ( .A1(n7036), .A2(n6477), .B1(n6406), .B2(n6390), .ZN(n4843)
         );
  AOI21_X1 U5986 ( .B1(n6522), .B2(n5137), .A(n4843), .ZN(n4844) );
  OAI211_X1 U5987 ( .C1(n5140), .C2(n5250), .A(n4845), .B(n4844), .ZN(U3070)
         );
  NOR2_X1 U5988 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4846), .ZN(n5095)
         );
  INV_X1 U5989 ( .A(n6413), .ZN(n6509) );
  INV_X1 U5990 ( .A(n6409), .ZN(n4847) );
  OR2_X1 U5991 ( .A1(n6410), .A2(n4847), .ZN(n4851) );
  AOI21_X1 U5992 ( .B1(n4851), .B2(STATE2_REG_2__SCAN_IN), .A(n4957), .ZN(
        n4899) );
  OAI211_X1 U5993 ( .C1(n6693), .C2(n5095), .A(n6509), .B(n4899), .ZN(n4850)
         );
  NAND3_X1 U5994 ( .A1(n5091), .A2(n6456), .A3(n6562), .ZN(n4848) );
  AOI21_X1 U5995 ( .B1(n4848), .B2(n5801), .A(n4852), .ZN(n4849) );
  NOR2_X1 U5996 ( .A1(n5091), .A2(n6390), .ZN(n4854) );
  INV_X1 U5997 ( .A(n4851), .ZN(n4905) );
  AOI22_X1 U5998 ( .A1(n4852), .A2(n6456), .B1(n5806), .B2(n4905), .ZN(n5092)
         );
  OAI22_X1 U5999 ( .A1(n5065), .A2(n5092), .B1(n6477), .B2(n6562), .ZN(n4853)
         );
  AOI211_X1 U6000 ( .C1(n5095), .C2(n6521), .A(n4854), .B(n4853), .ZN(n4855)
         );
  OAI21_X1 U6001 ( .B1(n5098), .B2(n6787), .A(n4855), .ZN(U3022) );
  OAI22_X1 U6002 ( .A1(n6562), .A2(n7038), .B1(n5092), .B2(n7044), .ZN(n4857)
         );
  NOR2_X1 U6003 ( .A1(n5091), .A2(n7035), .ZN(n4856) );
  AOI211_X1 U6004 ( .C1(n5095), .C2(n7041), .A(n4857), .B(n4856), .ZN(n4858)
         );
  OAI21_X1 U6005 ( .B1(n5098), .B2(n4859), .A(n4858), .ZN(U3027) );
  INV_X1 U6006 ( .A(n4861), .ZN(n4862) );
  AOI21_X1 U6007 ( .B1(n4863), .B2(n4860), .A(n4862), .ZN(n5085) );
  INV_X1 U6008 ( .A(n5085), .ZN(n5276) );
  OAI21_X1 U6009 ( .B1(n4866), .B2(n4865), .A(n4864), .ZN(n4867) );
  AND2_X1 U6010 ( .A1(n5121), .A2(n4867), .ZN(n6248) );
  AOI22_X1 U6011 ( .A1(n6159), .A2(n6248), .B1(EBX_REG_8__SCAN_IN), .B2(n5529), 
        .ZN(n4868) );
  OAI21_X1 U6012 ( .B1(n5276), .B2(n5531), .A(n4868), .ZN(U2851) );
  NAND2_X1 U6013 ( .A1(n7034), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4872) );
  NAND2_X1 U6014 ( .A1(n6226), .A2(DATAI_30_), .ZN(n6491) );
  NAND2_X1 U6015 ( .A1(n6226), .A2(DATAI_22_), .ZN(n6352) );
  OAI22_X1 U6016 ( .A1(n6491), .A2(n7037), .B1(n7036), .B2(n6352), .ZN(n4870)
         );
  AOI21_X1 U6017 ( .B1(n6544), .B2(n7040), .A(n4870), .ZN(n4871) );
  OAI211_X1 U6018 ( .C1(n7045), .C2(n5217), .A(n4872), .B(n4871), .ZN(U3066)
         );
  NAND2_X1 U6019 ( .A1(n5135), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4875) );
  OAI22_X1 U6020 ( .A1(n6406), .A2(n6480), .B1(n5041), .B2(n5236), .ZN(n4873)
         );
  AOI21_X1 U6021 ( .B1(n6530), .B2(n5043), .A(n4873), .ZN(n4874) );
  OAI211_X1 U6022 ( .C1(n5140), .C2(n5242), .A(n4875), .B(n4874), .ZN(U3071)
         );
  OAI22_X1 U6023 ( .A1(n6562), .A2(n6426), .B1(n5092), .B2(n5222), .ZN(n4877)
         );
  NOR2_X1 U6024 ( .A1(n5091), .A2(n6474), .ZN(n4876) );
  AOI211_X1 U6025 ( .C1(n5095), .C2(n6515), .A(n4877), .B(n4876), .ZN(n4878)
         );
  OAI21_X1 U6026 ( .B1(n5098), .B2(n6968), .A(n4878), .ZN(U3021) );
  INV_X1 U6027 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4882) );
  OAI22_X1 U6028 ( .A1(n6562), .A2(n6431), .B1(n5092), .B2(n5236), .ZN(n4880)
         );
  NOR2_X1 U6029 ( .A1(n5091), .A2(n6480), .ZN(n4879) );
  AOI211_X1 U6030 ( .C1(n5095), .C2(n6529), .A(n4880), .B(n4879), .ZN(n4881)
         );
  OAI21_X1 U6031 ( .B1(n5098), .B2(n4882), .A(n4881), .ZN(U3023) );
  INV_X1 U6032 ( .A(DATAI_8_), .ZN(n7014) );
  OAI222_X1 U6033 ( .A1(n5276), .A2(n5924), .B1(n5324), .B2(n7014), .C1(n5379), 
        .C2(n6184), .ZN(U2883) );
  NAND2_X1 U6034 ( .A1(n5135), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U6035 ( .A1(n6406), .A2(n6474), .B1(n5041), .B2(n5222), .ZN(n4883)
         );
  AOI21_X1 U6036 ( .B1(n6516), .B2(n5043), .A(n4883), .ZN(n4884) );
  OAI211_X1 U6037 ( .C1(n5140), .C2(n5226), .A(n4885), .B(n4884), .ZN(U3069)
         );
  INV_X1 U6038 ( .A(n6535), .ZN(n5231) );
  NAND2_X1 U6039 ( .A1(n7034), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6040 ( .A1(n6226), .A2(DATAI_28_), .ZN(n6434) );
  NAND2_X1 U6041 ( .A1(n6226), .A2(DATAI_20_), .ZN(n6485) );
  OAI22_X1 U6042 ( .A1(n6434), .A2(n7037), .B1(n7036), .B2(n6485), .ZN(n4887)
         );
  AOI21_X1 U6043 ( .B1(n6536), .B2(n7040), .A(n4887), .ZN(n4888) );
  OAI211_X1 U6044 ( .C1(n7045), .C2(n5231), .A(n4889), .B(n4888), .ZN(U3064)
         );
  INV_X1 U6045 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4893) );
  OAI22_X1 U6046 ( .A1(n6562), .A2(n6474), .B1(n5145), .B2(n5222), .ZN(n4891)
         );
  NOR2_X1 U6047 ( .A1(n5226), .A2(n5146), .ZN(n4890) );
  AOI211_X1 U6048 ( .C1(n6572), .C2(n6516), .A(n4891), .B(n4890), .ZN(n4892)
         );
  OAI21_X1 U6049 ( .B1(n6577), .B2(n4893), .A(n4892), .ZN(U3141) );
  INV_X1 U6050 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4897) );
  OAI22_X1 U6051 ( .A1(n6562), .A2(n6480), .B1(n5145), .B2(n5236), .ZN(n4895)
         );
  NOR2_X1 U6052 ( .A1(n5242), .A2(n5146), .ZN(n4894) );
  AOI211_X1 U6053 ( .C1(n6572), .C2(n6530), .A(n4895), .B(n4894), .ZN(n4896)
         );
  OAI21_X1 U6054 ( .B1(n6577), .B2(n4897), .A(n4896), .ZN(U3143) );
  NOR2_X1 U6055 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4898), .ZN(n6364)
         );
  INV_X1 U6056 ( .A(n6364), .ZN(n5037) );
  INV_X1 U6057 ( .A(n5806), .ZN(n6504) );
  OAI211_X1 U6058 ( .C1(n6693), .C2(n6364), .A(n6504), .B(n4899), .ZN(n4904)
         );
  NAND2_X1 U6059 ( .A1(n4754), .A2(n6372), .ZN(n4900) );
  AOI21_X1 U6060 ( .B1(n6370), .B2(n7037), .A(n6033), .ZN(n4902) );
  NOR3_X1 U6061 ( .A1(n4902), .A2(n4901), .A3(n6499), .ZN(n4903) );
  NAND2_X1 U6062 ( .A1(n6367), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4910) );
  NAND3_X1 U6063 ( .A1(n6418), .A2(n6456), .A3(n6500), .ZN(n4907) );
  NAND2_X1 U6064 ( .A1(n4905), .A2(n6413), .ZN(n4906) );
  AND2_X1 U6065 ( .A1(n4907), .A2(n4906), .ZN(n5033) );
  OAI22_X1 U6066 ( .A1(n7037), .A2(n6480), .B1(n5033), .B2(n5236), .ZN(n4908)
         );
  AOI21_X1 U6067 ( .B1(n6530), .B2(n6353), .A(n4908), .ZN(n4909) );
  OAI211_X1 U6068 ( .C1(n5037), .C2(n5242), .A(n4910), .B(n4909), .ZN(U3055)
         );
  NAND2_X1 U6069 ( .A1(n6367), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4913) );
  OAI22_X1 U6070 ( .A1(n7037), .A2(n7035), .B1(n5033), .B2(n7044), .ZN(n4911)
         );
  AOI21_X1 U6071 ( .B1(n6552), .B2(n6353), .A(n4911), .ZN(n4912) );
  OAI211_X1 U6072 ( .C1(n5037), .C2(n5216), .A(n4913), .B(n4912), .ZN(U3059)
         );
  NAND2_X1 U6073 ( .A1(n6367), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4916) );
  OAI22_X1 U6074 ( .A1(n7037), .A2(n6474), .B1(n5033), .B2(n5222), .ZN(n4914)
         );
  AOI21_X1 U6075 ( .B1(n6516), .B2(n6353), .A(n4914), .ZN(n4915) );
  OAI211_X1 U6076 ( .C1(n5226), .C2(n5037), .A(n4916), .B(n4915), .ZN(U3053)
         );
  INV_X1 U6077 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6035) );
  NAND2_X1 U6078 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6035), .ZN(n4955) );
  INV_X1 U6079 ( .A(n4955), .ZN(n4950) );
  INV_X1 U6080 ( .A(n4917), .ZN(n5353) );
  NAND2_X1 U6081 ( .A1(n6580), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4918) );
  OAI21_X1 U6082 ( .B1(n4939), .B2(n5353), .A(n4918), .ZN(n4924) );
  NOR2_X1 U6083 ( .A1(n4920), .A2(n4919), .ZN(n4925) );
  MUX2_X1 U6084 ( .A(n4939), .B(n4925), .S(n4917), .Z(n4922) );
  NAND2_X1 U6085 ( .A1(n6580), .A2(n4921), .ZN(n5357) );
  NAND2_X1 U6086 ( .A1(n4922), .A2(n5357), .ZN(n4923) );
  MUX2_X1 U6087 ( .A(n4924), .B(n4923), .S(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .Z(n4928) );
  INV_X1 U6088 ( .A(n4925), .ZN(n4944) );
  NOR2_X1 U6089 ( .A1(n4917), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4926)
         );
  NAND2_X1 U6090 ( .A1(n4944), .A2(n4926), .ZN(n4946) );
  OAI21_X1 U6091 ( .B1(n4751), .B2(n5358), .A(n4946), .ZN(n4927) );
  NOR2_X1 U6092 ( .A1(n4928), .A2(n4927), .ZN(n5345) );
  MUX2_X1 U6093 ( .A(n3217), .B(n5345), .S(n6581), .Z(n6578) );
  INV_X1 U6094 ( .A(n5358), .ZN(n4948) );
  INV_X1 U6095 ( .A(n4933), .ZN(n4931) );
  OAI21_X1 U6096 ( .B1(n5353), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n4931), 
        .ZN(n4943) );
  NAND2_X1 U6097 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4932) );
  AOI22_X1 U6098 ( .A1(n4933), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n4932), .ZN(n4940) );
  INV_X1 U6099 ( .A(n4934), .ZN(n4936) );
  NAND2_X1 U6100 ( .A1(n5353), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6101 ( .A1(n4936), .A2(n4935), .ZN(n4938) );
  NOR2_X1 U6102 ( .A1(n4938), .A2(n4937), .ZN(n5796) );
  OAI22_X1 U6103 ( .A1(n4941), .A2(n4940), .B1(n5796), .B2(n4939), .ZN(n4942)
         );
  AOI21_X1 U6104 ( .B1(n4944), .B2(n4943), .A(n4942), .ZN(n4945) );
  OAI21_X1 U6105 ( .B1(n4946), .B2(n4929), .A(n4945), .ZN(n4947) );
  AOI21_X1 U6106 ( .B1(n4749), .B2(n4948), .A(n4947), .ZN(n5798) );
  MUX2_X1 U6107 ( .A(n4929), .B(n5798), .S(n6581), .Z(n6590) );
  NOR3_X1 U6108 ( .A1(n6578), .A2(STATE2_REG_1__SCAN_IN), .A3(n6590), .ZN(
        n4949) );
  AOI21_X1 U6109 ( .B1(n4951), .B2(n4950), .A(n4949), .ZN(n6599) );
  NOR2_X1 U6110 ( .A1(n6599), .A2(n4952), .ZN(n4960) );
  XNOR2_X1 U6111 ( .A(n4953), .B(n6024), .ZN(n6128) );
  INV_X1 U6112 ( .A(n4219), .ZN(n6021) );
  INV_X1 U6113 ( .A(n6581), .ZN(n4954) );
  AOI22_X1 U6114 ( .A1(n6128), .A2(n6021), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4954), .ZN(n4956) );
  OAI22_X1 U6115 ( .A1(n4956), .A2(STATE2_REG_1__SCAN_IN), .B1(n4955), .B2(
        n6024), .ZN(n6592) );
  NOR3_X1 U6116 ( .A1(n4960), .A2(n6592), .A3(FLUSH_REG_SCAN_IN), .ZN(n4958)
         );
  NOR3_X1 U6117 ( .A1(n4960), .A2(n4959), .A3(n6592), .ZN(n6610) );
  NOR2_X1 U6118 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5351), .ZN(n5792) );
  OAI22_X1 U6119 ( .A1(n3745), .A2(n6499), .B1(n6378), .B2(n5792), .ZN(n4961)
         );
  OAI21_X1 U6120 ( .B1(n6610), .B2(n4961), .A(n6322), .ZN(n4962) );
  OAI21_X1 U6121 ( .B1(n6322), .B2(n6978), .A(n4962), .ZN(U3465) );
  OAI22_X1 U6122 ( .A1(n6562), .A2(n6491), .B1(n5092), .B2(n5217), .ZN(n4964)
         );
  NOR2_X1 U6123 ( .A1(n5091), .A2(n6352), .ZN(n4963) );
  AOI211_X1 U6124 ( .C1(n5095), .C2(n6544), .A(n4964), .B(n4963), .ZN(n4965)
         );
  OAI21_X1 U6125 ( .B1(n5098), .B2(n6750), .A(n4965), .ZN(U3026) );
  OAI22_X1 U6126 ( .A1(n6562), .A2(n6434), .B1(n5092), .B2(n5231), .ZN(n4967)
         );
  NOR2_X1 U6127 ( .A1(n5091), .A2(n6485), .ZN(n4966) );
  AOI211_X1 U6128 ( .C1(n5095), .C2(n6536), .A(n4967), .B(n4966), .ZN(n4968)
         );
  OAI21_X1 U6129 ( .B1(n5098), .B2(n4969), .A(n4968), .ZN(U3024) );
  NAND2_X1 U6130 ( .A1(n6521), .A2(n6364), .ZN(n4971) );
  INV_X1 U6131 ( .A(n5033), .ZN(n6365) );
  INV_X1 U6132 ( .A(n7037), .ZN(n6366) );
  AOI22_X1 U6133 ( .A1(n6522), .A2(n6365), .B1(n6524), .B2(n6366), .ZN(n4970)
         );
  OAI211_X1 U6134 ( .C1(n6370), .C2(n6477), .A(n4971), .B(n4970), .ZN(n4972)
         );
  AOI21_X1 U6135 ( .B1(n6367), .B2(INSTQUEUE_REG_4__2__SCAN_IN), .A(n4972), 
        .ZN(n4973) );
  INV_X1 U6136 ( .A(n4973), .ZN(U3054) );
  OAI22_X1 U6137 ( .A1(n6562), .A2(n6471), .B1(n5092), .B2(n5208), .ZN(n4974)
         );
  AOI21_X1 U6138 ( .B1(n6564), .B2(n5109), .A(n4974), .ZN(n4976) );
  NAND2_X1 U6139 ( .A1(n6561), .A2(n5095), .ZN(n4975) );
  OAI211_X1 U6140 ( .C1(n5098), .C2(n4977), .A(n4976), .B(n4975), .ZN(U3020)
         );
  NAND2_X1 U6141 ( .A1(n5135), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4980) );
  OAI22_X1 U6142 ( .A1(n6406), .A2(n5810), .B1(n5041), .B2(n5208), .ZN(n4978)
         );
  AOI21_X1 U6143 ( .B1(n6563), .B2(n5043), .A(n4978), .ZN(n4979) );
  OAI211_X1 U6144 ( .C1(n5212), .C2(n5140), .A(n4980), .B(n4979), .ZN(U3068)
         );
  AOI21_X1 U6145 ( .B1(n4983), .B2(n4861), .A(n4982), .ZN(n4984) );
  INV_X1 U6146 ( .A(n4984), .ZN(n5260) );
  XNOR2_X1 U6147 ( .A(n5121), .B(n5123), .ZN(n6241) );
  INV_X1 U6148 ( .A(n6241), .ZN(n4985) );
  OAI222_X1 U6149 ( .A1(n5260), .A2(n5531), .B1(n4986), .B2(n6163), .C1(n6155), 
        .C2(n4985), .ZN(U2850) );
  INV_X1 U6150 ( .A(DATAI_9_), .ZN(n6996) );
  OAI222_X1 U6151 ( .A1(n5260), .A2(n5924), .B1(n5324), .B2(n6996), .C1(n5379), 
        .C2(n6182), .ZN(U2882) );
  AOI22_X1 U6152 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5108), .B1(n6543), 
        .B2(n5107), .ZN(n4988) );
  INV_X1 U6153 ( .A(n6491), .ZN(n6545) );
  INV_X1 U6154 ( .A(n6352), .ZN(n6546) );
  AOI22_X1 U6155 ( .A1(n6545), .A2(n5109), .B1(n5840), .B2(n6546), .ZN(n4987)
         );
  OAI211_X1 U6156 ( .C1(n5221), .C2(n5112), .A(n4988), .B(n4987), .ZN(U3034)
         );
  NAND3_X1 U6157 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6584), .ZN(n6498) );
  OR2_X1 U6158 ( .A1(n6978), .A2(n6498), .ZN(n5117) );
  NAND2_X1 U6159 ( .A1(n4989), .A2(n6455), .ZN(n4996) );
  INV_X1 U6160 ( .A(n4996), .ZN(n4997) );
  NAND2_X1 U6161 ( .A1(n4997), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5791) );
  NAND2_X1 U6162 ( .A1(n6456), .A2(n5791), .ZN(n4994) );
  NAND2_X1 U6163 ( .A1(n4990), .A2(n6500), .ZN(n4991) );
  AND2_X1 U6164 ( .A1(n4991), .A2(n5117), .ZN(n4995) );
  INV_X1 U6165 ( .A(n4995), .ZN(n4993) );
  AOI21_X1 U6166 ( .B1(n6499), .B2(n6498), .A(n6462), .ZN(n4992) );
  OAI21_X1 U6167 ( .B1(n4994), .B2(n4993), .A(n4992), .ZN(n5114) );
  OAI22_X1 U6168 ( .A1(n4995), .A2(n4994), .B1(n5022), .B2(n6498), .ZN(n5113)
         );
  AOI22_X1 U6169 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n5114), .B1(n6550), 
        .B2(n5113), .ZN(n4999) );
  NOR2_X2 U6170 ( .A1(n4996), .A2(n3745), .ZN(n5239) );
  AOI22_X1 U6171 ( .A1(n5239), .A2(n6555), .B1(n6554), .B2(n6552), .ZN(n4998)
         );
  OAI211_X1 U6172 ( .C1(n5216), .C2(n5117), .A(n4999), .B(n4998), .ZN(U3131)
         );
  AOI22_X1 U6173 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n5114), .B1(n6522), 
        .B2(n5113), .ZN(n5001) );
  AOI22_X1 U6174 ( .A1(n5239), .A2(n6524), .B1(n6554), .B2(n6523), .ZN(n5000)
         );
  OAI211_X1 U6175 ( .C1(n5250), .C2(n5117), .A(n5001), .B(n5000), .ZN(U3126)
         );
  AOI22_X1 U6176 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n5114), .B1(n6560), 
        .B2(n5113), .ZN(n5003) );
  AOI22_X1 U6177 ( .A1(n5239), .A2(n6564), .B1(n6554), .B2(n6563), .ZN(n5002)
         );
  OAI211_X1 U6178 ( .C1(n5212), .C2(n5117), .A(n5003), .B(n5002), .ZN(U3124)
         );
  AOI22_X1 U6179 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n5114), .B1(n6528), 
        .B2(n5113), .ZN(n5005) );
  AOI22_X1 U6180 ( .A1(n5239), .A2(n6531), .B1(n6554), .B2(n6530), .ZN(n5004)
         );
  OAI211_X1 U6181 ( .C1(n5242), .C2(n5117), .A(n5005), .B(n5004), .ZN(U3127)
         );
  AOI22_X1 U6182 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n5114), .B1(n6514), 
        .B2(n5113), .ZN(n5007) );
  AOI22_X1 U6183 ( .A1(n5239), .A2(n6517), .B1(n6554), .B2(n6516), .ZN(n5006)
         );
  OAI211_X1 U6184 ( .C1(n5226), .C2(n5117), .A(n5007), .B(n5006), .ZN(U3125)
         );
  AOI22_X1 U6185 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n5114), .B1(n6543), 
        .B2(n5113), .ZN(n5009) );
  AOI22_X1 U6186 ( .A1(n5239), .A2(n6546), .B1(n6554), .B2(n6545), .ZN(n5008)
         );
  OAI211_X1 U6187 ( .C1(n5221), .C2(n5117), .A(n5009), .B(n5008), .ZN(U3130)
         );
  INV_X1 U6188 ( .A(n6536), .ZN(n5235) );
  AOI22_X1 U6189 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5108), .B1(n6535), 
        .B2(n5107), .ZN(n5011) );
  INV_X1 U6190 ( .A(n6434), .ZN(n6537) );
  INV_X1 U6191 ( .A(n6485), .ZN(n6538) );
  AOI22_X1 U6192 ( .A1(n6537), .A2(n5109), .B1(n5840), .B2(n6538), .ZN(n5010)
         );
  OAI211_X1 U6193 ( .C1(n5235), .C2(n5112), .A(n5011), .B(n5010), .ZN(U3032)
         );
  AOI22_X1 U6194 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5114), .B1(n6535), 
        .B2(n5113), .ZN(n5013) );
  AOI22_X1 U6195 ( .A1(n5239), .A2(n6538), .B1(n6554), .B2(n6537), .ZN(n5012)
         );
  OAI211_X1 U6196 ( .C1(n5235), .C2(n5117), .A(n5013), .B(n5012), .ZN(U3128)
         );
  NAND3_X1 U6197 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6589), .A3(n6584), .ZN(n6407) );
  INV_X1 U6198 ( .A(n6407), .ZN(n5014) );
  NAND2_X1 U6199 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5014), .ZN(n5016) );
  INV_X1 U6200 ( .A(n5016), .ZN(n6448) );
  AOI22_X1 U6201 ( .A1(n6544), .A2(n6448), .B1(n6449), .B2(n6546), .ZN(n5024)
         );
  AOI21_X1 U6202 ( .B1(n5015), .B2(n6456), .A(n6502), .ZN(n5018) );
  OAI21_X1 U6203 ( .B1(n5017), .B2(n6417), .A(n5016), .ZN(n5020) );
  NOR2_X1 U6204 ( .A1(n5018), .A2(n5020), .ZN(n5019) );
  AOI211_X1 U6205 ( .C1(n6499), .C2(n6407), .A(n5019), .B(n6462), .ZN(n6453)
         );
  INV_X1 U6206 ( .A(n6453), .ZN(n5088) );
  NAND2_X1 U6207 ( .A1(n5020), .A2(n6456), .ZN(n5021) );
  OAI21_X1 U6208 ( .B1(n5022), .B2(n6407), .A(n5021), .ZN(n6450) );
  AOI22_X1 U6209 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5088), .B1(n6543), 
        .B2(n6450), .ZN(n5023) );
  OAI211_X1 U6210 ( .C1(n6491), .C2(n6415), .A(n5024), .B(n5023), .ZN(U3098)
         );
  AOI22_X1 U6211 ( .A1(n6529), .A2(n6448), .B1(n6449), .B2(n6531), .ZN(n5026)
         );
  AOI22_X1 U6212 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5088), .B1(n6528), 
        .B2(n6450), .ZN(n5025) );
  OAI211_X1 U6213 ( .C1(n6431), .C2(n6415), .A(n5026), .B(n5025), .ZN(U3095)
         );
  AOI22_X1 U6214 ( .A1(n6515), .A2(n6448), .B1(n6449), .B2(n6517), .ZN(n5028)
         );
  AOI22_X1 U6215 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5088), .B1(n6514), 
        .B2(n6450), .ZN(n5027) );
  OAI211_X1 U6216 ( .C1(n6426), .C2(n6415), .A(n5028), .B(n5027), .ZN(U3093)
         );
  AOI22_X1 U6217 ( .A1(n6521), .A2(n6448), .B1(n6449), .B2(n6524), .ZN(n5030)
         );
  AOI22_X1 U6218 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5088), .B1(n6522), 
        .B2(n6450), .ZN(n5029) );
  OAI211_X1 U6219 ( .C1(n6477), .C2(n6415), .A(n5030), .B(n5029), .ZN(U3094)
         );
  AOI22_X1 U6220 ( .A1(n7041), .A2(n6448), .B1(n6449), .B2(n6555), .ZN(n5032)
         );
  AOI22_X1 U6221 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5088), .B1(n6550), 
        .B2(n6450), .ZN(n5031) );
  OAI211_X1 U6222 ( .C1(n7038), .C2(n6415), .A(n5032), .B(n5031), .ZN(U3099)
         );
  NAND2_X1 U6223 ( .A1(n6367), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5036) );
  OAI22_X1 U6224 ( .A1(n7037), .A2(n6352), .B1(n5033), .B2(n5217), .ZN(n5034)
         );
  AOI21_X1 U6225 ( .B1(n6545), .B2(n6353), .A(n5034), .ZN(n5035) );
  OAI211_X1 U6226 ( .C1(n5037), .C2(n5221), .A(n5036), .B(n5035), .ZN(U3058)
         );
  NAND2_X1 U6227 ( .A1(n5135), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5040) );
  OAI22_X1 U6228 ( .A1(n6406), .A2(n6352), .B1(n5041), .B2(n5217), .ZN(n5038)
         );
  AOI21_X1 U6229 ( .B1(n6545), .B2(n5043), .A(n5038), .ZN(n5039) );
  OAI211_X1 U6230 ( .C1(n5140), .C2(n5221), .A(n5040), .B(n5039), .ZN(U3074)
         );
  NAND2_X1 U6231 ( .A1(n5135), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5045) );
  OAI22_X1 U6232 ( .A1(n6406), .A2(n6485), .B1(n5041), .B2(n5231), .ZN(n5042)
         );
  AOI21_X1 U6233 ( .B1(n6537), .B2(n5043), .A(n5042), .ZN(n5044) );
  OAI211_X1 U6234 ( .C1(n5140), .C2(n5235), .A(n5045), .B(n5044), .ZN(U3072)
         );
  NAND2_X1 U6235 ( .A1(n5100), .A2(n6497), .ZN(n5046) );
  AOI21_X1 U6236 ( .B1(n5046), .B2(STATEBS16_REG_SCAN_IN), .A(n6499), .ZN(
        n5051) );
  AND2_X1 U6237 ( .A1(n4750), .A2(n4751), .ZN(n5802) );
  AND2_X1 U6238 ( .A1(n5802), .A2(n4749), .ZN(n6459) );
  NAND2_X1 U6239 ( .A1(n5051), .A2(n6459), .ZN(n5048) );
  NAND3_X1 U6240 ( .A1(n5806), .A2(n6410), .A3(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5047) );
  NOR2_X1 U6241 ( .A1(n6413), .A2(n5200), .ZN(n5804) );
  INV_X1 U6242 ( .A(n6459), .ZN(n5050) );
  NAND2_X1 U6243 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5800), .ZN(n6466) );
  NOR2_X1 U6244 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6466), .ZN(n5102)
         );
  INV_X1 U6245 ( .A(n5102), .ZN(n5049) );
  AOI22_X1 U6246 ( .A1(n5051), .A2(n5050), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5049), .ZN(n5052) );
  OAI211_X1 U6247 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6465), .A(n5804), .B(n5052), .ZN(n5099) );
  NAND2_X1 U6248 ( .A1(n5099), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5055)
         );
  OAI22_X1 U6249 ( .A1(n5100), .A2(n6426), .B1(n6497), .B2(n6474), .ZN(n5053)
         );
  AOI21_X1 U6250 ( .B1(n5102), .B2(n6515), .A(n5053), .ZN(n5054) );
  OAI211_X1 U6251 ( .C1(n5106), .C2(n5222), .A(n5055), .B(n5054), .ZN(U3101)
         );
  NAND2_X1 U6252 ( .A1(n5099), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5058)
         );
  OAI22_X1 U6253 ( .A1(n5100), .A2(n6491), .B1(n6497), .B2(n6352), .ZN(n5056)
         );
  AOI21_X1 U6254 ( .B1(n5102), .B2(n6544), .A(n5056), .ZN(n5057) );
  OAI211_X1 U6255 ( .C1(n5106), .C2(n5217), .A(n5058), .B(n5057), .ZN(U3106)
         );
  NAND2_X1 U6256 ( .A1(n5099), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5061)
         );
  OAI22_X1 U6257 ( .A1(n5100), .A2(n7038), .B1(n6497), .B2(n7035), .ZN(n5059)
         );
  AOI21_X1 U6258 ( .B1(n5102), .B2(n7041), .A(n5059), .ZN(n5060) );
  OAI211_X1 U6259 ( .C1(n5106), .C2(n7044), .A(n5061), .B(n5060), .ZN(U3107)
         );
  NAND2_X1 U6260 ( .A1(n5099), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5064)
         );
  OAI22_X1 U6261 ( .A1(n5100), .A2(n6477), .B1(n6497), .B2(n6390), .ZN(n5062)
         );
  AOI21_X1 U6262 ( .B1(n5102), .B2(n6521), .A(n5062), .ZN(n5063) );
  OAI211_X1 U6263 ( .C1(n5106), .C2(n5065), .A(n5064), .B(n5063), .ZN(U3102)
         );
  NAND2_X1 U6264 ( .A1(n5099), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5068)
         );
  OAI22_X1 U6265 ( .A1(n5100), .A2(n6434), .B1(n6497), .B2(n6485), .ZN(n5066)
         );
  AOI21_X1 U6266 ( .B1(n5102), .B2(n6536), .A(n5066), .ZN(n5067) );
  OAI211_X1 U6267 ( .C1(n5106), .C2(n5231), .A(n5068), .B(n5067), .ZN(U3104)
         );
  NAND2_X1 U6268 ( .A1(n5099), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5071)
         );
  OAI22_X1 U6269 ( .A1(n5100), .A2(n6431), .B1(n6497), .B2(n6480), .ZN(n5069)
         );
  AOI21_X1 U6270 ( .B1(n5102), .B2(n6529), .A(n5069), .ZN(n5070) );
  OAI211_X1 U6271 ( .C1(n5106), .C2(n5236), .A(n5071), .B(n5070), .ZN(U3103)
         );
  NAND2_X1 U6272 ( .A1(n5099), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5074)
         );
  OAI22_X1 U6273 ( .A1(n5100), .A2(n6471), .B1(n6497), .B2(n5810), .ZN(n5072)
         );
  AOI21_X1 U6274 ( .B1(n6561), .B2(n5102), .A(n5072), .ZN(n5073) );
  OAI211_X1 U6275 ( .C1(n5106), .C2(n5208), .A(n5074), .B(n5073), .ZN(U3100)
         );
  INV_X1 U6276 ( .A(n6570), .ZN(n5105) );
  NAND2_X1 U6277 ( .A1(n7034), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5078) );
  NOR2_X2 U6278 ( .A1(n5075), .A2(n3360), .ZN(n6568) );
  NAND2_X1 U6279 ( .A1(n6226), .A2(DATAI_29_), .ZN(n6488) );
  NAND2_X1 U6280 ( .A1(n6226), .A2(DATAI_21_), .ZN(n6398) );
  OAI22_X1 U6281 ( .A1(n6488), .A2(n7037), .B1(n7036), .B2(n6398), .ZN(n5076)
         );
  AOI21_X1 U6282 ( .B1(n6568), .B2(n7040), .A(n5076), .ZN(n5077) );
  OAI211_X1 U6283 ( .C1(n7045), .C2(n5105), .A(n5078), .B(n5077), .ZN(U3065)
         );
  OAI21_X1 U6284 ( .B1(n5081), .B2(n5080), .A(n5079), .ZN(n6249) );
  INV_X1 U6285 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U6286 ( .A1(n6232), .A2(n5082), .ZN(n6247) );
  AND2_X1 U6287 ( .A1(n6222), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5083)
         );
  AOI211_X1 U6288 ( .C1(n5084), .C2(n5966), .A(n6247), .B(n5083), .ZN(n5087)
         );
  NAND2_X1 U6289 ( .A1(n5085), .A2(n6226), .ZN(n5086) );
  OAI211_X1 U6290 ( .C1(n6249), .C2(n6034), .A(n5087), .B(n5086), .ZN(U2978)
         );
  INV_X1 U6291 ( .A(n6398), .ZN(n6573) );
  AOI22_X1 U6292 ( .A1(n6568), .A2(n6448), .B1(n6449), .B2(n6573), .ZN(n5090)
         );
  AOI22_X1 U6293 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5088), .B1(n6570), 
        .B2(n6450), .ZN(n5089) );
  OAI211_X1 U6294 ( .C1(n6488), .C2(n6415), .A(n5090), .B(n5089), .ZN(U3097)
         );
  NOR2_X1 U6295 ( .A1(n5091), .A2(n6398), .ZN(n5094) );
  OAI22_X1 U6296 ( .A1(n5105), .A2(n5092), .B1(n6488), .B2(n6562), .ZN(n5093)
         );
  AOI211_X1 U6297 ( .C1(n5095), .C2(n6568), .A(n5094), .B(n5093), .ZN(n5096)
         );
  OAI21_X1 U6298 ( .B1(n5098), .B2(n5097), .A(n5096), .ZN(U3025) );
  NAND2_X1 U6299 ( .A1(n5099), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5104)
         );
  OAI22_X1 U6300 ( .A1(n5100), .A2(n6488), .B1(n6497), .B2(n6398), .ZN(n5101)
         );
  AOI21_X1 U6301 ( .B1(n5102), .B2(n6568), .A(n5101), .ZN(n5103) );
  OAI211_X1 U6302 ( .C1(n5106), .C2(n5105), .A(n5104), .B(n5103), .ZN(U3105)
         );
  INV_X1 U6303 ( .A(n6568), .ZN(n5230) );
  AOI22_X1 U6304 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5108), .B1(n6570), 
        .B2(n5107), .ZN(n5111) );
  INV_X1 U6305 ( .A(n6488), .ZN(n6571) );
  AOI22_X1 U6306 ( .A1(n6571), .A2(n5109), .B1(n5840), .B2(n6573), .ZN(n5110)
         );
  OAI211_X1 U6307 ( .C1(n5230), .C2(n5112), .A(n5111), .B(n5110), .ZN(U3033)
         );
  AOI22_X1 U6308 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n5114), .B1(n6570), 
        .B2(n5113), .ZN(n5116) );
  AOI22_X1 U6309 ( .A1(n5239), .A2(n6573), .B1(n6554), .B2(n6571), .ZN(n5115)
         );
  OAI211_X1 U6310 ( .C1(n5230), .C2(n5117), .A(n5116), .B(n5115), .ZN(U3129)
         );
  NOR2_X1 U6311 ( .A1(n4982), .A2(n5119), .ZN(n5120) );
  OR2_X1 U6312 ( .A1(n5118), .A2(n5120), .ZN(n6081) );
  INV_X1 U6313 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5126) );
  INV_X1 U6314 ( .A(n5121), .ZN(n5124) );
  AOI21_X1 U6315 ( .B1(n5124), .B2(n5123), .A(n5122), .ZN(n5125) );
  OR2_X1 U6316 ( .A1(n5125), .A2(n5131), .ZN(n6078) );
  OAI222_X1 U6317 ( .A1(n6081), .A2(n5531), .B1(n5126), .B2(n6163), .C1(n6155), 
        .C2(n6078), .ZN(U2849) );
  INV_X1 U6318 ( .A(DATAI_10_), .ZN(n6816) );
  OAI222_X1 U6319 ( .A1(n6081), .A2(n5924), .B1(n5324), .B2(n6816), .C1(n5379), 
        .C2(n6180), .ZN(U2881) );
  OR2_X1 U6320 ( .A1(n5118), .A2(n5128), .ZN(n5129) );
  NAND2_X1 U6321 ( .A1(n5127), .A2(n5129), .ZN(n6068) );
  OAI21_X1 U6322 ( .B1(n5131), .B2(n5130), .A(n5196), .ZN(n6234) );
  INV_X1 U6323 ( .A(n6234), .ZN(n5132) );
  AOI22_X1 U6324 ( .A1(n5132), .A2(n6159), .B1(EBX_REG_11__SCAN_IN), .B2(n5529), .ZN(n5133) );
  OAI21_X1 U6325 ( .B1(n6068), .B2(n5531), .A(n5133), .ZN(U2848) );
  AOI22_X1 U6326 ( .A1(n5547), .A2(DATAI_11_), .B1(n6167), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5134) );
  OAI21_X1 U6327 ( .B1(n6068), .B2(n5924), .A(n5134), .ZN(U2880) );
  NAND2_X1 U6328 ( .A1(n5135), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5139) );
  OAI22_X1 U6329 ( .A1(n7036), .A2(n6488), .B1(n6406), .B2(n6398), .ZN(n5136)
         );
  AOI21_X1 U6330 ( .B1(n6570), .B2(n5137), .A(n5136), .ZN(n5138) );
  OAI211_X1 U6331 ( .C1(n5140), .C2(n5230), .A(n5139), .B(n5138), .ZN(U3073)
         );
  INV_X1 U6332 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5144) );
  OAI22_X1 U6333 ( .A1(n6562), .A2(n6352), .B1(n5145), .B2(n5217), .ZN(n5142)
         );
  NOR2_X1 U6334 ( .A1(n5221), .A2(n5146), .ZN(n5141) );
  AOI211_X1 U6335 ( .C1(n6572), .C2(n6545), .A(n5142), .B(n5141), .ZN(n5143)
         );
  OAI21_X1 U6336 ( .B1(n6577), .B2(n5144), .A(n5143), .ZN(U3146) );
  INV_X1 U6337 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5150) );
  OAI22_X1 U6338 ( .A1(n6562), .A2(n6485), .B1(n5145), .B2(n5231), .ZN(n5148)
         );
  NOR2_X1 U6339 ( .A1(n5235), .A2(n5146), .ZN(n5147) );
  AOI211_X1 U6340 ( .C1(n6572), .C2(n6537), .A(n5148), .B(n5147), .ZN(n5149)
         );
  OAI21_X1 U6341 ( .B1(n6577), .B2(n5150), .A(n5149), .ZN(U3144) );
  INV_X1 U6342 ( .A(n3388), .ZN(n5151) );
  OAI21_X1 U6343 ( .B1(n5152), .B2(n5151), .A(n6105), .ZN(n6124) );
  INV_X1 U6344 ( .A(n6124), .ZN(n6147) );
  NOR2_X1 U6345 ( .A1(n5152), .A2(n3367), .ZN(n6127) );
  NOR2_X1 U6346 ( .A1(n6098), .A2(REIP_REG_1__SCAN_IN), .ZN(n5164) );
  INV_X1 U6347 ( .A(n5164), .ZN(n5160) );
  OAI22_X1 U6348 ( .A1(n5153), .A2(n6140), .B1(n6096), .B2(n6815), .ZN(n5154)
         );
  AOI21_X1 U6349 ( .B1(n6142), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5154), 
        .ZN(n5159) );
  NAND2_X1 U6350 ( .A1(n6108), .A2(n5155), .ZN(n5158) );
  NAND2_X1 U6351 ( .A1(n6143), .A2(n5156), .ZN(n5157) );
  NAND4_X1 U6352 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n5161)
         );
  AOI21_X1 U6353 ( .B1(n4750), .B2(n6127), .A(n5161), .ZN(n5162) );
  OAI21_X1 U6354 ( .B1(n5163), .B2(n6147), .A(n5162), .ZN(U2826) );
  NOR2_X1 U6355 ( .A1(n5164), .A2(n6131), .ZN(n6141) );
  INV_X1 U6356 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6357 ( .A1(n6227), .A2(n6124), .ZN(n5176) );
  INV_X1 U6358 ( .A(n4751), .ZN(n5174) );
  NAND2_X1 U6359 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  AND2_X1 U6360 ( .A1(n5168), .A2(n5167), .ZN(n6309) );
  AOI22_X1 U6361 ( .A1(n3126), .A2(EBX_REG_2__SCAN_IN), .B1(n6143), .B2(n6309), 
        .ZN(n5172) );
  INV_X1 U6362 ( .A(n6230), .ZN(n5169) );
  AOI22_X1 U6363 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6142), .B1(n6108), 
        .B2(n5169), .ZN(n5171) );
  NAND3_X1 U6364 ( .A1(n6121), .A2(REIP_REG_1__SCAN_IN), .A3(n5177), .ZN(n5170) );
  NAND3_X1 U6365 ( .A1(n5172), .A2(n5171), .A3(n5170), .ZN(n5173) );
  AOI21_X1 U6366 ( .B1(n5174), .B2(n6127), .A(n5173), .ZN(n5175) );
  OAI211_X1 U6367 ( .C1(n6141), .C2(n5177), .A(n5176), .B(n5175), .ZN(U2825)
         );
  NAND2_X1 U6368 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  XNOR2_X1 U6369 ( .A(n5181), .B(n5180), .ZN(n6243) );
  NAND2_X1 U6370 ( .A1(n6243), .A2(n4529), .ZN(n5185) );
  INV_X1 U6371 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5182) );
  NOR2_X1 U6372 ( .A1(n6232), .A2(n5182), .ZN(n6240) );
  NOR2_X1 U6373 ( .A1(n6231), .A2(n5254), .ZN(n5183) );
  AOI211_X1 U6374 ( .C1(n6222), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6240), 
        .B(n5183), .ZN(n5184) );
  OAI211_X1 U6375 ( .C1(n5955), .C2(n5260), .A(n5185), .B(n5184), .ZN(U2977)
         );
  INV_X1 U6376 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6377 ( .A1(n6143), .A2(n5187), .ZN(n5189) );
  OAI21_X1 U6378 ( .B1(n6142), .B2(n6108), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5188) );
  NAND2_X1 U6379 ( .A1(n5189), .A2(n5188), .ZN(n5191) );
  INV_X1 U6380 ( .A(n6129), .ZN(n5433) );
  INV_X1 U6381 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6699) );
  INV_X1 U6382 ( .A(n6127), .ZN(n6145) );
  OAI22_X1 U6383 ( .A1(n5433), .A2(n6699), .B1(n6378), .B2(n6145), .ZN(n5190)
         );
  AOI211_X1 U6384 ( .C1(EBX_REG_0__SCAN_IN), .C2(n3126), .A(n5191), .B(n5190), 
        .ZN(n5192) );
  OAI21_X1 U6385 ( .B1(n6147), .B2(n5193), .A(n5192), .ZN(U2827) );
  AOI21_X1 U6386 ( .B1(n5194), .B2(n5127), .A(n3137), .ZN(n6061) );
  INV_X1 U6387 ( .A(n6061), .ZN(n5252) );
  NAND2_X1 U6388 ( .A1(n5196), .A2(n5195), .ZN(n5197) );
  AND2_X1 U6389 ( .A1(n3127), .A2(n5197), .ZN(n6053) );
  AOI22_X1 U6390 ( .A1(n6053), .A2(n6159), .B1(EBX_REG_12__SCAN_IN), .B2(n5529), .ZN(n5198) );
  OAI21_X1 U6391 ( .B1(n5252), .B2(n5531), .A(n5198), .ZN(U2847) );
  NOR2_X1 U6392 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5199), .ZN(n5205)
         );
  INV_X1 U6393 ( .A(n5205), .ZN(n5251) );
  NOR3_X1 U6394 ( .A1(n5200), .A2(n6325), .A3(n5806), .ZN(n5204) );
  INV_X1 U6395 ( .A(n5207), .ZN(n5202) );
  OAI21_X1 U6396 ( .B1(n5239), .B2(n6572), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5201) );
  NAND3_X1 U6397 ( .A1(n5202), .A2(n6456), .A3(n5201), .ZN(n5203) );
  NAND2_X1 U6398 ( .A1(n5243), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5211)
         );
  NOR2_X1 U6399 ( .A1(n6418), .A2(n6499), .ZN(n6408) );
  NOR2_X1 U6400 ( .A1(n6509), .A2(n6325), .ZN(n5206) );
  AOI22_X1 U6401 ( .A1(n6408), .A2(n5207), .B1(n6410), .B2(n5206), .ZN(n5237)
         );
  OAI22_X1 U6402 ( .A1(n5244), .A2(n5810), .B1(n5237), .B2(n5208), .ZN(n5209)
         );
  AOI21_X1 U6403 ( .B1(n6563), .B2(n5239), .A(n5209), .ZN(n5210) );
  OAI211_X1 U6404 ( .C1(n5212), .C2(n5251), .A(n5211), .B(n5210), .ZN(U3132)
         );
  NAND2_X1 U6405 ( .A1(n5243), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5215)
         );
  OAI22_X1 U6406 ( .A1(n5244), .A2(n7035), .B1(n5237), .B2(n7044), .ZN(n5213)
         );
  AOI21_X1 U6407 ( .B1(n6552), .B2(n5239), .A(n5213), .ZN(n5214) );
  OAI211_X1 U6408 ( .C1(n5251), .C2(n5216), .A(n5215), .B(n5214), .ZN(U3139)
         );
  NAND2_X1 U6409 ( .A1(n5243), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5220)
         );
  OAI22_X1 U6410 ( .A1(n5244), .A2(n6352), .B1(n5237), .B2(n5217), .ZN(n5218)
         );
  AOI21_X1 U6411 ( .B1(n6545), .B2(n5239), .A(n5218), .ZN(n5219) );
  OAI211_X1 U6412 ( .C1(n5251), .C2(n5221), .A(n5220), .B(n5219), .ZN(U3138)
         );
  NAND2_X1 U6413 ( .A1(n5243), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5225)
         );
  OAI22_X1 U6414 ( .A1(n5244), .A2(n6474), .B1(n5237), .B2(n5222), .ZN(n5223)
         );
  AOI21_X1 U6415 ( .B1(n6516), .B2(n5239), .A(n5223), .ZN(n5224) );
  OAI211_X1 U6416 ( .C1(n5251), .C2(n5226), .A(n5225), .B(n5224), .ZN(U3133)
         );
  NAND2_X1 U6417 ( .A1(n5243), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5229)
         );
  INV_X1 U6418 ( .A(n5237), .ZN(n5247) );
  INV_X1 U6419 ( .A(n5239), .ZN(n5245) );
  OAI22_X1 U6420 ( .A1(n6488), .A2(n5245), .B1(n5244), .B2(n6398), .ZN(n5227)
         );
  AOI21_X1 U6421 ( .B1(n6570), .B2(n5247), .A(n5227), .ZN(n5228) );
  OAI211_X1 U6422 ( .C1(n5251), .C2(n5230), .A(n5229), .B(n5228), .ZN(U3137)
         );
  NAND2_X1 U6423 ( .A1(n5243), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5234)
         );
  OAI22_X1 U6424 ( .A1(n5244), .A2(n6485), .B1(n5237), .B2(n5231), .ZN(n5232)
         );
  AOI21_X1 U6425 ( .B1(n6537), .B2(n5239), .A(n5232), .ZN(n5233) );
  OAI211_X1 U6426 ( .C1(n5251), .C2(n5235), .A(n5234), .B(n5233), .ZN(U3136)
         );
  NAND2_X1 U6427 ( .A1(n5243), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5241)
         );
  OAI22_X1 U6428 ( .A1(n5244), .A2(n6480), .B1(n5237), .B2(n5236), .ZN(n5238)
         );
  AOI21_X1 U6429 ( .B1(n6530), .B2(n5239), .A(n5238), .ZN(n5240) );
  OAI211_X1 U6430 ( .C1(n5251), .C2(n5242), .A(n5241), .B(n5240), .ZN(U3135)
         );
  NAND2_X1 U6431 ( .A1(n5243), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5249)
         );
  OAI22_X1 U6432 ( .A1(n6477), .A2(n5245), .B1(n5244), .B2(n6390), .ZN(n5246)
         );
  AOI21_X1 U6433 ( .B1(n6522), .B2(n5247), .A(n5246), .ZN(n5248) );
  OAI211_X1 U6434 ( .C1(n5251), .C2(n5250), .A(n5249), .B(n5248), .ZN(U3134)
         );
  INV_X1 U6435 ( .A(DATAI_12_), .ZN(n7003) );
  OAI222_X1 U6436 ( .A1(n5252), .A2(n5924), .B1(n5324), .B2(n7003), .C1(n5379), 
        .C2(n6176), .ZN(U2879) );
  INV_X1 U6437 ( .A(n5255), .ZN(n6074) );
  NAND3_X1 U6438 ( .A1(n6121), .A2(n5182), .A3(n6074), .ZN(n5253) );
  OAI21_X1 U6439 ( .B1(n6146), .B2(n5254), .A(n5253), .ZN(n5258) );
  NAND2_X1 U6440 ( .A1(n6121), .A2(n5255), .ZN(n5271) );
  NAND2_X1 U6441 ( .A1(n6096), .A2(n5271), .ZN(n6080) );
  AOI22_X1 U6442 ( .A1(EBX_REG_9__SCAN_IN), .A2(n3126), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6080), .ZN(n5256) );
  OAI211_X1 U6443 ( .C1(n6117), .C2(n6950), .A(n5256), .B(n6232), .ZN(n5257)
         );
  AOI211_X1 U6444 ( .C1(n6143), .C2(n6241), .A(n5258), .B(n5257), .ZN(n5259)
         );
  OAI21_X1 U6445 ( .B1(n6105), .B2(n5260), .A(n5259), .ZN(U2818) );
  NAND2_X1 U6446 ( .A1(n5289), .A2(n5261), .ZN(n5263) );
  XOR2_X1 U6447 ( .A(n5263), .B(n5262), .Z(n5288) );
  INV_X1 U6448 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5264) );
  NAND2_X1 U6449 ( .A1(n6308), .A2(REIP_REG_10__SCAN_IN), .ZN(n5283) );
  OAI21_X1 U6450 ( .B1(n5969), .B2(n5264), .A(n5283), .ZN(n5266) );
  NOR2_X1 U6451 ( .A1(n6081), .A2(n5955), .ZN(n5265) );
  AOI211_X1 U6452 ( .C1(n5966), .C2(n6082), .A(n5266), .B(n5265), .ZN(n5267)
         );
  OAI21_X1 U6453 ( .B1(n5288), .B2(n6034), .A(n5267), .ZN(U2976) );
  INV_X1 U6454 ( .A(n5268), .ZN(n5270) );
  OAI22_X1 U6455 ( .A1(n5271), .A2(n5270), .B1(n6146), .B2(n5269), .ZN(n5274)
         );
  AOI22_X1 U6456 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6142), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6080), .ZN(n5272) );
  OAI211_X1 U6457 ( .C1(n6140), .C2(n6828), .A(n5272), .B(n6232), .ZN(n5273)
         );
  AOI211_X1 U6458 ( .C1(n6143), .C2(n6248), .A(n5274), .B(n5273), .ZN(n5275)
         );
  OAI21_X1 U6459 ( .B1(n6105), .B2(n5276), .A(n5275), .ZN(U2819) );
  INV_X1 U6460 ( .A(n5280), .ZN(n5277) );
  OAI21_X1 U6461 ( .B1(n5277), .B2(n6291), .A(n6267), .ZN(n5278) );
  AOI21_X1 U6462 ( .B1(n6269), .B2(n5279), .A(n5278), .ZN(n6263) );
  OAI21_X1 U6463 ( .B1(n6250), .B2(n6270), .A(n6263), .ZN(n6242) );
  AOI21_X1 U6464 ( .B1(n6317), .B2(n6284), .A(n6311), .ZN(n6288) );
  NOR2_X1 U6465 ( .A1(n6288), .A2(n5280), .ZN(n6258) );
  NAND2_X1 U6466 ( .A1(n6250), .A2(n6258), .ZN(n6246) );
  AOI221_X1 U6467 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n5281), .C2(n3635), .A(n6246), 
        .ZN(n5282) );
  AOI21_X1 U6468 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6242), .A(n5282), 
        .ZN(n5287) );
  INV_X1 U6469 ( .A(n6078), .ZN(n5285) );
  INV_X1 U6470 ( .A(n5283), .ZN(n5284) );
  AOI21_X1 U6471 ( .B1(n5285), .B2(n6310), .A(n5284), .ZN(n5286) );
  OAI211_X1 U6472 ( .C1(n5288), .C2(n5992), .A(n5287), .B(n5286), .ZN(U3008)
         );
  NAND2_X1 U6473 ( .A1(n5290), .A2(n5289), .ZN(n5292) );
  XNOR2_X1 U6474 ( .A(n5633), .B(n6970), .ZN(n5291) );
  XNOR2_X1 U6475 ( .A(n5292), .B(n5291), .ZN(n6236) );
  NAND2_X1 U6476 ( .A1(n6236), .A2(n4529), .ZN(n5297) );
  INV_X1 U6477 ( .A(n6067), .ZN(n5295) );
  INV_X1 U6478 ( .A(REIP_REG_11__SCAN_IN), .ZN(n5293) );
  OAI22_X1 U6479 ( .A1(n5969), .A2(n6746), .B1(n6232), .B2(n5293), .ZN(n5294)
         );
  AOI21_X1 U6480 ( .B1(n5966), .B2(n5295), .A(n5294), .ZN(n5296) );
  OAI211_X1 U6481 ( .C1(n5955), .C2(n6068), .A(n5297), .B(n5296), .ZN(U2975)
         );
  OAI21_X1 U6482 ( .B1(n5298), .B2(n5300), .A(n5299), .ZN(n5656) );
  AND2_X1 U6483 ( .A1(n3127), .A2(n5301), .ZN(n5302) );
  NOR2_X1 U6484 ( .A1(n5332), .A2(n5302), .ZN(n5772) );
  NOR2_X1 U6485 ( .A1(n6163), .A2(n5313), .ZN(n5303) );
  AOI21_X1 U6486 ( .B1(n5772), .B2(n6159), .A(n5303), .ZN(n5304) );
  OAI21_X1 U6487 ( .B1(n5656), .B2(n5531), .A(n5304), .ZN(U2846) );
  OAI21_X1 U6488 ( .B1(n6131), .B2(n6055), .A(n6129), .ZN(n6072) );
  INV_X1 U6489 ( .A(n6072), .ZN(n5305) );
  NOR2_X1 U6490 ( .A1(n6098), .A2(REIP_REG_12__SCAN_IN), .ZN(n6054) );
  OAI21_X1 U6491 ( .B1(n5305), .B2(n6054), .A(REIP_REG_13__SCAN_IN), .ZN(n5312) );
  INV_X1 U6492 ( .A(n5652), .ZN(n5310) );
  INV_X1 U6493 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6749) );
  NAND3_X1 U6494 ( .A1(n6121), .A2(n6749), .A3(n5306), .ZN(n5307) );
  OAI211_X1 U6495 ( .C1(n6117), .C2(n5308), .A(n6232), .B(n5307), .ZN(n5309)
         );
  AOI21_X1 U6496 ( .B1(n6108), .B2(n5310), .A(n5309), .ZN(n5311) );
  OAI211_X1 U6497 ( .C1(n5313), .C2(n6140), .A(n5312), .B(n5311), .ZN(n5314)
         );
  AOI21_X1 U6498 ( .B1(n5772), .B2(n6143), .A(n5314), .ZN(n5315) );
  OAI21_X1 U6499 ( .B1(n5656), .B2(n6105), .A(n5315), .ZN(U2814) );
  NOR2_X1 U6500 ( .A1(n5317), .A2(n3154), .ZN(n5318) );
  XNOR2_X1 U6501 ( .A(n5316), .B(n5318), .ZN(n5785) );
  INV_X1 U6502 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5320) );
  NAND2_X1 U6503 ( .A1(n5966), .A2(n6060), .ZN(n5319) );
  NAND2_X1 U6504 ( .A1(n6308), .A2(REIP_REG_12__SCAN_IN), .ZN(n5775) );
  OAI211_X1 U6505 ( .C1(n5969), .C2(n5320), .A(n5319), .B(n5775), .ZN(n5321)
         );
  AOI21_X1 U6506 ( .B1(n6061), .B2(n6226), .A(n5321), .ZN(n5322) );
  OAI21_X1 U6507 ( .B1(n5785), .B2(n6034), .A(n5322), .ZN(U2974) );
  INV_X1 U6508 ( .A(DATAI_13_), .ZN(n5323) );
  OAI222_X1 U6509 ( .A1(n5656), .A2(n5924), .B1(n5324), .B2(n5323), .C1(n6716), 
        .C2(n5379), .ZN(U2878) );
  INV_X1 U6510 ( .A(n5325), .ZN(n5329) );
  NAND3_X1 U6511 ( .A1(n5299), .A2(n5327), .A3(n5326), .ZN(n5328) );
  NAND2_X1 U6512 ( .A1(n5329), .A2(n5328), .ZN(n5649) );
  AOI22_X1 U6513 ( .A1(n5547), .A2(DATAI_14_), .B1(n6167), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5330) );
  OAI21_X1 U6514 ( .B1(n5649), .B2(n5924), .A(n5330), .ZN(U2877) );
  NOR2_X1 U6515 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  OR2_X1 U6516 ( .A1(n5472), .A2(n5333), .ZN(n5343) );
  INV_X1 U6517 ( .A(n5343), .ZN(n6009) );
  OAI21_X1 U6518 ( .B1(n6098), .B2(n5334), .A(n6096), .ZN(n5478) );
  INV_X1 U6519 ( .A(n5478), .ZN(n5335) );
  OAI22_X1 U6520 ( .A1(n5335), .A2(n4490), .B1(n5645), .B2(n6146), .ZN(n5341)
         );
  NAND2_X1 U6521 ( .A1(n6121), .A2(n5336), .ZN(n5338) );
  AOI22_X1 U6522 ( .A1(EBX_REG_14__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n6142), .ZN(n5337) );
  OAI211_X1 U6523 ( .C1(n5339), .C2(n5338), .A(n5337), .B(n6232), .ZN(n5340)
         );
  AOI211_X1 U6524 ( .C1(n6009), .C2(n6143), .A(n5341), .B(n5340), .ZN(n5342)
         );
  OAI21_X1 U6525 ( .B1(n5649), .B2(n6105), .A(n5342), .ZN(U2813) );
  INV_X1 U6526 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5344) );
  OAI222_X1 U6527 ( .A1(n5649), .A2(n5531), .B1(n5344), .B2(n6163), .C1(n6155), 
        .C2(n5343), .ZN(U2845) );
  INV_X1 U6528 ( .A(n5345), .ZN(n5348) );
  AOI22_X1 U6529 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n3189), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6313), .ZN(n5360) );
  NOR3_X1 U6530 ( .A1(n5351), .A2(n6306), .A3(n5360), .ZN(n5347) );
  NOR3_X1 U6531 ( .A1(n5353), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6612), 
        .ZN(n5346) );
  AOI211_X1 U6532 ( .C1(n5348), .C2(n6022), .A(n5347), .B(n5346), .ZN(n5350)
         );
  INV_X1 U6533 ( .A(n6025), .ZN(n5365) );
  AOI21_X1 U6534 ( .B1(n5353), .B2(n5362), .A(n5365), .ZN(n5349) );
  OAI22_X1 U6535 ( .A1(n5350), .A2(n5365), .B1(n5349), .B2(n3217), .ZN(U3459)
         );
  NOR2_X1 U6536 ( .A1(n5351), .A2(n6306), .ZN(n5359) );
  INV_X1 U6537 ( .A(n5352), .ZN(n5355) );
  INV_X1 U6538 ( .A(n4952), .ZN(n5354) );
  NAND3_X1 U6539 ( .A1(n5355), .A2(n5354), .A3(n5353), .ZN(n5356) );
  OAI211_X1 U6540 ( .C1(n5787), .C2(n5358), .A(n5357), .B(n5356), .ZN(n6582)
         );
  AOI222_X1 U6541 ( .A1(n5362), .A2(n5361), .B1(n5360), .B2(n5359), .C1(n6582), 
        .C2(n6022), .ZN(n5366) );
  INV_X1 U6542 ( .A(n5363), .ZN(n5364) );
  OAI22_X1 U6543 ( .A1(n5366), .A2(n5365), .B1(n4921), .B2(n5364), .ZN(U3460)
         );
  AOI22_X1 U6544 ( .A1(n6164), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6167), .ZN(n5370) );
  AND2_X1 U6545 ( .A1(n3360), .A2(n3389), .ZN(n5368) );
  NAND2_X1 U6546 ( .A1(n6168), .A2(DATAI_14_), .ZN(n5369) );
  OAI211_X1 U6547 ( .C1(n5378), .C2(n5924), .A(n5370), .B(n5369), .ZN(U2861)
         );
  AOI22_X1 U6548 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6142), .B1(n6108), 
        .B2(n5552), .ZN(n5371) );
  OAI21_X1 U6549 ( .B1(n6140), .B2(n5372), .A(n5371), .ZN(n5376) );
  NAND2_X1 U6550 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5387) );
  AOI21_X1 U6551 ( .B1(n5386), .B2(n5387), .A(n5373), .ZN(n5393) );
  AOI21_X1 U6552 ( .B1(n5386), .B2(REIP_REG_29__SCAN_IN), .A(
        REIP_REG_30__SCAN_IN), .ZN(n5374) );
  NOR2_X1 U6553 ( .A1(n5393), .A2(n5374), .ZN(n5375) );
  AOI211_X1 U6554 ( .C1(n6143), .C2(n5664), .A(n5376), .B(n5375), .ZN(n5377)
         );
  OAI21_X1 U6555 ( .B1(n5378), .B2(n6105), .A(n5377), .ZN(U2797) );
  NAND3_X1 U6556 ( .A1(n5382), .A2(n4453), .A3(n5379), .ZN(n5381) );
  AOI22_X1 U6557 ( .A1(n6164), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6167), .ZN(n5380) );
  NAND2_X1 U6558 ( .A1(n5381), .A2(n5380), .ZN(U2860) );
  NAND2_X1 U6559 ( .A1(n5382), .A2(n6094), .ZN(n5392) );
  NAND4_X1 U6560 ( .A1(n6702), .A2(n5383), .A3(EBX_REG_31__SCAN_IN), .A4(n6608), .ZN(n5384) );
  OAI21_X1 U6561 ( .B1(n6117), .B2(n5385), .A(n5384), .ZN(n5390) );
  INV_X1 U6562 ( .A(n5386), .ZN(n5388) );
  NOR3_X1 U6563 ( .A1(n5388), .A2(REIP_REG_31__SCAN_IN), .A3(n5387), .ZN(n5389) );
  AOI211_X1 U6564 ( .C1(n5486), .C2(n6143), .A(n5390), .B(n5389), .ZN(n5391)
         );
  OAI211_X1 U6565 ( .C1(n5393), .C2(n6917), .A(n5392), .B(n5391), .ZN(U2796)
         );
  NAND2_X1 U6567 ( .A1(n5396), .A2(n5397), .ZN(n5398) );
  AND2_X1 U6568 ( .A1(n5394), .A2(n5398), .ZN(n5947) );
  INV_X1 U6569 ( .A(n5947), .ZN(n5413) );
  NOR2_X1 U6570 ( .A1(n5433), .A2(n5399), .ZN(n5872) );
  INV_X1 U6571 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6572 ( .A1(n5401), .A2(n5400), .ZN(n5867) );
  INV_X1 U6573 ( .A(n5867), .ZN(n5402) );
  OAI21_X1 U6574 ( .B1(n5872), .B2(n5402), .A(REIP_REG_25__SCAN_IN), .ZN(n5412) );
  INV_X1 U6575 ( .A(n5403), .ZN(n5410) );
  INV_X1 U6576 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5409) );
  NOR2_X1 U6577 ( .A1(n5508), .A2(n5404), .ZN(n5405) );
  OR2_X1 U6578 ( .A1(n5497), .A2(n5405), .ZN(n5693) );
  OAI22_X1 U6579 ( .A1(n4114), .A2(n6117), .B1(n6146), .B2(n5950), .ZN(n5406)
         );
  AOI21_X1 U6580 ( .B1(n3126), .B2(EBX_REG_25__SCAN_IN), .A(n5406), .ZN(n5407)
         );
  OAI21_X1 U6581 ( .B1(n5693), .B2(n6115), .A(n5407), .ZN(n5408) );
  AOI21_X1 U6582 ( .B1(n5410), .B2(n5409), .A(n5408), .ZN(n5411) );
  OAI211_X1 U6583 ( .C1(n5413), .C2(n6105), .A(n5412), .B(n5411), .ZN(U2802)
         );
  NAND2_X1 U6584 ( .A1(n5415), .A2(n5416), .ZN(n5417) );
  NAND2_X1 U6585 ( .A1(n5414), .A2(n5417), .ZN(n5939) );
  NAND2_X1 U6586 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  NAND2_X1 U6587 ( .A1(n5514), .A2(n5420), .ZN(n5731) );
  INV_X1 U6588 ( .A(n5731), .ZN(n5425) );
  AOI22_X1 U6589 ( .A1(EBX_REG_21__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6142), .ZN(n5421) );
  OAI21_X1 U6590 ( .B1(n6146), .B2(n5607), .A(n5421), .ZN(n5424) );
  AND2_X1 U6591 ( .A1(n6129), .A2(n5422), .ZN(n5894) );
  AND2_X1 U6592 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5894), .ZN(n5423) );
  AOI211_X1 U6593 ( .C1(n6143), .C2(n5425), .A(n5424), .B(n5423), .ZN(n5427)
         );
  NOR2_X1 U6594 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5871), .ZN(n5883) );
  INV_X1 U6595 ( .A(n5883), .ZN(n5426) );
  OAI211_X1 U6596 ( .C1(n5939), .C2(n6105), .A(n5427), .B(n5426), .ZN(U2806)
         );
  INV_X1 U6597 ( .A(n5912), .ZN(n5889) );
  INV_X1 U6598 ( .A(n5428), .ZN(n5431) );
  OAI21_X1 U6599 ( .B1(n5431), .B2(n3155), .A(n5430), .ZN(n5624) );
  INV_X1 U6600 ( .A(n5624), .ZN(n5432) );
  NAND2_X1 U6601 ( .A1(n5432), .A2(n6094), .ZN(n5444) );
  NOR2_X1 U6602 ( .A1(n5434), .A2(n5433), .ZN(n5901) );
  AOI22_X1 U6603 ( .A1(n5622), .A2(n6108), .B1(REIP_REG_18__SCAN_IN), .B2(
        n5901), .ZN(n5435) );
  OAI211_X1 U6604 ( .C1(n6117), .C2(n5436), .A(n5435), .B(n6232), .ZN(n5442)
         );
  MUX2_X1 U6605 ( .A(n5520), .B(n5438), .S(n3132), .Z(n5439) );
  INV_X1 U6606 ( .A(n5439), .ZN(n5905) );
  XNOR2_X1 U6607 ( .A(n5906), .B(n5905), .ZN(n5750) );
  OAI22_X1 U6608 ( .A1(n5750), .A2(n6115), .B1(n5440), .B2(n6140), .ZN(n5441)
         );
  NOR2_X1 U6609 ( .A1(n5442), .A2(n5441), .ZN(n5443) );
  OAI211_X1 U6610 ( .C1(REIP_REG_18__SCAN_IN), .C2(n5889), .A(n5444), .B(n5443), .ZN(U2809) );
  NAND2_X1 U6611 ( .A1(n5445), .A2(n5446), .ZN(n5447) );
  AND2_X1 U6612 ( .A1(n5428), .A2(n5447), .ZN(n6166) );
  INV_X1 U6613 ( .A(n6166), .ZN(n5456) );
  NAND2_X1 U6614 ( .A1(n6798), .A2(n5448), .ZN(n5454) );
  AND2_X1 U6615 ( .A1(n5458), .A2(n5449), .ZN(n5450) );
  OR2_X1 U6616 ( .A1(n5450), .A2(n5906), .ZN(n5991) );
  AOI21_X1 U6617 ( .B1(n3126), .B2(EBX_REG_17__SCAN_IN), .A(n6308), .ZN(n5451)
         );
  OAI21_X1 U6618 ( .B1(n5991), .B2(n6115), .A(n5451), .ZN(n5453) );
  INV_X1 U6619 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6900) );
  OAI22_X1 U6620 ( .A1(n6900), .A2(n6117), .B1(n5965), .B2(n6146), .ZN(n5452)
         );
  AOI211_X1 U6621 ( .C1(n5454), .C2(n5901), .A(n5453), .B(n5452), .ZN(n5455)
         );
  OAI21_X1 U6622 ( .B1(n5456), .B2(n6105), .A(n5455), .ZN(U2810) );
  OAI21_X1 U6623 ( .B1(n3149), .B2(n5457), .A(n5445), .ZN(n5631) );
  INV_X1 U6624 ( .A(n5458), .ZN(n5459) );
  AOI21_X1 U6625 ( .B1(n5460), .B2(n5474), .A(n5459), .ZN(n6000) );
  AOI21_X1 U6626 ( .B1(n6142), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6308), 
        .ZN(n5461) );
  OAI21_X1 U6627 ( .B1(n5627), .B2(n6146), .A(n5461), .ZN(n5469) );
  INV_X1 U6628 ( .A(n5462), .ZN(n5465) );
  NOR2_X1 U6629 ( .A1(n5463), .A2(REIP_REG_15__SCAN_IN), .ZN(n5483) );
  NOR2_X1 U6630 ( .A1(n5483), .A2(n5478), .ZN(n5464) );
  MUX2_X1 U6631 ( .A(n5465), .B(n5464), .S(REIP_REG_16__SCAN_IN), .Z(n5466) );
  OAI21_X1 U6632 ( .B1(n5467), .B2(n6140), .A(n5466), .ZN(n5468) );
  AOI211_X1 U6633 ( .C1(n6000), .C2(n6143), .A(n5469), .B(n5468), .ZN(n5470)
         );
  OAI21_X1 U6634 ( .B1(n5631), .B2(n6105), .A(n5470), .ZN(U2811) );
  OR2_X1 U6635 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U6636 ( .A1(n5474), .A2(n5473), .ZN(n5757) );
  NOR2_X1 U6637 ( .A1(n5325), .A2(n5475), .ZN(n5476) );
  OR2_X1 U6638 ( .A1(n3149), .A2(n5476), .ZN(n5637) );
  INV_X1 U6639 ( .A(n5637), .ZN(n5477) );
  NAND2_X1 U6640 ( .A1(n5477), .A2(n6094), .ZN(n5485) );
  NAND2_X1 U6641 ( .A1(n6108), .A2(n5636), .ZN(n5481) );
  NAND2_X1 U6642 ( .A1(n6142), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5480)
         );
  AOI22_X1 U6643 ( .A1(EBX_REG_15__SCAN_IN), .A2(n3126), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5478), .ZN(n5479) );
  NAND4_X1 U6644 ( .A1(n5481), .A2(n5480), .A3(n5479), .A4(n6232), .ZN(n5482)
         );
  NOR2_X1 U6645 ( .A1(n5483), .A2(n5482), .ZN(n5484) );
  OAI211_X1 U6646 ( .C1(n5757), .C2(n6115), .A(n5485), .B(n5484), .ZN(U2812)
         );
  INV_X1 U6647 ( .A(n5486), .ZN(n5488) );
  OAI22_X1 U6648 ( .A1(n5488), .A2(n6155), .B1(n6163), .B2(n5487), .ZN(U2828)
         );
  OAI222_X1 U6649 ( .A1(n5531), .A2(n5534), .B1(n5490), .B2(n6163), .C1(n5489), 
        .C2(n6155), .ZN(U2830) );
  INV_X1 U6650 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5491) );
  OAI222_X1 U6651 ( .A1(n5531), .A2(n5537), .B1(n5491), .B2(n6163), .C1(n5674), 
        .C2(n6155), .ZN(U2831) );
  BUF_X1 U6652 ( .A(n5492), .Z(n5493) );
  NAND2_X1 U6653 ( .A1(n5394), .A2(n5494), .ZN(n5495) );
  NOR2_X1 U6654 ( .A1(n5497), .A2(n5496), .ZN(n5498) );
  OR2_X1 U6655 ( .A1(n5680), .A2(n5498), .ZN(n5972) );
  OAI22_X1 U6656 ( .A1(n5972), .A2(n6155), .B1(n5863), .B2(n6163), .ZN(n5499)
         );
  AOI21_X1 U6657 ( .B1(n5860), .B2(n6160), .A(n5499), .ZN(n5500) );
  INV_X1 U6658 ( .A(n5500), .ZN(U2833) );
  OAI22_X1 U6659 ( .A1(n5693), .A2(n6155), .B1(n5501), .B2(n6163), .ZN(n5502)
         );
  AOI21_X1 U6660 ( .B1(n5947), .B2(n6160), .A(n5502), .ZN(n5503) );
  INV_X1 U6661 ( .A(n5503), .ZN(U2834) );
  OR2_X1 U6662 ( .A1(n5504), .A2(n5505), .ZN(n5506) );
  NAND2_X1 U6663 ( .A1(n5396), .A2(n5506), .ZN(n5865) );
  INV_X1 U6664 ( .A(n5706), .ZN(n5513) );
  AOI21_X1 U6665 ( .B1(n5513), .B2(n5705), .A(n5507), .ZN(n5509) );
  NOR2_X1 U6666 ( .A1(n5509), .A2(n5508), .ZN(n5866) );
  AOI22_X1 U6667 ( .A1(n5866), .A2(n6159), .B1(EBX_REG_24__SCAN_IN), .B2(n5529), .ZN(n5510) );
  OAI21_X1 U6668 ( .B1(n5865), .B2(n5531), .A(n5510), .ZN(U2835) );
  AOI21_X1 U6669 ( .B1(n5512), .B2(n5414), .A(n5511), .ZN(n5936) );
  INV_X1 U6670 ( .A(n5936), .ZN(n5517) );
  AOI21_X1 U6671 ( .B1(n5515), .B2(n5514), .A(n5513), .ZN(n5882) );
  AOI22_X1 U6672 ( .A1(n5882), .A2(n6159), .B1(EBX_REG_22__SCAN_IN), .B2(n5529), .ZN(n5516) );
  OAI21_X1 U6673 ( .B1(n5517), .B2(n5531), .A(n5516), .ZN(U2837) );
  OAI222_X1 U6674 ( .A1(n5939), .A2(n5531), .B1(n5518), .B2(n6163), .C1(n6155), 
        .C2(n5731), .ZN(U2838) );
  MUX2_X1 U6675 ( .A(n3128), .B(n5520), .S(n5519), .Z(n5522) );
  XNOR2_X1 U6676 ( .A(n5522), .B(n5521), .ZN(n5737) );
  INV_X1 U6677 ( .A(n5737), .ZN(n5890) );
  INV_X1 U6678 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5525) );
  OAI21_X1 U6679 ( .B1(n5523), .B2(n5524), .A(n5415), .ZN(n5891) );
  OAI222_X1 U6680 ( .A1(n5890), .A2(n6155), .B1(n6163), .B2(n5525), .C1(n5891), 
        .C2(n5531), .ZN(U2839) );
  OAI222_X1 U6681 ( .A1(n5750), .A2(n6155), .B1(n6163), .B2(n5440), .C1(n5624), 
        .C2(n5531), .ZN(U2841) );
  OAI22_X1 U6682 ( .A1(n5991), .A2(n6155), .B1(n5526), .B2(n6163), .ZN(n5527)
         );
  AOI21_X1 U6683 ( .B1(n6166), .B2(n6160), .A(n5527), .ZN(n5528) );
  INV_X1 U6684 ( .A(n5528), .ZN(U2842) );
  AOI22_X1 U6685 ( .A1(n6000), .A2(n6159), .B1(EBX_REG_16__SCAN_IN), .B2(n5529), .ZN(n5530) );
  OAI21_X1 U6686 ( .B1(n5631), .B2(n5531), .A(n5530), .ZN(U2843) );
  INV_X1 U6687 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6962) );
  OAI222_X1 U6688 ( .A1(n5637), .A2(n5531), .B1(n6163), .B2(n6962), .C1(n5757), 
        .C2(n6155), .ZN(U2844) );
  AOI22_X1 U6689 ( .A1(n6168), .A2(DATAI_13_), .B1(n6167), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U6690 ( .A1(n6164), .A2(DATAI_29_), .ZN(n5532) );
  OAI211_X1 U6691 ( .C1(n5534), .C2(n5924), .A(n5533), .B(n5532), .ZN(U2862)
         );
  AOI22_X1 U6692 ( .A1(n6168), .A2(DATAI_12_), .B1(n6167), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5536) );
  NAND2_X1 U6693 ( .A1(n6164), .A2(DATAI_28_), .ZN(n5535) );
  OAI211_X1 U6694 ( .C1(n5537), .C2(n5924), .A(n5536), .B(n5535), .ZN(U2863)
         );
  INV_X1 U6695 ( .A(n5860), .ZN(n5540) );
  AOI22_X1 U6696 ( .A1(n6168), .A2(DATAI_10_), .B1(n6167), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U6697 ( .A1(n6164), .A2(DATAI_26_), .ZN(n5538) );
  OAI211_X1 U6698 ( .C1(n5540), .C2(n5924), .A(n5539), .B(n5538), .ZN(U2865)
         );
  AOI22_X1 U6699 ( .A1(n6168), .A2(DATAI_4_), .B1(n6167), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6700 ( .A1(n6164), .A2(DATAI_20_), .ZN(n5541) );
  OAI211_X1 U6701 ( .C1(n5891), .C2(n5924), .A(n5542), .B(n5541), .ZN(U2871)
         );
  AOI22_X1 U6702 ( .A1(n6164), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6167), .ZN(n5544) );
  NAND2_X1 U6703 ( .A1(n6168), .A2(DATAI_2_), .ZN(n5543) );
  OAI211_X1 U6704 ( .C1(n5624), .C2(n5924), .A(n5544), .B(n5543), .ZN(U2873)
         );
  AOI22_X1 U6705 ( .A1(n6164), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6167), .ZN(n5546) );
  NAND2_X1 U6706 ( .A1(n6168), .A2(DATAI_0_), .ZN(n5545) );
  OAI211_X1 U6707 ( .C1(n5631), .C2(n5924), .A(n5546), .B(n5545), .ZN(U2875)
         );
  AOI22_X1 U6708 ( .A1(n5547), .A2(DATAI_15_), .B1(n6167), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5548) );
  OAI21_X1 U6709 ( .B1(n5637), .B2(n5924), .A(n5548), .ZN(U2876) );
  MUX2_X2 U6710 ( .A(n5550), .B(n5549), .S(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .Z(n5551) );
  XNOR2_X1 U6711 ( .A(n5551), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5666)
         );
  NAND2_X1 U6712 ( .A1(n5966), .A2(n5552), .ZN(n5553) );
  NAND2_X1 U6713 ( .A1(n6308), .A2(REIP_REG_30__SCAN_IN), .ZN(n5661) );
  OAI211_X1 U6714 ( .C1(n5554), .C2(n5969), .A(n5553), .B(n5661), .ZN(n5555)
         );
  AOI21_X1 U6715 ( .B1(n5556), .B2(n6226), .A(n5555), .ZN(n5557) );
  OAI21_X1 U6716 ( .B1(n5666), .B2(n6034), .A(n5557), .ZN(U2956) );
  NAND2_X1 U6717 ( .A1(n5559), .A2(n5558), .ZN(n5560) );
  XNOR2_X1 U6718 ( .A(n5560), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5689)
         );
  NOR2_X1 U6719 ( .A1(n6232), .A2(n6676), .ZN(n5681) );
  AOI21_X1 U6720 ( .B1(n6222), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5681), 
        .ZN(n5563) );
  OAI21_X1 U6721 ( .B1(n5848), .B2(n6231), .A(n5563), .ZN(n5564) );
  AOI21_X1 U6722 ( .B1(n5925), .B2(n6226), .A(n5564), .ZN(n5565) );
  OAI21_X1 U6723 ( .B1(n5689), .B2(n6034), .A(n5565), .ZN(U2959) );
  NOR2_X1 U6724 ( .A1(n5567), .A2(n5566), .ZN(n5569) );
  XOR2_X1 U6725 ( .A(n5569), .B(n5568), .Z(n5971) );
  NAND2_X1 U6726 ( .A1(n5860), .A2(n6226), .ZN(n5574) );
  INV_X1 U6727 ( .A(REIP_REG_26__SCAN_IN), .ZN(n5570) );
  OAI22_X1 U6728 ( .A1(n5969), .A2(n5571), .B1(n6232), .B2(n5570), .ZN(n5572)
         );
  AOI21_X1 U6729 ( .B1(n5966), .B2(n5855), .A(n5572), .ZN(n5573) );
  OAI211_X1 U6730 ( .C1(n5971), .C2(n6034), .A(n5574), .B(n5573), .ZN(U2960)
         );
  XNOR2_X1 U6731 ( .A(n5633), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5951)
         );
  NAND2_X1 U6732 ( .A1(n5952), .A2(n5951), .ZN(n5953) );
  OR2_X1 U6733 ( .A1(n5584), .A2(n6971), .ZN(n5575) );
  NAND2_X1 U6734 ( .A1(n5584), .A2(n5576), .ZN(n5578) );
  NOR2_X1 U6735 ( .A1(n5633), .A2(n5576), .ZN(n5577) );
  AOI21_X1 U6736 ( .B1(n5612), .B2(n5578), .A(n5577), .ZN(n5604) );
  XNOR2_X1 U6737 ( .A(n5633), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5605)
         );
  AND2_X2 U6738 ( .A1(n5604), .A2(n5605), .ZN(n5602) );
  NOR2_X1 U6739 ( .A1(n5633), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5595)
         );
  NAND2_X1 U6740 ( .A1(n5602), .A2(n5595), .ZN(n5585) );
  NAND4_X1 U6741 ( .A1(n5596), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n5584), .ZN(n5579) );
  OAI21_X1 U6742 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5585), .A(n5579), 
        .ZN(n5580) );
  XNOR2_X1 U6743 ( .A(n5580), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5704)
         );
  NAND2_X1 U6744 ( .A1(n6308), .A2(REIP_REG_24__SCAN_IN), .ZN(n5697) );
  OAI21_X1 U6745 ( .B1(n5969), .B2(n6808), .A(n5697), .ZN(n5582) );
  NOR2_X1 U6746 ( .A1(n5865), .A2(n5955), .ZN(n5581) );
  AOI211_X1 U6747 ( .C1(n5966), .C2(n5864), .A(n5582), .B(n5581), .ZN(n5583)
         );
  OAI21_X1 U6748 ( .B1(n5704), .B2(n6034), .A(n5583), .ZN(U2962) );
  NAND3_X1 U6749 ( .A1(n5584), .A2(n5734), .A3(n5718), .ZN(n5586) );
  OAI21_X1 U6750 ( .B1(n5587), .B2(n5586), .A(n5585), .ZN(n5588) );
  XNOR2_X1 U6751 ( .A(n5588), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5714)
         );
  INV_X1 U6752 ( .A(n5589), .ZN(n5591) );
  INV_X1 U6753 ( .A(n5511), .ZN(n5590) );
  AOI21_X1 U6754 ( .B1(n5591), .B2(n5590), .A(n5504), .ZN(n5933) );
  NAND2_X1 U6755 ( .A1(n6308), .A2(REIP_REG_23__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U6756 ( .A1(n6222), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5592)
         );
  OAI211_X1 U6757 ( .C1(n6231), .C2(n5873), .A(n5709), .B(n5592), .ZN(n5593)
         );
  AOI21_X1 U6758 ( .B1(n5933), .B2(n6226), .A(n5593), .ZN(n5594) );
  OAI21_X1 U6759 ( .B1(n5714), .B2(n6034), .A(n5594), .ZN(U2963) );
  AOI21_X1 U6760 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5633), .A(n5595), 
        .ZN(n5597) );
  XOR2_X1 U6761 ( .A(n5597), .B(n5596), .Z(n5723) );
  INV_X1 U6762 ( .A(n5881), .ZN(n5599) );
  NAND2_X1 U6763 ( .A1(n6308), .A2(REIP_REG_22__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U6764 ( .A1(n6222), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5598)
         );
  OAI211_X1 U6765 ( .C1(n6231), .C2(n5599), .A(n5715), .B(n5598), .ZN(n5600)
         );
  AOI21_X1 U6766 ( .B1(n5936), .B2(n6226), .A(n5600), .ZN(n5601) );
  OAI21_X1 U6767 ( .B1(n5723), .B2(n6034), .A(n5601), .ZN(U2964) );
  INV_X1 U6768 ( .A(n5602), .ZN(n5603) );
  OAI21_X1 U6769 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5724) );
  NAND2_X1 U6770 ( .A1(n5724), .A2(n4529), .ZN(n5610) );
  INV_X1 U6771 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5606) );
  NOR2_X1 U6772 ( .A1(n6232), .A2(n5606), .ZN(n5727) );
  NOR2_X1 U6773 ( .A1(n6231), .A2(n5607), .ZN(n5608) );
  AOI211_X1 U6774 ( .C1(n6222), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5727), 
        .B(n5608), .ZN(n5609) );
  OAI211_X1 U6775 ( .C1(n5955), .C2(n5939), .A(n5610), .B(n5609), .ZN(U2965)
         );
  XNOR2_X1 U6776 ( .A(n5633), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5611)
         );
  XNOR2_X1 U6777 ( .A(n5612), .B(n5611), .ZN(n5742) );
  NAND2_X1 U6778 ( .A1(n6308), .A2(REIP_REG_20__SCAN_IN), .ZN(n5732) );
  OAI21_X1 U6779 ( .B1(n5969), .B2(n5897), .A(n5732), .ZN(n5614) );
  NOR2_X1 U6780 ( .A1(n5891), .A2(n5955), .ZN(n5613) );
  AOI211_X1 U6781 ( .C1(n5966), .C2(n5888), .A(n5614), .B(n5613), .ZN(n5615)
         );
  OAI21_X1 U6782 ( .B1(n5742), .B2(n6034), .A(n5615), .ZN(U2966) );
  NOR2_X1 U6783 ( .A1(n3138), .A2(n6947), .ZN(n5962) );
  NAND2_X1 U6784 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5962), .ZN(n5618) );
  NOR2_X1 U6785 ( .A1(n5633), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5961)
         );
  NAND3_X1 U6786 ( .A1(n5961), .A2(n5963), .A3(n5616), .ZN(n5617) );
  OAI21_X1 U6787 ( .B1(n5618), .B2(n5616), .A(n5617), .ZN(n5619) );
  XNOR2_X1 U6788 ( .A(n5743), .B(n5619), .ZN(n5747) );
  AOI22_X1 U6789 ( .A1(n4529), .A2(n5747), .B1(n6308), .B2(
        REIP_REG_18__SCAN_IN), .ZN(n5620) );
  OAI21_X1 U6790 ( .B1(n5436), .B2(n5969), .A(n5620), .ZN(n5621) );
  AOI21_X1 U6791 ( .B1(n5966), .B2(n5622), .A(n5621), .ZN(n5623) );
  OAI21_X1 U6792 ( .B1(n5624), .B2(n5955), .A(n5623), .ZN(U2968) );
  NOR2_X1 U6793 ( .A1(n5962), .A2(n5961), .ZN(n5625) );
  XOR2_X1 U6794 ( .A(n5625), .B(n5616), .Z(n6002) );
  NAND2_X1 U6795 ( .A1(n6002), .A2(n4529), .ZN(n5630) );
  INV_X1 U6796 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5626) );
  NOR2_X1 U6797 ( .A1(n6232), .A2(n5626), .ZN(n5999) );
  NOR2_X1 U6798 ( .A1(n5627), .A2(n6231), .ZN(n5628) );
  AOI211_X1 U6799 ( .C1(n6222), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5999), 
        .B(n5628), .ZN(n5629) );
  OAI211_X1 U6800 ( .C1(n5955), .C2(n5631), .A(n5630), .B(n5629), .ZN(U2970)
         );
  XNOR2_X1 U6801 ( .A(n5633), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5634)
         );
  XNOR2_X1 U6802 ( .A(n5632), .B(n5634), .ZN(n5762) );
  OAI22_X1 U6803 ( .A1(n5969), .A2(n3923), .B1(n6232), .B2(n6659), .ZN(n5635)
         );
  AOI21_X1 U6804 ( .B1(n5636), .B2(n5966), .A(n5635), .ZN(n5639) );
  OR2_X1 U6805 ( .A1(n5637), .A2(n5955), .ZN(n5638) );
  OAI211_X1 U6806 ( .C1(n5762), .C2(n6034), .A(n5639), .B(n5638), .ZN(U2971)
         );
  INV_X1 U6807 ( .A(n5641), .ZN(n5643) );
  NOR2_X1 U6808 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  XNOR2_X1 U6809 ( .A(n5640), .B(n5644), .ZN(n6016) );
  NAND2_X1 U6810 ( .A1(n6016), .A2(n4529), .ZN(n5648) );
  NOR2_X1 U6811 ( .A1(n6232), .A2(n4490), .ZN(n6008) );
  NOR2_X1 U6812 ( .A1(n6231), .A2(n5645), .ZN(n5646) );
  AOI211_X1 U6813 ( .C1(n6222), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6008), 
        .B(n5646), .ZN(n5647) );
  OAI211_X1 U6814 ( .C1(n5955), .C2(n5649), .A(n5648), .B(n5647), .ZN(U2972)
         );
  XNOR2_X1 U6815 ( .A(n5651), .B(n5650), .ZN(n5763) );
  NAND2_X1 U6816 ( .A1(n5763), .A2(n4529), .ZN(n5655) );
  AND2_X1 U6817 ( .A1(n6308), .A2(REIP_REG_13__SCAN_IN), .ZN(n5771) );
  NOR2_X1 U6818 ( .A1(n6231), .A2(n5652), .ZN(n5653) );
  AOI211_X1 U6819 ( .C1(n6222), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5771), 
        .B(n5653), .ZN(n5654) );
  OAI211_X1 U6820 ( .C1(n5955), .C2(n5656), .A(n5655), .B(n5654), .ZN(U2973)
         );
  OAI211_X1 U6821 ( .C1(n5657), .C2(n6830), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5686), .ZN(n5662) );
  NAND3_X1 U6822 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5658), .ZN(n5660) );
  NAND3_X1 U6823 ( .A1(n5662), .A2(n5661), .A3(n5660), .ZN(n5663) );
  AOI21_X1 U6824 ( .B1(n5664), .B2(n6310), .A(n5663), .ZN(n5665) );
  OAI21_X1 U6825 ( .B1(n5666), .B2(n5992), .A(n5665), .ZN(U2988) );
  INV_X1 U6826 ( .A(n5686), .ZN(n5668) );
  OR2_X1 U6827 ( .A1(n5669), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5683)
         );
  OAI21_X1 U6828 ( .B1(n5668), .B2(n5667), .A(n5683), .ZN(n5676) );
  INV_X1 U6829 ( .A(n5669), .ZN(n5671) );
  INV_X1 U6830 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5670) );
  NAND3_X1 U6831 ( .A1(n5671), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5670), .ZN(n5672) );
  OAI211_X1 U6832 ( .C1(n5674), .C2(n6233), .A(n5673), .B(n5672), .ZN(n5675)
         );
  AOI21_X1 U6833 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5676), .A(n5675), 
        .ZN(n5677) );
  OAI21_X1 U6834 ( .B1(n5678), .B2(n5992), .A(n5677), .ZN(U2990) );
  XNOR2_X1 U6835 ( .A(n5680), .B(n5679), .ZN(n5916) );
  INV_X1 U6836 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U6837 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  AOI21_X1 U6838 ( .B1(n5916), .B2(n6310), .A(n5684), .ZN(n5688) );
  NAND3_X1 U6839 ( .A1(n5686), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5685), .ZN(n5687) );
  OAI211_X1 U6840 ( .C1(n5689), .C2(n5992), .A(n5688), .B(n5687), .ZN(U2991)
         );
  NAND2_X1 U6841 ( .A1(n3656), .A2(n5690), .ZN(n5691) );
  NAND2_X1 U6842 ( .A1(n4190), .A2(n5691), .ZN(n5946) );
  NOR2_X1 U6843 ( .A1(n5699), .A2(n5976), .ZN(n5695) );
  AOI22_X1 U6844 ( .A1(n5975), .A2(n5976), .B1(REIP_REG_25__SCAN_IN), .B2(
        n6308), .ZN(n5692) );
  OAI21_X1 U6845 ( .B1(n5693), .B2(n6233), .A(n5692), .ZN(n5694) );
  AOI211_X1 U6846 ( .C1(n5946), .C2(n6315), .A(n5695), .B(n5694), .ZN(n5696)
         );
  INV_X1 U6847 ( .A(n5696), .ZN(U2993) );
  INV_X1 U6848 ( .A(n5697), .ZN(n5698) );
  AOI21_X1 U6849 ( .B1(n5866), .B2(n6310), .A(n5698), .ZN(n5703) );
  INV_X1 U6850 ( .A(n5699), .ZN(n5970) );
  INV_X1 U6851 ( .A(n5700), .ZN(n5701) );
  OAI211_X1 U6852 ( .C1(INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n5707), .A(n5970), .B(n5701), .ZN(n5702) );
  OAI211_X1 U6853 ( .C1(n5704), .C2(n5992), .A(n5703), .B(n5702), .ZN(U2994)
         );
  XNOR2_X1 U6854 ( .A(n5706), .B(n5705), .ZN(n5919) );
  INV_X1 U6855 ( .A(n5707), .ZN(n5711) );
  NAND2_X1 U6856 ( .A1(n5708), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5710) );
  OAI211_X1 U6857 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5711), .A(n5710), .B(n5709), .ZN(n5712) );
  AOI21_X1 U6858 ( .B1(n5919), .B2(n6310), .A(n5712), .ZN(n5713) );
  OAI21_X1 U6859 ( .B1(n5714), .B2(n5992), .A(n5713), .ZN(U2995) );
  INV_X1 U6860 ( .A(n5715), .ZN(n5720) );
  INV_X1 U6861 ( .A(n5716), .ZN(n5725) );
  NOR3_X1 U6862 ( .A1(n5725), .A2(n5718), .A3(n5717), .ZN(n5719) );
  AOI211_X1 U6863 ( .C1(n5728), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5720), .B(n5719), .ZN(n5722) );
  NAND2_X1 U6864 ( .A1(n5882), .A2(n6310), .ZN(n5721) );
  OAI211_X1 U6865 ( .C1(n5723), .C2(n5992), .A(n5722), .B(n5721), .ZN(U2996)
         );
  NAND2_X1 U6866 ( .A1(n5724), .A2(n6315), .ZN(n5730) );
  NOR2_X1 U6867 ( .A1(n5725), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5726)
         );
  AOI211_X1 U6868 ( .C1(n5728), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5727), .B(n5726), .ZN(n5729) );
  OAI211_X1 U6869 ( .C1(n6233), .C2(n5731), .A(n5730), .B(n5729), .ZN(U2997)
         );
  INV_X1 U6870 ( .A(n5732), .ZN(n5736) );
  NOR3_X1 U6871 ( .A1(n5734), .A2(n5733), .A3(n5988), .ZN(n5735) );
  AOI211_X1 U6872 ( .C1(n5737), .C2(n6310), .A(n5736), .B(n5735), .ZN(n5741)
         );
  OAI221_X1 U6873 ( .B1(n6291), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n6291), .C2(n5739), .A(n5738), .ZN(n5996) );
  AOI21_X1 U6874 ( .B1(n6317), .B2(n5963), .A(n5996), .ZN(n5744) );
  OAI21_X1 U6875 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6270), .A(n5744), 
        .ZN(n5984) );
  NAND2_X1 U6876 ( .A1(n5984), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5740) );
  OAI211_X1 U6877 ( .C1(n5742), .C2(n5992), .A(n5741), .B(n5740), .ZN(U2998)
         );
  INV_X1 U6878 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6664) );
  OAI22_X1 U6879 ( .A1(n5744), .A2(n5743), .B1(n6232), .B2(n6664), .ZN(n5745)
         );
  INV_X1 U6880 ( .A(n5745), .ZN(n5749) );
  NOR3_X1 U6881 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5963), .A3(n5998), 
        .ZN(n5746) );
  AOI21_X1 U6882 ( .B1(n6315), .B2(n5747), .A(n5746), .ZN(n5748) );
  OAI211_X1 U6883 ( .C1(n5750), .C2(n6233), .A(n5749), .B(n5748), .ZN(U3000)
         );
  INV_X1 U6884 ( .A(n5751), .ZN(n5756) );
  NOR2_X1 U6885 ( .A1(n5753), .A2(n5752), .ZN(n5754) );
  AOI221_X1 U6886 ( .B1(n6311), .B2(n6011), .C1(n5755), .C2(n6011), .A(n5754), 
        .ZN(n6238) );
  OAI21_X1 U6887 ( .B1(n6270), .B2(n5756), .A(n6238), .ZN(n6001) );
  OAI22_X1 U6888 ( .A1(n5757), .A2(n6233), .B1(n6659), .B2(n6232), .ZN(n5758)
         );
  AOI21_X1 U6889 ( .B1(n6001), .B2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5758), 
        .ZN(n5761) );
  NAND2_X1 U6890 ( .A1(n6004), .A2(n5759), .ZN(n5760) );
  OAI211_X1 U6891 ( .C1(n5762), .C2(n5992), .A(n5761), .B(n5760), .ZN(U3003)
         );
  INV_X1 U6892 ( .A(n5763), .ZN(n5774) );
  INV_X1 U6893 ( .A(n5764), .ZN(n6239) );
  INV_X1 U6894 ( .A(n5769), .ZN(n5777) );
  NAND2_X1 U6895 ( .A1(n5777), .A2(n4318), .ZN(n6014) );
  OAI21_X1 U6896 ( .B1(n5766), .B2(n5765), .A(n6238), .ZN(n5767) );
  AOI21_X1 U6897 ( .B1(n5769), .B2(n5768), .A(n5767), .ZN(n6012) );
  OAI22_X1 U6898 ( .A1(n6239), .A2(n6014), .B1(n6012), .B2(n4318), .ZN(n5770)
         );
  AOI211_X1 U6899 ( .C1(n6310), .C2(n5772), .A(n5771), .B(n5770), .ZN(n5773)
         );
  OAI21_X1 U6900 ( .B1(n5774), .B2(n5992), .A(n5773), .ZN(U3005) );
  INV_X1 U6901 ( .A(n5775), .ZN(n5776) );
  AOI21_X1 U6902 ( .B1(n6053), .B2(n6310), .A(n5776), .ZN(n5784) );
  INV_X1 U6903 ( .A(n6238), .ZN(n5782) );
  AOI21_X1 U6904 ( .B1(n6291), .B2(n5778), .A(n5777), .ZN(n5781) );
  INV_X1 U6905 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6970) );
  OAI21_X1 U6906 ( .B1(n6239), .B2(n6970), .A(n5779), .ZN(n5780) );
  OAI21_X1 U6907 ( .B1(n5782), .B2(n5781), .A(n5780), .ZN(n5783) );
  OAI211_X1 U6908 ( .C1(n5785), .C2(n5992), .A(n5784), .B(n5783), .ZN(U3006)
         );
  NOR2_X1 U6909 ( .A1(n6455), .A2(n6033), .ZN(n6326) );
  INV_X1 U6910 ( .A(n6326), .ZN(n6458) );
  OAI211_X1 U6911 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6372), .A(n6458), .B(
        n6456), .ZN(n5786) );
  OAI21_X1 U6912 ( .B1(n5792), .B2(n5787), .A(n5786), .ZN(n5788) );
  MUX2_X1 U6913 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5788), .S(n6322), 
        .Z(U3464) );
  XNOR2_X1 U6914 ( .A(n6458), .B(n4754), .ZN(n5789) );
  OAI22_X1 U6915 ( .A1(n5789), .A2(n6499), .B1(n4751), .B2(n5792), .ZN(n5790)
         );
  MUX2_X1 U6916 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5790), .S(n6322), 
        .Z(U3463) );
  INV_X1 U6917 ( .A(n4792), .ZN(n5794) );
  NAND2_X1 U6918 ( .A1(n5791), .A2(n6457), .ZN(n6328) );
  NOR2_X1 U6919 ( .A1(n6458), .A2(n6371), .ZN(n6383) );
  NOR2_X1 U6920 ( .A1(n6328), .A2(n6383), .ZN(n5793) );
  OAI222_X1 U6921 ( .A1(n5801), .A2(n5794), .B1(n6499), .B2(n5793), .C1(n5792), 
        .C2(n6418), .ZN(n5795) );
  MUX2_X1 U6922 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5795), .S(n6322), 
        .Z(U3462) );
  INV_X1 U6923 ( .A(n6022), .ZN(n5797) );
  OAI22_X1 U6924 ( .A1(n5798), .A2(n5797), .B1(n5796), .B2(n6612), .ZN(n5799)
         );
  MUX2_X1 U6925 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5799), .S(n6025), 
        .Z(U3456) );
  NAND2_X1 U6926 ( .A1(n5800), .A2(n6325), .ZN(n6334) );
  NOR2_X1 U6927 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6334), .ZN(n5843)
         );
  INV_X1 U6928 ( .A(n6359), .ZN(n6349) );
  OAI21_X1 U6929 ( .B1(n6349), .B2(n5840), .A(n5801), .ZN(n5803) );
  NAND2_X1 U6930 ( .A1(n6418), .A2(n5802), .ZN(n6329) );
  NAND2_X1 U6931 ( .A1(n5803), .A2(n6329), .ZN(n5805) );
  OAI221_X1 U6932 ( .B1(n5843), .B2(n6693), .C1(n5843), .C2(n5805), .A(n5804), 
        .ZN(n5833) );
  INV_X1 U6933 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5813) );
  OR2_X1 U6934 ( .A1(n6329), .A2(n6499), .ZN(n5808) );
  NAND3_X1 U6935 ( .A1(n5806), .A2(n6410), .A3(n6325), .ZN(n5807) );
  NAND2_X1 U6936 ( .A1(n5808), .A2(n5807), .ZN(n5839) );
  AOI22_X1 U6937 ( .A1(n5840), .A2(n6563), .B1(n6560), .B2(n5839), .ZN(n5809)
         );
  OAI21_X1 U6938 ( .B1(n5810), .B2(n6359), .A(n5809), .ZN(n5811) );
  AOI21_X1 U6939 ( .B1(n6561), .B2(n5843), .A(n5811), .ZN(n5812) );
  OAI21_X1 U6940 ( .B1(n5846), .B2(n5813), .A(n5812), .ZN(U3036) );
  INV_X1 U6941 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5817) );
  AOI22_X1 U6942 ( .A1(n5840), .A2(n6516), .B1(n6514), .B2(n5839), .ZN(n5814)
         );
  OAI21_X1 U6943 ( .B1(n6474), .B2(n6359), .A(n5814), .ZN(n5815) );
  AOI21_X1 U6944 ( .B1(n6515), .B2(n5843), .A(n5815), .ZN(n5816) );
  OAI21_X1 U6945 ( .B1(n5846), .B2(n5817), .A(n5816), .ZN(U3037) );
  NAND2_X1 U6946 ( .A1(n6521), .A2(n5843), .ZN(n5819) );
  AOI22_X1 U6947 ( .A1(n6522), .A2(n5839), .B1(n6523), .B2(n5840), .ZN(n5818)
         );
  OAI211_X1 U6948 ( .C1(n6359), .C2(n6390), .A(n5819), .B(n5818), .ZN(n5820)
         );
  AOI21_X1 U6949 ( .B1(n5833), .B2(INSTQUEUE_REG_2__2__SCAN_IN), .A(n5820), 
        .ZN(n5821) );
  INV_X1 U6950 ( .A(n5821), .ZN(U3038) );
  INV_X1 U6951 ( .A(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5825) );
  AOI22_X1 U6952 ( .A1(n5840), .A2(n6530), .B1(n6528), .B2(n5839), .ZN(n5822)
         );
  OAI21_X1 U6953 ( .B1(n6480), .B2(n6359), .A(n5822), .ZN(n5823) );
  AOI21_X1 U6954 ( .B1(n6529), .B2(n5843), .A(n5823), .ZN(n5824) );
  OAI21_X1 U6955 ( .B1(n5846), .B2(n5825), .A(n5824), .ZN(U3039) );
  INV_X1 U6956 ( .A(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5829) );
  AOI22_X1 U6957 ( .A1(n5840), .A2(n6537), .B1(n6535), .B2(n5839), .ZN(n5826)
         );
  OAI21_X1 U6958 ( .B1(n6485), .B2(n6359), .A(n5826), .ZN(n5827) );
  AOI21_X1 U6959 ( .B1(n6536), .B2(n5843), .A(n5827), .ZN(n5828) );
  OAI21_X1 U6960 ( .B1(n5846), .B2(n5829), .A(n5828), .ZN(U3040) );
  NAND2_X1 U6961 ( .A1(n6568), .A2(n5843), .ZN(n5831) );
  AOI22_X1 U6962 ( .A1(n6570), .A2(n5839), .B1(n6571), .B2(n5840), .ZN(n5830)
         );
  OAI211_X1 U6963 ( .C1(n6359), .C2(n6398), .A(n5831), .B(n5830), .ZN(n5832)
         );
  AOI21_X1 U6964 ( .B1(n5833), .B2(INSTQUEUE_REG_2__5__SCAN_IN), .A(n5832), 
        .ZN(n5834) );
  INV_X1 U6965 ( .A(n5834), .ZN(U3041) );
  INV_X1 U6966 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5838) );
  AOI22_X1 U6967 ( .A1(n5840), .A2(n6545), .B1(n6543), .B2(n5839), .ZN(n5835)
         );
  OAI21_X1 U6968 ( .B1(n6352), .B2(n6359), .A(n5835), .ZN(n5836) );
  AOI21_X1 U6969 ( .B1(n6544), .B2(n5843), .A(n5836), .ZN(n5837) );
  OAI21_X1 U6970 ( .B1(n5846), .B2(n5838), .A(n5837), .ZN(U3042) );
  INV_X1 U6971 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5845) );
  AOI22_X1 U6972 ( .A1(n5840), .A2(n6552), .B1(n6550), .B2(n5839), .ZN(n5841)
         );
  OAI21_X1 U6973 ( .B1(n7035), .B2(n6359), .A(n5841), .ZN(n5842) );
  AOI21_X1 U6974 ( .B1(n7041), .B2(n5843), .A(n5842), .ZN(n5844) );
  OAI21_X1 U6975 ( .B1(n5846), .B2(n5845), .A(n5844), .ZN(U3043) );
  AND2_X1 U6976 ( .A1(DATAO_REG_31__SCAN_IN), .A2(n5847), .ZN(U2892) );
  NOR2_X1 U6977 ( .A1(n5848), .A2(n6146), .ZN(n5851) );
  OAI22_X1 U6978 ( .A1(n5849), .A2(n6117), .B1(n6676), .B2(n5857), .ZN(n5850)
         );
  AOI211_X1 U6979 ( .C1(n3126), .C2(EBX_REG_27__SCAN_IN), .A(n5851), .B(n5850), 
        .ZN(n5853) );
  AOI22_X1 U6980 ( .A1(n5925), .A2(n6094), .B1(n6143), .B2(n5916), .ZN(n5852)
         );
  OAI211_X1 U6981 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5854), .A(n5853), .B(n5852), .ZN(U2800) );
  AOI22_X1 U6982 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6142), .B1(n5855), 
        .B2(n6108), .ZN(n5862) );
  NOR2_X1 U6983 ( .A1(REIP_REG_26__SCAN_IN), .A2(n5856), .ZN(n5858) );
  OAI22_X1 U6984 ( .A1(n5858), .A2(n5857), .B1(n6115), .B2(n5972), .ZN(n5859)
         );
  AOI21_X1 U6985 ( .B1(n5860), .B2(n6094), .A(n5859), .ZN(n5861) );
  OAI211_X1 U6986 ( .C1(n5863), .C2(n6140), .A(n5862), .B(n5861), .ZN(U2801)
         );
  AOI22_X1 U6987 ( .A1(EBX_REG_24__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6142), .ZN(n5870) );
  AOI22_X1 U6988 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5872), .B1(n5864), .B2(
        n6108), .ZN(n5869) );
  INV_X1 U6989 ( .A(n5865), .ZN(n5930) );
  AOI22_X1 U6990 ( .A1(n5930), .A2(n6094), .B1(n5866), .B2(n6143), .ZN(n5868)
         );
  NAND4_X1 U6991 ( .A1(n5870), .A2(n5869), .A3(n5868), .A4(n5867), .ZN(U2803)
         );
  NOR2_X1 U6992 ( .A1(n5606), .A2(n5871), .ZN(n5880) );
  AOI21_X1 U6993 ( .B1(REIP_REG_22__SCAN_IN), .B2(n5880), .A(
        REIP_REG_23__SCAN_IN), .ZN(n5879) );
  INV_X1 U6994 ( .A(n5872), .ZN(n5878) );
  INV_X1 U6995 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5874) );
  OAI22_X1 U6996 ( .A1(n5874), .A2(n6117), .B1(n5873), .B2(n6146), .ZN(n5875)
         );
  AOI21_X1 U6997 ( .B1(EBX_REG_23__SCAN_IN), .B2(n3126), .A(n5875), .ZN(n5877)
         );
  AOI22_X1 U6998 ( .A1(n5933), .A2(n6094), .B1(n6143), .B2(n5919), .ZN(n5876)
         );
  OAI211_X1 U6999 ( .C1(n5879), .C2(n5878), .A(n5877), .B(n5876), .ZN(U2804)
         );
  AOI22_X1 U7000 ( .A1(EBX_REG_22__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6142), .ZN(n5887) );
  INV_X1 U7001 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6669) );
  AOI22_X1 U7002 ( .A1(n5881), .A2(n6108), .B1(n5880), .B2(n6669), .ZN(n5886)
         );
  AOI22_X1 U7003 ( .A1(n5936), .A2(n6094), .B1(n5882), .B2(n6143), .ZN(n5885)
         );
  OAI21_X1 U7004 ( .B1(n5894), .B2(n5883), .A(REIP_REG_22__SCAN_IN), .ZN(n5884) );
  NAND4_X1 U7005 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(U2805)
         );
  AOI22_X1 U7006 ( .A1(EBX_REG_20__SCAN_IN), .A2(n3126), .B1(n5888), .B2(n6108), .ZN(n5896) );
  NAND2_X1 U7007 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5911) );
  INV_X1 U7008 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U7009 ( .B1(n5911), .B2(n5889), .A(n6667), .ZN(n5893) );
  OAI22_X1 U7010 ( .A1(n5891), .A2(n6105), .B1(n6115), .B2(n5890), .ZN(n5892)
         );
  AOI21_X1 U7011 ( .B1(n5894), .B2(n5893), .A(n5892), .ZN(n5895) );
  OAI211_X1 U7012 ( .C1(n5897), .C2(n6117), .A(n5896), .B(n5895), .ZN(U2807)
         );
  INV_X1 U7013 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5898) );
  OAI21_X1 U7014 ( .B1(n6117), .B2(n5898), .A(n6232), .ZN(n5900) );
  OAI22_X1 U7015 ( .A1(n5923), .A2(n6140), .B1(n5960), .B2(n6146), .ZN(n5899)
         );
  AOI211_X1 U7016 ( .C1(REIP_REG_19__SCAN_IN), .C2(n5901), .A(n5900), .B(n5899), .ZN(n5915) );
  INV_X1 U7017 ( .A(n5523), .ZN(n5904) );
  NAND2_X1 U7018 ( .A1(n5430), .A2(n5902), .ZN(n5903) );
  NAND2_X1 U7019 ( .A1(n5904), .A2(n5903), .ZN(n5956) );
  NAND2_X1 U7020 ( .A1(n5906), .A2(n5905), .ZN(n5909) );
  INV_X1 U7021 ( .A(n5907), .ZN(n5908) );
  XNOR2_X1 U7022 ( .A(n5909), .B(n5908), .ZN(n5982) );
  OAI22_X1 U7023 ( .A1(n5956), .A2(n6105), .B1(n6115), .B2(n5982), .ZN(n5910)
         );
  INV_X1 U7024 ( .A(n5910), .ZN(n5914) );
  OAI211_X1 U7025 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5912), .B(n5911), .ZN(n5913) );
  NAND3_X1 U7026 ( .A1(n5915), .A2(n5914), .A3(n5913), .ZN(U2808) );
  AOI22_X1 U7027 ( .A1(n5925), .A2(n6160), .B1(n6159), .B2(n5916), .ZN(n5917)
         );
  OAI21_X1 U7028 ( .B1(n6163), .B2(n5918), .A(n5917), .ZN(U2832) );
  AOI22_X1 U7029 ( .A1(n5933), .A2(n6160), .B1(n6159), .B2(n5919), .ZN(n5920)
         );
  OAI21_X1 U7030 ( .B1(n6163), .B2(n6717), .A(n5920), .ZN(U2836) );
  OAI22_X1 U7031 ( .A1(n5956), .A2(n5531), .B1(n6155), .B2(n5982), .ZN(n5921)
         );
  INV_X1 U7032 ( .A(n5921), .ZN(n5922) );
  OAI21_X1 U7033 ( .B1(n6163), .B2(n5923), .A(n5922), .ZN(U2840) );
  AOI22_X1 U7034 ( .A1(n5925), .A2(n6165), .B1(n6164), .B2(DATAI_27_), .ZN(
        n5927) );
  AOI22_X1 U7035 ( .A1(n6168), .A2(DATAI_11_), .B1(n6167), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7036 ( .A1(n5927), .A2(n5926), .ZN(U2864) );
  AOI22_X1 U7037 ( .A1(n5947), .A2(n6165), .B1(n6164), .B2(DATAI_25_), .ZN(
        n5929) );
  AOI22_X1 U7038 ( .A1(n6168), .A2(DATAI_9_), .B1(n6167), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7039 ( .A1(n5929), .A2(n5928), .ZN(U2866) );
  AOI22_X1 U7040 ( .A1(n5930), .A2(n6165), .B1(n6164), .B2(DATAI_24_), .ZN(
        n5932) );
  AOI22_X1 U7041 ( .A1(n6168), .A2(DATAI_8_), .B1(n6167), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7042 ( .A1(n5932), .A2(n5931), .ZN(U2867) );
  AOI22_X1 U7043 ( .A1(n5933), .A2(n6165), .B1(n6164), .B2(DATAI_23_), .ZN(
        n5935) );
  AOI22_X1 U7044 ( .A1(n6168), .A2(DATAI_7_), .B1(n6167), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7045 ( .A1(n5935), .A2(n5934), .ZN(U2868) );
  AOI22_X1 U7046 ( .A1(n5936), .A2(n6165), .B1(n6164), .B2(DATAI_22_), .ZN(
        n5938) );
  AOI22_X1 U7047 ( .A1(n6168), .A2(DATAI_6_), .B1(n6167), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7048 ( .A1(n5938), .A2(n5937), .ZN(U2869) );
  INV_X1 U7049 ( .A(n5939), .ZN(n5940) );
  AOI22_X1 U7050 ( .A1(n5940), .A2(n6165), .B1(n6164), .B2(DATAI_21_), .ZN(
        n5942) );
  AOI22_X1 U7051 ( .A1(n6168), .A2(DATAI_5_), .B1(n6167), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7052 ( .A1(n5942), .A2(n5941), .ZN(U2870) );
  INV_X1 U7053 ( .A(n5956), .ZN(n5943) );
  AOI22_X1 U7054 ( .A1(n5943), .A2(n6165), .B1(n6164), .B2(DATAI_19_), .ZN(
        n5945) );
  AOI22_X1 U7055 ( .A1(n6168), .A2(DATAI_3_), .B1(n6167), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7056 ( .A1(n5945), .A2(n5944), .ZN(U2872) );
  AOI22_X1 U7057 ( .A1(n6308), .A2(REIP_REG_25__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5949) );
  AOI22_X1 U7058 ( .A1(n5947), .A2(n6226), .B1(n4529), .B2(n5946), .ZN(n5948)
         );
  OAI211_X1 U7059 ( .C1(n6231), .C2(n5950), .A(n5949), .B(n5948), .ZN(U2961)
         );
  AOI22_X1 U7060 ( .A1(n6308), .A2(REIP_REG_19__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7061 ( .A1(n5952), .A2(n5951), .ZN(n5954) );
  AND2_X1 U7062 ( .A1(n5954), .A2(n5953), .ZN(n5985) );
  NOR2_X1 U7063 ( .A1(n5956), .A2(n5955), .ZN(n5957) );
  AOI21_X1 U7064 ( .B1(n5985), .B2(n4529), .A(n5957), .ZN(n5958) );
  OAI211_X1 U7065 ( .C1(n6231), .C2(n5960), .A(n5959), .B(n5958), .ZN(U2967)
         );
  MUX2_X1 U7066 ( .A(n5962), .B(n5961), .S(n5616), .Z(n5964) );
  XNOR2_X1 U7067 ( .A(n5964), .B(n5963), .ZN(n5990) );
  INV_X1 U7068 ( .A(n5965), .ZN(n5967) );
  AOI222_X1 U7069 ( .A1(n5990), .A2(n4529), .B1(n6226), .B2(n6166), .C1(n5967), 
        .C2(n5966), .ZN(n5968) );
  NAND2_X1 U7070 ( .A1(n6308), .A2(REIP_REG_17__SCAN_IN), .ZN(n5989) );
  OAI211_X1 U7071 ( .C1(n6900), .C2(n5969), .A(n5968), .B(n5989), .ZN(U2969)
         );
  AOI22_X1 U7072 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n5970), .B1(n6308), .B2(REIP_REG_26__SCAN_IN), .ZN(n5980) );
  INV_X1 U7073 ( .A(n5971), .ZN(n5974) );
  INV_X1 U7074 ( .A(n5972), .ZN(n5973) );
  AOI22_X1 U7075 ( .A1(n5974), .A2(n6315), .B1(n6310), .B2(n5973), .ZN(n5979)
         );
  OAI221_X1 U7076 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .C1(n5977), .C2(n5976), .A(n5975), 
        .ZN(n5978) );
  NAND3_X1 U7077 ( .A1(n5980), .A2(n5979), .A3(n5978), .ZN(U2992) );
  INV_X1 U7078 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5981) );
  OAI22_X1 U7079 ( .A1(n5982), .A2(n6233), .B1(n6232), .B2(n5981), .ZN(n5983)
         );
  INV_X1 U7080 ( .A(n5983), .ZN(n5987) );
  AOI22_X1 U7081 ( .A1(n5985), .A2(n6315), .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5984), .ZN(n5986) );
  OAI211_X1 U7082 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5988), .A(n5987), .B(n5986), .ZN(U2999) );
  INV_X1 U7083 ( .A(n5989), .ZN(n5995) );
  INV_X1 U7084 ( .A(n5990), .ZN(n5993) );
  OAI22_X1 U7085 ( .A1(n5993), .A2(n5992), .B1(n6233), .B2(n5991), .ZN(n5994)
         );
  AOI211_X1 U7086 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5996), .A(n5995), .B(n5994), .ZN(n5997) );
  OAI21_X1 U7087 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5998), .A(n5997), 
        .ZN(U3001) );
  AOI21_X1 U7088 ( .B1(n6000), .B2(n6310), .A(n5999), .ZN(n6007) );
  AOI22_X1 U7089 ( .A1(n6002), .A2(n6315), .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6001), .ZN(n6006) );
  OAI211_X1 U7090 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n6004), .B(n6003), .ZN(n6005) );
  NAND3_X1 U7091 ( .A1(n6007), .A2(n6006), .A3(n6005), .ZN(U3002) );
  AOI21_X1 U7092 ( .B1(n6009), .B2(n6310), .A(n6008), .ZN(n6018) );
  AND2_X1 U7093 ( .A1(n6011), .A2(n6010), .ZN(n6013) );
  OAI21_X1 U7094 ( .B1(n6014), .B2(n6013), .A(n6012), .ZN(n6015) );
  AOI22_X1 U7095 ( .A1(n6016), .A2(n6315), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6015), .ZN(n6017) );
  OAI211_X1 U7096 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6019), .A(n6018), .B(n6017), .ZN(U3004) );
  NAND4_X1 U7097 ( .A1(n6128), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n6023)
         );
  OAI21_X1 U7098 ( .B1(n6025), .B2(n6024), .A(n6023), .ZN(U3455) );
  INV_X1 U7099 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6952) );
  OAI21_X1 U7100 ( .B1(n6952), .B2(STATE_REG_2__SCAN_IN), .A(
        STATE_REG_0__SCAN_IN), .ZN(n6031) );
  NOR2_X2 U7101 ( .A1(STATE_REG_0__SCAN_IN), .A2(n6952), .ZN(n6712) );
  INV_X2 U7102 ( .A(n6712), .ZN(n6685) );
  OAI21_X1 U7103 ( .B1(n6031), .B2(ADS_N_REG_SCAN_IN), .A(n6685), .ZN(n6026)
         );
  INV_X1 U7104 ( .A(n6026), .ZN(U2789) );
  OAI21_X1 U7105 ( .B1(n6027), .B2(n6617), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6028) );
  OAI21_X1 U7106 ( .B1(n6029), .B2(n6611), .A(n6028), .ZN(U2790) );
  NOR2_X1 U7107 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n6032) );
  OAI21_X1 U7108 ( .B1(D_C_N_REG_SCAN_IN), .B2(n6032), .A(n6685), .ZN(n6030)
         );
  OAI21_X1 U7109 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6685), .A(n6030), .ZN(
        U2791) );
  NAND2_X1 U7110 ( .A1(n6685), .A2(n6031), .ZN(n6627) );
  INV_X1 U7111 ( .A(n6627), .ZN(n6690) );
  OAI21_X1 U7112 ( .B1(n6032), .B2(BS16_N), .A(n6690), .ZN(n6688) );
  OAI21_X1 U7113 ( .B1(n6690), .B2(n6033), .A(n6688), .ZN(U2792) );
  OAI21_X1 U7114 ( .B1(n6036), .B2(n6035), .A(n6034), .ZN(U2793) );
  NOR4_X1 U7115 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_3__SCAN_IN), .ZN(n6046) );
  NOR4_X1 U7116 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(
        n6045) );
  AOI211_X1 U7117 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_24__SCAN_IN), .B(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6037) );
  INV_X1 U7118 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6896) );
  INV_X1 U7119 ( .A(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6626) );
  NAND3_X1 U7120 ( .A1(n6037), .A2(n6896), .A3(n6626), .ZN(n6043) );
  NOR4_X1 U7121 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAWIDTH_REG_19__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U7122 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAWIDTH_REG_11__SCAN_IN), .ZN(
        n6040) );
  NOR4_X1 U7123 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6039) );
  NOR4_X1 U7124 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6038) );
  NAND4_X1 U7125 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n6042)
         );
  NOR4_X1 U7126 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(n6043), .A4(n6042), .ZN(n6044) );
  NAND3_X1 U7127 ( .A1(n6046), .A2(n6045), .A3(n6044), .ZN(n6700) );
  INV_X1 U7128 ( .A(n6700), .ZN(n6697) );
  INV_X1 U7129 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6689) );
  NAND2_X1 U7130 ( .A1(n6697), .A2(n6689), .ZN(n6050) );
  NOR3_X1 U7131 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(n6050), .ZN(n6047) );
  AOI21_X1 U7132 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6700), .A(n6047), .ZN(
        n6048) );
  OAI21_X1 U7133 ( .B1(n6815), .B2(n6700), .A(n6048), .ZN(U2794) );
  INV_X1 U7134 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6052) );
  NOR2_X1 U7135 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .ZN(n6049) );
  NOR2_X1 U7136 ( .A1(n6049), .A2(n6815), .ZN(n6051) );
  OAI22_X1 U7137 ( .A1(n6697), .A2(n6052), .B1(n6051), .B2(n6050), .ZN(U2795)
         );
  AOI22_X1 U7138 ( .A1(n6053), .A2(n6143), .B1(PHYADDRPOINTER_REG_12__SCAN_IN), 
        .B2(n6142), .ZN(n6064) );
  INV_X1 U7139 ( .A(n6054), .ZN(n6056) );
  NOR2_X1 U7140 ( .A1(n6056), .A2(n6055), .ZN(n6059) );
  NOR2_X1 U7141 ( .A1(n6057), .A2(n6072), .ZN(n6058) );
  AOI211_X1 U7142 ( .C1(n3126), .C2(EBX_REG_12__SCAN_IN), .A(n6059), .B(n6058), 
        .ZN(n6063) );
  AOI22_X1 U7143 ( .A1(n6061), .A2(n6094), .B1(n6108), .B2(n6060), .ZN(n6062)
         );
  NAND4_X1 U7144 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6232), .ZN(U2815)
         );
  AOI21_X1 U7145 ( .B1(n6121), .B2(n6065), .A(REIP_REG_11__SCAN_IN), .ZN(n6073) );
  OAI22_X1 U7146 ( .A1(n6234), .A2(n6115), .B1(n6746), .B2(n6117), .ZN(n6066)
         );
  AOI211_X1 U7147 ( .C1(n3126), .C2(EBX_REG_11__SCAN_IN), .A(n6308), .B(n6066), 
        .ZN(n6071) );
  OAI22_X1 U7148 ( .A1(n6068), .A2(n6105), .B1(n6067), .B2(n6146), .ZN(n6069)
         );
  INV_X1 U7149 ( .A(n6069), .ZN(n6070) );
  OAI211_X1 U7150 ( .C1(n6073), .C2(n6072), .A(n6071), .B(n6070), .ZN(U2816)
         );
  INV_X1 U7151 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6730) );
  NAND2_X1 U7152 ( .A1(n5182), .A2(n6730), .ZN(n6075) );
  NAND4_X1 U7153 ( .A1(n6121), .A2(n6076), .A3(n6075), .A4(n6074), .ZN(n6077)
         );
  OAI21_X1 U7154 ( .B1(n6078), .B2(n6115), .A(n6077), .ZN(n6079) );
  INV_X1 U7155 ( .A(n6079), .ZN(n6087) );
  AOI22_X1 U7156 ( .A1(EBX_REG_10__SCAN_IN), .A2(n3126), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6142), .ZN(n6086) );
  AOI21_X1 U7157 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6080), .A(n6308), .ZN(n6085) );
  INV_X1 U7158 ( .A(n6081), .ZN(n6083) );
  AOI22_X1 U7159 ( .A1(n6083), .A2(n6094), .B1(n6108), .B2(n6082), .ZN(n6084)
         );
  NAND4_X1 U7160 ( .A1(n6087), .A2(n6086), .A3(n6085), .A4(n6084), .ZN(U2817)
         );
  INV_X1 U7161 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7162 ( .B1(n6117), .B2(n6088), .A(n6232), .ZN(n6091) );
  NOR3_X1 U7163 ( .A1(n6098), .A2(REIP_REG_7__SCAN_IN), .A3(n6089), .ZN(n6090)
         );
  AOI211_X1 U7164 ( .C1(EBX_REG_7__SCAN_IN), .C2(n3126), .A(n6091), .B(n6090), 
        .ZN(n6092) );
  OAI21_X1 U7165 ( .B1(n6256), .B2(n6115), .A(n6092), .ZN(n6093) );
  AOI21_X1 U7166 ( .B1(n6202), .B2(n6094), .A(n6093), .ZN(n6100) );
  INV_X1 U7167 ( .A(n6097), .ZN(n6095) );
  NOR3_X1 U7168 ( .A1(n6098), .A2(REIP_REG_6__SCAN_IN), .A3(n6095), .ZN(n6101)
         );
  OAI21_X1 U7169 ( .B1(n6098), .B2(n6097), .A(n6096), .ZN(n6123) );
  OAI21_X1 U7170 ( .B1(n6101), .B2(n6123), .A(REIP_REG_7__SCAN_IN), .ZN(n6099)
         );
  OAI211_X1 U7171 ( .C1(n6146), .C2(n6205), .A(n6100), .B(n6099), .ZN(U2820)
         );
  AOI21_X1 U7172 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6123), .A(n6101), .ZN(n6111)
         );
  NOR2_X1 U7173 ( .A1(n6115), .A2(n6102), .ZN(n6103) );
  AOI211_X1 U7174 ( .C1(n6142), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6308), 
        .B(n6103), .ZN(n6104) );
  OAI21_X1 U7175 ( .B1(n6106), .B2(n6105), .A(n6104), .ZN(n6107) );
  AOI21_X1 U7176 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(n6110) );
  OAI211_X1 U7177 ( .C1(n6112), .C2(n6140), .A(n6111), .B(n6110), .ZN(U2821)
         );
  XNOR2_X1 U7178 ( .A(n6114), .B(n6113), .ZN(n6277) );
  NOR2_X1 U7179 ( .A1(n6115), .A2(n6277), .ZN(n6119) );
  INV_X1 U7180 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U7181 ( .A1(n3126), .A2(EBX_REG_5__SCAN_IN), .ZN(n6116) );
  OAI211_X1 U7182 ( .C1(n6987), .C2(n6117), .A(n6116), .B(n6232), .ZN(n6118)
         );
  NOR2_X1 U7183 ( .A1(n6119), .A2(n6118), .ZN(n6126) );
  INV_X1 U7184 ( .A(n6130), .ZN(n6120) );
  NAND2_X1 U7185 ( .A1(n6121), .A2(n6120), .ZN(n6132) );
  OAI21_X1 U7186 ( .B1(n6132), .B2(n6934), .A(n6648), .ZN(n6122) );
  AOI22_X1 U7187 ( .A1(n6210), .A2(n6124), .B1(n6123), .B2(n6122), .ZN(n6125)
         );
  OAI211_X1 U7188 ( .C1(n6213), .C2(n6146), .A(n6126), .B(n6125), .ZN(U2822)
         );
  AOI22_X1 U7189 ( .A1(n6128), .A2(n6127), .B1(n6143), .B2(n6290), .ZN(n6139)
         );
  OAI21_X1 U7190 ( .B1(n6131), .B2(n6130), .A(n6129), .ZN(n6154) );
  OAI221_X1 U7191 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6132), .C1(n6934), .C2(
        n6154), .A(n6232), .ZN(n6137) );
  INV_X1 U7192 ( .A(n6133), .ZN(n6134) );
  OAI22_X1 U7193 ( .A1(n6135), .A2(n6147), .B1(n6134), .B2(n6146), .ZN(n6136)
         );
  AOI211_X1 U7194 ( .C1(PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n6142), .A(n6137), 
        .B(n6136), .ZN(n6138) );
  OAI211_X1 U7195 ( .C1(n6827), .C2(n6140), .A(n6139), .B(n6138), .ZN(U2823)
         );
  INV_X1 U7196 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6928) );
  NAND2_X1 U7197 ( .A1(n6141), .A2(REIP_REG_2__SCAN_IN), .ZN(n6153) );
  AOI22_X1 U7198 ( .A1(n6143), .A2(n6299), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6142), .ZN(n6144) );
  OAI21_X1 U7199 ( .B1(n6418), .B2(n6145), .A(n6144), .ZN(n6150) );
  OAI22_X1 U7200 ( .A1(n6148), .A2(n6147), .B1(n6221), .B2(n6146), .ZN(n6149)
         );
  AOI211_X1 U7201 ( .C1(EBX_REG_3__SCAN_IN), .C2(n3126), .A(n6150), .B(n6149), 
        .ZN(n6152) );
  OAI221_X1 U7202 ( .B1(n6154), .B2(n6928), .C1(n6154), .C2(n6153), .A(n6152), 
        .ZN(U2824) );
  NOR2_X1 U7203 ( .A1(n6155), .A2(n6277), .ZN(n6156) );
  AOI21_X1 U7204 ( .B1(n6210), .B2(n6160), .A(n6156), .ZN(n6157) );
  OAI21_X1 U7205 ( .B1(n6163), .B2(n6158), .A(n6157), .ZN(U2854) );
  AOI22_X1 U7206 ( .A1(n6227), .A2(n6160), .B1(n6159), .B2(n6309), .ZN(n6161)
         );
  OAI21_X1 U7207 ( .B1(n6163), .B2(n6162), .A(n6161), .ZN(U2857) );
  AOI22_X1 U7208 ( .A1(n6166), .A2(n6165), .B1(n6164), .B2(DATAI_17_), .ZN(
        n6170) );
  AOI22_X1 U7209 ( .A1(n6168), .A2(DATAI_1_), .B1(n6167), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7210 ( .A1(n6170), .A2(n6169), .ZN(U2874) );
  AOI22_X1 U7211 ( .A1(n6195), .A2(LWORD_REG_15__SCAN_IN), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n5847), .ZN(n6171) );
  OAI21_X1 U7212 ( .B1(n6172), .B2(n6197), .A(n6171), .ZN(U2908) );
  AOI22_X1 U7213 ( .A1(n6195), .A2(LWORD_REG_14__SCAN_IN), .B1(
        DATAO_REG_14__SCAN_IN), .B2(n5847), .ZN(n6173) );
  OAI21_X1 U7214 ( .B1(n6795), .B2(n6197), .A(n6173), .ZN(U2909) );
  AOI22_X1 U7215 ( .A1(n6195), .A2(LWORD_REG_13__SCAN_IN), .B1(
        DATAO_REG_13__SCAN_IN), .B2(n5847), .ZN(n6174) );
  OAI21_X1 U7216 ( .B1(n6716), .B2(n6197), .A(n6174), .ZN(U2910) );
  AOI22_X1 U7217 ( .A1(n6195), .A2(LWORD_REG_12__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6175) );
  OAI21_X1 U7218 ( .B1(n6176), .B2(n6197), .A(n6175), .ZN(U2911) );
  AOI22_X1 U7219 ( .A1(n6195), .A2(LWORD_REG_11__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6177) );
  OAI21_X1 U7220 ( .B1(n6178), .B2(n6197), .A(n6177), .ZN(U2912) );
  AOI22_X1 U7221 ( .A1(n6195), .A2(LWORD_REG_10__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U7222 ( .B1(n6180), .B2(n6197), .A(n6179), .ZN(U2913) );
  AOI22_X1 U7223 ( .A1(n6195), .A2(LWORD_REG_9__SCAN_IN), .B1(
        DATAO_REG_9__SCAN_IN), .B2(n5847), .ZN(n6181) );
  OAI21_X1 U7224 ( .B1(n6182), .B2(n6197), .A(n6181), .ZN(U2914) );
  AOI22_X1 U7225 ( .A1(n6195), .A2(LWORD_REG_8__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6183) );
  OAI21_X1 U7226 ( .B1(n6184), .B2(n6197), .A(n6183), .ZN(U2915) );
  INV_X1 U7227 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7228 ( .A1(EAX_REG_7__SCAN_IN), .A2(n6185), .B1(n5847), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U7229 ( .B1(n6604), .B2(n6753), .A(n6186), .ZN(U2916) );
  AOI22_X1 U7230 ( .A1(n6195), .A2(LWORD_REG_6__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6187) );
  OAI21_X1 U7231 ( .B1(n3735), .B2(n6197), .A(n6187), .ZN(U2917) );
  AOI22_X1 U7232 ( .A1(n6195), .A2(LWORD_REG_5__SCAN_IN), .B1(
        DATAO_REG_5__SCAN_IN), .B2(n5847), .ZN(n6188) );
  OAI21_X1 U7233 ( .B1(n4766), .B2(n6197), .A(n6188), .ZN(U2918) );
  AOI22_X1 U7234 ( .A1(n6195), .A2(LWORD_REG_4__SCAN_IN), .B1(
        DATAO_REG_4__SCAN_IN), .B2(n5847), .ZN(n6189) );
  OAI21_X1 U7235 ( .B1(n6190), .B2(n6197), .A(n6189), .ZN(U2919) );
  AOI22_X1 U7236 ( .A1(n6195), .A2(LWORD_REG_3__SCAN_IN), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n5847), .ZN(n6191) );
  OAI21_X1 U7237 ( .B1(n3776), .B2(n6197), .A(n6191), .ZN(U2920) );
  AOI22_X1 U7238 ( .A1(n6195), .A2(LWORD_REG_2__SCAN_IN), .B1(n5847), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6192) );
  OAI21_X1 U7239 ( .B1(n6193), .B2(n6197), .A(n6192), .ZN(U2921) );
  AOI22_X1 U7240 ( .A1(n6195), .A2(LWORD_REG_1__SCAN_IN), .B1(
        DATAO_REG_1__SCAN_IN), .B2(n5847), .ZN(n6194) );
  OAI21_X1 U7241 ( .B1(n3741), .B2(n6197), .A(n6194), .ZN(U2922) );
  AOI22_X1 U7242 ( .A1(n6195), .A2(LWORD_REG_0__SCAN_IN), .B1(
        DATAO_REG_0__SCAN_IN), .B2(n5847), .ZN(n6196) );
  OAI21_X1 U7243 ( .B1(n3748), .B2(n6197), .A(n6196), .ZN(U2923) );
  AOI22_X1 U7244 ( .A1(n6308), .A2(REIP_REG_7__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6204) );
  OAI21_X1 U7245 ( .B1(n6200), .B2(n6199), .A(n6198), .ZN(n6201) );
  INV_X1 U7246 ( .A(n6201), .ZN(n6259) );
  AOI22_X1 U7247 ( .A1(n6259), .A2(n4529), .B1(n6226), .B2(n6202), .ZN(n6203)
         );
  OAI211_X1 U7248 ( .C1(n6231), .C2(n6205), .A(n6204), .B(n6203), .ZN(U2979)
         );
  AOI22_X1 U7249 ( .A1(n6308), .A2(REIP_REG_5__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6212) );
  OR2_X1 U7250 ( .A1(n6207), .A2(n6206), .ZN(n6208) );
  AND2_X1 U7251 ( .A1(n6209), .A2(n6208), .ZN(n6280) );
  AOI22_X1 U7252 ( .A1(n6280), .A2(n4529), .B1(n6226), .B2(n6210), .ZN(n6211)
         );
  OAI211_X1 U7253 ( .C1(n6231), .C2(n6213), .A(n6212), .B(n6211), .ZN(U2981)
         );
  AOI22_X1 U7254 ( .A1(n6308), .A2(REIP_REG_3__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6220) );
  OR2_X1 U7255 ( .A1(n6215), .A2(n6214), .ZN(n6217) );
  AND2_X1 U7256 ( .A1(n6217), .A2(n6216), .ZN(n6300) );
  AOI22_X1 U7257 ( .A1(n6218), .A2(n6226), .B1(n4529), .B2(n6300), .ZN(n6219)
         );
  OAI211_X1 U7258 ( .C1(n6231), .C2(n6221), .A(n6220), .B(n6219), .ZN(U2983)
         );
  AOI22_X1 U7259 ( .A1(n6308), .A2(REIP_REG_2__SCAN_IN), .B1(n6222), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6229) );
  XOR2_X1 U7260 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(n6223), .Z(n6224) );
  XNOR2_X1 U7261 ( .A(n6225), .B(n6224), .ZN(n6314) );
  AOI22_X1 U7262 ( .A1(n6314), .A2(n4529), .B1(n6227), .B2(n6226), .ZN(n6228)
         );
  OAI211_X1 U7263 ( .C1(n6231), .C2(n6230), .A(n6229), .B(n6228), .ZN(U2984)
         );
  OAI22_X1 U7264 ( .A1(n6234), .A2(n6233), .B1(n5293), .B2(n6232), .ZN(n6235)
         );
  AOI21_X1 U7265 ( .B1(n6315), .B2(n6236), .A(n6235), .ZN(n6237) );
  OAI221_X1 U7266 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n6239), .C1(
        n6970), .C2(n6238), .A(n6237), .ZN(U3007) );
  AOI21_X1 U7267 ( .B1(n6241), .B2(n6310), .A(n6240), .ZN(n6245) );
  AOI22_X1 U7268 ( .A1(n6243), .A2(n6315), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6242), .ZN(n6244) );
  OAI211_X1 U7269 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6246), .A(n6245), 
        .B(n6244), .ZN(U3009) );
  AOI21_X1 U7270 ( .B1(n6248), .B2(n6310), .A(n6247), .ZN(n6254) );
  INV_X1 U7271 ( .A(n6249), .ZN(n6252) );
  AOI21_X1 U7272 ( .B1(n6262), .B2(n6255), .A(n6250), .ZN(n6251) );
  AOI22_X1 U7273 ( .A1(n6252), .A2(n6315), .B1(n6258), .B2(n6251), .ZN(n6253)
         );
  OAI211_X1 U7274 ( .C1(n6263), .C2(n6255), .A(n6254), .B(n6253), .ZN(U3010)
         );
  INV_X1 U7275 ( .A(n6256), .ZN(n6257) );
  AOI22_X1 U7276 ( .A1(n6257), .A2(n6310), .B1(n6308), .B2(REIP_REG_7__SCAN_IN), .ZN(n6261) );
  AOI22_X1 U7277 ( .A1(n6259), .A2(n6315), .B1(n6258), .B2(n6262), .ZN(n6260)
         );
  OAI211_X1 U7278 ( .C1(n6263), .C2(n6262), .A(n6261), .B(n6260), .ZN(U3011)
         );
  NAND2_X1 U7279 ( .A1(n6271), .A2(n6264), .ZN(n6276) );
  AOI21_X1 U7280 ( .B1(n6266), .B2(n6310), .A(n6265), .ZN(n6275) );
  INV_X1 U7281 ( .A(n6284), .ZN(n6307) );
  INV_X1 U7282 ( .A(n6267), .ZN(n6268) );
  AOI21_X1 U7283 ( .B1(n6269), .B2(n6307), .A(n6268), .ZN(n6321) );
  OAI21_X1 U7284 ( .B1(n6271), .B2(n6270), .A(n6321), .ZN(n6282) );
  INV_X1 U7285 ( .A(n6272), .ZN(n6273) );
  AOI22_X1 U7286 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n6282), .B1(n6273), 
        .B2(n6315), .ZN(n6274) );
  OAI211_X1 U7287 ( .C1(n6288), .C2(n6276), .A(n6275), .B(n6274), .ZN(U3012)
         );
  INV_X1 U7288 ( .A(n6277), .ZN(n6278) );
  AOI22_X1 U7289 ( .A1(n6278), .A2(n6310), .B1(n6308), .B2(REIP_REG_5__SCAN_IN), .ZN(n6287) );
  OAI21_X1 U7290 ( .B1(n6291), .B2(n6279), .A(n6283), .ZN(n6281) );
  AOI22_X1 U7291 ( .A1(n6282), .A2(n6281), .B1(n6315), .B2(n6280), .ZN(n6286)
         );
  NAND4_X1 U7292 ( .A1(n6297), .A2(n6317), .A3(n6284), .A4(n6283), .ZN(n6285)
         );
  NAND3_X1 U7293 ( .A1(n6287), .A2(n6286), .A3(n6285), .ZN(U3013) );
  INV_X1 U7294 ( .A(n6288), .ZN(n6298) );
  OAI211_X1 U7295 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n6298), .B(n6305), .ZN(n6296) );
  AOI21_X1 U7296 ( .B1(n6290), .B2(n6310), .A(n6289), .ZN(n6295) );
  OAI21_X1 U7297 ( .B1(n6305), .B2(n6291), .A(n6321), .ZN(n6301) );
  INV_X1 U7298 ( .A(n6292), .ZN(n6293) );
  AOI22_X1 U7299 ( .A1(n6301), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n6315), 
        .B2(n6293), .ZN(n6294) );
  OAI211_X1 U7300 ( .C1(n6297), .C2(n6296), .A(n6295), .B(n6294), .ZN(U3014)
         );
  NAND2_X1 U7301 ( .A1(n6305), .A2(n6298), .ZN(n6304) );
  AOI22_X1 U7302 ( .A1(n6299), .A2(n6310), .B1(n6308), .B2(REIP_REG_3__SCAN_IN), .ZN(n6303) );
  AOI22_X1 U7303 ( .A1(n6301), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6315), 
        .B2(n6300), .ZN(n6302) );
  OAI211_X1 U7304 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n6304), .A(n6303), 
        .B(n6302), .ZN(U3015) );
  OAI21_X1 U7305 ( .B1(n6307), .B2(n6306), .A(n6305), .ZN(n6312) );
  AOI222_X1 U7306 ( .A1(n6312), .A2(n6311), .B1(n6310), .B2(n6309), .C1(
        REIP_REG_2__SCAN_IN), .C2(n6308), .ZN(n6319) );
  NOR2_X1 U7307 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6313), .ZN(n6316)
         );
  AOI22_X1 U7308 ( .A1(n6317), .A2(n6316), .B1(n6315), .B2(n6314), .ZN(n6318)
         );
  OAI211_X1 U7309 ( .C1(n6321), .C2(n6320), .A(n6319), .B(n6318), .ZN(U3016)
         );
  NOR2_X1 U7310 ( .A1(n6323), .A2(n6322), .ZN(U3019) );
  INV_X1 U7311 ( .A(n6324), .ZN(n6454) );
  NAND2_X1 U7312 ( .A1(n6454), .A2(n6325), .ZN(n6330) );
  INV_X1 U7313 ( .A(n6330), .ZN(n6354) );
  AOI22_X1 U7314 ( .A1(n6561), .A2(n6354), .B1(n6564), .B2(n6353), .ZN(n6338)
         );
  NAND2_X1 U7315 ( .A1(n6326), .A2(n4754), .ZN(n6327) );
  OAI21_X1 U7316 ( .B1(n6328), .B2(n6327), .A(n6456), .ZN(n6336) );
  OR2_X1 U7317 ( .A1(n6329), .A2(n6378), .ZN(n6331) );
  NAND2_X1 U7318 ( .A1(n6331), .A2(n6330), .ZN(n6333) );
  AOI21_X1 U7319 ( .B1(n6334), .B2(n6499), .A(n6462), .ZN(n6332) );
  OAI21_X1 U7320 ( .B1(n6336), .B2(n6333), .A(n6332), .ZN(n6356) );
  INV_X1 U7321 ( .A(n6333), .ZN(n6335) );
  OAI22_X1 U7322 ( .A1(n6336), .A2(n6335), .B1(n6334), .B2(n6465), .ZN(n6355)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6356), .B1(n6560), 
        .B2(n6355), .ZN(n6337) );
  OAI211_X1 U7324 ( .C1(n6471), .C2(n6359), .A(n6338), .B(n6337), .ZN(U3044)
         );
  AOI22_X1 U7325 ( .A1(n6515), .A2(n6354), .B1(n6517), .B2(n6353), .ZN(n6340)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6356), .B1(n6514), 
        .B2(n6355), .ZN(n6339) );
  OAI211_X1 U7327 ( .C1(n6359), .C2(n6426), .A(n6340), .B(n6339), .ZN(U3045)
         );
  AOI22_X1 U7328 ( .A1(n6521), .A2(n6354), .B1(n6524), .B2(n6353), .ZN(n6342)
         );
  AOI22_X1 U7329 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6356), .B1(n6522), 
        .B2(n6355), .ZN(n6341) );
  OAI211_X1 U7330 ( .C1(n6359), .C2(n6477), .A(n6342), .B(n6341), .ZN(U3046)
         );
  AOI22_X1 U7331 ( .A1(n6529), .A2(n6354), .B1(n6530), .B2(n6349), .ZN(n6344)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6356), .B1(n6528), 
        .B2(n6355), .ZN(n6343) );
  OAI211_X1 U7333 ( .C1(n6480), .C2(n6370), .A(n6344), .B(n6343), .ZN(U3047)
         );
  AOI22_X1 U7334 ( .A1(n6536), .A2(n6354), .B1(n6538), .B2(n6353), .ZN(n6346)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6356), .B1(n6535), 
        .B2(n6355), .ZN(n6345) );
  OAI211_X1 U7336 ( .C1(n6359), .C2(n6434), .A(n6346), .B(n6345), .ZN(U3048)
         );
  AOI22_X1 U7337 ( .A1(n6568), .A2(n6354), .B1(n6573), .B2(n6353), .ZN(n6348)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6356), .B1(n6570), 
        .B2(n6355), .ZN(n6347) );
  OAI211_X1 U7339 ( .C1(n6359), .C2(n6488), .A(n6348), .B(n6347), .ZN(U3049)
         );
  AOI22_X1 U7340 ( .A1(n6544), .A2(n6354), .B1(n6545), .B2(n6349), .ZN(n6351)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6356), .B1(n6543), 
        .B2(n6355), .ZN(n6350) );
  OAI211_X1 U7342 ( .C1(n6352), .C2(n6370), .A(n6351), .B(n6350), .ZN(U3050)
         );
  AOI22_X1 U7343 ( .A1(n7041), .A2(n6354), .B1(n6555), .B2(n6353), .ZN(n6358)
         );
  AOI22_X1 U7344 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6356), .B1(n6550), 
        .B2(n6355), .ZN(n6357) );
  OAI211_X1 U7345 ( .C1(n6359), .C2(n7038), .A(n6358), .B(n6357), .ZN(U3051)
         );
  AOI22_X1 U7346 ( .A1(n6561), .A2(n6364), .B1(n6560), .B2(n6365), .ZN(n6361)
         );
  AOI22_X1 U7347 ( .A1(n6367), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n6564), 
        .B2(n6366), .ZN(n6360) );
  OAI211_X1 U7348 ( .C1(n6471), .C2(n6370), .A(n6361), .B(n6360), .ZN(U3052)
         );
  AOI22_X1 U7349 ( .A1(n6536), .A2(n6364), .B1(n6535), .B2(n6365), .ZN(n6363)
         );
  AOI22_X1 U7350 ( .A1(n6367), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n6538), 
        .B2(n6366), .ZN(n6362) );
  OAI211_X1 U7351 ( .C1(n6434), .C2(n6370), .A(n6363), .B(n6362), .ZN(U3056)
         );
  AOI22_X1 U7352 ( .A1(n6570), .A2(n6365), .B1(n6568), .B2(n6364), .ZN(n6369)
         );
  AOI22_X1 U7353 ( .A1(n6367), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n6573), 
        .B2(n6366), .ZN(n6368) );
  OAI211_X1 U7354 ( .C1(n6488), .C2(n6370), .A(n6369), .B(n6368), .ZN(U3057)
         );
  INV_X1 U7355 ( .A(n6377), .ZN(n6401) );
  NOR2_X1 U7356 ( .A1(n6371), .A2(n3745), .ZN(n6373) );
  AOI22_X1 U7357 ( .A1(n6561), .A2(n6401), .B1(n6564), .B2(n6416), .ZN(n6385)
         );
  NAND2_X1 U7358 ( .A1(n6456), .A2(n6383), .ZN(n6374) );
  NAND2_X1 U7359 ( .A1(n6374), .A2(n6381), .ZN(n6375) );
  NAND2_X1 U7360 ( .A1(n6376), .A2(n6375), .ZN(n6403) );
  OAI21_X1 U7361 ( .B1(n6379), .B2(n6378), .A(n6377), .ZN(n6380) );
  NAND2_X1 U7362 ( .A1(n6380), .A2(n6456), .ZN(n6382) );
  OAI22_X1 U7363 ( .A1(n6383), .A2(n6382), .B1(n6381), .B2(n6465), .ZN(n6402)
         );
  AOI22_X1 U7364 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6403), .B1(n6560), 
        .B2(n6402), .ZN(n6384) );
  OAI211_X1 U7365 ( .C1(n6471), .C2(n6406), .A(n6385), .B(n6384), .ZN(U3076)
         );
  AOI22_X1 U7366 ( .A1(n6515), .A2(n6401), .B1(n6517), .B2(n6416), .ZN(n6387)
         );
  AOI22_X1 U7367 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6403), .B1(n6514), 
        .B2(n6402), .ZN(n6386) );
  OAI211_X1 U7368 ( .C1(n6426), .C2(n6406), .A(n6387), .B(n6386), .ZN(U3077)
         );
  INV_X1 U7369 ( .A(n6406), .ZN(n6395) );
  AOI22_X1 U7370 ( .A1(n6521), .A2(n6401), .B1(n6523), .B2(n6395), .ZN(n6389)
         );
  AOI22_X1 U7371 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6403), .B1(n6522), 
        .B2(n6402), .ZN(n6388) );
  OAI211_X1 U7372 ( .C1(n6390), .C2(n6444), .A(n6389), .B(n6388), .ZN(U3078)
         );
  AOI22_X1 U7373 ( .A1(n6529), .A2(n6401), .B1(n6531), .B2(n6416), .ZN(n6392)
         );
  AOI22_X1 U7374 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6403), .B1(n6528), 
        .B2(n6402), .ZN(n6391) );
  OAI211_X1 U7375 ( .C1(n6431), .C2(n6406), .A(n6392), .B(n6391), .ZN(U3079)
         );
  AOI22_X1 U7376 ( .A1(n6536), .A2(n6401), .B1(n6537), .B2(n6395), .ZN(n6394)
         );
  AOI22_X1 U7377 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6403), .B1(n6535), 
        .B2(n6402), .ZN(n6393) );
  OAI211_X1 U7378 ( .C1(n6485), .C2(n6444), .A(n6394), .B(n6393), .ZN(U3080)
         );
  AOI22_X1 U7379 ( .A1(n6568), .A2(n6401), .B1(n6571), .B2(n6395), .ZN(n6397)
         );
  AOI22_X1 U7380 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6403), .B1(n6570), 
        .B2(n6402), .ZN(n6396) );
  OAI211_X1 U7381 ( .C1(n6398), .C2(n6444), .A(n6397), .B(n6396), .ZN(U3081)
         );
  AOI22_X1 U7382 ( .A1(n6544), .A2(n6401), .B1(n6546), .B2(n6416), .ZN(n6400)
         );
  AOI22_X1 U7383 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6403), .B1(n6543), 
        .B2(n6402), .ZN(n6399) );
  OAI211_X1 U7384 ( .C1(n6491), .C2(n6406), .A(n6400), .B(n6399), .ZN(U3082)
         );
  AOI22_X1 U7385 ( .A1(n7041), .A2(n6401), .B1(n6555), .B2(n6416), .ZN(n6405)
         );
  AOI22_X1 U7386 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6403), .B1(n6550), 
        .B2(n6402), .ZN(n6404) );
  OAI211_X1 U7387 ( .C1(n7038), .C2(n6406), .A(n6405), .B(n6404), .ZN(U3083)
         );
  NOR2_X1 U7388 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6407), .ZN(n6440)
         );
  INV_X1 U7389 ( .A(n6408), .ZN(n6511) );
  OR2_X1 U7390 ( .A1(n6410), .A2(n6409), .ZN(n6508) );
  OAI22_X1 U7391 ( .A1(n6511), .A2(n6417), .B1(n6504), .B2(n6508), .ZN(n6439)
         );
  AOI22_X1 U7392 ( .A1(n6561), .A2(n6440), .B1(n6560), .B2(n6439), .ZN(n6423)
         );
  INV_X1 U7393 ( .A(n6440), .ZN(n6414) );
  INV_X1 U7394 ( .A(n6508), .ZN(n6412) );
  OAI21_X1 U7395 ( .B1(n6412), .B2(n5022), .A(n6411), .ZN(n6507) );
  AOI211_X1 U7396 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6414), .A(n6413), .B(
        n6507), .ZN(n6421) );
  NOR3_X1 U7397 ( .A1(n6447), .A2(n6416), .A3(n6499), .ZN(n6419) );
  OAI22_X1 U7398 ( .A1(n6419), .A2(n6502), .B1(n6418), .B2(n6417), .ZN(n6420)
         );
  NAND2_X1 U7399 ( .A1(n6421), .A2(n6420), .ZN(n6441) );
  AOI22_X1 U7400 ( .A1(n6441), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6564), 
        .B2(n6447), .ZN(n6422) );
  OAI211_X1 U7401 ( .C1(n6471), .C2(n6444), .A(n6423), .B(n6422), .ZN(U3084)
         );
  AOI22_X1 U7402 ( .A1(n6515), .A2(n6440), .B1(n6514), .B2(n6439), .ZN(n6425)
         );
  AOI22_X1 U7403 ( .A1(n6441), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6517), 
        .B2(n6447), .ZN(n6424) );
  OAI211_X1 U7404 ( .C1(n6426), .C2(n6444), .A(n6425), .B(n6424), .ZN(U3085)
         );
  AOI22_X1 U7405 ( .A1(n6522), .A2(n6439), .B1(n6521), .B2(n6440), .ZN(n6428)
         );
  AOI22_X1 U7406 ( .A1(n6441), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6524), 
        .B2(n6447), .ZN(n6427) );
  OAI211_X1 U7407 ( .C1(n6477), .C2(n6444), .A(n6428), .B(n6427), .ZN(U3086)
         );
  AOI22_X1 U7408 ( .A1(n6529), .A2(n6440), .B1(n6528), .B2(n6439), .ZN(n6430)
         );
  AOI22_X1 U7409 ( .A1(n6441), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6531), 
        .B2(n6447), .ZN(n6429) );
  OAI211_X1 U7410 ( .C1(n6431), .C2(n6444), .A(n6430), .B(n6429), .ZN(U3087)
         );
  AOI22_X1 U7411 ( .A1(n6536), .A2(n6440), .B1(n6535), .B2(n6439), .ZN(n6433)
         );
  AOI22_X1 U7412 ( .A1(n6441), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6538), 
        .B2(n6447), .ZN(n6432) );
  OAI211_X1 U7413 ( .C1(n6434), .C2(n6444), .A(n6433), .B(n6432), .ZN(U3088)
         );
  AOI22_X1 U7414 ( .A1(n6570), .A2(n6439), .B1(n6568), .B2(n6440), .ZN(n6436)
         );
  AOI22_X1 U7415 ( .A1(n6441), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6573), 
        .B2(n6447), .ZN(n6435) );
  OAI211_X1 U7416 ( .C1(n6488), .C2(n6444), .A(n6436), .B(n6435), .ZN(U3089)
         );
  AOI22_X1 U7417 ( .A1(n6544), .A2(n6440), .B1(n6543), .B2(n6439), .ZN(n6438)
         );
  AOI22_X1 U7418 ( .A1(n6441), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6546), 
        .B2(n6447), .ZN(n6437) );
  OAI211_X1 U7419 ( .C1(n6491), .C2(n6444), .A(n6438), .B(n6437), .ZN(U3090)
         );
  AOI22_X1 U7420 ( .A1(n7041), .A2(n6440), .B1(n6550), .B2(n6439), .ZN(n6443)
         );
  AOI22_X1 U7421 ( .A1(n6441), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6555), 
        .B2(n6447), .ZN(n6442) );
  OAI211_X1 U7422 ( .C1(n7038), .C2(n6444), .A(n6443), .B(n6442), .ZN(U3091)
         );
  INV_X1 U7423 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7424 ( .A1(n6561), .A2(n6448), .B1(n6447), .B2(n6563), .ZN(n6446)
         );
  AOI22_X1 U7425 ( .A1(n6450), .A2(n6560), .B1(n6449), .B2(n6564), .ZN(n6445)
         );
  OAI211_X1 U7426 ( .C1(n6453), .C2(n6756), .A(n6446), .B(n6445), .ZN(U3092)
         );
  INV_X1 U7427 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6729) );
  AOI22_X1 U7428 ( .A1(n6536), .A2(n6448), .B1(n6447), .B2(n6537), .ZN(n6452)
         );
  AOI22_X1 U7429 ( .A1(n6450), .A2(n6535), .B1(n6449), .B2(n6538), .ZN(n6451)
         );
  OAI211_X1 U7430 ( .C1(n6453), .C2(n6729), .A(n6452), .B(n6451), .ZN(U3096)
         );
  NAND2_X1 U7431 ( .A1(n6454), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6460) );
  INV_X1 U7432 ( .A(n6460), .ZN(n6492) );
  AOI22_X1 U7433 ( .A1(n6561), .A2(n6492), .B1(n6564), .B2(n6553), .ZN(n6470)
         );
  OAI21_X1 U7434 ( .B1(n6458), .B2(n6457), .A(n6456), .ZN(n6468) );
  NAND2_X1 U7435 ( .A1(n6459), .A2(n3134), .ZN(n6461) );
  NAND2_X1 U7436 ( .A1(n6461), .A2(n6460), .ZN(n6464) );
  AOI21_X1 U7437 ( .B1(n6466), .B2(n6499), .A(n6462), .ZN(n6463) );
  OAI21_X1 U7438 ( .B1(n6468), .B2(n6464), .A(n6463), .ZN(n6494) );
  INV_X1 U7439 ( .A(n6464), .ZN(n6467) );
  OAI22_X1 U7440 ( .A1(n6468), .A2(n6467), .B1(n6466), .B2(n6465), .ZN(n6493)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6494), .B1(n6560), 
        .B2(n6493), .ZN(n6469) );
  OAI211_X1 U7442 ( .C1(n6471), .C2(n6497), .A(n6470), .B(n6469), .ZN(U3108)
         );
  INV_X1 U7443 ( .A(n6497), .ZN(n6481) );
  AOI22_X1 U7444 ( .A1(n6515), .A2(n6492), .B1(n6481), .B2(n6516), .ZN(n6473)
         );
  AOI22_X1 U7445 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6494), .B1(n6514), 
        .B2(n6493), .ZN(n6472) );
  OAI211_X1 U7446 ( .C1(n6474), .C2(n6484), .A(n6473), .B(n6472), .ZN(U3109)
         );
  AOI22_X1 U7447 ( .A1(n6521), .A2(n6492), .B1(n6524), .B2(n6553), .ZN(n6476)
         );
  AOI22_X1 U7448 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6494), .B1(n6522), 
        .B2(n6493), .ZN(n6475) );
  OAI211_X1 U7449 ( .C1(n6477), .C2(n6497), .A(n6476), .B(n6475), .ZN(U3110)
         );
  AOI22_X1 U7450 ( .A1(n6529), .A2(n6492), .B1(n6481), .B2(n6530), .ZN(n6479)
         );
  AOI22_X1 U7451 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6494), .B1(n6528), 
        .B2(n6493), .ZN(n6478) );
  OAI211_X1 U7452 ( .C1(n6480), .C2(n6484), .A(n6479), .B(n6478), .ZN(U3111)
         );
  AOI22_X1 U7453 ( .A1(n6536), .A2(n6492), .B1(n6481), .B2(n6537), .ZN(n6483)
         );
  AOI22_X1 U7454 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6494), .B1(n6535), 
        .B2(n6493), .ZN(n6482) );
  OAI211_X1 U7455 ( .C1(n6485), .C2(n6484), .A(n6483), .B(n6482), .ZN(U3112)
         );
  AOI22_X1 U7456 ( .A1(n6568), .A2(n6492), .B1(n6573), .B2(n6553), .ZN(n6487)
         );
  AOI22_X1 U7457 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6494), .B1(n6570), 
        .B2(n6493), .ZN(n6486) );
  OAI211_X1 U7458 ( .C1(n6488), .C2(n6497), .A(n6487), .B(n6486), .ZN(U3113)
         );
  AOI22_X1 U7459 ( .A1(n6544), .A2(n6492), .B1(n6546), .B2(n6553), .ZN(n6490)
         );
  AOI22_X1 U7460 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6494), .B1(n6543), 
        .B2(n6493), .ZN(n6489) );
  OAI211_X1 U7461 ( .C1(n6491), .C2(n6497), .A(n6490), .B(n6489), .ZN(U3114)
         );
  AOI22_X1 U7462 ( .A1(n7041), .A2(n6492), .B1(n6555), .B2(n6553), .ZN(n6496)
         );
  AOI22_X1 U7463 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6494), .B1(n6550), 
        .B2(n6493), .ZN(n6495) );
  OAI211_X1 U7464 ( .C1(n7038), .C2(n6497), .A(n6496), .B(n6495), .ZN(U3115)
         );
  NOR2_X1 U7465 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6498), .ZN(n6551)
         );
  NOR3_X1 U7466 ( .A1(n6554), .A2(n6553), .A3(n6499), .ZN(n6503) );
  INV_X1 U7467 ( .A(n6500), .ZN(n6510) );
  OAI22_X1 U7468 ( .A1(n6503), .A2(n6502), .B1(n6501), .B2(n6510), .ZN(n6505)
         );
  OAI211_X1 U7469 ( .C1(n6551), .C2(n6693), .A(n6505), .B(n6504), .ZN(n6506)
         );
  INV_X1 U7470 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n7017) );
  OAI22_X1 U7471 ( .A1(n6511), .A2(n6510), .B1(n6509), .B2(n6508), .ZN(n6549)
         );
  AOI22_X1 U7472 ( .A1(n6561), .A2(n6551), .B1(n6560), .B2(n6549), .ZN(n6513)
         );
  AOI22_X1 U7473 ( .A1(n6564), .A2(n6554), .B1(n6553), .B2(n6563), .ZN(n6512)
         );
  OAI211_X1 U7474 ( .C1(n6559), .C2(n7017), .A(n6513), .B(n6512), .ZN(U3116)
         );
  INV_X1 U7475 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n6520) );
  AOI22_X1 U7476 ( .A1(n6515), .A2(n6551), .B1(n6514), .B2(n6549), .ZN(n6519)
         );
  AOI22_X1 U7477 ( .A1(n6517), .A2(n6554), .B1(n6553), .B2(n6516), .ZN(n6518)
         );
  OAI211_X1 U7478 ( .C1(n6559), .C2(n6520), .A(n6519), .B(n6518), .ZN(U3117)
         );
  INV_X1 U7479 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6527) );
  AOI22_X1 U7480 ( .A1(n6522), .A2(n6549), .B1(n6521), .B2(n6551), .ZN(n6526)
         );
  AOI22_X1 U7481 ( .A1(n6524), .A2(n6554), .B1(n6553), .B2(n6523), .ZN(n6525)
         );
  OAI211_X1 U7482 ( .C1(n6559), .C2(n6527), .A(n6526), .B(n6525), .ZN(U3118)
         );
  INV_X1 U7483 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n6534) );
  AOI22_X1 U7484 ( .A1(n6529), .A2(n6551), .B1(n6528), .B2(n6549), .ZN(n6533)
         );
  AOI22_X1 U7485 ( .A1(n6531), .A2(n6554), .B1(n6553), .B2(n6530), .ZN(n6532)
         );
  OAI211_X1 U7486 ( .C1(n6559), .C2(n6534), .A(n6533), .B(n6532), .ZN(U3119)
         );
  INV_X1 U7487 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n7002) );
  AOI22_X1 U7488 ( .A1(n6536), .A2(n6551), .B1(n6535), .B2(n6549), .ZN(n6540)
         );
  AOI22_X1 U7489 ( .A1(n6538), .A2(n6554), .B1(n6553), .B2(n6537), .ZN(n6539)
         );
  OAI211_X1 U7490 ( .C1(n6559), .C2(n7002), .A(n6540), .B(n6539), .ZN(U3120)
         );
  INV_X1 U7491 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n7000) );
  AOI22_X1 U7492 ( .A1(n6570), .A2(n6549), .B1(n6568), .B2(n6551), .ZN(n6542)
         );
  AOI22_X1 U7493 ( .A1(n6573), .A2(n6554), .B1(n6553), .B2(n6571), .ZN(n6541)
         );
  OAI211_X1 U7494 ( .C1(n6559), .C2(n7000), .A(n6542), .B(n6541), .ZN(U3121)
         );
  INV_X1 U7495 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6994) );
  AOI22_X1 U7496 ( .A1(n6544), .A2(n6551), .B1(n6543), .B2(n6549), .ZN(n6548)
         );
  AOI22_X1 U7497 ( .A1(n6546), .A2(n6554), .B1(n6553), .B2(n6545), .ZN(n6547)
         );
  OAI211_X1 U7498 ( .C1(n6559), .C2(n6994), .A(n6548), .B(n6547), .ZN(U3122)
         );
  INV_X1 U7499 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6558) );
  AOI22_X1 U7500 ( .A1(n7041), .A2(n6551), .B1(n6550), .B2(n6549), .ZN(n6557)
         );
  AOI22_X1 U7501 ( .A1(n6555), .A2(n6554), .B1(n6553), .B2(n6552), .ZN(n6556)
         );
  OAI211_X1 U7502 ( .C1(n6559), .C2(n6558), .A(n6557), .B(n6556), .ZN(U3123)
         );
  INV_X1 U7503 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7504 ( .A1(n6561), .A2(n6567), .B1(n6560), .B2(n6569), .ZN(n6566)
         );
  INV_X1 U7505 ( .A(n6562), .ZN(n6574) );
  AOI22_X1 U7506 ( .A1(n6574), .A2(n6564), .B1(n6572), .B2(n6563), .ZN(n6565)
         );
  OAI211_X1 U7507 ( .C1(n6577), .C2(n6747), .A(n6566), .B(n6565), .ZN(U3140)
         );
  INV_X1 U7508 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7509 ( .A1(n6570), .A2(n6569), .B1(n6568), .B2(n6567), .ZN(n6576)
         );
  AOI22_X1 U7510 ( .A1(n6574), .A2(n6573), .B1(n6572), .B2(n6571), .ZN(n6575)
         );
  OAI211_X1 U7511 ( .C1(n6577), .C2(n6772), .A(n6576), .B(n6575), .ZN(U3145)
         );
  INV_X1 U7512 ( .A(n6578), .ZN(n6588) );
  AOI211_X1 U7513 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6580), .A(n6978), .B(n6579), .ZN(n6586) );
  INV_X1 U7514 ( .A(n6586), .ZN(n6583) );
  OAI211_X1 U7515 ( .C1(n6584), .C2(n6583), .A(n6582), .B(n6581), .ZN(n6585)
         );
  OAI21_X1 U7516 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6586), .A(n6585), 
        .ZN(n6587) );
  AOI222_X1 U7517 ( .A1(n6589), .A2(n6588), .B1(n6589), .B2(n6587), .C1(n6588), 
        .C2(n6587), .ZN(n6591) );
  AOI21_X1 U7518 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6591), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6603) );
  OAI21_X1 U7519 ( .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6591), .A(n6590), 
        .ZN(n6602) );
  INV_X1 U7520 ( .A(n6592), .ZN(n6598) );
  INV_X1 U7521 ( .A(n6593), .ZN(n6596) );
  OAI21_X1 U7522 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6594), 
        .ZN(n6595) );
  NAND4_X1 U7523 ( .A1(n6598), .A2(n6597), .A3(n6596), .A4(n6595), .ZN(n6601)
         );
  INV_X1 U7524 ( .A(n6599), .ZN(n6600) );
  AOI211_X1 U7525 ( .C1(n6603), .C2(n6602), .A(n6601), .B(n6600), .ZN(n6615)
         );
  INV_X1 U7526 ( .A(n6615), .ZN(n6605) );
  OAI22_X1 U7527 ( .A1(n6605), .A2(n6617), .B1(n6604), .B2(n6704), .ZN(n6606)
         );
  OAI21_X1 U7528 ( .B1(n6608), .B2(n6607), .A(n6606), .ZN(n6692) );
  OAI21_X1 U7529 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6704), .A(n6692), .ZN(
        n6616) );
  AOI221_X1 U7530 ( .B1(n6610), .B2(STATE2_REG_0__SCAN_IN), .C1(n6616), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6609), .ZN(n6614) );
  OAI211_X1 U7531 ( .C1(n6623), .C2(n6612), .A(n6611), .B(n6692), .ZN(n6613)
         );
  OAI211_X1 U7532 ( .C1(n6615), .C2(n6617), .A(n6614), .B(n6613), .ZN(U3148)
         );
  OAI211_X1 U7533 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6616), .ZN(n6622) );
  OAI21_X1 U7534 ( .B1(READY_N), .B2(n6618), .A(n6617), .ZN(n6620) );
  AOI21_X1 U7535 ( .B1(n6620), .B2(n6692), .A(n6619), .ZN(n6621) );
  NAND2_X1 U7536 ( .A1(n6622), .A2(n6621), .ZN(U3149) );
  INV_X1 U7537 ( .A(n6623), .ZN(n6707) );
  OAI221_X1 U7538 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n6704), .A(n6691), .ZN(n6625) );
  OAI21_X1 U7539 ( .B1(n6707), .B2(n6625), .A(n6624), .ZN(U3150) );
  AND2_X1 U7540 ( .A1(n6627), .A2(DATAWIDTH_REG_31__SCAN_IN), .ZN(U3151) );
  AND2_X1 U7541 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6627), .ZN(U3152) );
  AND2_X1 U7542 ( .A1(n6627), .A2(DATAWIDTH_REG_29__SCAN_IN), .ZN(U3153) );
  AND2_X1 U7543 ( .A1(n6627), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U7544 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6627), .ZN(U3155) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6627), .ZN(U3156) );
  AND2_X1 U7546 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6627), .ZN(U3157) );
  AND2_X1 U7547 ( .A1(n6627), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6627), .ZN(U3159) );
  AND2_X1 U7549 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6627), .ZN(U3160) );
  AND2_X1 U7550 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6627), .ZN(U3161) );
  AND2_X1 U7551 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6627), .ZN(U3162) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6627), .ZN(U3163) );
  AND2_X1 U7553 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6627), .ZN(U3164) );
  AND2_X1 U7554 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6627), .ZN(U3165) );
  AND2_X1 U7555 ( .A1(n6627), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U7556 ( .A1(n6627), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  NOR2_X1 U7557 ( .A1(n6690), .A2(n6896), .ZN(U3168) );
  AND2_X1 U7558 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6627), .ZN(U3169) );
  AND2_X1 U7559 ( .A1(n6627), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6627), .ZN(U3171) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6627), .ZN(U3172) );
  AND2_X1 U7562 ( .A1(n6627), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U7563 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6627), .ZN(U3174) );
  AND2_X1 U7564 ( .A1(n6627), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  AND2_X1 U7565 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6627), .ZN(U3176) );
  AND2_X1 U7566 ( .A1(n6627), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  NOR2_X1 U7567 ( .A1(n6690), .A2(n6626), .ZN(U3178) );
  AND2_X1 U7568 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6627), .ZN(U3179) );
  AND2_X1 U7569 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6627), .ZN(U3180) );
  NAND2_X1 U7570 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6630) );
  AND2_X1 U7571 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6634) );
  NAND2_X1 U7572 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6635) );
  INV_X1 U7573 ( .A(n6635), .ZN(n6639) );
  INV_X1 U7574 ( .A(NA_N), .ZN(n6628) );
  AOI221_X1 U7575 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6628), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6641) );
  AOI221_X1 U7576 ( .B1(n6634), .B2(n6636), .C1(n6639), .C2(n6636), .A(n6641), 
        .ZN(n6629) );
  OAI221_X1 U7577 ( .B1(n6712), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6712), 
        .C2(n6630), .A(n6629), .ZN(U3181) );
  INV_X1 U7578 ( .A(n6630), .ZN(n6631) );
  AOI21_X1 U7579 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_0__SCAN_IN), 
        .A(n6631), .ZN(n6633) );
  OAI211_X1 U7580 ( .C1(n6634), .C2(n6633), .A(n6632), .B(n6635), .ZN(U3182)
         );
  AOI221_X1 U7581 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6704), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6638) );
  OAI21_X1 U7582 ( .B1(n6636), .B2(n6635), .A(STATE_REG_0__SCAN_IN), .ZN(n6637) );
  AOI221_X1 U7583 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6638), .C2(HOLD), .A(n6637), .ZN(n6642) );
  NAND3_X1 U7584 ( .A1(STATE_REG_0__SCAN_IN), .A2(REQUESTPENDING_REG_SCAN_IN), 
        .A3(n6639), .ZN(n6640) );
  OAI22_X1 U7585 ( .A1(n6642), .A2(n6641), .B1(NA_N), .B2(n6640), .ZN(U3183)
         );
  NAND2_X1 U7586 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6712), .ZN(n6680) );
  NOR2_X2 U7587 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6685), .ZN(n6678) );
  AOI22_X1 U7588 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6685), .ZN(n6643) );
  OAI21_X1 U7589 ( .B1(n6815), .B2(n6680), .A(n6643), .ZN(U3184) );
  AOI22_X1 U7590 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6685), .ZN(n6644) );
  OAI21_X1 U7591 ( .B1(n5177), .B2(n6680), .A(n6644), .ZN(U3185) );
  AOI22_X1 U7592 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6685), .ZN(n6645) );
  OAI21_X1 U7593 ( .B1(n6928), .B2(n6680), .A(n6645), .ZN(U3186) );
  AOI22_X1 U7594 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6685), .ZN(n6646) );
  OAI21_X1 U7595 ( .B1(n6934), .B2(n6680), .A(n6646), .ZN(U3187) );
  AOI22_X1 U7596 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6685), .ZN(n6647) );
  OAI21_X1 U7597 ( .B1(n6648), .B2(n6680), .A(n6647), .ZN(U3188) );
  INV_X1 U7598 ( .A(n6680), .ZN(n6682) );
  AOI22_X1 U7599 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6685), .ZN(n6649) );
  OAI21_X1 U7600 ( .B1(n6651), .B2(n6684), .A(n6649), .ZN(U3189) );
  AOI22_X1 U7601 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6685), .ZN(n6650) );
  OAI21_X1 U7602 ( .B1(n6651), .B2(n6680), .A(n6650), .ZN(U3190) );
  INV_X1 U7603 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6652) );
  OAI222_X1 U7604 ( .A1(n6684), .A2(n5182), .B1(n6652), .B2(n6712), .C1(n5082), 
        .C2(n6680), .ZN(U3191) );
  AOI22_X1 U7605 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6685), .ZN(n6653) );
  OAI21_X1 U7606 ( .B1(n6730), .B2(n6684), .A(n6653), .ZN(U3192) );
  AOI22_X1 U7607 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6685), .ZN(n6654) );
  OAI21_X1 U7608 ( .B1(n6730), .B2(n6680), .A(n6654), .ZN(U3193) );
  AOI22_X1 U7609 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6685), .ZN(n6655) );
  OAI21_X1 U7610 ( .B1(n5293), .B2(n6680), .A(n6655), .ZN(U3194) );
  AOI22_X1 U7611 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6685), .ZN(n6656) );
  OAI21_X1 U7612 ( .B1(n6749), .B2(n6684), .A(n6656), .ZN(U3195) );
  AOI222_X1 U7613 ( .A1(n6682), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6685), .C1(REIP_REG_14__SCAN_IN), .C2(
        n6678), .ZN(n6657) );
  INV_X1 U7614 ( .A(n6657), .ZN(U3196) );
  AOI22_X1 U7615 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6685), .ZN(n6658) );
  OAI21_X1 U7616 ( .B1(n6659), .B2(n6684), .A(n6658), .ZN(U3197) );
  AOI22_X1 U7617 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6685), .ZN(n6660) );
  OAI21_X1 U7618 ( .B1(n5626), .B2(n6684), .A(n6660), .ZN(U3198) );
  AOI22_X1 U7619 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6685), .ZN(n6661) );
  OAI21_X1 U7620 ( .B1(n5626), .B2(n6680), .A(n6661), .ZN(U3199) );
  AOI22_X1 U7621 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6685), .ZN(n6662) );
  OAI21_X1 U7622 ( .B1(n6798), .B2(n6680), .A(n6662), .ZN(U3200) );
  AOI22_X1 U7623 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6685), .ZN(n6663) );
  OAI21_X1 U7624 ( .B1(n6664), .B2(n6680), .A(n6663), .ZN(U3201) );
  AOI22_X1 U7625 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6685), .ZN(n6665) );
  OAI21_X1 U7626 ( .B1(n6667), .B2(n6684), .A(n6665), .ZN(U3202) );
  AOI22_X1 U7627 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6685), .ZN(n6666) );
  OAI21_X1 U7628 ( .B1(n6667), .B2(n6680), .A(n6666), .ZN(U3203) );
  AOI22_X1 U7629 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6685), .ZN(n6668) );
  OAI21_X1 U7630 ( .B1(n6669), .B2(n6684), .A(n6668), .ZN(U3204) );
  INV_X1 U7631 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6762) );
  AOI22_X1 U7632 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6685), .ZN(n6670) );
  OAI21_X1 U7633 ( .B1(n6762), .B2(n6684), .A(n6670), .ZN(U3205) );
  AOI22_X1 U7634 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6685), .ZN(n6671) );
  OAI21_X1 U7635 ( .B1(n6762), .B2(n6680), .A(n6671), .ZN(U3206) );
  AOI22_X1 U7636 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6685), .ZN(n6672) );
  OAI21_X1 U7637 ( .B1(n5409), .B2(n6684), .A(n6672), .ZN(U3207) );
  INV_X1 U7638 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6673) );
  OAI222_X1 U7639 ( .A1(n6680), .A2(n5409), .B1(n6673), .B2(n6712), .C1(n5570), 
        .C2(n6684), .ZN(U3208) );
  AOI22_X1 U7640 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6685), .ZN(n6674) );
  OAI21_X1 U7641 ( .B1(n6676), .B2(n6684), .A(n6674), .ZN(U3209) );
  AOI22_X1 U7642 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6685), .ZN(n6675) );
  OAI21_X1 U7643 ( .B1(n6676), .B2(n6680), .A(n6675), .ZN(U3210) );
  AOI22_X1 U7644 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6685), .ZN(n6677) );
  OAI21_X1 U7645 ( .B1(n6681), .B2(n6684), .A(n6677), .ZN(U3211) );
  AOI22_X1 U7646 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6678), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6685), .ZN(n6679) );
  OAI21_X1 U7647 ( .B1(n6681), .B2(n6680), .A(n6679), .ZN(U3212) );
  AOI22_X1 U7648 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6682), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6685), .ZN(n6683) );
  OAI21_X1 U7649 ( .B1(n6917), .B2(n6684), .A(n6683), .ZN(U3213) );
  MUX2_X1 U7650 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6712), .Z(U3445) );
  MUX2_X1 U7651 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6712), .Z(U3446) );
  OAI22_X1 U7652 ( .A1(n6685), .A2(BYTEENABLE_REG_1__SCAN_IN), .B1(
        BE_N_REG_1__SCAN_IN), .B2(n6712), .ZN(n6686) );
  INV_X1 U7653 ( .A(n6686), .ZN(U3447) );
  MUX2_X1 U7654 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6712), .Z(U3448) );
  OAI21_X1 U7655 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6690), .A(n6688), .ZN(
        n6687) );
  INV_X1 U7656 ( .A(n6687), .ZN(U3451) );
  OAI21_X1 U7657 ( .B1(n6690), .B2(n6689), .A(n6688), .ZN(U3452) );
  OAI221_X1 U7658 ( .B1(n6693), .B2(STATE2_REG_0__SCAN_IN), .C1(n6693), .C2(
        n6692), .A(n6691), .ZN(U3453) );
  INV_X1 U7659 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6696) );
  AOI21_X1 U7660 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6694) );
  OAI221_X1 U7661 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6694), .C1(n6815), .C2(
        REIP_REG_0__SCAN_IN), .A(n6697), .ZN(n6695) );
  OAI21_X1 U7662 ( .B1(n6697), .B2(n6696), .A(n6695), .ZN(U3468) );
  INV_X1 U7663 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6897) );
  NOR2_X1 U7664 ( .A1(n6700), .A2(REIP_REG_1__SCAN_IN), .ZN(n6698) );
  AOI22_X1 U7665 ( .A1(n6897), .A2(n6700), .B1(n6699), .B2(n6698), .ZN(U3469)
         );
  NAND2_X1 U7666 ( .A1(n6685), .A2(W_R_N_REG_SCAN_IN), .ZN(n6701) );
  OAI21_X1 U7667 ( .B1(n6685), .B2(READREQUEST_REG_SCAN_IN), .A(n6701), .ZN(
        U3470) );
  AOI211_X1 U7668 ( .C1(n6195), .C2(n6704), .A(n6703), .B(n6702), .ZN(n6711)
         );
  OAI211_X1 U7669 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6706), .A(n6705), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6708) );
  AOI21_X1 U7670 ( .B1(n6708), .B2(STATE2_REG_0__SCAN_IN), .A(n6707), .ZN(
        n6710) );
  NAND2_X1 U7671 ( .A1(n6711), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6709) );
  OAI21_X1 U7672 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(U3472) );
  MUX2_X1 U7673 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6712), .Z(U3473) );
  INV_X1 U7674 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6714) );
  AOI22_X1 U7675 ( .A1(n4766), .A2(keyinput74), .B1(n6714), .B2(keyinput41), 
        .ZN(n6713) );
  OAI221_X1 U7676 ( .B1(n4766), .B2(keyinput74), .C1(n6714), .C2(keyinput41), 
        .A(n6713), .ZN(n6727) );
  AOI22_X1 U7677 ( .A1(n6717), .A2(keyinput117), .B1(keyinput79), .B2(n6716), 
        .ZN(n6715) );
  OAI221_X1 U7678 ( .B1(n6717), .B2(keyinput117), .C1(n6716), .C2(keyinput79), 
        .A(n6715), .ZN(n6726) );
  INV_X1 U7679 ( .A(keyinput45), .ZN(n6720) );
  INV_X1 U7680 ( .A(keyinput81), .ZN(n6719) );
  AOI22_X1 U7681 ( .A1(n6720), .A2(DATAO_REG_15__SCAN_IN), .B1(
        DATAWIDTH_REG_31__SCAN_IN), .B2(n6719), .ZN(n6718) );
  OAI221_X1 U7682 ( .B1(n6720), .B2(DATAO_REG_15__SCAN_IN), .C1(n6719), .C2(
        DATAWIDTH_REG_31__SCAN_IN), .A(n6718), .ZN(n6725) );
  INV_X1 U7683 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6723) );
  INV_X1 U7684 ( .A(keyinput23), .ZN(n6722) );
  AOI22_X1 U7685 ( .A1(n6723), .A2(keyinput107), .B1(ADDRESS_REG_1__SCAN_IN), 
        .B2(n6722), .ZN(n6721) );
  OAI221_X1 U7686 ( .B1(n6723), .B2(keyinput107), .C1(n6722), .C2(
        ADDRESS_REG_1__SCAN_IN), .A(n6721), .ZN(n6724) );
  NOR4_X1 U7687 ( .A1(n6727), .A2(n6726), .A3(n6725), .A4(n6724), .ZN(n7033)
         );
  AOI22_X1 U7688 ( .A1(n6730), .A2(keyinput33), .B1(n6729), .B2(keyinput89), 
        .ZN(n6728) );
  OAI221_X1 U7689 ( .B1(n6730), .B2(keyinput33), .C1(n6729), .C2(keyinput89), 
        .A(n6728), .ZN(n6744) );
  INV_X1 U7690 ( .A(keyinput104), .ZN(n6733) );
  INV_X1 U7691 ( .A(keyinput1), .ZN(n6732) );
  AOI22_X1 U7692 ( .A1(n6733), .A2(DATAO_REG_31__SCAN_IN), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6732), .ZN(n6731) );
  OAI221_X1 U7693 ( .B1(n6733), .B2(DATAO_REG_31__SCAN_IN), .C1(n6732), .C2(
        ADDRESS_REG_29__SCAN_IN), .A(n6731), .ZN(n6743) );
  INV_X1 U7694 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6736) );
  INV_X1 U7695 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7696 ( .A1(n6736), .A2(keyinput32), .B1(n6735), .B2(keyinput108), 
        .ZN(n6734) );
  OAI221_X1 U7697 ( .B1(n6736), .B2(keyinput32), .C1(n6735), .C2(keyinput108), 
        .A(n6734), .ZN(n6742) );
  INV_X1 U7698 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6737) );
  XOR2_X1 U7699 ( .A(n6737), .B(keyinput5), .Z(n6740) );
  XNOR2_X1 U7700 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput2), .ZN(
        n6739) );
  NAND2_X1 U7701 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  NOR4_X1 U7702 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n7032)
         );
  OAI22_X1 U7703 ( .A1(n6750), .A2(keyinput69), .B1(n6749), .B2(keyinput7), 
        .ZN(n6748) );
  AOI221_X1 U7704 ( .B1(n6750), .B2(keyinput69), .C1(keyinput7), .C2(n6749), 
        .A(n6748), .ZN(n6759) );
  INV_X1 U7705 ( .A(keyinput34), .ZN(n6752) );
  OAI22_X1 U7706 ( .A1(keyinput63), .A2(n6753), .B1(n6752), .B2(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6751) );
  AOI221_X1 U7707 ( .B1(n6753), .B2(keyinput63), .C1(n6752), .C2(
        DATAWIDTH_REG_16__SCAN_IN), .A(n6751), .ZN(n6758) );
  INV_X1 U7708 ( .A(keyinput44), .ZN(n6755) );
  OAI22_X1 U7709 ( .A1(n6756), .A2(keyinput19), .B1(n6755), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6754) );
  AOI221_X1 U7710 ( .B1(n6756), .B2(keyinput19), .C1(DATAO_REG_3__SCAN_IN), 
        .C2(n6755), .A(n6754), .ZN(n6757) );
  NAND4_X1 U7711 ( .A1(n6760), .A2(n6759), .A3(n6758), .A4(n6757), .ZN(n6842)
         );
  INV_X1 U7712 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n6763) );
  OAI22_X1 U7713 ( .A1(n6763), .A2(keyinput65), .B1(n6762), .B2(keyinput72), 
        .ZN(n6761) );
  AOI221_X1 U7714 ( .B1(n6763), .B2(keyinput65), .C1(keyinput72), .C2(n6762), 
        .A(n6761), .ZN(n6776) );
  INV_X1 U7715 ( .A(keyinput85), .ZN(n6765) );
  OAI22_X1 U7716 ( .A1(n6766), .A2(keyinput58), .B1(n6765), .B2(
        M_IO_N_REG_SCAN_IN), .ZN(n6764) );
  AOI221_X1 U7717 ( .B1(n6766), .B2(keyinput58), .C1(M_IO_N_REG_SCAN_IN), .C2(
        n6765), .A(n6764), .ZN(n6775) );
  INV_X1 U7718 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6769) );
  INV_X1 U7719 ( .A(keyinput84), .ZN(n6768) );
  OAI22_X1 U7720 ( .A1(n6769), .A2(keyinput115), .B1(n6768), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6767) );
  AOI221_X1 U7721 ( .B1(n6769), .B2(keyinput115), .C1(DATAO_REG_13__SCAN_IN), 
        .C2(n6768), .A(n6767), .ZN(n6774) );
  INV_X1 U7722 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6771) );
  OAI22_X1 U7723 ( .A1(n6772), .A2(keyinput98), .B1(n6771), .B2(keyinput80), 
        .ZN(n6770) );
  AOI221_X1 U7724 ( .B1(n6772), .B2(keyinput98), .C1(keyinput80), .C2(n6771), 
        .A(n6770), .ZN(n6773) );
  NAND4_X1 U7725 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6841)
         );
  INV_X1 U7726 ( .A(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n6779) );
  AOI22_X1 U7727 ( .A1(n6779), .A2(keyinput92), .B1(keyinput121), .B2(n6778), 
        .ZN(n6777) );
  OAI221_X1 U7728 ( .B1(n6779), .B2(keyinput92), .C1(n6778), .C2(keyinput121), 
        .A(n6777), .ZN(n6791) );
  INV_X1 U7729 ( .A(keyinput77), .ZN(n6781) );
  AOI22_X1 U7730 ( .A1(n5385), .A2(keyinput25), .B1(ADDRESS_REG_24__SCAN_IN), 
        .B2(n6781), .ZN(n6780) );
  OAI221_X1 U7731 ( .B1(n5385), .B2(keyinput25), .C1(n6781), .C2(
        ADDRESS_REG_24__SCAN_IN), .A(n6780), .ZN(n6790) );
  INV_X1 U7732 ( .A(keyinput68), .ZN(n6784) );
  INV_X1 U7733 ( .A(keyinput30), .ZN(n6783) );
  AOI22_X1 U7734 ( .A1(n6784), .A2(ADDRESS_REG_3__SCAN_IN), .B1(
        DATAWIDTH_REG_24__SCAN_IN), .B2(n6783), .ZN(n6782) );
  OAI221_X1 U7735 ( .B1(n6784), .B2(ADDRESS_REG_3__SCAN_IN), .C1(n6783), .C2(
        DATAWIDTH_REG_24__SCAN_IN), .A(n6782), .ZN(n6789) );
  INV_X1 U7736 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6786) );
  AOI22_X1 U7737 ( .A1(n6787), .A2(keyinput4), .B1(n6786), .B2(keyinput20), 
        .ZN(n6785) );
  OAI221_X1 U7738 ( .B1(n6787), .B2(keyinput4), .C1(n6786), .C2(keyinput20), 
        .A(n6785), .ZN(n6788) );
  NOR4_X1 U7739 ( .A1(n6791), .A2(n6790), .A3(n6789), .A4(n6788), .ZN(n6839)
         );
  INV_X1 U7740 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6793) );
  INV_X1 U7741 ( .A(keyinput122), .ZN(n6867) );
  AOI22_X1 U7742 ( .A1(n6793), .A2(keyinput37), .B1(REQUESTPENDING_REG_SCAN_IN), .B2(n6867), .ZN(n6792) );
  OAI221_X1 U7743 ( .B1(n6793), .B2(keyinput37), .C1(n6867), .C2(
        REQUESTPENDING_REG_SCAN_IN), .A(n6792), .ZN(n6805) );
  AOI22_X1 U7744 ( .A1(n5182), .A2(keyinput27), .B1(n6795), .B2(keyinput31), 
        .ZN(n6794) );
  OAI221_X1 U7745 ( .B1(n5182), .B2(keyinput27), .C1(n6795), .C2(keyinput31), 
        .A(n6794), .ZN(n6804) );
  INV_X1 U7746 ( .A(keyinput75), .ZN(n6797) );
  AOI22_X1 U7747 ( .A1(n6798), .A2(keyinput18), .B1(DATAO_REG_1__SCAN_IN), 
        .B2(n6797), .ZN(n6796) );
  OAI221_X1 U7748 ( .B1(n6798), .B2(keyinput18), .C1(n6797), .C2(
        DATAO_REG_1__SCAN_IN), .A(n6796), .ZN(n6803) );
  INV_X1 U7749 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6801) );
  INV_X1 U7750 ( .A(keyinput125), .ZN(n6800) );
  AOI22_X1 U7751 ( .A1(n6801), .A2(keyinput55), .B1(DATAWIDTH_REG_12__SCAN_IN), 
        .B2(n6800), .ZN(n6799) );
  OAI221_X1 U7752 ( .B1(n6801), .B2(keyinput55), .C1(n6800), .C2(
        DATAWIDTH_REG_12__SCAN_IN), .A(n6799), .ZN(n6802) );
  NOR4_X1 U7753 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n6838)
         );
  INV_X1 U7754 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6807) );
  AOI22_X1 U7755 ( .A1(n6808), .A2(keyinput101), .B1(n6807), .B2(keyinput38), 
        .ZN(n6806) );
  OAI221_X1 U7756 ( .B1(n6808), .B2(keyinput101), .C1(n6807), .C2(keyinput38), 
        .A(n6806), .ZN(n6820) );
  INV_X1 U7757 ( .A(keyinput99), .ZN(n6810) );
  AOI22_X1 U7758 ( .A1(n4829), .A2(keyinput124), .B1(DATAWIDTH_REG_4__SCAN_IN), 
        .B2(n6810), .ZN(n6809) );
  OAI221_X1 U7759 ( .B1(n4829), .B2(keyinput124), .C1(n6810), .C2(
        DATAWIDTH_REG_4__SCAN_IN), .A(n6809), .ZN(n6819) );
  INV_X1 U7760 ( .A(keyinput96), .ZN(n6812) );
  AOI22_X1 U7761 ( .A1(n6813), .A2(keyinput76), .B1(DATAO_REG_4__SCAN_IN), 
        .B2(n6812), .ZN(n6811) );
  OAI221_X1 U7762 ( .B1(n6813), .B2(keyinput76), .C1(n6812), .C2(
        DATAO_REG_4__SCAN_IN), .A(n6811), .ZN(n6818) );
  AOI22_X1 U7763 ( .A1(n6816), .A2(keyinput105), .B1(n6815), .B2(keyinput100), 
        .ZN(n6814) );
  OAI221_X1 U7764 ( .B1(n6816), .B2(keyinput105), .C1(n6815), .C2(keyinput100), 
        .A(n6814), .ZN(n6817) );
  NOR4_X1 U7765 ( .A1(n6820), .A2(n6819), .A3(n6818), .A4(n6817), .ZN(n6837)
         );
  INV_X1 U7766 ( .A(keyinput102), .ZN(n6823) );
  INV_X1 U7767 ( .A(keyinput15), .ZN(n6822) );
  AOI22_X1 U7768 ( .A1(n6823), .A2(DATAO_REG_27__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6822), .ZN(n6821) );
  OAI221_X1 U7769 ( .B1(n6823), .B2(DATAO_REG_27__SCAN_IN), .C1(n6822), .C2(
        ADDRESS_REG_5__SCAN_IN), .A(n6821), .ZN(n6835) );
  INV_X1 U7770 ( .A(DATAI_23_), .ZN(n6825) );
  AOI22_X1 U7771 ( .A1(n6825), .A2(keyinput97), .B1(n5126), .B2(keyinput49), 
        .ZN(n6824) );
  OAI221_X1 U7772 ( .B1(n6825), .B2(keyinput97), .C1(n5126), .C2(keyinput49), 
        .A(n6824), .ZN(n6834) );
  AOI22_X1 U7773 ( .A1(n6828), .A2(keyinput82), .B1(n6827), .B2(keyinput9), 
        .ZN(n6826) );
  OAI221_X1 U7774 ( .B1(n6828), .B2(keyinput82), .C1(n6827), .C2(keyinput9), 
        .A(n6826), .ZN(n6833) );
  AOI22_X1 U7775 ( .A1(n6831), .A2(keyinput91), .B1(keyinput39), .B2(n6830), 
        .ZN(n6829) );
  OAI221_X1 U7776 ( .B1(n6831), .B2(keyinput91), .C1(n6830), .C2(keyinput39), 
        .A(n6829), .ZN(n6832) );
  NOR4_X1 U7777 ( .A1(n6835), .A2(n6834), .A3(n6833), .A4(n6832), .ZN(n6836)
         );
  NAND4_X1 U7778 ( .A1(n6839), .A2(n6838), .A3(n6837), .A4(n6836), .ZN(n6840)
         );
  NOR3_X1 U7779 ( .A1(n6842), .A2(n6841), .A3(n6840), .ZN(n7031) );
  INV_X1 U7780 ( .A(keyinput105), .ZN(n6843) );
  NAND4_X1 U7781 ( .A1(keyinput100), .A2(keyinput96), .A3(keyinput76), .A4(
        n6843), .ZN(n6844) );
  NOR3_X1 U7782 ( .A1(keyinput101), .A2(keyinput38), .A3(n6844), .ZN(n6858) );
  NAND2_X1 U7783 ( .A1(keyinput19), .A2(keyinput120), .ZN(n6845) );
  NOR3_X1 U7784 ( .A1(keyinput7), .A2(keyinput34), .A3(n6845), .ZN(n6846) );
  NAND3_X1 U7785 ( .A1(keyinput44), .A2(keyinput63), .A3(n6846), .ZN(n6856) );
  NAND2_X1 U7786 ( .A1(keyinput115), .A2(keyinput98), .ZN(n6847) );
  NOR3_X1 U7787 ( .A1(keyinput84), .A2(keyinput80), .A3(n6847), .ZN(n6854) );
  INV_X1 U7788 ( .A(keyinput58), .ZN(n6848) );
  NOR4_X1 U7789 ( .A1(keyinput65), .A2(keyinput85), .A3(keyinput72), .A4(n6848), .ZN(n6853) );
  NAND2_X1 U7790 ( .A1(keyinput9), .A2(keyinput91), .ZN(n6849) );
  NOR3_X1 U7791 ( .A1(keyinput82), .A2(keyinput39), .A3(n6849), .ZN(n6852) );
  NAND2_X1 U7792 ( .A1(keyinput102), .A2(keyinput49), .ZN(n6850) );
  NOR3_X1 U7793 ( .A1(keyinput97), .A2(keyinput15), .A3(n6850), .ZN(n6851) );
  NAND4_X1 U7794 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6855)
         );
  NOR4_X1 U7795 ( .A1(keyinput69), .A2(keyinput51), .A3(n6856), .A4(n6855), 
        .ZN(n6857) );
  NAND4_X1 U7796 ( .A1(keyinput99), .A2(keyinput124), .A3(n6858), .A4(n6857), 
        .ZN(n6894) );
  NOR4_X1 U7797 ( .A1(keyinput28), .A2(keyinput29), .A3(keyinput36), .A4(
        keyinput56), .ZN(n6862) );
  NOR4_X1 U7798 ( .A1(keyinput14), .A2(keyinput35), .A3(keyinput22), .A4(
        keyinput26), .ZN(n6861) );
  NOR4_X1 U7799 ( .A1(keyinput24), .A2(keyinput93), .A3(keyinput109), .A4(
        keyinput113), .ZN(n6860) );
  NOR4_X1 U7800 ( .A1(keyinput0), .A2(keyinput8), .A3(keyinput13), .A4(
        keyinput21), .ZN(n6859) );
  NAND4_X1 U7801 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6893)
         );
  NOR4_X1 U7802 ( .A1(keyinput71), .A2(keyinput70), .A3(keyinput119), .A4(
        keyinput118), .ZN(n6866) );
  NOR4_X1 U7803 ( .A1(keyinput10), .A2(keyinput103), .A3(keyinput106), .A4(
        keyinput66), .ZN(n6865) );
  NOR4_X1 U7804 ( .A1(keyinput110), .A2(keyinput54), .A3(keyinput62), .A4(
        keyinput50), .ZN(n6864) );
  NOR4_X1 U7805 ( .A1(keyinput123), .A2(keyinput86), .A3(keyinput78), .A4(
        keyinput111), .ZN(n6863) );
  NAND4_X1 U7806 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6892)
         );
  NAND4_X1 U7807 ( .A1(keyinput55), .A2(keyinput125), .A3(keyinput75), .A4(
        keyinput18), .ZN(n6871) );
  NAND4_X1 U7808 ( .A1(keyinput31), .A2(keyinput27), .A3(keyinput37), .A4(
        n6867), .ZN(n6870) );
  NAND4_X1 U7809 ( .A1(keyinput92), .A2(keyinput121), .A3(keyinput68), .A4(
        keyinput30), .ZN(n6869) );
  OR4_X1 U7810 ( .A1(keyinput77), .A2(keyinput25), .A3(keyinput4), .A4(
        keyinput20), .ZN(n6868) );
  NOR4_X1 U7811 ( .A1(n6871), .A2(n6870), .A3(n6869), .A4(n6868), .ZN(n6890)
         );
  NOR3_X1 U7812 ( .A1(keyinput5), .A2(keyinput108), .A3(keyinput32), .ZN(n6872) );
  NAND2_X1 U7813 ( .A1(keyinput2), .A2(n6872), .ZN(n6877) );
  NAND4_X1 U7814 ( .A1(keyinput104), .A2(keyinput1), .A3(keyinput33), .A4(
        keyinput89), .ZN(n6876) );
  NOR3_X1 U7815 ( .A1(keyinput45), .A2(keyinput81), .A3(keyinput41), .ZN(n6873) );
  NAND2_X1 U7816 ( .A1(keyinput74), .A2(n6873), .ZN(n6875) );
  NAND4_X1 U7817 ( .A1(keyinput117), .A2(keyinput79), .A3(keyinput107), .A4(
        keyinput23), .ZN(n6874) );
  NOR4_X1 U7818 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6889)
         );
  NAND4_X1 U7819 ( .A1(keyinput60), .A2(keyinput52), .A3(keyinput40), .A4(
        keyinput53), .ZN(n6881) );
  NAND4_X1 U7820 ( .A1(keyinput17), .A2(keyinput12), .A3(keyinput57), .A4(
        keyinput48), .ZN(n6880) );
  NAND4_X1 U7821 ( .A1(keyinput47), .A2(keyinput42), .A3(keyinput46), .A4(
        keyinput11), .ZN(n6879) );
  NAND4_X1 U7822 ( .A1(keyinput59), .A2(keyinput3), .A3(keyinput43), .A4(
        keyinput6), .ZN(n6878) );
  NOR4_X1 U7823 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6888)
         );
  NAND4_X1 U7824 ( .A1(keyinput114), .A2(keyinput83), .A3(keyinput126), .A4(
        keyinput95), .ZN(n6886) );
  INV_X1 U7825 ( .A(keyinput61), .ZN(n6882) );
  NAND4_X1 U7826 ( .A1(keyinput87), .A2(keyinput67), .A3(keyinput127), .A4(
        n6882), .ZN(n6885) );
  NAND4_X1 U7827 ( .A1(keyinput64), .A2(keyinput112), .A3(keyinput116), .A4(
        keyinput16), .ZN(n6884) );
  NAND4_X1 U7828 ( .A1(keyinput90), .A2(keyinput94), .A3(keyinput88), .A4(
        keyinput73), .ZN(n6883) );
  NOR4_X1 U7829 ( .A1(n6886), .A2(n6885), .A3(n6884), .A4(n6883), .ZN(n6887)
         );
  NAND4_X1 U7830 ( .A1(n6890), .A2(n6889), .A3(n6888), .A4(n6887), .ZN(n6891)
         );
  NOR4_X1 U7831 ( .A1(n6894), .A2(n6893), .A3(n6892), .A4(n6891), .ZN(n7029)
         );
  OAI22_X1 U7832 ( .A1(keyinput54), .A2(n6897), .B1(n6896), .B2(keyinput61), 
        .ZN(n6895) );
  AOI221_X1 U7833 ( .B1(n6897), .B2(keyinput54), .C1(n6896), .C2(keyinput61), 
        .A(n6895), .ZN(n6909) );
  OAI22_X1 U7834 ( .A1(n6900), .A2(keyinput29), .B1(n6899), .B2(keyinput88), 
        .ZN(n6898) );
  AOI221_X1 U7835 ( .B1(n6900), .B2(keyinput29), .C1(keyinput88), .C2(n6899), 
        .A(n6898), .ZN(n6908) );
  INV_X1 U7836 ( .A(keyinput13), .ZN(n6902) );
  OAI22_X1 U7837 ( .A1(n5082), .A2(keyinput119), .B1(n6902), .B2(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6901) );
  AOI221_X1 U7838 ( .B1(n5082), .B2(keyinput119), .C1(DATAWIDTH_REG_5__SCAN_IN), .C2(n6902), .A(n6901), .ZN(n6907) );
  INV_X1 U7839 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n6905) );
  INV_X1 U7840 ( .A(keyinput111), .ZN(n6904) );
  OAI22_X1 U7841 ( .A1(n6905), .A2(keyinput70), .B1(n6904), .B2(
        DATAWIDTH_REG_9__SCAN_IN), .ZN(n6903) );
  AOI221_X1 U7842 ( .B1(n6905), .B2(keyinput70), .C1(DATAWIDTH_REG_9__SCAN_IN), 
        .C2(n6904), .A(n6903), .ZN(n6906) );
  NAND4_X1 U7843 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n7028)
         );
  INV_X1 U7844 ( .A(keyinput95), .ZN(n6911) );
  AOI22_X1 U7845 ( .A1(n6912), .A2(keyinput112), .B1(UWORD_REG_12__SCAN_IN), 
        .B2(n6911), .ZN(n6910) );
  OAI221_X1 U7846 ( .B1(n6912), .B2(keyinput112), .C1(n6911), .C2(
        UWORD_REG_12__SCAN_IN), .A(n6910), .ZN(n6925) );
  INV_X1 U7847 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6915) );
  INV_X1 U7848 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U7849 ( .A1(n6915), .A2(keyinput87), .B1(n6914), .B2(keyinput127), 
        .ZN(n6913) );
  OAI221_X1 U7850 ( .B1(n6915), .B2(keyinput87), .C1(n6914), .C2(keyinput127), 
        .A(n6913), .ZN(n6924) );
  INV_X1 U7851 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n6918) );
  AOI22_X1 U7852 ( .A1(n6918), .A2(keyinput67), .B1(keyinput48), .B2(n6917), 
        .ZN(n6916) );
  OAI221_X1 U7853 ( .B1(n6918), .B2(keyinput67), .C1(n6917), .C2(keyinput48), 
        .A(n6916), .ZN(n6923) );
  INV_X1 U7854 ( .A(keyinput62), .ZN(n6920) );
  AOI22_X1 U7855 ( .A1(n6921), .A2(keyinput26), .B1(UWORD_REG_1__SCAN_IN), 
        .B2(n6920), .ZN(n6919) );
  OAI221_X1 U7856 ( .B1(n6921), .B2(keyinput26), .C1(n6920), .C2(
        UWORD_REG_1__SCAN_IN), .A(n6919), .ZN(n6922) );
  NOR4_X1 U7857 ( .A1(n6925), .A2(n6924), .A3(n6923), .A4(n6922), .ZN(n6959)
         );
  INV_X1 U7858 ( .A(keyinput60), .ZN(n6927) );
  AOI22_X1 U7859 ( .A1(n6928), .A2(keyinput71), .B1(UWORD_REG_2__SCAN_IN), 
        .B2(n6927), .ZN(n6926) );
  OAI221_X1 U7860 ( .B1(n6928), .B2(keyinput71), .C1(n6927), .C2(
        UWORD_REG_2__SCAN_IN), .A(n6926), .ZN(n6941) );
  INV_X1 U7861 ( .A(keyinput114), .ZN(n6931) );
  INV_X1 U7862 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7863 ( .A1(n6931), .A2(DATAO_REG_0__SCAN_IN), .B1(keyinput57), 
        .B2(n6930), .ZN(n6929) );
  OAI221_X1 U7864 ( .B1(n6931), .B2(DATAO_REG_0__SCAN_IN), .C1(n6930), .C2(
        keyinput57), .A(n6929), .ZN(n6940) );
  INV_X1 U7865 ( .A(keyinput10), .ZN(n6933) );
  AOI22_X1 U7866 ( .A1(n6934), .A2(keyinput0), .B1(BE_N_REG_1__SCAN_IN), .B2(
        n6933), .ZN(n6932) );
  OAI221_X1 U7867 ( .B1(n6934), .B2(keyinput0), .C1(n6933), .C2(
        BE_N_REG_1__SCAN_IN), .A(n6932), .ZN(n6939) );
  INV_X1 U7868 ( .A(DATAI_18_), .ZN(n6937) );
  INV_X1 U7869 ( .A(keyinput64), .ZN(n6936) );
  AOI22_X1 U7870 ( .A1(n6937), .A2(keyinput118), .B1(ADDRESS_REG_12__SCAN_IN), 
        .B2(n6936), .ZN(n6935) );
  OAI221_X1 U7871 ( .B1(n6937), .B2(keyinput118), .C1(n6936), .C2(
        ADDRESS_REG_12__SCAN_IN), .A(n6935), .ZN(n6938) );
  NOR4_X1 U7872 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n6958)
         );
  INV_X1 U7873 ( .A(LWORD_REG_12__SCAN_IN), .ZN(n6944) );
  INV_X1 U7874 ( .A(keyinput109), .ZN(n6943) );
  OAI22_X1 U7875 ( .A1(keyinput35), .A2(n6944), .B1(n6943), .B2(
        DATAWIDTH_REG_7__SCAN_IN), .ZN(n6942) );
  AOI221_X1 U7876 ( .B1(n6944), .B2(keyinput35), .C1(n6943), .C2(
        DATAWIDTH_REG_7__SCAN_IN), .A(n6942), .ZN(n6957) );
  INV_X1 U7877 ( .A(keyinput73), .ZN(n6946) );
  AOI22_X1 U7878 ( .A1(n6947), .A2(keyinput53), .B1(ADDRESS_REG_7__SCAN_IN), 
        .B2(n6946), .ZN(n6945) );
  OAI221_X1 U7879 ( .B1(n6947), .B2(keyinput53), .C1(n6946), .C2(
        ADDRESS_REG_7__SCAN_IN), .A(n6945), .ZN(n6955) );
  AOI22_X1 U7880 ( .A1(n6950), .A2(keyinput123), .B1(n6949), .B2(keyinput11), 
        .ZN(n6948) );
  OAI221_X1 U7881 ( .B1(n6950), .B2(keyinput123), .C1(n6949), .C2(keyinput11), 
        .A(n6948), .ZN(n6954) );
  AOI22_X1 U7882 ( .A1(n6952), .A2(keyinput78), .B1(keyinput110), .B2(n5570), 
        .ZN(n6951) );
  OAI221_X1 U7883 ( .B1(n6952), .B2(keyinput78), .C1(n5570), .C2(keyinput110), 
        .A(n6951), .ZN(n6953) );
  NOR3_X1 U7884 ( .A1(n6955), .A2(n6954), .A3(n6953), .ZN(n6956) );
  NAND4_X1 U7885 ( .A1(n6959), .A2(n6958), .A3(n6957), .A4(n6956), .ZN(n7027)
         );
  INV_X1 U7886 ( .A(keyinput86), .ZN(n6961) );
  AOI22_X1 U7887 ( .A1(n6962), .A2(keyinput103), .B1(DATAWIDTH_REG_15__SCAN_IN), .B2(n6961), .ZN(n6960) );
  OAI221_X1 U7888 ( .B1(n6962), .B2(keyinput103), .C1(n6961), .C2(
        DATAWIDTH_REG_15__SCAN_IN), .A(n6960), .ZN(n6975) );
  INV_X1 U7889 ( .A(keyinput16), .ZN(n6965) );
  INV_X1 U7890 ( .A(keyinput42), .ZN(n6964) );
  AOI22_X1 U7891 ( .A1(n6965), .A2(DATAO_REG_14__SCAN_IN), .B1(
        BYTEENABLE_REG_1__SCAN_IN), .B2(n6964), .ZN(n6963) );
  OAI221_X1 U7892 ( .B1(n6965), .B2(DATAO_REG_14__SCAN_IN), .C1(n6964), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6963), .ZN(n6974) );
  INV_X1 U7893 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7894 ( .A1(n6968), .A2(keyinput83), .B1(keyinput59), .B2(n6967), 
        .ZN(n6966) );
  OAI221_X1 U7895 ( .B1(n6968), .B2(keyinput83), .C1(n6967), .C2(keyinput59), 
        .A(n6966), .ZN(n6973) );
  AOI22_X1 U7896 ( .A1(n6971), .A2(keyinput113), .B1(n6970), .B2(keyinput90), 
        .ZN(n6969) );
  OAI221_X1 U7897 ( .B1(n6971), .B2(keyinput113), .C1(n6970), .C2(keyinput90), 
        .A(n6969), .ZN(n6972) );
  NOR4_X1 U7898 ( .A1(n6975), .A2(n6974), .A3(n6973), .A4(n6972), .ZN(n7025)
         );
  AOI22_X1 U7899 ( .A1(n6978), .A2(keyinput21), .B1(keyinput24), .B2(n6977), 
        .ZN(n6976) );
  OAI221_X1 U7900 ( .B1(n6978), .B2(keyinput21), .C1(n6977), .C2(keyinput24), 
        .A(n6976), .ZN(n6991) );
  INV_X1 U7901 ( .A(DATAI_29_), .ZN(n6981) );
  INV_X1 U7902 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7903 ( .A1(n6981), .A2(keyinput12), .B1(n6980), .B2(keyinput40), 
        .ZN(n6979) );
  OAI221_X1 U7904 ( .B1(n6981), .B2(keyinput12), .C1(n6980), .C2(keyinput40), 
        .A(n6979), .ZN(n6990) );
  INV_X1 U7905 ( .A(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n6984) );
  INV_X1 U7906 ( .A(keyinput47), .ZN(n6983) );
  AOI22_X1 U7907 ( .A1(n6984), .A2(keyinput3), .B1(DATAWIDTH_REG_28__SCAN_IN), 
        .B2(n6983), .ZN(n6982) );
  OAI221_X1 U7908 ( .B1(n6984), .B2(keyinput3), .C1(n6983), .C2(
        DATAWIDTH_REG_28__SCAN_IN), .A(n6982), .ZN(n6989) );
  INV_X1 U7909 ( .A(keyinput93), .ZN(n6986) );
  AOI22_X1 U7910 ( .A1(n6987), .A2(keyinput36), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n6986), .ZN(n6985) );
  OAI221_X1 U7911 ( .B1(n6987), .B2(keyinput36), .C1(n6986), .C2(
        DATAO_REG_9__SCAN_IN), .A(n6985), .ZN(n6988) );
  NOR4_X1 U7912 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n7024)
         );
  INV_X1 U7913 ( .A(keyinput28), .ZN(n6993) );
  AOI22_X1 U7914 ( .A1(n6994), .A2(keyinput43), .B1(DATAWIDTH_REG_29__SCAN_IN), 
        .B2(n6993), .ZN(n6992) );
  OAI221_X1 U7915 ( .B1(n6994), .B2(keyinput43), .C1(n6993), .C2(
        DATAWIDTH_REG_29__SCAN_IN), .A(n6992), .ZN(n7007) );
  INV_X1 U7916 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U7917 ( .A1(n6997), .A2(keyinput50), .B1(keyinput94), .B2(n6996), 
        .ZN(n6995) );
  OAI221_X1 U7918 ( .B1(n6997), .B2(keyinput50), .C1(n6996), .C2(keyinput94), 
        .A(n6995), .ZN(n7006) );
  INV_X1 U7919 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6999) );
  AOI22_X1 U7920 ( .A1(n7000), .A2(keyinput56), .B1(keyinput46), .B2(n6999), 
        .ZN(n6998) );
  OAI221_X1 U7921 ( .B1(n7000), .B2(keyinput56), .C1(n6999), .C2(keyinput46), 
        .A(n6998), .ZN(n7005) );
  AOI22_X1 U7922 ( .A1(n7003), .A2(keyinput22), .B1(n7002), .B2(keyinput116), 
        .ZN(n7001) );
  OAI221_X1 U7923 ( .B1(n7003), .B2(keyinput22), .C1(n7002), .C2(keyinput116), 
        .A(n7001), .ZN(n7004) );
  NOR4_X1 U7924 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n7023)
         );
  INV_X1 U7925 ( .A(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n7010) );
  INV_X1 U7926 ( .A(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n7009) );
  AOI22_X1 U7927 ( .A1(n7010), .A2(keyinput14), .B1(keyinput17), .B2(n7009), 
        .ZN(n7008) );
  OAI221_X1 U7928 ( .B1(n7010), .B2(keyinput14), .C1(n7009), .C2(keyinput17), 
        .A(n7008), .ZN(n7021) );
  INV_X1 U7929 ( .A(keyinput52), .ZN(n7012) );
  AOI22_X1 U7930 ( .A1(n4508), .A2(keyinput126), .B1(DATAO_REG_5__SCAN_IN), 
        .B2(n7012), .ZN(n7011) );
  OAI221_X1 U7931 ( .B1(n4508), .B2(keyinput126), .C1(n7012), .C2(
        DATAO_REG_5__SCAN_IN), .A(n7011), .ZN(n7020) );
  AOI22_X1 U7932 ( .A1(n7014), .A2(keyinput66), .B1(n4114), .B2(keyinput6), 
        .ZN(n7013) );
  OAI221_X1 U7933 ( .B1(n7014), .B2(keyinput66), .C1(n4114), .C2(keyinput6), 
        .A(n7013), .ZN(n7019) );
  INV_X1 U7934 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n7016) );
  AOI22_X1 U7935 ( .A1(n7017), .A2(keyinput106), .B1(keyinput8), .B2(n7016), 
        .ZN(n7015) );
  OAI221_X1 U7936 ( .B1(n7017), .B2(keyinput106), .C1(n7016), .C2(keyinput8), 
        .A(n7015), .ZN(n7018) );
  NOR4_X1 U7937 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7022)
         );
  NAND4_X1 U7938 ( .A1(n7025), .A2(n7024), .A3(n7023), .A4(n7022), .ZN(n7026)
         );
  NOR4_X1 U7939 ( .A1(n7029), .A2(n7028), .A3(n7027), .A4(n7026), .ZN(n7030)
         );
  NAND4_X1 U7940 ( .A1(n7033), .A2(n7032), .A3(n7031), .A4(n7030), .ZN(n7047)
         );
  NAND2_X1 U7941 ( .A1(n7034), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n7043) );
  OAI22_X1 U7942 ( .A1(n7038), .A2(n7037), .B1(n7036), .B2(n7035), .ZN(n7039)
         );
  AOI21_X1 U7943 ( .B1(n7041), .B2(n7040), .A(n7039), .ZN(n7042) );
  OAI211_X1 U7944 ( .C1(n7045), .C2(n7044), .A(n7043), .B(n7042), .ZN(n7046)
         );
  XNOR2_X1 U7945 ( .A(n7047), .B(n7046), .ZN(U3067) );
  CLKBUF_X1 U3599 ( .A(n3336), .Z(n4434) );
  CLKBUF_X2 U3603 ( .A(n5437), .Z(n3132) );
  CLKBUF_X1 U3623 ( .A(n3746), .Z(n3134) );
  CLKBUF_X1 U3665 ( .A(n5395), .Z(n5396) );
endmodule

