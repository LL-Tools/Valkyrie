

module b20_C_SARLock_k_128_1 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362;

  INV_X4 U4920 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  XNOR2_X1 U4921 ( .A(n6995), .B(n6996), .ZN(n6861) );
  INV_X2 U4922 ( .A(n9204), .ZN(n9140) );
  INV_X1 U4923 ( .A(n6752), .ZN(n9207) );
  OR2_X1 U4924 ( .A1(n6445), .A2(n6444), .ZN(n6454) );
  CLKBUF_X2 U4925 ( .A(n5186), .Z(n7854) );
  OAI21_X1 U4926 ( .B1(n5709), .B2(n5697), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5698) );
  NAND2_X1 U4927 ( .A1(n5595), .A2(n5596), .ZN(n5181) );
  OAI22_X1 U4929 ( .A1(n6646), .A2(n4839), .B1(n4445), .B2(n10154), .ZN(n10153) );
  NAND2_X1 U4930 ( .A1(n8264), .A2(n8076), .ZN(n8256) );
  INV_X1 U4931 ( .A(n7613), .ZN(n7527) );
  INV_X1 U4933 ( .A(n8256), .ZN(n8249) );
  NAND2_X1 U4934 ( .A1(n8724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5053) );
  INV_X1 U4936 ( .A(n7592), .ZN(n6082) );
  NAND2_X1 U4937 ( .A1(n7722), .A2(n7755), .ZN(n6326) );
  NOR2_X2 U4938 ( .A1(n6316), .A2(n6498), .ZN(n6526) );
  XNOR2_X1 U4939 ( .A(n6980), .B(n6996), .ZN(n6844) );
  NAND2_X1 U4940 ( .A1(n5721), .A2(n5725), .ZN(n7534) );
  OAI21_X1 U4941 ( .B1(n9543), .B2(n7809), .A(n7808), .ZN(n9521) );
  INV_X1 U4942 ( .A(n5179), .ZN(n5939) );
  XNOR2_X1 U4943 ( .A(n5225), .B(n5224), .ZN(n6655) );
  NAND2_X4 U4944 ( .A1(n5759), .A2(n5918), .ZN(n9201) );
  XNOR2_X2 U4945 ( .A(n8071), .B(n4758), .ZN(n7864) );
  NAND2_X2 U4946 ( .A1(n7852), .A2(n7851), .ZN(n8071) );
  NAND2_X4 U4947 ( .A1(n5728), .A2(n5727), .ZN(n6231) );
  NAND4_X2 U4948 ( .A1(n6086), .A2(n6085), .A3(n6084), .A4(n6083), .ZN(n9395)
         );
  OAI21_X2 U4949 ( .B1(n5587), .B2(n4730), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5653) );
  XNOR2_X1 U4950 ( .A(n9397), .B(n6672), .ZN(n7698) );
  NAND4_X2 U4951 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n9397)
         );
  BUF_X8 U4952 ( .A(n5200), .Z(n4414) );
  AOI21_X2 U4953 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10171), .A(n10169), .ZN(
        n7305) );
  AOI21_X2 U4954 ( .B1(n5888), .B2(n5887), .A(n6363), .ZN(n6362) );
  XNOR2_X2 U4955 ( .A(n5156), .B(n5155), .ZN(n5596) );
  NAND2_X4 U4956 ( .A1(n4527), .A2(n4526), .ZN(n5179) );
  NAND3_X2 U4957 ( .A1(n4604), .A2(n4603), .A3(n4602), .ZN(n4527) );
  INV_X1 U4958 ( .A(n7896), .ZN(n7932) );
  INV_X2 U4959 ( .A(n6076), .ZN(n9082) );
  NAND4_X4 U4960 ( .A1(n5204), .A2(n5203), .A3(n5202), .A4(n5201), .ZN(n8283)
         );
  NOR2_X2 U4961 ( .A1(n6454), .A2(n6453), .ZN(n6615) );
  XNOR2_X2 U4962 ( .A(n5053), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8729) );
  XNOR2_X2 U4963 ( .A(n5299), .B(n5019), .ZN(n9023) );
  XNOR2_X2 U4964 ( .A(n9399), .B(n7642), .ZN(n6238) );
  XNOR2_X2 U4965 ( .A(n6841), .B(n6847), .ZN(n6646) );
  CLKBUF_X1 U4966 ( .A(n9946), .Z(n4416) );
  XNOR2_X2 U4967 ( .A(n8372), .B(n8373), .ZN(n8352) );
  NOR2_X2 U4968 ( .A1(n8350), .A2(n4498), .ZN(n8372) );
  AOI21_X2 U4969 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n10155), .A(n10153), .ZN(
        n6980) );
  OR4_X1 U4970 ( .A1(n9211), .A2(n9217), .A3(n9218), .A4(n9370), .ZN(n9222) );
  OAI21_X1 U4971 ( .B1(n9288), .B2(n4912), .A(n4423), .ZN(n9160) );
  NAND2_X1 U4972 ( .A1(n9116), .A2(n9115), .ZN(n9189) );
  NAND2_X1 U4973 ( .A1(n9223), .A2(n4488), .ZN(n9117) );
  NAND2_X1 U4974 ( .A1(n9224), .A2(n9225), .ZN(n9223) );
  NAND2_X1 U4975 ( .A1(n9292), .A2(n9103), .ZN(n9224) );
  INV_X1 U4976 ( .A(n7606), .ZN(n7688) );
  INV_X1 U4977 ( .A(n6957), .ZN(n10272) );
  NOR2_X1 U4978 ( .A1(n6488), .A2(n9394), .ZN(n7465) );
  NAND2_X1 U4979 ( .A1(n6074), .A2(n9201), .ZN(n4417) );
  NAND2_X1 U4980 ( .A1(n5182), .A2(n6211), .ZN(n5601) );
  CLKBUF_X3 U4981 ( .A(n5185), .Z(n5432) );
  INV_X2 U4982 ( .A(n7589), .ZN(n5836) );
  OAI21_X1 U4983 ( .B1(n7724), .B2(n7755), .A(n5012), .ZN(n4967) );
  NAND2_X1 U4984 ( .A1(n9185), .A2(n9286), .ZN(n4641) );
  NAND2_X1 U4985 ( .A1(n4642), .A2(n9187), .ZN(n9185) );
  NAND2_X1 U4986 ( .A1(n9189), .A2(n4863), .ZN(n4642) );
  CLKBUF_X1 U4987 ( .A(n9603), .Z(n4509) );
  NOR2_X1 U4988 ( .A1(n7726), .A2(n5757), .ZN(n5012) );
  NAND2_X1 U4989 ( .A1(n5615), .A2(n8192), .ZN(n8531) );
  AND3_X1 U4990 ( .A1(n4848), .A2(n4850), .A3(n8417), .ZN(n8420) );
  OR2_X1 U4991 ( .A1(n9724), .A2(n9353), .ZN(n7675) );
  OR2_X1 U4992 ( .A1(n7340), .A2(n7339), .ZN(n8298) );
  XNOR2_X1 U4993 ( .A(n6759), .B(n4515), .ZN(n6781) );
  NAND2_X1 U4994 ( .A1(n4671), .A2(n6750), .ZN(n6759) );
  OR2_X1 U4995 ( .A1(n7362), .A2(n7309), .ZN(n4838) );
  OR2_X1 U4996 ( .A1(n6590), .A2(n4740), .ZN(n4737) );
  NAND2_X1 U4997 ( .A1(n8140), .A2(n8141), .ZN(n8134) );
  NAND2_X1 U4998 ( .A1(n5311), .A2(n5310), .ZN(n7181) );
  NAND2_X2 U4999 ( .A1(n6331), .A2(n10042), .ZN(n10067) );
  AND2_X1 U5000 ( .A1(n7700), .A2(n4510), .ZN(n4865) );
  CLKBUF_X3 U5001 ( .A(n6073), .Z(n4514) );
  NAND2_X1 U5002 ( .A1(n5758), .A2(n5756), .ZN(n5759) );
  NAND2_X1 U5003 ( .A1(n4988), .A2(n4987), .ZN(n10205) );
  OR2_X1 U5004 ( .A1(n7546), .A2(n9299), .ZN(n7561) );
  AND4_X1 U5005 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n6962)
         );
  NAND2_X1 U5006 ( .A1(n5755), .A2(n5918), .ZN(n6074) );
  NAND2_X1 U5007 ( .A1(n5757), .A2(n7755), .ZN(n7684) );
  OR2_X1 U5008 ( .A1(n5850), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U5009 ( .A1(n5995), .A2(n5994), .ZN(n6672) );
  CLKBUF_X2 U5010 ( .A(n7835), .Z(n4418) );
  AND2_X1 U5011 ( .A1(n8729), .A2(n8731), .ZN(n5185) );
  CLKBUF_X1 U5012 ( .A(n5056), .Z(n8731) );
  INV_X2 U5013 ( .A(n5426), .ZN(n8060) );
  INV_X2 U5014 ( .A(n7521), .ZN(n7612) );
  CLKBUF_X1 U5015 ( .A(n5288), .Z(n8061) );
  NAND2_X1 U5016 ( .A1(n4465), .A2(n4594), .ZN(n7642) );
  XNOR2_X1 U5017 ( .A(n5754), .B(P1_IR_REG_19__SCAN_IN), .ZN(n7835) );
  XNOR2_X1 U5018 ( .A(n5055), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5056) );
  NAND2_X2 U5019 ( .A1(n9865), .A2(n9870), .ZN(n7592) );
  NAND2_X1 U5020 ( .A1(n5753), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U5021 ( .A1(n5630), .A2(n5629), .ZN(n7143) );
  AND2_X2 U5022 ( .A1(n5725), .A2(n9870), .ZN(n7589) );
  NAND2_X2 U5023 ( .A1(n6253), .A2(n5939), .ZN(n7613) );
  NOR2_X1 U5024 ( .A1(n6366), .A2(n6376), .ZN(n6367) );
  NAND2_X1 U5025 ( .A1(n5630), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5626) );
  NAND2_X1 U5026 ( .A1(n5735), .A2(n5734), .ZN(n7755) );
  INV_X1 U5027 ( .A(n5721), .ZN(n9870) );
  NAND2_X1 U5028 ( .A1(n5054), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5055) );
  XNOR2_X1 U5029 ( .A(n4673), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7722) );
  AND2_X1 U5030 ( .A1(n10124), .A2(n10123), .ZN(n10129) );
  INV_X1 U5031 ( .A(n5725), .ZN(n9865) );
  XNOR2_X1 U5032 ( .A(n5743), .B(n5742), .ZN(n7769) );
  AND2_X1 U5033 ( .A1(n5731), .A2(n5696), .ZN(n5729) );
  XNOR2_X1 U5034 ( .A(n4836), .B(n5744), .ZN(n9946) );
  XNOR2_X1 U5035 ( .A(n5717), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5725) );
  OR2_X1 U5036 ( .A1(n6710), .A2(n6709), .ZN(n6802) );
  NAND2_X1 U5037 ( .A1(n5749), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U5038 ( .A1(n5704), .A2(n4679), .ZN(n5716) );
  NOR2_X2 U5039 ( .A1(n5859), .A2(n5692), .ZN(n5704) );
  INV_X2 U5040 ( .A(n5939), .ZN(n5534) );
  NAND2_X2 U5041 ( .A1(n5939), .A2(P1_U3086), .ZN(n9868) );
  INV_X1 U5042 ( .A(n5427), .ZN(n5049) );
  NOR2_X2 U5043 ( .A1(n5190), .A2(n5209), .ZN(n6375) );
  OR2_X1 U5044 ( .A1(n6306), .A2(n6305), .ZN(n6445) );
  NAND2_X1 U5045 ( .A1(n4842), .A2(n5166), .ZN(n6356) );
  AND2_X1 U5046 ( .A1(n5189), .A2(n4993), .ZN(n4716) );
  CLKBUF_X1 U5047 ( .A(n5779), .Z(n5797) );
  AND2_X1 U5048 ( .A1(n10112), .A2(n4785), .ZN(n5894) );
  AND4_X1 U5049 ( .A1(n5044), .A2(n5043), .A3(n5257), .A4(n5224), .ZN(n5045)
         );
  AND4_X1 U5050 ( .A1(n5047), .A2(n4784), .A3(n4783), .A4(n4782), .ZN(n5048)
         );
  INV_X1 U5051 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5224) );
  INV_X1 U5052 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5750) );
  INV_X1 U5053 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5627) );
  INV_X4 U5054 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5055 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5652) );
  NOR2_X1 U5056 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5044) );
  INV_X1 U5057 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5625) );
  NOR2_X1 U5058 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5689) );
  NOR2_X1 U5059 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5690) );
  NOR2_X1 U5060 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n4639) );
  NAND2_X1 U5061 ( .A1(n6074), .A2(n9201), .ZN(n6073) );
  NAND2_X2 U5062 ( .A1(n5546), .A2(n5545), .ZN(n8475) );
  NOR2_X2 U5063 ( .A1(n7561), .A2(n9230), .ZN(n7573) );
  NAND2_X2 U5064 ( .A1(n7450), .A2(n7828), .ZN(n7829) );
  OR2_X1 U5065 ( .A1(n8445), .A2(n7938), .ZN(n8244) );
  INV_X1 U5066 ( .A(n5362), .ZN(n5119) );
  INV_X1 U5067 ( .A(SI_14_), .ZN(n5118) );
  OR2_X1 U5068 ( .A1(n5618), .A2(n8501), .ZN(n8217) );
  OR2_X1 U5069 ( .A1(n8556), .A2(n8566), .ZN(n8194) );
  NAND2_X1 U5070 ( .A1(n7805), .A2(n4519), .ZN(n9603) );
  OR2_X1 U5071 ( .A1(n9627), .A2(n9380), .ZN(n4519) );
  NAND2_X1 U5072 ( .A1(n9681), .A2(n9340), .ZN(n4894) );
  NAND2_X1 U5073 ( .A1(n4696), .A2(n4458), .ZN(n4693) );
  NOR2_X1 U5074 ( .A1(n4946), .A2(n5113), .ZN(n4944) );
  INV_X1 U5075 ( .A(n5337), .ZN(n5113) );
  NAND2_X1 U5076 ( .A1(n8243), .A2(n8256), .ZN(n4537) );
  OAI21_X1 U5077 ( .B1(n5511), .B2(n4962), .A(n5530), .ZN(n4961) );
  NOR2_X1 U5078 ( .A1(n4997), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4996) );
  INV_X1 U5079 ( .A(n4729), .ZN(n4728) );
  OAI21_X1 U5080 ( .B1(n8511), .B2(n7913), .A(n7951), .ZN(n4729) );
  NAND2_X1 U5081 ( .A1(n4541), .A2(n8249), .ZN(n4538) );
  NAND2_X1 U5082 ( .A1(n5050), .A2(n4998), .ZN(n4997) );
  INV_X1 U5083 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5050) );
  INV_X1 U5084 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4998) );
  INV_X1 U5085 ( .A(n5056), .ZN(n5159) );
  OR2_X1 U5086 ( .A1(n6893), .A2(n5304), .ZN(n4793) );
  OR2_X1 U5087 ( .A1(n5850), .A2(n5648), .ZN(n5669) );
  AND2_X1 U5088 ( .A1(n5637), .A2(n5636), .ZN(n6162) );
  OR2_X1 U5089 ( .A1(n5850), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5637) );
  INV_X1 U5090 ( .A(n8684), .ZN(n5490) );
  AND2_X1 U5091 ( .A1(n8684), .A2(n8525), .ZN(n8202) );
  OR2_X1 U5092 ( .A1(n7274), .A2(n7243), .ZN(n8171) );
  NOR2_X1 U5093 ( .A1(n4995), .A2(n4790), .ZN(n4789) );
  NAND2_X1 U5094 ( .A1(n5013), .A2(n4791), .ZN(n4790) );
  INV_X1 U5095 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4791) );
  INV_X1 U5096 ( .A(n9049), .ZN(n4875) );
  OR2_X1 U5097 ( .A1(n10091), .A2(n6763), .ZN(n7477) );
  NAND2_X1 U5098 ( .A1(n6261), .A2(n7647), .ZN(n7458) );
  INV_X1 U5099 ( .A(n6241), .ZN(n4824) );
  INV_X1 U5100 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5101 ( .B1(n7698), .B2(n4824), .A(n7640), .ZN(n4823) );
  NAND2_X1 U5102 ( .A1(n7814), .A2(n9212), .ZN(n7687) );
  NAND2_X1 U5103 ( .A1(n7391), .A2(n7390), .ZN(n7611) );
  OR2_X1 U5104 ( .A1(n7389), .A2(n7388), .ZN(n7390) );
  OR2_X1 U5105 ( .A1(n7405), .A2(n7387), .ZN(n7391) );
  NAND2_X1 U5106 ( .A1(n5552), .A2(n5551), .ZN(n5571) );
  NAND2_X1 U5107 ( .A1(n5550), .A2(n5549), .ZN(n5552) );
  INV_X1 U5108 ( .A(n5481), .ZN(n4545) );
  AOI21_X1 U5109 ( .B1(n4938), .B2(n4935), .A(n4464), .ZN(n4934) );
  INV_X1 U5110 ( .A(n5139), .ZN(n4935) );
  XNOR2_X1 U5111 ( .A(n5141), .B(SI_20_), .ZN(n5456) );
  AOI21_X1 U5112 ( .B1(n4568), .B2(n4566), .A(n4469), .ZN(n4565) );
  INV_X1 U5113 ( .A(n4440), .ZN(n4566) );
  NAND2_X1 U5114 ( .A1(n5117), .A2(n5116), .ZN(n5364) );
  XNOR2_X1 U5115 ( .A(n5111), .B(SI_12_), .ZN(n5337) );
  AND3_X1 U5116 ( .A1(n4640), .A2(n4639), .A3(n4638), .ZN(n5687) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4640) );
  NAND2_X1 U5118 ( .A1(n4596), .A2(n5075), .ZN(n5251) );
  NAND3_X1 U5119 ( .A1(n4601), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4526) );
  INV_X1 U5120 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4601) );
  INV_X1 U5121 ( .A(n6744), .ZN(n4736) );
  NAND2_X1 U5122 ( .A1(n4712), .A2(n4711), .ZN(n6572) );
  INV_X1 U5123 ( .A(n6479), .ZN(n4711) );
  AND2_X1 U5124 ( .A1(n6150), .A2(n5851), .ZN(n4741) );
  NAND2_X1 U5125 ( .A1(n7962), .A2(n7881), .ZN(n8004) );
  INV_X1 U5126 ( .A(n5184), .ZN(n7857) );
  AND2_X2 U5127 ( .A1(n8729), .A2(n5159), .ZN(n5186) );
  OAI21_X1 U5128 ( .B1(n6657), .B2(n6656), .A(n4442), .ZN(n6658) );
  OR2_X1 U5129 ( .A1(n6861), .A2(n10313), .ZN(n4812) );
  XNOR2_X1 U5130 ( .A(n8239), .B(n8455), .ZN(n8058) );
  INV_X1 U5131 ( .A(n8224), .ZN(n4970) );
  NAND2_X1 U5132 ( .A1(n4781), .A2(n4778), .ZN(n8532) );
  AND2_X1 U5133 ( .A1(n8533), .A2(n4448), .ZN(n4778) );
  INV_X1 U5134 ( .A(n8431), .ZN(n8409) );
  AOI21_X1 U5135 ( .B1(n8175), .B2(n4761), .A(n4459), .ZN(n4760) );
  NAND2_X1 U5136 ( .A1(n8175), .A2(n4763), .ZN(n4762) );
  AND2_X1 U5137 ( .A1(n8180), .A2(n8177), .ZN(n4985) );
  NAND2_X1 U5138 ( .A1(n5181), .A2(n5939), .ZN(n5426) );
  INV_X1 U5139 ( .A(n5181), .ZN(n5256) );
  OR2_X1 U5140 ( .A1(n5490), .A2(n8525), .ZN(n4771) );
  AND2_X1 U5141 ( .A1(n8194), .A2(n8186), .ZN(n4994) );
  OR2_X1 U5142 ( .A1(n8571), .A2(n7967), .ZN(n8186) );
  NAND2_X1 U5144 ( .A1(n5049), .A2(n4789), .ZN(n5634) );
  NAND2_X1 U5145 ( .A1(n5628), .A2(n5627), .ZN(n5630) );
  INV_X1 U5146 ( .A(n7754), .ZN(n7721) );
  AND2_X1 U5147 ( .A1(n9708), .A2(n9384), .ZN(n4516) );
  NAND2_X1 U5148 ( .A1(n7801), .A2(n9068), .ZN(n4517) );
  OAI21_X1 U5149 ( .B1(n9386), .B2(n9309), .A(n7161), .ZN(n7208) );
  NAND2_X1 U5150 ( .A1(n6723), .A2(n6722), .ZN(n6724) );
  OR2_X1 U5151 ( .A1(n10091), .A2(n9390), .ZN(n6722) );
  OR2_X1 U5152 ( .A1(n9729), .A2(n9375), .ZN(n7810) );
  OAI21_X1 U5153 ( .B1(n9603), .B2(n4901), .A(n4899), .ZN(n9554) );
  AOI21_X1 U5154 ( .B1(n4900), .B2(n4902), .A(n4484), .ZN(n4899) );
  NAND2_X1 U5155 ( .A1(n4902), .A2(n4436), .ZN(n4901) );
  NAND2_X1 U5156 ( .A1(n9651), .A2(n5018), .ZN(n9640) );
  AND2_X1 U5157 ( .A1(n4600), .A2(n4894), .ZN(n4891) );
  AND2_X1 U5158 ( .A1(n9840), .A2(n9382), .ZN(n4895) );
  INV_X1 U5159 ( .A(n6253), .ZN(n7526) );
  NAND2_X1 U5160 ( .A1(n6253), .A2(n5534), .ZN(n7521) );
  NAND2_X2 U5161 ( .A1(n7769), .A2(n9946), .ZN(n6253) );
  NAND2_X1 U5162 ( .A1(n4923), .A2(n5718), .ZN(n4922) );
  OR2_X1 U5163 ( .A1(n5729), .A2(n5864), .ZN(n4673) );
  NOR2_X1 U5164 ( .A1(n7462), .A2(n7468), .ZN(n4686) );
  AOI21_X1 U5165 ( .B1(n7472), .B2(n7471), .A(n7470), .ZN(n4688) );
  NOR2_X1 U5166 ( .A1(n7693), .A2(n7666), .ZN(n4690) );
  OR2_X1 U5167 ( .A1(n8208), .A2(n8213), .ZN(n4576) );
  NAND2_X1 U5168 ( .A1(n4699), .A2(n4697), .ZN(n7621) );
  AND2_X1 U5169 ( .A1(n4477), .A2(n4698), .ZN(n4697) );
  NAND2_X1 U5170 ( .A1(n4700), .A2(n4704), .ZN(n4698) );
  AND2_X1 U5171 ( .A1(n7477), .A2(n6700), .ZN(n7474) );
  INV_X1 U5172 ( .A(n4954), .ZN(n4953) );
  OAI21_X1 U5173 ( .B1(n5570), .B2(n4955), .A(n7381), .ZN(n4954) );
  INV_X1 U5174 ( .A(n5572), .ZN(n4955) );
  INV_X1 U5175 ( .A(n5513), .ZN(n4962) );
  NOR2_X1 U5176 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4782) );
  AND3_X1 U5177 ( .A1(n10112), .A2(n4785), .A3(n5046), .ZN(n5189) );
  INV_X1 U5178 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5046) );
  INV_X1 U5179 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4785) );
  NAND2_X1 U5180 ( .A1(n7621), .A2(n9937), .ZN(n4969) );
  NAND2_X1 U5181 ( .A1(n9487), .A2(n4677), .ZN(n4968) );
  AND2_X1 U5182 ( .A1(n9846), .A2(n7802), .ZN(n7665) );
  NOR2_X1 U5183 ( .A1(n9644), .A2(n9648), .ZN(n9624) );
  NOR2_X1 U5184 ( .A1(n4962), .A2(n4958), .ZN(n4957) );
  INV_X1 U5185 ( .A(n5503), .ZN(n4958) );
  AOI21_X1 U5186 ( .B1(n5440), .B2(n5139), .A(n4939), .ZN(n4938) );
  INV_X1 U5187 ( .A(n5456), .ZN(n4939) );
  INV_X1 U5188 ( .A(n5382), .ZN(n5122) );
  NAND2_X1 U5189 ( .A1(n7955), .A2(n4724), .ZN(n7903) );
  OR2_X1 U5190 ( .A1(n7900), .A2(n8272), .ZN(n4724) );
  NAND2_X1 U5191 ( .A1(n4534), .A2(n4537), .ZN(n4533) );
  NAND2_X1 U5192 ( .A1(n4419), .A2(n4429), .ZN(n4534) );
  OR2_X1 U5193 ( .A1(n8245), .A2(n4536), .ZN(n4535) );
  NAND2_X1 U5194 ( .A1(n4537), .A2(n8249), .ZN(n4536) );
  OR2_X1 U5195 ( .A1(n8254), .A2(n4532), .ZN(n4531) );
  NAND2_X1 U5196 ( .A1(n4537), .A2(n7908), .ZN(n4532) );
  AOI21_X1 U5197 ( .B1(n4419), .B2(n4428), .A(n4446), .ZN(n4530) );
  AOI21_X1 U5198 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10116), .A(n10113), .ZN(
        n6377) );
  AND2_X1 U5199 ( .A1(n8298), .A2(n8297), .ZN(n8326) );
  OR2_X1 U5200 ( .A1(n8706), .A2(n8565), .ZN(n8180) );
  INV_X1 U5201 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7286) );
  OR2_X1 U5202 ( .A1(n5328), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5342) );
  OR2_X1 U5203 ( .A1(n5312), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5328) );
  INV_X1 U5204 ( .A(n6211), .ZN(n5183) );
  NAND2_X1 U5205 ( .A1(n8089), .A2(n8090), .ZN(n8036) );
  OR2_X1 U5206 ( .A1(n8667), .A2(n8486), .ZN(n8224) );
  OR2_X1 U5207 ( .A1(n8632), .A2(n7946), .ZN(n8196) );
  OR2_X1 U5208 ( .A1(n8154), .A2(n8274), .ZN(n8158) );
  AND2_X1 U5209 ( .A1(n4789), .A2(n5155), .ZN(n4786) );
  NAND2_X1 U5210 ( .A1(n4996), .A2(n4449), .ZN(n4995) );
  NAND4_X1 U5211 ( .A1(n4716), .A2(n5048), .A3(n5045), .A4(n4715), .ZN(n5427)
         );
  INV_X1 U5212 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4715) );
  INV_X1 U5213 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5685) );
  AND2_X1 U5214 ( .A1(n5017), .A2(n6502), .ZN(n4921) );
  NAND2_X1 U5215 ( .A1(n6631), .A2(n6501), .ZN(n6502) );
  INV_X1 U5216 ( .A(n9194), .ZN(n4652) );
  XNOR2_X1 U5217 ( .A(n5998), .B(n6074), .ZN(n4648) );
  INV_X1 U5218 ( .A(n4617), .ZN(n4616) );
  NOR2_X1 U5219 ( .A1(n7733), .A2(n4618), .ZN(n4617) );
  INV_X1 U5220 ( .A(n7817), .ZN(n4618) );
  NOR2_X1 U5221 ( .A1(n9690), .A2(n9840), .ZN(n9662) );
  NOR2_X1 U5222 ( .A1(n9241), .A2(n9309), .ZN(n4589) );
  INV_X1 U5223 ( .A(n5014), .ZN(n4868) );
  OR2_X1 U5224 ( .A1(n4869), .A2(n7703), .ZN(n4510) );
  NAND2_X1 U5225 ( .A1(n4605), .A2(n4835), .ZN(n9561) );
  NOR2_X1 U5226 ( .A1(n9559), .A2(n9560), .ZN(n4835) );
  XNOR2_X1 U5227 ( .A(n7389), .B(n7388), .ZN(n7405) );
  AND2_X1 U5228 ( .A1(n5532), .A2(n5517), .ZN(n5530) );
  AND2_X1 U5229 ( .A1(n5513), .A2(n5507), .ZN(n5511) );
  INV_X1 U5230 ( .A(n4938), .ZN(n4936) );
  NOR2_X1 U5231 ( .A1(n5749), .A2(n5695), .ZN(n5731) );
  OAI21_X1 U5232 ( .B1(n5364), .B2(n4564), .A(n4466), .ZN(n5410) );
  NAND2_X1 U5233 ( .A1(n4565), .A2(n4482), .ZN(n4564) );
  XNOR2_X1 U5234 ( .A(n5128), .B(SI_17_), .ZN(n5409) );
  XNOR2_X1 U5235 ( .A(n5115), .B(SI_13_), .ZN(n5349) );
  NAND2_X1 U5236 ( .A1(n4550), .A2(n4551), .ZN(n5350) );
  AOI21_X1 U5237 ( .B1(n4553), .B2(n4559), .A(n4552), .ZN(n4551) );
  NOR2_X1 U5238 ( .A1(n4942), .A2(n4554), .ZN(n4553) );
  OAI21_X1 U5239 ( .B1(n5179), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4528), .ZN(
        n5062) );
  NAND2_X1 U5240 ( .A1(n5179), .A2(n5940), .ZN(n4528) );
  AOI21_X1 U5241 ( .B1(n6577), .B2(n4739), .A(n4460), .ZN(n4738) );
  INV_X1 U5242 ( .A(n6591), .ZN(n4739) );
  INV_X1 U5243 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5244 ( .B1(n7889), .B2(n4723), .A(n7943), .ZN(n4722) );
  INV_X1 U5245 ( .A(n10205), .ZN(n5198) );
  AND2_X1 U5246 ( .A1(n8262), .A2(n5882), .ZN(n6142) );
  INV_X1 U5247 ( .A(n8475), .ZN(n8015) );
  NOR2_X1 U5248 ( .A1(n4735), .A2(n4468), .ZN(n4734) );
  INV_X1 U5249 ( .A(n7129), .ZN(n4735) );
  INV_X1 U5250 ( .A(n7189), .ZN(n4733) );
  AND2_X1 U5251 ( .A1(n5196), .A2(n5193), .ZN(n4987) );
  NAND2_X1 U5252 ( .A1(n5184), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5196) );
  AND2_X1 U5253 ( .A1(n5195), .A2(n5194), .ZN(n4988) );
  XNOR2_X1 U5254 ( .A(n6375), .B(n6374), .ZN(n10115) );
  NAND2_X1 U5255 ( .A1(n4861), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4859) );
  OR2_X1 U5256 ( .A1(n6645), .A2(n6644), .ZN(n6841) );
  INV_X1 U5257 ( .A(n6658), .ZN(n4802) );
  NAND2_X1 U5258 ( .A1(n4838), .A2(n4837), .ZN(n8288) );
  INV_X1 U5259 ( .A(n7312), .ZN(n4837) );
  OR2_X1 U5260 ( .A1(n5351), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5352) );
  XNOR2_X1 U5261 ( .A(n8326), .B(n4511), .ZN(n8299) );
  NOR2_X1 U5262 ( .A1(n8299), .A2(n8300), .ZN(n8328) );
  AND2_X1 U5263 ( .A1(n8288), .A2(n8287), .ZN(n8310) );
  INV_X1 U5264 ( .A(n8362), .ZN(n4847) );
  INV_X1 U5265 ( .A(n8412), .ZN(n8413) );
  NAND2_X1 U5266 ( .A1(n4849), .A2(n4421), .ZN(n4848) );
  NAND2_X1 U5267 ( .A1(n4747), .A2(n10207), .ZN(n4745) );
  NAND2_X1 U5268 ( .A1(n4748), .A2(n4752), .ZN(n4747) );
  NAND2_X1 U5269 ( .A1(n7853), .A2(n4753), .ZN(n4752) );
  NOR2_X1 U5270 ( .A1(n4746), .A2(n10225), .ZN(n4744) );
  AND2_X1 U5271 ( .A1(n4748), .A2(n4479), .ZN(n4746) );
  OR2_X1 U5272 ( .A1(n8667), .A2(n8272), .ZN(n5529) );
  NAND2_X1 U5273 ( .A1(n5520), .A2(n8831), .ZN(n5540) );
  NOR2_X1 U5274 ( .A1(n8687), .A2(n8536), .ZN(n5480) );
  OR2_X1 U5275 ( .A1(n5460), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5475) );
  OR2_X1 U5276 ( .A1(n5430), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5450) );
  OR2_X1 U5277 ( .A1(n5403), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5415) );
  OR2_X1 U5278 ( .A1(n5373), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5389) );
  AND4_X1 U5279 ( .A1(n5378), .A2(n5377), .A3(n5376), .A4(n5375), .ZN(n7243)
         );
  NAND2_X1 U5280 ( .A1(n5032), .A2(n7286), .ZN(n5355) );
  INV_X1 U5281 ( .A(n5342), .ZN(n5032) );
  AOI21_X1 U5282 ( .B1(n8045), .B2(n8137), .A(n4982), .ZN(n4981) );
  INV_X1 U5283 ( .A(n8141), .ZN(n4982) );
  AOI21_X1 U5284 ( .B1(n7051), .B2(n5336), .A(n4444), .ZN(n7101) );
  NAND2_X1 U5285 ( .A1(n4971), .A2(n4974), .ZN(n6890) );
  AOI21_X1 U5286 ( .B1(n4976), .B2(n8130), .A(n4975), .ZN(n4974) );
  INV_X1 U5287 ( .A(n8126), .ZN(n4975) );
  OR2_X1 U5288 ( .A1(n5278), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U5289 ( .A1(n5027), .A2(n5026), .ZN(n5244) );
  INV_X1 U5290 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5026) );
  NAND2_X1 U5291 ( .A1(n5197), .A2(n8036), .ZN(n10227) );
  AND2_X1 U5292 ( .A1(n8409), .A2(n8260), .ZN(n6194) );
  AND3_X1 U5293 ( .A1(n6141), .A2(n5622), .A3(n10282), .ZN(n10230) );
  NOR2_X1 U5294 ( .A1(n5164), .A2(n5534), .ZN(n4742) );
  NAND2_X1 U5295 ( .A1(n6164), .A2(n6163), .ZN(n6170) );
  NAND2_X1 U5296 ( .A1(n5539), .A2(n5538), .ZN(n8012) );
  NAND2_X1 U5297 ( .A1(n4990), .A2(n8206), .ZN(n4989) );
  INV_X1 U5298 ( .A(n8512), .ZN(n4768) );
  NAND2_X1 U5299 ( .A1(n5597), .A2(n8249), .ZN(n10220) );
  INV_X1 U5300 ( .A(n10202), .ZN(n10221) );
  NAND2_X1 U5301 ( .A1(n8513), .A2(n8207), .ZN(n4992) );
  NOR2_X1 U5302 ( .A1(n8546), .A2(n4780), .ZN(n4779) );
  INV_X1 U5303 ( .A(n5438), .ZN(n4780) );
  NAND2_X1 U5304 ( .A1(n5614), .A2(n5613), .ZN(n8561) );
  AND2_X1 U5305 ( .A1(n8194), .A2(n8192), .ZN(n8546) );
  NOR2_X1 U5306 ( .A1(n7300), .A2(n7875), .ZN(n4761) );
  NAND2_X1 U5307 ( .A1(n8584), .A2(n8179), .ZN(n4986) );
  OR2_X1 U5308 ( .A1(n8712), .A2(n7875), .ZN(n8177) );
  NOR2_X1 U5309 ( .A1(n8050), .A2(n4777), .ZN(n4776) );
  INV_X1 U5310 ( .A(n5381), .ZN(n4777) );
  OR2_X1 U5311 ( .A1(n8051), .A2(n8050), .ZN(n8596) );
  AND2_X1 U5312 ( .A1(n8171), .A2(n8163), .ZN(n8165) );
  INV_X1 U5313 ( .A(n10220), .ZN(n10204) );
  AND2_X1 U5314 ( .A1(n6048), .A2(n6059), .ZN(n6144) );
  NAND2_X1 U5315 ( .A1(n5635), .A2(n5856), .ZN(n5850) );
  NAND2_X1 U5316 ( .A1(n5634), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5156) );
  NOR2_X1 U5317 ( .A1(n4995), .A2(n4788), .ZN(n4787) );
  INV_X1 U5318 ( .A(n5013), .ZN(n4788) );
  NAND2_X1 U5319 ( .A1(n5624), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5628) );
  AND2_X1 U5320 ( .A1(n5586), .A2(n4430), .ZN(n8076) );
  INV_X1 U5321 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5445) );
  INV_X1 U5322 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5442) );
  INV_X1 U5323 ( .A(n5894), .ZN(n4842) );
  NAND3_X1 U5324 ( .A1(n4918), .A2(n4920), .A3(n4672), .ZN(n4671) );
  INV_X1 U5325 ( .A(n6508), .ZN(n4672) );
  AND2_X1 U5326 ( .A1(n4870), .A2(n4669), .ZN(n4668) );
  NAND2_X1 U5327 ( .A1(n4872), .A2(n4670), .ZN(n4669) );
  AOI21_X1 U5328 ( .B1(n4872), .B2(n4875), .A(n4489), .ZN(n4870) );
  NAND2_X1 U5329 ( .A1(n9117), .A2(n4864), .ZN(n4863) );
  INV_X1 U5330 ( .A(n9314), .ZN(n4864) );
  AOI21_X1 U5331 ( .B1(n4463), .B2(n4661), .A(n4658), .ZN(n4657) );
  INV_X1 U5332 ( .A(n9337), .ZN(n4658) );
  AND2_X1 U5333 ( .A1(n5761), .A2(n5760), .ZN(n5936) );
  AND2_X1 U5334 ( .A1(n9132), .A2(n9131), .ZN(n9284) );
  AND2_X1 U5335 ( .A1(n5767), .A2(n5766), .ZN(n5937) );
  AOI21_X1 U5336 ( .B1(n4662), .B2(n9078), .A(n4499), .ZN(n4661) );
  INV_X1 U5337 ( .A(n9246), .ZN(n4912) );
  NAND2_X1 U5338 ( .A1(n9246), .A2(n4911), .ZN(n4910) );
  INV_X1 U5339 ( .A(n9132), .ZN(n4911) );
  OR2_X1 U5340 ( .A1(n7779), .A2(n4418), .ZN(n5756) );
  AND4_X1 U5341 ( .A1(n7444), .A2(n7443), .A3(n7442), .A4(n7441), .ZN(n9351)
         );
  AND4_X1 U5342 ( .A1(n7156), .A2(n7155), .A3(n7154), .A4(n7153), .ZN(n9068)
         );
  AND4_X1 U5343 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n9042)
         );
  AND4_X1 U5344 ( .A1(n6451), .A2(n6450), .A3(n6449), .A4(n6448), .ZN(n6753)
         );
  OR2_X1 U5345 ( .A1(n7440), .A2(n10101), .ZN(n5930) );
  INV_X1 U5346 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5752) );
  NOR2_X1 U5347 ( .A1(n9487), .A2(n4584), .ZN(n4582) );
  INV_X1 U5348 ( .A(n4582), .ZN(n4579) );
  NOR2_X1 U5349 ( .A1(n4452), .A2(n4433), .ZN(n4622) );
  OR2_X1 U5350 ( .A1(n9511), .A2(n4627), .ZN(n4623) );
  NAND2_X1 U5351 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  OR2_X1 U5352 ( .A1(n9808), .A2(n9351), .ZN(n9522) );
  NAND2_X1 U5353 ( .A1(n9561), .A2(n7823), .ZN(n9538) );
  NAND2_X1 U5354 ( .A1(n9538), .A2(n9542), .ZN(n9537) );
  NOR2_X1 U5355 ( .A1(n9597), .A2(n9742), .ZN(n9580) );
  NAND2_X1 U5356 ( .A1(n7821), .A2(n7820), .ZN(n9572) );
  AND2_X1 U5357 ( .A1(n9648), .A2(n9381), .ZN(n7803) );
  NAND2_X1 U5358 ( .A1(n9676), .A2(n4818), .ZN(n9657) );
  NOR2_X1 U5359 ( .A1(n9654), .A2(n7666), .ZN(n4818) );
  OAI21_X1 U5360 ( .B1(n7730), .B2(n4600), .A(n4598), .ZN(n9674) );
  INV_X1 U5361 ( .A(n4599), .ZN(n4598) );
  OAI21_X1 U5362 ( .B1(n4600), .B2(n7729), .A(n7731), .ZN(n4599) );
  NOR2_X1 U5363 ( .A1(n6812), .A2(n9333), .ZN(n6919) );
  NAND2_X1 U5364 ( .A1(n6918), .A2(n4878), .ZN(n7090) );
  OR2_X1 U5365 ( .A1(n9333), .A2(n9388), .ZN(n4878) );
  OR2_X1 U5366 ( .A1(n6916), .A2(n9038), .ZN(n5006) );
  NAND2_X1 U5367 ( .A1(n6256), .A2(n7648), .ZN(n7700) );
  NAND2_X1 U5368 ( .A1(n4822), .A2(n4824), .ZN(n4820) );
  NAND2_X1 U5369 ( .A1(n6292), .A2(n7698), .ZN(n6291) );
  OR2_X1 U5370 ( .A1(n6398), .A2(n6672), .ZN(n6288) );
  OR2_X1 U5371 ( .A1(n6095), .A2(n6098), .ZN(n9664) );
  NOR2_X1 U5372 ( .A1(n5938), .A2(n5939), .ZN(n4593) );
  NAND2_X1 U5373 ( .A1(n7423), .A2(n7422), .ZN(n9724) );
  NAND2_X1 U5374 ( .A1(n7427), .A2(n7426), .ZN(n9729) );
  AOI21_X1 U5375 ( .B1(n4904), .B2(n4903), .A(n4491), .ZN(n4902) );
  INV_X1 U5376 ( .A(n4481), .ZN(n4903) );
  INV_X1 U5377 ( .A(n9600), .ZN(n9747) );
  NAND2_X1 U5378 ( .A1(n7560), .A2(n7559), .ZN(n9752) );
  NAND2_X1 U5379 ( .A1(n4885), .A2(n4887), .ZN(n9651) );
  AND2_X1 U5380 ( .A1(n9654), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U5381 ( .A1(n4889), .A2(n4890), .ZN(n4888) );
  OR2_X1 U5382 ( .A1(n4588), .A2(n9057), .ZN(n5007) );
  AND2_X1 U5383 ( .A1(n7508), .A2(n7729), .ZN(n7714) );
  INV_X1 U5384 ( .A(n7642), .ZN(n10080) );
  OR2_X1 U5385 ( .A1(n5926), .A2(n6095), .ZN(n10094) );
  OR3_X1 U5386 ( .A1(n6325), .A2(n6323), .A3(n6094), .ZN(n6432) );
  NAND2_X1 U5387 ( .A1(n5905), .A2(n5904), .ZN(n9854) );
  XNOR2_X1 U5388 ( .A(n7400), .B(n7399), .ZN(n8723) );
  OAI21_X1 U5389 ( .B1(n7611), .B2(n7610), .A(n7397), .ZN(n7400) );
  XNOR2_X1 U5390 ( .A(n7611), .B(n7610), .ZN(n8728) );
  NAND2_X1 U5391 ( .A1(n9857), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5719) );
  XNOR2_X1 U5392 ( .A(n7405), .B(SI_29_), .ZN(n7848) );
  XNOR2_X1 U5393 ( .A(n5571), .B(n5570), .ZN(n7421) );
  AND2_X1 U5394 ( .A1(n5703), .A2(n4680), .ZN(n4679) );
  INV_X1 U5395 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4680) );
  XNOR2_X1 U5396 ( .A(n5531), .B(n5530), .ZN(n7435) );
  NAND2_X1 U5397 ( .A1(n4959), .A2(n5513), .ZN(n5531) );
  NAND2_X1 U5398 ( .A1(n5512), .A2(n5511), .ZN(n4959) );
  XNOR2_X1 U5399 ( .A(n5512), .B(n5511), .ZN(n7598) );
  NAND2_X1 U5400 ( .A1(n4542), .A2(n4543), .ZN(n5502) );
  AOI21_X1 U5401 ( .B1(n4422), .B2(n4932), .A(n4544), .ZN(n4543) );
  INV_X1 U5402 ( .A(n5148), .ZN(n4544) );
  NAND2_X1 U5403 ( .A1(n4546), .A2(n4441), .ZN(n5482) );
  NAND2_X1 U5404 ( .A1(n4547), .A2(n4931), .ZN(n4546) );
  INV_X1 U5405 ( .A(n5425), .ZN(n4547) );
  NAND2_X1 U5406 ( .A1(n4937), .A2(n5139), .ZN(n5457) );
  OR2_X1 U5407 ( .A1(n5441), .A2(n5440), .ZN(n4937) );
  NAND2_X1 U5408 ( .A1(n5751), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U5409 ( .A1(n4562), .A2(n4565), .ZN(n5398) );
  NAND2_X1 U5410 ( .A1(n5364), .A2(n4568), .ZN(n4562) );
  NAND2_X1 U5411 ( .A1(n4570), .A2(n5120), .ZN(n5384) );
  NAND2_X1 U5412 ( .A1(n4571), .A2(n4440), .ZN(n4570) );
  NAND2_X1 U5413 ( .A1(n4945), .A2(n4943), .ZN(n5338) );
  INV_X1 U5414 ( .A(n4946), .ZN(n4943) );
  NAND2_X1 U5415 ( .A1(n5307), .A2(n4948), .ZN(n4945) );
  OAI21_X1 U5416 ( .B1(n5307), .B2(n5105), .A(n5104), .ZN(n5319) );
  INV_X1 U5417 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U5418 ( .A1(n4597), .A2(n5072), .ZN(n5223) );
  NAND2_X1 U5419 ( .A1(n5857), .A2(n5651), .ZN(n5879) );
  NAND2_X1 U5420 ( .A1(n8003), .A2(n7884), .ZN(n7987) );
  NAND2_X1 U5421 ( .A1(n4710), .A2(n7877), .ZN(n7964) );
  AND3_X1 U5422 ( .A1(n5059), .A2(n5058), .A3(n5057), .ZN(n8511) );
  NAND2_X1 U5423 ( .A1(n6473), .A2(n6472), .ZN(n4714) );
  INV_X1 U5424 ( .A(n8277), .ZN(n7114) );
  AND4_X1 U5425 ( .A1(n5455), .A2(n5454), .A3(n5453), .A4(n5452), .ZN(n8566)
         );
  AND2_X1 U5426 ( .A1(n8032), .A2(n5594), .ZN(n7938) );
  OAI211_X1 U5427 ( .C1(n7857), .C2(n8682), .A(n5489), .B(n5488), .ZN(n8525)
         );
  INV_X1 U5428 ( .A(n7875), .ZN(n8599) );
  NAND4_X1 U5429 ( .A1(n5221), .A2(n5220), .A3(n5219), .A4(n5218), .ZN(n10203)
         );
  INV_X1 U5430 ( .A(n4812), .ZN(n6997) );
  XNOR2_X1 U5431 ( .A(n8310), .B(n4511), .ZN(n8289) );
  OR2_X1 U5432 ( .A1(n8340), .A2(n8341), .ZN(n4846) );
  NOR2_X1 U5433 ( .A1(n8428), .A2(n8427), .ZN(n9890) );
  NAND2_X1 U5434 ( .A1(n5429), .A2(n5428), .ZN(n8571) );
  OR2_X1 U5435 ( .A1(n7522), .A2(n5426), .ZN(n5429) );
  INV_X1 U5436 ( .A(n8652), .ZN(n8606) );
  NAND2_X1 U5437 ( .A1(n5574), .A2(n5573), .ZN(n8239) );
  OR2_X1 U5438 ( .A1(n5623), .A2(n10294), .ZN(n5009) );
  INV_X1 U5439 ( .A(n8012), .ZN(n8665) );
  INV_X1 U5440 ( .A(n6488), .ZN(n6428) );
  NAND2_X1 U5441 ( .A1(n4967), .A2(n4965), .ZN(n4964) );
  AOI21_X1 U5442 ( .B1(n7761), .B2(n7762), .A(n4966), .ZN(n4965) );
  INV_X1 U5443 ( .A(n7779), .ZN(n7766) );
  INV_X1 U5444 ( .A(n9729), .ZN(n9534) );
  NAND2_X1 U5445 ( .A1(n9023), .A2(n7612), .ZN(n6606) );
  INV_X1 U5446 ( .A(n6342), .ZN(n6669) );
  AOI21_X1 U5447 ( .B1(n4426), .B2(n4420), .A(n4880), .ZN(n4879) );
  OR2_X1 U5448 ( .A1(n10100), .A2(n7832), .ZN(n4636) );
  NAND2_X1 U5449 ( .A1(n4828), .A2(n4832), .ZN(n4827) );
  NOR2_X1 U5450 ( .A1(n7836), .A2(n4833), .ZN(n4832) );
  INV_X1 U5451 ( .A(n7843), .ZN(n4828) );
  AND2_X1 U5452 ( .A1(n7814), .A2(n9767), .ZN(n4833) );
  NAND2_X1 U5453 ( .A1(n10100), .A2(n10096), .ZN(n9842) );
  NAND2_X1 U5454 ( .A1(n5748), .A2(n5747), .ZN(n7779) );
  OR2_X1 U5455 ( .A1(n5746), .A2(n5745), .ZN(n5747) );
  NOR2_X1 U5456 ( .A1(n7037), .A2(n7036), .ZN(n10341) );
  NOR2_X1 U5457 ( .A1(n10343), .A2(n10342), .ZN(n7036) );
  NAND2_X1 U5458 ( .A1(n4676), .A2(n4678), .ZN(n7466) );
  NAND2_X1 U5459 ( .A1(n7458), .A2(n4453), .ZN(n4678) );
  NAND2_X1 U5460 ( .A1(n7471), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5461 ( .A1(n4696), .A2(n4427), .ZN(n4689) );
  NAND2_X1 U5462 ( .A1(n4696), .A2(n4432), .ZN(n4694) );
  NOR2_X1 U5463 ( .A1(n8491), .A2(n4576), .ZN(n4575) );
  INV_X1 U5464 ( .A(n8209), .ZN(n4577) );
  NAND2_X1 U5465 ( .A1(n8211), .A2(n8210), .ZN(n4574) );
  NAND2_X1 U5466 ( .A1(n7602), .A2(n9559), .ZN(n4705) );
  AND2_X1 U5467 ( .A1(n4707), .A2(n4701), .ZN(n4700) );
  NAND2_X1 U5468 ( .A1(n4703), .A2(n4702), .ZN(n4701) );
  INV_X1 U5469 ( .A(n7609), .ZN(n4707) );
  INV_X1 U5470 ( .A(n7602), .ZN(n4702) );
  OR2_X1 U5471 ( .A1(n7456), .A2(n7678), .ZN(n4706) );
  INV_X1 U5472 ( .A(n5019), .ZN(n4561) );
  NAND2_X1 U5473 ( .A1(n10205), .A2(n10219), .ZN(n8089) );
  INV_X1 U5474 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5257) );
  NAND2_X1 U5475 ( .A1(n7470), .A2(n7474), .ZN(n6696) );
  OR2_X1 U5476 ( .A1(n9719), .A2(n9208), .ZN(n7450) );
  AND2_X1 U5477 ( .A1(n9534), .A2(n9375), .ZN(n7606) );
  NAND2_X1 U5478 ( .A1(n4951), .A2(n4950), .ZN(n7389) );
  AOI21_X1 U5479 ( .B1(n4953), .B2(n4955), .A(n4503), .ZN(n4950) );
  NAND2_X1 U5480 ( .A1(n5571), .A2(n4953), .ZN(n4951) );
  INV_X1 U5481 ( .A(n5396), .ZN(n5125) );
  INV_X1 U5482 ( .A(SI_16_), .ZN(n5124) );
  INV_X1 U5483 ( .A(n4944), .ZN(n4942) );
  INV_X1 U5484 ( .A(n4556), .ZN(n4554) );
  INV_X1 U5485 ( .A(n4940), .ZN(n4552) );
  AOI21_X1 U5486 ( .B1(n4944), .B2(n4941), .A(n4470), .ZN(n4940) );
  INV_X1 U5487 ( .A(n4948), .ZN(n4941) );
  INV_X1 U5488 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5489 ( .A1(n5107), .A2(n8826), .ZN(n5110) );
  AOI21_X1 U5490 ( .B1(n4560), .B2(n4558), .A(n4557), .ZN(n4556) );
  INV_X1 U5491 ( .A(n5101), .ZN(n4557) );
  INV_X1 U5492 ( .A(n5096), .ZN(n4558) );
  NOR2_X1 U5493 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4638) );
  OR2_X1 U5494 ( .A1(n5078), .A2(n5077), .ZN(n5080) );
  INV_X1 U5495 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4602) );
  INV_X1 U5496 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4604) );
  NOR2_X1 U5497 ( .A1(n10162), .A2(n4522), .ZN(n7330) );
  NOR2_X1 U5498 ( .A1(n6999), .A2(n10315), .ZN(n4522) );
  AND3_X1 U5499 ( .A1(n4805), .A2(n4495), .A3(n4803), .ZN(n7335) );
  INV_X1 U5500 ( .A(n4754), .ZN(n4753) );
  OAI22_X1 U5501 ( .A1(n7846), .A2(n4755), .B1(n8242), .B2(n7908), .ZN(n4754)
         );
  NAND2_X1 U5502 ( .A1(n5569), .A2(n5568), .ZN(n4755) );
  NOR2_X1 U5503 ( .A1(n7846), .A2(n4757), .ZN(n4756) );
  INV_X1 U5504 ( .A(n5568), .ZN(n4757) );
  OAI21_X1 U5505 ( .B1(n4758), .B2(n4750), .A(n4749), .ZN(n4748) );
  NAND2_X1 U5506 ( .A1(n4758), .A2(n4753), .ZN(n4749) );
  AND2_X1 U5507 ( .A1(n4753), .A2(n4751), .ZN(n4750) );
  INV_X1 U5508 ( .A(n4756), .ZN(n4751) );
  OR2_X1 U5509 ( .A1(n8034), .A2(n8228), .ZN(n8223) );
  INV_X1 U5510 ( .A(n8585), .ZN(n4763) );
  NOR2_X1 U5511 ( .A1(n8134), .A2(n4980), .ZN(n4979) );
  INV_X1 U5512 ( .A(n8129), .ZN(n4980) );
  NOR2_X1 U5513 ( .A1(n4977), .A2(n4973), .ZN(n4972) );
  INV_X1 U5514 ( .A(n8130), .ZN(n4977) );
  NAND2_X1 U5515 ( .A1(n6822), .A2(n5291), .ZN(n6904) );
  NAND2_X1 U5516 ( .A1(n5605), .A2(n8114), .ZN(n6819) );
  INV_X1 U5517 ( .A(n5199), .ZN(n4775) );
  NAND2_X1 U5518 ( .A1(n5174), .A2(n5183), .ZN(n8080) );
  OR2_X1 U5519 ( .A1(n8012), .A2(n8015), .ZN(n8230) );
  AND2_X1 U5520 ( .A1(n8012), .A2(n8015), .ZN(n8228) );
  NOR2_X1 U5521 ( .A1(n8658), .A2(n8463), .ZN(n8233) );
  OR2_X1 U5522 ( .A1(n8687), .A2(n8510), .ZN(n8199) );
  INV_X1 U5523 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4993) );
  NOR2_X1 U5524 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5047) );
  NOR2_X1 U5525 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4784) );
  NOR2_X1 U5526 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4783) );
  OR2_X1 U5527 ( .A1(n5308), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5320) );
  INV_X1 U5528 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5155) );
  INV_X1 U5529 ( .A(SI_9_), .ZN(n8798) );
  INV_X1 U5530 ( .A(SI_11_), .ZN(n8826) );
  INV_X1 U5531 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5208) );
  OR2_X1 U5532 ( .A1(n9235), .A2(n4875), .ZN(n4874) );
  INV_X1 U5533 ( .A(n9327), .ZN(n4670) );
  NAND2_X1 U5534 ( .A1(n4969), .A2(n4968), .ZN(n7620) );
  AND2_X1 U5535 ( .A1(n7428), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n7407) );
  OAI21_X1 U5536 ( .B1(n4629), .B2(n7830), .A(n4625), .ZN(n4624) );
  NAND2_X1 U5537 ( .A1(n4629), .A2(n4626), .ZN(n4625) );
  NAND2_X1 U5538 ( .A1(n4632), .A2(n4628), .ZN(n4626) );
  INV_X1 U5539 ( .A(n7830), .ZN(n4628) );
  AOI21_X1 U5540 ( .B1(n4631), .B2(n4633), .A(n4630), .ZN(n4629) );
  INV_X1 U5541 ( .A(n7828), .ZN(n4630) );
  NAND2_X1 U5542 ( .A1(n9572), .A2(n9570), .ZN(n4605) );
  NAND2_X1 U5543 ( .A1(n9635), .A2(n9636), .ZN(n4619) );
  INV_X1 U5544 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6453) );
  NOR2_X1 U5545 ( .A1(n6757), .A2(n6532), .ZN(n4592) );
  INV_X1 U5546 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6305) );
  AND2_X1 U5547 ( .A1(n6699), .A2(n6695), .ZN(n7471) );
  AND2_X1 U5548 ( .A1(n7766), .A2(n7722), .ZN(n7752) );
  AND2_X1 U5549 ( .A1(n4905), .A2(n4436), .ZN(n4900) );
  NAND2_X1 U5550 ( .A1(n9610), .A2(n9747), .ZN(n9597) );
  NOR2_X1 U5551 ( .A1(n9625), .A2(n9752), .ZN(n9610) );
  NAND2_X1 U5552 ( .A1(n9624), .A2(n9828), .ZN(n9625) );
  INV_X1 U5553 ( .A(n4891), .ZN(n4889) );
  AND2_X1 U5554 ( .A1(n6919), .A2(n4585), .ZN(n9691) );
  NOR2_X1 U5555 ( .A1(n9708), .A2(n4587), .ZN(n4585) );
  NAND2_X1 U5556 ( .A1(n10080), .A2(n10061), .ZN(n6398) );
  AND2_X1 U5557 ( .A1(n5907), .A2(n9855), .ZN(n6325) );
  NAND2_X1 U5558 ( .A1(n4925), .A2(n5742), .ZN(n4924) );
  INV_X1 U5559 ( .A(n4926), .ZN(n4925) );
  INV_X1 U5560 ( .A(n4924), .ZN(n4923) );
  NAND2_X1 U5561 ( .A1(n5533), .A2(n5532), .ZN(n5550) );
  NAND2_X1 U5562 ( .A1(n4956), .A2(n4960), .ZN(n5533) );
  INV_X1 U5563 ( .A(n4961), .ZN(n4960) );
  AND2_X1 U5564 ( .A1(n5551), .A2(n5537), .ZN(n5549) );
  NAND2_X1 U5565 ( .A1(n4931), .A2(n4549), .ZN(n4548) );
  AOI21_X1 U5566 ( .B1(n4931), .B2(n4936), .A(n4492), .ZN(n4930) );
  INV_X1 U5567 ( .A(n5136), .ZN(n4549) );
  INV_X1 U5568 ( .A(n5120), .ZN(n4569) );
  INV_X1 U5569 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n5121) );
  INV_X1 U5570 ( .A(n5364), .ZN(n4571) );
  NOR2_X1 U5571 ( .A1(n5318), .A2(n4949), .ZN(n4948) );
  INV_X1 U5572 ( .A(n5104), .ZN(n4949) );
  OAI21_X1 U5573 ( .B1(n5318), .B2(n4947), .A(n5110), .ZN(n4946) );
  NAND2_X1 U5574 ( .A1(n5105), .A2(n5104), .ZN(n4947) );
  NAND2_X1 U5575 ( .A1(n4555), .A2(n4556), .ZN(n5307) );
  OR2_X1 U5576 ( .A1(n5287), .A2(n4559), .ZN(n4555) );
  INV_X1 U5577 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5087) );
  NAND3_X1 U5578 ( .A1(n5685), .A2(n4675), .A3(n4674), .ZN(n5779) );
  INV_X1 U5579 ( .A(n4996), .ZN(n4730) );
  INV_X1 U5580 ( .A(n6577), .ZN(n4740) );
  XNOR2_X1 U5581 ( .A(n7061), .B(n7059), .ZN(n6958) );
  NAND2_X1 U5582 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  AND2_X1 U5583 ( .A1(n7899), .A2(n7952), .ZN(n4726) );
  INV_X1 U5584 ( .A(n7965), .ZN(n4708) );
  INV_X1 U5585 ( .A(n7964), .ZN(n4709) );
  NAND2_X1 U5586 ( .A1(n5031), .A2(n5030), .ZN(n5312) );
  INV_X1 U5587 ( .A(n5293), .ZN(n5031) );
  NAND2_X1 U5588 ( .A1(n4720), .A2(n4718), .ZN(n7994) );
  AOI21_X1 U5589 ( .B1(n4721), .B2(n4723), .A(n4719), .ZN(n4718) );
  INV_X1 U5590 ( .A(n7893), .ZN(n4719) );
  NAND2_X1 U5591 ( .A1(n7192), .A2(n7189), .ZN(n7247) );
  AND2_X1 U5592 ( .A1(n5650), .A2(n5674), .ZN(n6048) );
  NAND2_X1 U5593 ( .A1(n4530), .A2(n4529), .ZN(n4539) );
  AOI21_X1 U5594 ( .B1(n8606), .B2(n8243), .A(n6939), .ZN(n5002) );
  AND4_X1 U5595 ( .A1(n5249), .A2(n5248), .A3(n5247), .A4(n5246), .ZN(n6824)
         );
  AND4_X1 U5596 ( .A1(n5173), .A2(n5170), .A3(n5172), .A4(n5171), .ZN(n5182)
         );
  NAND2_X1 U5597 ( .A1(n4841), .A2(n6371), .ZN(n5895) );
  AND2_X1 U5598 ( .A1(n4859), .A2(n4860), .ZN(n6381) );
  AOI21_X1 U5599 ( .B1(n6650), .B2(n6655), .A(n6649), .ZN(n6651) );
  NOR2_X1 U5600 ( .A1(n6651), .A2(n6652), .ZN(n6846) );
  AND3_X1 U5601 ( .A1(n4800), .A2(n6857), .A3(P2_REG1_REG_5__SCAN_IN), .ZN(
        n6859) );
  AOI21_X1 U5602 ( .B1(n6848), .B2(n6847), .A(n6846), .ZN(n10151) );
  OR2_X1 U5603 ( .A1(n10154), .A2(n6647), .ZN(n4839) );
  OR2_X1 U5604 ( .A1(n6646), .A2(n6647), .ZN(n4840) );
  OAI21_X1 U5605 ( .B1(n6844), .B2(n4854), .A(n4853), .ZN(n10169) );
  NAND2_X1 U5606 ( .A1(n4855), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4854) );
  NAND2_X1 U5607 ( .A1(n6982), .A2(n4855), .ZN(n4853) );
  INV_X1 U5608 ( .A(n10170), .ZN(n4855) );
  XNOR2_X1 U5609 ( .A(n7330), .B(n9021), .ZN(n7000) );
  AOI21_X1 U5610 ( .B1(n7317), .B2(n7316), .A(n7315), .ZN(n10188) );
  NOR2_X1 U5611 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  OAI21_X1 U5612 ( .B1(n6983), .B2(n4857), .A(n4856), .ZN(n10189) );
  NAND2_X1 U5613 ( .A1(n4858), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5614 ( .A1(n7307), .A2(n4858), .ZN(n4856) );
  INV_X1 U5615 ( .A(n10190), .ZN(n4858) );
  OR2_X1 U5616 ( .A1(n7000), .A2(n4806), .ZN(n4805) );
  OR2_X1 U5617 ( .A1(n10181), .A2(n10317), .ZN(n4806) );
  NAND2_X1 U5618 ( .A1(n7332), .A2(n4804), .ZN(n4803) );
  INV_X1 U5619 ( .A(n10181), .ZN(n4804) );
  NOR2_X1 U5620 ( .A1(n7320), .A2(n10186), .ZN(n7370) );
  NOR2_X1 U5621 ( .A1(n7370), .A2(n7371), .ZN(n7369) );
  XNOR2_X1 U5622 ( .A(n7335), .B(n7334), .ZN(n7365) );
  NOR2_X1 U5623 ( .A1(n7323), .A2(n7369), .ZN(n8293) );
  NOR2_X1 U5624 ( .A1(n8328), .A2(n8329), .ZN(n8332) );
  OAI21_X1 U5625 ( .B1(n8352), .B2(n4815), .A(n4814), .ZN(n8396) );
  NAND2_X1 U5626 ( .A1(n4816), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4815) );
  NAND2_X1 U5627 ( .A1(n8375), .A2(n4816), .ZN(n4814) );
  INV_X1 U5628 ( .A(n8377), .ZN(n4816) );
  NOR2_X1 U5629 ( .A1(n8352), .A2(n8892), .ZN(n8374) );
  AOI21_X1 U5630 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8397), .A(n8396), .ZN(
        n8405) );
  OR2_X1 U5631 ( .A1(n9878), .A2(n9877), .ZN(n9875) );
  AOI21_X1 U5632 ( .B1(n8453), .B2(n8033), .A(n8233), .ZN(n5620) );
  NAND2_X1 U5633 ( .A1(n8473), .A2(n8472), .ZN(n4772) );
  NAND2_X1 U5634 ( .A1(n5493), .A2(n5492), .ZN(n5521) );
  INV_X1 U5635 ( .A(n5494), .ZN(n5493) );
  OR2_X1 U5636 ( .A1(n5487), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5494) );
  NAND2_X1 U5637 ( .A1(n5041), .A2(n5040), .ZN(n5485) );
  INV_X1 U5638 ( .A(n5475), .ZN(n5041) );
  NAND2_X1 U5639 ( .A1(n5039), .A2(n8977), .ZN(n5460) );
  INV_X1 U5640 ( .A(n5450), .ZN(n5039) );
  NAND2_X1 U5641 ( .A1(n5038), .A2(n5037), .ZN(n5430) );
  INV_X1 U5642 ( .A(n5415), .ZN(n5038) );
  NAND2_X1 U5643 ( .A1(n5036), .A2(n5035), .ZN(n5403) );
  INV_X1 U5644 ( .A(n5389), .ZN(n5036) );
  NAND2_X1 U5645 ( .A1(n5034), .A2(n5033), .ZN(n5373) );
  INV_X1 U5646 ( .A(n5355), .ZN(n5034) );
  INV_X1 U5647 ( .A(n8152), .ZN(n5606) );
  NAND2_X1 U5648 ( .A1(n4437), .A2(n5606), .ZN(n7100) );
  AND4_X1 U5649 ( .A1(n5333), .A2(n5332), .A3(n5331), .A4(n5330), .ZN(n7124)
         );
  NAND2_X1 U5650 ( .A1(n4793), .A2(n4792), .ZN(n7051) );
  AND2_X1 U5651 ( .A1(n5022), .A2(n5305), .ZN(n4792) );
  AND2_X1 U5652 ( .A1(n8139), .A2(n8136), .ZN(n8044) );
  NAND2_X1 U5653 ( .A1(n4793), .A2(n5305), .ZN(n6944) );
  NAND2_X1 U5654 ( .A1(n6819), .A2(n8122), .ZN(n6902) );
  NAND2_X1 U5655 ( .A1(n5029), .A2(n5028), .ZN(n5278) );
  INV_X1 U5656 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5028) );
  INV_X1 U5657 ( .A(n5266), .ZN(n5029) );
  AND3_X1 U5658 ( .A1(n5242), .A2(n5241), .A3(n5240), .ZN(n6573) );
  OAI21_X1 U5659 ( .B1(n6544), .B2(n5230), .A(n5229), .ZN(n6678) );
  AND4_X1 U5660 ( .A1(n5236), .A2(n5235), .A3(n5234), .A4(n5233), .ZN(n6575)
         );
  AND2_X1 U5661 ( .A1(n5671), .A2(n5670), .ZN(n6164) );
  NAND2_X1 U5662 ( .A1(n8224), .A2(n8225), .ZN(n8472) );
  NAND2_X1 U5663 ( .A1(n4572), .A2(n5508), .ZN(n5618) );
  NAND2_X1 U5664 ( .A1(n7598), .A2(n8060), .ZN(n4572) );
  NOR2_X1 U5665 ( .A1(n4455), .A2(n4766), .ZN(n4765) );
  NAND2_X1 U5666 ( .A1(n4768), .A2(n4770), .ZN(n4764) );
  INV_X1 U5667 ( .A(n4771), .ZN(n4766) );
  NAND2_X1 U5668 ( .A1(n5466), .A2(n7946), .ZN(n5467) );
  NAND2_X1 U5669 ( .A1(n5439), .A2(n5438), .ZN(n8547) );
  AND2_X1 U5670 ( .A1(n8158), .A2(n8155), .ZN(n8047) );
  NOR2_X1 U5671 ( .A1(n10230), .A2(n10255), .ZN(n10294) );
  OAI22_X1 U5672 ( .A1(n5894), .A2(n4817), .B1(P2_IR_REG_2__SCAN_IN), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U5673 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4817) );
  NAND2_X1 U5674 ( .A1(n4919), .A2(n4921), .ZN(n4918) );
  AOI21_X1 U5675 ( .B1(n6628), .B2(n6500), .A(n6629), .ZN(n6503) );
  INV_X1 U5676 ( .A(n9030), .ZN(n4917) );
  INV_X1 U5677 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6801) );
  NOR2_X1 U5678 ( .A1(n6123), .A2(n6425), .ZN(n6264) );
  NAND2_X1 U5679 ( .A1(n7588), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6205) );
  INV_X1 U5680 ( .A(n6758), .ZN(n4515) );
  NAND2_X1 U5681 ( .A1(n4649), .A2(n4650), .ZN(n9293) );
  AOI21_X1 U5682 ( .B1(n4651), .B2(n4659), .A(n4500), .ZN(n4650) );
  OR2_X1 U5683 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  INV_X1 U5684 ( .A(n4863), .ZN(n4862) );
  AND2_X1 U5685 ( .A1(n4648), .A2(n6079), .ZN(n4644) );
  NAND2_X1 U5686 ( .A1(n4647), .A2(n4646), .ZN(n4645) );
  INV_X1 U5687 ( .A(n6079), .ZN(n4646) );
  INV_X1 U5688 ( .A(n4648), .ZN(n4647) );
  AOI21_X1 U5689 ( .B1(n4664), .B2(n4663), .A(n9270), .ZN(n4662) );
  INV_X1 U5690 ( .A(n9079), .ZN(n4663) );
  NAND2_X1 U5691 ( .A1(n6417), .A2(n5015), .ZN(n6627) );
  NAND2_X1 U5692 ( .A1(n7760), .A2(n4451), .ZN(n4966) );
  AND4_X1 U5693 ( .A1(n7411), .A2(n7410), .A3(n7409), .A4(n7408), .ZN(n9212)
         );
  AND2_X1 U5694 ( .A1(n7580), .A2(n7579), .ZN(n9180) );
  AND2_X1 U5695 ( .A1(n7553), .A2(n7552), .ZN(n9227) );
  AND3_X1 U5696 ( .A1(n7537), .A2(n7536), .A3(n7535), .ZN(n9341) );
  INV_X1 U5697 ( .A(n7534), .ZN(n7594) );
  AND4_X1 U5698 ( .A1(n7085), .A2(n7084), .A3(n7083), .A4(n7082), .ZN(n9057)
         );
  AND4_X1 U5699 ( .A1(n6931), .A2(n6930), .A3(n6929), .A4(n6928), .ZN(n9050)
         );
  AND4_X1 U5700 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n9038)
         );
  INV_X1 U5701 ( .A(n7440), .ZN(n7616) );
  AND4_X1 U5702 ( .A1(n6460), .A2(n6459), .A3(n6458), .A4(n6457), .ZN(n6763)
         );
  AND4_X1 U5703 ( .A1(n6312), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n6504)
         );
  AND4_X1 U5704 ( .A1(n6270), .A2(n6269), .A3(n6268), .A4(n6267), .ZN(n6510)
         );
  NOR2_X1 U5705 ( .A1(n9208), .A2(n9350), .ZN(n4831) );
  INV_X1 U5706 ( .A(n7827), .ZN(n4633) );
  NAND2_X1 U5707 ( .A1(n9537), .A2(n4834), .ZN(n7826) );
  AND2_X1 U5708 ( .A1(n9523), .A2(n9522), .ZN(n4834) );
  INV_X1 U5709 ( .A(n9283), .ZN(n9556) );
  INV_X1 U5710 ( .A(n4605), .ZN(n9573) );
  NAND2_X1 U5711 ( .A1(n4612), .A2(n4610), .ZN(n9589) );
  AOI21_X1 U5712 ( .B1(n4614), .B2(n4616), .A(n4611), .ZN(n4610) );
  INV_X1 U5713 ( .A(n7818), .ZN(n4611) );
  AND2_X1 U5714 ( .A1(n4620), .A2(n4615), .ZN(n4614) );
  AND2_X1 U5715 ( .A1(n9604), .A2(n9606), .ZN(n4620) );
  NAND2_X1 U5716 ( .A1(n9639), .A2(n4617), .ZN(n4615) );
  OR2_X1 U5717 ( .A1(n9635), .A2(n4616), .ZN(n4613) );
  NAND2_X1 U5718 ( .A1(n4619), .A2(n4617), .ZN(n9605) );
  AND2_X1 U5719 ( .A1(n4619), .A2(n7695), .ZN(n9620) );
  OR2_X1 U5720 ( .A1(n7532), .A2(n6015), .ZN(n7546) );
  NAND2_X1 U5721 ( .A1(n9657), .A2(n7732), .ZN(n9635) );
  NAND2_X1 U5722 ( .A1(n4819), .A2(n4696), .ZN(n9676) );
  NOR2_X1 U5723 ( .A1(n7218), .A2(n7217), .ZN(n7516) );
  NAND2_X1 U5724 ( .A1(n7080), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7151) );
  OR2_X1 U5725 ( .A1(n7151), .A2(n7150), .ZN(n7218) );
  NAND2_X1 U5726 ( .A1(n7091), .A2(n9042), .ZN(n4876) );
  AND2_X1 U5727 ( .A1(n7637), .A2(n4609), .ZN(n4606) );
  NAND2_X1 U5728 ( .A1(n7654), .A2(n7655), .ZN(n4609) );
  NAND2_X1 U5729 ( .A1(n6919), .A2(n4589), .ZN(n7162) );
  NAND2_X1 U5730 ( .A1(n6919), .A2(n7091), .ZN(n7093) );
  NAND2_X1 U5731 ( .A1(n6793), .A2(n6792), .ZN(n6917) );
  NAND2_X1 U5732 ( .A1(n9929), .A2(n6707), .ZN(n6792) );
  NAND2_X1 U5733 ( .A1(n4608), .A2(n7478), .ZN(n7079) );
  NAND2_X1 U5734 ( .A1(n6703), .A2(n7650), .ZN(n7653) );
  NAND2_X1 U5735 ( .A1(n6526), .A2(n4590), .ZN(n6812) );
  AND2_X1 U5736 ( .A1(n9929), .A2(n4425), .ZN(n4590) );
  NAND2_X1 U5737 ( .A1(n6526), .A2(n4425), .ZN(n6726) );
  OR2_X1 U5738 ( .A1(n9391), .A2(n6757), .ZN(n6609) );
  NAND2_X1 U5739 ( .A1(n6526), .A2(n4592), .ZN(n6614) );
  AND2_X1 U5740 ( .A1(n6526), .A2(n10087), .ZN(n6527) );
  OAI21_X1 U5741 ( .B1(n9393), .B2(n6498), .A(n6464), .ZN(n6525) );
  OAI21_X1 U5742 ( .B1(n6300), .B2(n7465), .A(n7648), .ZN(n6697) );
  NAND2_X1 U5743 ( .A1(n7458), .A2(n7463), .ZN(n6300) );
  NAND2_X1 U5744 ( .A1(n4867), .A2(n6275), .ZN(n4866) );
  NOR2_X1 U5745 ( .A1(n4869), .A2(n4868), .ZN(n4867) );
  OR2_X1 U5746 ( .A1(n6259), .A2(n6428), .ZN(n6316) );
  NAND2_X1 U5747 ( .A1(n6275), .A2(n5014), .ZN(n6235) );
  NAND2_X1 U5748 ( .A1(n6235), .A2(n7703), .ZN(n6251) );
  NOR2_X1 U5749 ( .A1(n6288), .A2(n6669), .ZN(n6277) );
  NOR2_X1 U5750 ( .A1(n9664), .A2(n5757), .ZN(n6094) );
  NOR2_X1 U5751 ( .A1(n9505), .A2(n9208), .ZN(n4880) );
  OR2_X1 U5752 ( .A1(n7613), .A2(n9869), .ZN(n4928) );
  NAND2_X1 U5753 ( .A1(n7848), .A2(n7612), .ZN(n4929) );
  AND2_X1 U5754 ( .A1(n4883), .A2(n7812), .ZN(n4882) );
  NAND2_X1 U5755 ( .A1(n9510), .A2(n4884), .ZN(n4883) );
  INV_X1 U5756 ( .A(n7810), .ZN(n4884) );
  NAND2_X1 U5757 ( .A1(n7545), .A2(n7544), .ZN(n9627) );
  INV_X1 U5758 ( .A(n10094), .ZN(n9767) );
  AND2_X1 U5759 ( .A1(n5906), .A2(n9856), .ZN(n6322) );
  NAND2_X1 U5760 ( .A1(n5744), .A2(n4927), .ZN(n4926) );
  INV_X1 U5761 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5742) );
  XNOR2_X1 U5762 ( .A(n7382), .B(n7381), .ZN(n7412) );
  NAND2_X1 U5763 ( .A1(n4952), .A2(n5572), .ZN(n7382) );
  INV_X1 U5764 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U5765 ( .A(n5550), .B(n5549), .ZN(n7424) );
  NOR2_X1 U5766 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NOR2_X1 U5767 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5699) );
  INV_X1 U5768 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5700) );
  INV_X1 U5769 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5710) );
  INV_X1 U5770 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U5771 ( .A1(n4933), .A2(n4934), .ZN(n5470) );
  OR2_X1 U5772 ( .A1(n5441), .A2(n4936), .ZN(n4933) );
  INV_X1 U5773 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U5774 ( .A1(n5065), .A2(n5064), .ZN(n4595) );
  XNOR2_X1 U5775 ( .A(n5062), .B(SI_1_), .ZN(n5163) );
  NOR2_X1 U5776 ( .A1(n10351), .A2(n7017), .ZN(n7018) );
  NOR2_X1 U5777 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10350), .ZN(n7017) );
  XNOR2_X1 U5778 ( .A(n5653), .B(n5652), .ZN(n5880) );
  AND4_X1 U5779 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n6959)
         );
  NAND2_X1 U5780 ( .A1(n4737), .A2(n4738), .ZN(n6743) );
  AND2_X1 U5781 ( .A1(n5559), .A2(n5558), .ZN(n7912) );
  OR2_X1 U5782 ( .A1(n7987), .A2(n4723), .ZN(n4717) );
  NAND2_X1 U5783 ( .A1(n7130), .A2(n7129), .ZN(n7283) );
  AND4_X1 U5784 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n8565)
         );
  NAND2_X1 U5785 ( .A1(n7130), .A2(n4734), .ZN(n7192) );
  INV_X1 U5786 ( .A(n8275), .ZN(n8148) );
  NAND2_X1 U5787 ( .A1(n6589), .A2(n6577), .ZN(n6741) );
  NAND2_X1 U5788 ( .A1(n6590), .A2(n6591), .ZN(n6589) );
  NAND2_X1 U5789 ( .A1(n6144), .A2(n6062), .ZN(n8020) );
  OAI21_X1 U5790 ( .B1(n7130), .B2(n4733), .A(n4731), .ZN(n7298) );
  NOR2_X1 U5791 ( .A1(n4732), .A2(n4461), .ZN(n4731) );
  NOR2_X1 U5792 ( .A1(n4734), .A2(n4733), .ZN(n4732) );
  INV_X1 U5793 ( .A(n7972), .ZN(n8016) );
  XNOR2_X1 U5794 ( .A(n5584), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8264) );
  INV_X1 U5795 ( .A(n8486), .ZN(n8272) );
  INV_X1 U5796 ( .A(n8511), .ZN(n8273) );
  INV_X1 U5797 ( .A(n6959), .ZN(n8279) );
  INV_X1 U5798 ( .A(n6824), .ZN(n8281) );
  INV_X1 U5799 ( .A(n6575), .ZN(n8282) );
  OR2_X1 U5800 ( .A1(n5879), .A2(n5855), .ZN(n8285) );
  NOR2_X1 U5801 ( .A1(n5875), .A2(n5874), .ZN(n6355) );
  NAND2_X1 U5802 ( .A1(n4795), .A2(n4794), .ZN(n10133) );
  NAND2_X1 U5803 ( .A1(n6366), .A2(n6376), .ZN(n4794) );
  NOR2_X1 U5804 ( .A1(n6378), .A2(n4859), .ZN(n10138) );
  NOR2_X1 U5805 ( .A1(n6360), .A2(n6361), .ZN(n6649) );
  INV_X1 U5806 ( .A(n6859), .ZN(n4797) );
  NOR2_X1 U5807 ( .A1(n10148), .A2(n10309), .ZN(n4799) );
  NOR2_X1 U5808 ( .A1(n6844), .A2(n6845), .ZN(n6981) );
  OAI21_X1 U5809 ( .B1(n6861), .B2(n4810), .A(n4809), .ZN(n10162) );
  NAND2_X1 U5810 ( .A1(n4813), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4810) );
  NAND2_X1 U5811 ( .A1(n6998), .A2(n4813), .ZN(n4809) );
  INV_X1 U5812 ( .A(n10163), .ZN(n4813) );
  INV_X1 U5813 ( .A(n6998), .ZN(n4811) );
  XNOR2_X1 U5814 ( .A(n7305), .B(n9021), .ZN(n6983) );
  NOR2_X1 U5815 ( .A1(n6983), .A2(n6984), .ZN(n7306) );
  OR2_X1 U5816 ( .A1(n7000), .A2(n10317), .ZN(n4808) );
  NAND2_X1 U5817 ( .A1(n4803), .A2(n4805), .ZN(n10180) );
  AND2_X1 U5818 ( .A1(n5885), .A2(n5884), .ZN(n10185) );
  INV_X1 U5819 ( .A(n4838), .ZN(n7313) );
  NOR2_X1 U5820 ( .A1(n8311), .A2(n8312), .ZN(n8315) );
  INV_X1 U5821 ( .A(n8361), .ZN(n4845) );
  NAND2_X1 U5822 ( .A1(n8361), .A2(n4847), .ZN(n4843) );
  OR2_X1 U5823 ( .A1(n8340), .A2(n4844), .ZN(n4521) );
  NAND2_X1 U5824 ( .A1(n4847), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4844) );
  OAI21_X1 U5825 ( .B1(n4852), .B2(n4851), .A(n4443), .ZN(n9886) );
  OR2_X1 U5826 ( .A1(n8415), .A2(n8416), .ZN(n4852) );
  NAND2_X1 U5827 ( .A1(n5892), .A2(n5886), .ZN(n10199) );
  INV_X1 U5828 ( .A(n8434), .ZN(n4524) );
  NAND2_X1 U5829 ( .A1(n4520), .A2(n10167), .ZN(n4525) );
  XNOR2_X1 U5830 ( .A(n8429), .B(n8430), .ZN(n4520) );
  AOI21_X1 U5831 ( .B1(n9888), .B2(n9887), .A(n9890), .ZN(n8429) );
  NAND2_X1 U5832 ( .A1(n7863), .A2(n4512), .ZN(n8444) );
  AND2_X1 U5833 ( .A1(n4743), .A2(n4513), .ZN(n4512) );
  OR2_X1 U5834 ( .A1(n4745), .A2(n8454), .ZN(n4513) );
  INV_X1 U5835 ( .A(n8058), .ZN(n5583) );
  AND2_X1 U5836 ( .A1(n4781), .A2(n4448), .ZN(n8534) );
  NAND2_X1 U5837 ( .A1(n5459), .A2(n5458), .ZN(n8632) );
  NAND2_X1 U5838 ( .A1(n5449), .A2(n5448), .ZN(n8556) );
  NAND2_X1 U5839 ( .A1(n5341), .A2(n5340), .ZN(n10298) );
  NAND2_X1 U5840 ( .A1(n4983), .A2(n8136), .ZN(n7049) );
  NAND2_X1 U5841 ( .A1(n6942), .A2(n8129), .ZN(n4983) );
  NAND2_X1 U5842 ( .A1(n5327), .A2(n5326), .ZN(n10292) );
  AND3_X1 U5843 ( .A1(n5262), .A2(n5261), .A3(n5260), .ZN(n6690) );
  NAND2_X1 U5844 ( .A1(n6171), .A2(n7262), .ZN(n8516) );
  AND2_X1 U5845 ( .A1(n8601), .A2(n6543), .ZN(n10213) );
  NAND2_X1 U5846 ( .A1(n10227), .A2(n5199), .ZN(n10201) );
  NAND2_X1 U5847 ( .A1(n6059), .A2(n6058), .ZN(n10217) );
  AND3_X2 U5848 ( .A1(n5169), .A2(n5168), .A3(n5167), .ZN(n6211) );
  NAND2_X1 U5849 ( .A1(n5181), .A2(n4742), .ZN(n5168) );
  AND2_X1 U5850 ( .A1(n6940), .A2(n6939), .ZN(n10299) );
  INV_X1 U5851 ( .A(n10217), .ZN(n10211) );
  AND2_X1 U5852 ( .A1(n8027), .A2(n8026), .ZN(n8652) );
  AND2_X1 U5853 ( .A1(n8063), .A2(n8062), .ZN(n8655) );
  NAND2_X1 U5854 ( .A1(n7850), .A2(n7849), .ZN(n8445) );
  NAND2_X1 U5855 ( .A1(n5519), .A2(n5518), .ZN(n8667) );
  INV_X1 U5856 ( .A(n5618), .ZN(n8672) );
  NAND2_X1 U5857 ( .A1(n4992), .A2(n4990), .ZN(n8490) );
  AND2_X1 U5858 ( .A1(n5158), .A2(n5157), .ZN(n8677) );
  NAND2_X1 U5859 ( .A1(n4767), .A2(n4771), .ZN(n8497) );
  NAND2_X1 U5860 ( .A1(n4769), .A2(n4768), .ZN(n4767) );
  NAND2_X1 U5861 ( .A1(n4992), .A2(n5617), .ZN(n8496) );
  AND2_X1 U5862 ( .A1(n5484), .A2(n5483), .ZN(n8684) );
  NAND2_X1 U5863 ( .A1(n8561), .A2(n8186), .ZN(n8545) );
  NAND2_X1 U5864 ( .A1(n5414), .A2(n5413), .ZN(n8706) );
  OAI21_X1 U5865 ( .B1(n8586), .B2(n8585), .A(n4759), .ZN(n8577) );
  INV_X1 U5866 ( .A(n4761), .ZN(n4759) );
  NAND2_X1 U5867 ( .A1(n4986), .A2(n8177), .ZN(n8575) );
  NAND2_X1 U5868 ( .A1(n5402), .A2(n5401), .ZN(n8712) );
  NAND2_X1 U5869 ( .A1(n5388), .A2(n5387), .ZN(n8718) );
  NAND2_X1 U5870 ( .A1(n7256), .A2(n5381), .ZN(n8597) );
  NAND2_X1 U5871 ( .A1(n5372), .A2(n5371), .ZN(n7274) );
  AND2_X1 U5872 ( .A1(n7260), .A2(n7259), .ZN(n7272) );
  NAND2_X1 U5873 ( .A1(n5354), .A2(n5353), .ZN(n8154) );
  INV_X1 U5874 ( .A(n7187), .ZN(n5857) );
  AND2_X1 U5875 ( .A1(n5880), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5853) );
  NAND2_X1 U5876 ( .A1(n5850), .A2(n6059), .ZN(n5862) );
  INV_X1 U5877 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8725) );
  NOR2_X1 U5878 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4984) );
  INV_X1 U5879 ( .A(n5596), .ZN(n7294) );
  NAND2_X1 U5880 ( .A1(n5634), .A2(n5633), .ZN(n7280) );
  INV_X1 U5881 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8865) );
  OR2_X1 U5882 ( .A1(n5628), .A2(n5627), .ZN(n5629) );
  INV_X1 U5883 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n6941) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6869) );
  XNOR2_X1 U5885 ( .A(n5589), .B(n5588), .ZN(n8260) );
  XNOR2_X1 U5886 ( .A(n5446), .B(n5445), .ZN(n8431) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n8967) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8800) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5867) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5849) );
  INV_X1 U5891 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5831) );
  INV_X1 U5892 ( .A(n6860), .ZN(n10155) );
  INV_X1 U5893 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n5818) );
  INV_X1 U5894 ( .A(n4671), .ZN(n6751) );
  NAND2_X1 U5895 ( .A1(n4920), .A2(n4918), .ZN(n6509) );
  AND2_X1 U5896 ( .A1(n4914), .A2(n4915), .ZN(n9921) );
  NAND2_X1 U5897 ( .A1(n4653), .A2(n4657), .ZN(n9196) );
  NAND2_X1 U5898 ( .A1(n4655), .A2(n4654), .ZN(n4653) );
  INV_X1 U5899 ( .A(n9257), .ZN(n4655) );
  INV_X1 U5900 ( .A(n4909), .ZN(n4908) );
  AOI21_X1 U5901 ( .B1(n4423), .B2(n4912), .A(n4474), .ZN(n4909) );
  AND2_X1 U5902 ( .A1(n9153), .A2(n9152), .ZN(n9217) );
  NOR2_X1 U5903 ( .A1(n5937), .A2(n5011), .ZN(n5990) );
  INV_X1 U5904 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U5905 ( .A1(n6122), .A2(n6121), .ZN(n6417) );
  NAND2_X1 U5906 ( .A1(n4871), .A2(n9049), .ZN(n9304) );
  NAND2_X1 U5907 ( .A1(n9234), .A2(n9235), .ZN(n4871) );
  NAND2_X1 U5908 ( .A1(n9117), .A2(n9189), .ZN(n9313) );
  NAND2_X1 U5909 ( .A1(n4643), .A2(n4645), .ZN(n6080) );
  INV_X1 U5910 ( .A(n4644), .ZN(n4643) );
  NAND2_X1 U5911 ( .A1(n4656), .A2(n4661), .ZN(n9339) );
  NAND2_X1 U5912 ( .A1(n9256), .A2(n4662), .ZN(n4656) );
  NAND2_X1 U5913 ( .A1(n7524), .A2(n7523), .ZN(n9766) );
  NAND2_X1 U5914 ( .A1(n9244), .A2(n4667), .ZN(n4666) );
  INV_X1 U5915 ( .A(n9348), .ZN(n4667) );
  NOR2_X2 U5916 ( .A1(n5925), .A2(n5924), .ZN(n9931) );
  INV_X1 U5917 ( .A(n9928), .ZN(n9368) );
  INV_X1 U5918 ( .A(n9931), .ZN(n9370) );
  INV_X1 U5919 ( .A(n9227), .ZN(n9380) );
  INV_X1 U5920 ( .A(n9042), .ZN(n9387) );
  OR2_X1 U5921 ( .A1(n7534), .A2(n6399), .ZN(n4681) );
  INV_X1 U5922 ( .A(P1_U3973), .ZN(n9398) );
  AND3_X1 U5923 ( .A1(n5724), .A2(n5723), .A3(n5722), .ZN(n5728) );
  OR2_X1 U5924 ( .A1(n5836), .A2(n5726), .ZN(n5727) );
  NOR2_X1 U5925 ( .A1(n9481), .A2(n9664), .ZN(n9714) );
  NAND2_X1 U5926 ( .A1(n4579), .A2(n9480), .ZN(n4578) );
  NAND2_X1 U5927 ( .A1(n4621), .A2(n4829), .ZN(n7843) );
  NOR2_X1 U5928 ( .A1(n4831), .A2(n4830), .ZN(n4829) );
  NAND2_X1 U5929 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  NOR2_X1 U5930 ( .A1(n7831), .A2(n9482), .ZN(n4830) );
  AND2_X1 U5931 ( .A1(n9541), .A2(n9540), .ZN(n9733) );
  NAND2_X1 U5932 ( .A1(n7585), .A2(n7584), .ZN(n9742) );
  NAND2_X1 U5933 ( .A1(n7572), .A2(n7571), .ZN(n9600) );
  NAND2_X1 U5934 ( .A1(n7529), .A2(n7528), .ZN(n9648) );
  NAND2_X1 U5935 ( .A1(n7730), .A2(n7729), .ZN(n9695) );
  INV_X1 U5936 ( .A(n10065), .ZN(n10042) );
  NAND2_X1 U5937 ( .A1(n10067), .A2(n6332), .ZN(n10062) );
  OR2_X1 U5938 ( .A1(n6331), .A2(n4418), .ZN(n10049) );
  INV_X1 U5939 ( .A(n9701), .ZN(n10053) );
  INV_X1 U5940 ( .A(n10049), .ZN(n9665) );
  NAND2_X1 U5941 ( .A1(n6291), .A2(n6241), .ZN(n6278) );
  OAI21_X1 U5942 ( .B1(n4593), .B2(n4431), .A(n6253), .ZN(n4594) );
  INV_X1 U5943 ( .A(n10062), .ZN(n10047) );
  AND2_X1 U5944 ( .A1(n9853), .A2(n6094), .ZN(n10065) );
  AND2_X1 U5945 ( .A1(n5993), .A2(n5020), .ZN(n5994) );
  OAI21_X1 U5946 ( .B1(n9521), .B2(n7811), .A(n7810), .ZN(n9509) );
  NAND2_X1 U5947 ( .A1(n7437), .A2(n7436), .ZN(n9808) );
  NAND2_X1 U5948 ( .A1(n7601), .A2(n7600), .ZN(n9813) );
  NAND2_X1 U5949 ( .A1(n4898), .A2(n4902), .ZN(n9571) );
  NAND2_X1 U5950 ( .A1(n4509), .A2(n4904), .ZN(n4898) );
  NAND2_X1 U5951 ( .A1(n4906), .A2(n4424), .ZN(n9593) );
  NAND2_X1 U5952 ( .A1(n4907), .A2(n4481), .ZN(n4906) );
  INV_X1 U5953 ( .A(n4509), .ZN(n4907) );
  INV_X1 U5954 ( .A(n9627), .ZN(n9828) );
  NAND2_X1 U5955 ( .A1(n4886), .A2(n4890), .ZN(n9652) );
  NAND2_X1 U5956 ( .A1(n4893), .A2(n4891), .ZN(n4886) );
  NAND2_X1 U5957 ( .A1(n7515), .A2(n7514), .ZN(n9840) );
  NAND2_X1 U5958 ( .A1(n4892), .A2(n4896), .ZN(n9672) );
  NAND2_X1 U5959 ( .A1(n4893), .A2(n4600), .ZN(n4892) );
  NAND2_X1 U5960 ( .A1(n7499), .A2(n7498), .ZN(n9846) );
  NAND2_X1 U5961 ( .A1(n7076), .A2(n7075), .ZN(n9309) );
  NAND2_X1 U5962 ( .A1(n6796), .A2(n6795), .ZN(n9333) );
  INV_X1 U5963 ( .A(n9852), .ZN(n9847) );
  AND2_X1 U5964 ( .A1(n6255), .A2(n6254), .ZN(n6488) );
  AND3_X1 U5965 ( .A1(n6119), .A2(n6118), .A3(n6117), .ZN(n6260) );
  AND3_X1 U5966 ( .A1(n6072), .A2(n6071), .A3(n6070), .ZN(n6342) );
  INV_X1 U5967 ( .A(n7848), .ZN(n9871) );
  XNOR2_X1 U5968 ( .A(n5705), .B(n4927), .ZN(n7255) );
  INV_X1 U5969 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U5970 ( .A(n5502), .B(n5501), .ZN(n7583) );
  INV_X1 U5971 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7781) );
  INV_X1 U5972 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8932) );
  INV_X1 U5973 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7543) );
  INV_X1 U5974 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6180) );
  INV_X1 U5975 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5865) );
  INV_X1 U5976 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8980) );
  OAI21_X1 U5977 ( .B1(n5287), .B2(n5286), .A(n5096), .ZN(n5299) );
  INV_X1 U5978 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8825) );
  OR3_X1 U5979 ( .A1(n5844), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .ZN(n5845) );
  INV_X1 U5980 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5823) );
  INV_X1 U5981 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6116) );
  INV_X1 U5982 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5991) );
  NOR2_X1 U5983 ( .A1(n7039), .A2(n7038), .ZN(n10339) );
  NOR2_X1 U5984 ( .A1(n10341), .A2(n10340), .ZN(n7038) );
  INV_X1 U5985 ( .A(n8285), .ZN(P2_U3893) );
  AND2_X1 U5986 ( .A1(n4714), .A2(n6479), .ZN(n4713) );
  INV_X1 U5987 ( .A(n4846), .ZN(n8360) );
  AND2_X1 U5988 ( .A1(n5683), .A2(n5682), .ZN(n5024) );
  MUX2_X1 U5989 ( .A(n8616), .B(n8662), .S(n10325), .Z(n8617) );
  MUX2_X1 U5990 ( .A(n8663), .B(n8662), .S(n10300), .Z(n8664) );
  NAND2_X1 U5991 ( .A1(n4963), .A2(n7767), .ZN(P1_U3242) );
  NAND2_X1 U5992 ( .A1(n4964), .A2(n5773), .ZN(n4963) );
  OAI21_X1 U5993 ( .B1(n4827), .B2(n4826), .A(n4825), .ZN(n7834) );
  OR2_X1 U5994 ( .A1(n10106), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4825) );
  NAND2_X1 U5995 ( .A1(n4827), .A2(n10100), .ZN(n4637) );
  OR2_X1 U5996 ( .A1(n8248), .A2(n8247), .ZN(n4419) );
  NAND2_X1 U5997 ( .A1(n4934), .A2(n4487), .ZN(n4932) );
  OR2_X1 U5998 ( .A1(n9508), .A2(n7811), .ZN(n4420) );
  AND2_X1 U5999 ( .A1(n4851), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4421) );
  AND2_X1 U6000 ( .A1(n4441), .A2(n4545), .ZN(n4422) );
  AND2_X1 U6001 ( .A1(n9144), .A2(n4910), .ZN(n4423) );
  NAND2_X1 U6002 ( .A1(n4929), .A2(n4928), .ZN(n7814) );
  OR2_X1 U6003 ( .A1(n9614), .A2(n9316), .ZN(n4424) );
  AND2_X1 U6004 ( .A1(n4592), .A2(n4591), .ZN(n4425) );
  AND2_X1 U6005 ( .A1(n4882), .A2(n4483), .ZN(n4426) );
  INV_X1 U6006 ( .A(n9510), .ZN(n9508) );
  OR2_X1 U6007 ( .A1(n7511), .A2(n7510), .ZN(n4427) );
  AND2_X1 U6008 ( .A1(n4538), .A2(n8256), .ZN(n4428) );
  AND2_X1 U6009 ( .A1(n4473), .A2(n8256), .ZN(n4429) );
  OR2_X1 U6010 ( .A1(n5587), .A2(n4997), .ZN(n4430) );
  INV_X1 U6011 ( .A(n10148), .ZN(n4801) );
  NAND2_X1 U6012 ( .A1(n7213), .A2(n7212), .ZN(n9708) );
  AND2_X1 U6013 ( .A1(n5939), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4431) );
  AND2_X1 U6014 ( .A1(n4462), .A2(n7512), .ZN(n4432) );
  INV_X1 U6015 ( .A(n4659), .ZN(n4654) );
  NAND2_X1 U6016 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  NAND2_X1 U6017 ( .A1(n4624), .A2(n9697), .ZN(n4433) );
  AND2_X1 U6018 ( .A1(n4976), .A2(n5264), .ZN(n4434) );
  AND2_X1 U6019 ( .A1(n8219), .A2(n4989), .ZN(n4435) );
  INV_X1 U6020 ( .A(n4932), .ZN(n4931) );
  AND3_X1 U6021 ( .A1(n5479), .A2(n5478), .A3(n5477), .ZN(n8510) );
  OR2_X1 U6022 ( .A1(n9742), .A2(n9377), .ZN(n4436) );
  AND2_X1 U6023 ( .A1(n4978), .A2(n4981), .ZN(n4437) );
  NOR2_X1 U6024 ( .A1(n8233), .A2(n8234), .ZN(n4438) );
  NOR2_X1 U6025 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5788) );
  AND2_X1 U6026 ( .A1(n7987), .A2(n7889), .ZN(n4439) );
  NAND2_X1 U6027 ( .A1(n4862), .A2(n9189), .ZN(n9186) );
  OR2_X1 U6028 ( .A1(n5119), .A2(n5118), .ZN(n4440) );
  AND2_X1 U6029 ( .A1(n4930), .A2(n4548), .ZN(n4441) );
  NAND2_X1 U6030 ( .A1(n6655), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4442) );
  AND2_X1 U6031 ( .A1(n4848), .A2(n4850), .ZN(n4443) );
  NOR2_X1 U6032 ( .A1(n5335), .A2(n8134), .ZN(n4444) );
  AND2_X1 U6033 ( .A1(n5045), .A2(n5209), .ZN(n5284) );
  NAND2_X1 U6034 ( .A1(n6841), .A2(n6847), .ZN(n4445) );
  AOI21_X1 U6035 ( .B1(n9257), .B2(n9079), .A(n9078), .ZN(n9269) );
  NAND2_X1 U6036 ( .A1(n4772), .A2(n5529), .ZN(n8461) );
  INV_X1 U6037 ( .A(n8114), .ZN(n4973) );
  INV_X1 U6038 ( .A(n7467), .ZN(n4685) );
  INV_X1 U6039 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5730) );
  OR2_X1 U6040 ( .A1(n8250), .A2(n8256), .ZN(n4446) );
  NAND2_X1 U6041 ( .A1(n5582), .A2(n5581), .ZN(n8455) );
  OR2_X1 U6042 ( .A1(n5587), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n4447) );
  NAND2_X1 U6043 ( .A1(n6915), .A2(n6914), .ZN(n9241) );
  NAND2_X1 U6044 ( .A1(n8556), .A2(n8535), .ZN(n4448) );
  AND3_X1 U6045 ( .A1(n5627), .A2(n5652), .A3(n5625), .ZN(n4449) );
  INV_X1 U6046 ( .A(n7829), .ZN(n9493) );
  AND2_X1 U6047 ( .A1(n4631), .A2(n7830), .ZN(n4450) );
  INV_X1 U6048 ( .A(n8463), .ZN(n8271) );
  AND2_X1 U6049 ( .A1(n5567), .A2(n5566), .ZN(n8463) );
  OR2_X1 U6050 ( .A1(n7725), .A2(n7684), .ZN(n4451) );
  AND2_X1 U6051 ( .A1(n9511), .A2(n4450), .ZN(n4452) );
  AND2_X1 U6052 ( .A1(n7463), .A2(n4677), .ZN(n4453) );
  NOR2_X1 U6053 ( .A1(n8374), .A2(n8375), .ZN(n4454) );
  INV_X1 U6054 ( .A(n8501), .ZN(n8474) );
  AND2_X1 U6055 ( .A1(n5500), .A2(n5499), .ZN(n8501) );
  AND2_X1 U6056 ( .A1(n8677), .A2(n8511), .ZN(n4455) );
  OR2_X1 U6057 ( .A1(n7661), .A2(n7506), .ZN(n4456) );
  AND2_X1 U6058 ( .A1(n5490), .A2(n8500), .ZN(n8206) );
  INV_X1 U6059 ( .A(n6648), .ZN(n6847) );
  INV_X1 U6060 ( .A(n7706), .ZN(n6797) );
  AND2_X1 U6061 ( .A1(n6708), .A2(n7478), .ZN(n7706) );
  AND2_X1 U6062 ( .A1(n4846), .A2(n4845), .ZN(n4457) );
  INV_X1 U6063 ( .A(n7655), .ZN(n7478) );
  AND2_X1 U6064 ( .A1(n9034), .A2(n6707), .ZN(n7655) );
  INV_X1 U6065 ( .A(n4560), .ZN(n4559) );
  AOI21_X1 U6066 ( .B1(n5286), .B2(n5096), .A(n4561), .ZN(n4560) );
  INV_X1 U6067 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5718) );
  NOR2_X1 U6068 ( .A1(n4456), .A2(n4695), .ZN(n4458) );
  AND2_X1 U6069 ( .A1(n8706), .A2(n8588), .ZN(n4459) );
  NOR2_X1 U6070 ( .A1(n6824), .A2(n6740), .ZN(n4460) );
  INV_X1 U6071 ( .A(n4704), .ZN(n4703) );
  NAND2_X1 U6072 ( .A1(n4705), .A2(n7688), .ZN(n4704) );
  NAND2_X1 U6073 ( .A1(n7248), .A2(n7246), .ZN(n4461) );
  NOR2_X1 U6074 ( .A1(n7665), .A2(n7625), .ZN(n4462) );
  NOR2_X1 U6075 ( .A1(n4662), .A2(n9336), .ZN(n4463) );
  AND2_X1 U6076 ( .A1(n8125), .A2(n6901), .ZN(n8122) );
  INV_X1 U6077 ( .A(n8122), .ZN(n4976) );
  AND2_X1 U6078 ( .A1(n5141), .A2(n5140), .ZN(n4464) );
  OR2_X1 U6079 ( .A1(n6253), .A2(n5941), .ZN(n4465) );
  AND2_X1 U6080 ( .A1(n4563), .A2(n5126), .ZN(n4466) );
  NAND2_X1 U6081 ( .A1(n5049), .A2(n4787), .ZN(n4467) );
  AOI21_X1 U6082 ( .B1(n9288), .B2(n4423), .A(n4908), .ZN(n9211) );
  NAND2_X1 U6083 ( .A1(n7135), .A2(n7134), .ZN(n4468) );
  INV_X1 U6084 ( .A(n4587), .ZN(n4586) );
  NAND2_X1 U6085 ( .A1(n4589), .A2(n4588), .ZN(n4587) );
  INV_X1 U6086 ( .A(n4873), .ZN(n4872) );
  NAND2_X1 U6087 ( .A1(n4874), .A2(n9303), .ZN(n4873) );
  AND2_X1 U6088 ( .A1(n5122), .A2(SI_15_), .ZN(n4469) );
  AND2_X1 U6089 ( .A1(n5112), .A2(SI_12_), .ZN(n4470) );
  AND2_X1 U6090 ( .A1(n4613), .A2(n4614), .ZN(n4471) );
  AND2_X1 U6091 ( .A1(n4717), .A2(n4721), .ZN(n4472) );
  INV_X1 U6092 ( .A(n4632), .ZN(n4631) );
  OAI21_X1 U6093 ( .B1(n4633), .B2(n9508), .A(n9493), .ZN(n4632) );
  INV_X1 U6094 ( .A(n7853), .ZN(n4758) );
  INV_X1 U6095 ( .A(n9078), .ZN(n4664) );
  AND2_X1 U6096 ( .A1(n8677), .A2(n8273), .ZN(n8213) );
  AND2_X1 U6097 ( .A1(n4538), .A2(n8253), .ZN(n4473) );
  AND2_X1 U6098 ( .A1(n8655), .A2(n8270), .ZN(n8243) );
  OR2_X1 U6099 ( .A1(n9159), .A2(n9158), .ZN(n4474) );
  INV_X1 U6100 ( .A(n9673), .ZN(n4696) );
  OR2_X1 U6101 ( .A1(n5893), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4475) );
  AND2_X1 U6102 ( .A1(n4738), .A2(n4736), .ZN(n4476) );
  AND2_X1 U6103 ( .A1(n4706), .A2(n7455), .ZN(n4477) );
  INV_X1 U6104 ( .A(n9929), .ZN(n9034) );
  AND2_X1 U6105 ( .A1(n6706), .A2(n6705), .ZN(n9929) );
  AND2_X1 U6106 ( .A1(n4689), .A2(n4690), .ZN(n4478) );
  NAND2_X1 U6107 ( .A1(n4758), .A2(n4756), .ZN(n4479) );
  AND2_X1 U6108 ( .A1(n5529), .A2(n5023), .ZN(n4480) );
  INV_X1 U6109 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5864) );
  AND2_X1 U6110 ( .A1(n4657), .A2(n4652), .ZN(n4651) );
  INV_X1 U6111 ( .A(n4991), .ZN(n4990) );
  NAND2_X1 U6112 ( .A1(n8214), .A2(n5617), .ZN(n4991) );
  INV_X1 U6113 ( .A(n5491), .ZN(n4770) );
  AND2_X1 U6114 ( .A1(n8505), .A2(n8273), .ZN(n5491) );
  NAND2_X1 U6115 ( .A1(n7146), .A2(n7145), .ZN(n9172) );
  INV_X1 U6116 ( .A(n9172), .ZN(n4588) );
  OR2_X1 U6117 ( .A1(n9752), .A2(n9379), .ZN(n4481) );
  AND2_X1 U6118 ( .A1(n7697), .A2(n7731), .ZN(n9694) );
  INV_X1 U6119 ( .A(n9694), .ZN(n4600) );
  NAND2_X1 U6120 ( .A1(n9323), .A2(n9327), .ZN(n9234) );
  OR2_X1 U6121 ( .A1(n5125), .A2(n5124), .ZN(n4482) );
  INV_X1 U6122 ( .A(n6999), .ZN(n10171) );
  NAND2_X1 U6123 ( .A1(n4424), .A2(n4485), .ZN(n4905) );
  INV_X1 U6124 ( .A(n7333), .ZN(n10184) );
  INV_X1 U6125 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4927) );
  NAND2_X1 U6126 ( .A1(n7615), .A2(n7614), .ZN(n9487) );
  NAND2_X1 U6127 ( .A1(n5380), .A2(n5379), .ZN(n7256) );
  OR2_X1 U6128 ( .A1(n9719), .A2(n9374), .ZN(n4483) );
  NAND2_X1 U6129 ( .A1(n5472), .A2(n5471), .ZN(n8687) );
  INV_X1 U6130 ( .A(n4568), .ZN(n4567) );
  NOR2_X1 U6131 ( .A1(n5123), .A2(n4569), .ZN(n4568) );
  AND2_X1 U6132 ( .A1(n9742), .A2(n9377), .ZN(n4484) );
  OR2_X1 U6133 ( .A1(n9747), .A2(n9180), .ZN(n4485) );
  NAND2_X1 U6134 ( .A1(n8571), .A2(n8578), .ZN(n4486) );
  NAND2_X1 U6135 ( .A1(n5468), .A2(n5142), .ZN(n4487) );
  AND2_X1 U6136 ( .A1(n9114), .A2(n9111), .ZN(n4488) );
  AND2_X1 U6137 ( .A1(n9056), .A2(n9055), .ZN(n4489) );
  AND2_X1 U6138 ( .A1(n9241), .A2(n9387), .ZN(n4490) );
  INV_X1 U6139 ( .A(n4905), .ZN(n4904) );
  AND2_X1 U6140 ( .A1(n7402), .A2(n7401), .ZN(n9793) );
  AND2_X1 U6141 ( .A1(n9747), .A2(n9180), .ZN(n4491) );
  INV_X1 U6142 ( .A(n4897), .ZN(n4896) );
  NOR2_X1 U6143 ( .A1(n9783), .A2(n7802), .ZN(n4897) );
  INV_X1 U6144 ( .A(n4584), .ZN(n4583) );
  OR2_X1 U6145 ( .A1(n7814), .A2(n9719), .ZN(n4584) );
  AND2_X1 U6146 ( .A1(n5143), .A2(SI_21_), .ZN(n4492) );
  NAND2_X1 U6147 ( .A1(n7414), .A2(n7413), .ZN(n9719) );
  OR2_X1 U6148 ( .A1(n4895), .A2(n4897), .ZN(n4493) );
  INV_X1 U6149 ( .A(n7334), .ZN(n7368) );
  AND2_X1 U6150 ( .A1(n5325), .A2(n5351), .ZN(n7334) );
  OR2_X1 U6151 ( .A1(n7160), .A2(n9050), .ZN(n4494) );
  NAND2_X1 U6152 ( .A1(n4493), .A2(n4894), .ZN(n4890) );
  OR2_X1 U6153 ( .A1(n7333), .A2(n10319), .ZN(n4495) );
  XNOR2_X1 U6154 ( .A(n5626), .B(n5625), .ZN(n7187) );
  AND2_X1 U6155 ( .A1(n6919), .A2(n4586), .ZN(n4496) );
  INV_X1 U6156 ( .A(n8316), .ZN(n4511) );
  AND2_X1 U6157 ( .A1(n5649), .A2(n5851), .ZN(n4497) );
  INV_X1 U6158 ( .A(n7942), .ZN(n4723) );
  AND2_X1 U6159 ( .A1(n8351), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4498) );
  AND2_X1 U6160 ( .A1(n9084), .A2(n9083), .ZN(n4499) );
  AND2_X1 U6161 ( .A1(n9098), .A2(n9097), .ZN(n4500) );
  NAND2_X1 U6162 ( .A1(n5265), .A2(n5264), .ZN(n6821) );
  NAND2_X1 U6163 ( .A1(n5048), .A2(n5284), .ZN(n5399) );
  NOR2_X1 U6164 ( .A1(n6981), .A2(n6982), .ZN(n4501) );
  NOR2_X1 U6165 ( .A1(n7306), .A2(n7307), .ZN(n4502) );
  INV_X1 U6166 ( .A(n9336), .ZN(n4660) );
  AND2_X1 U6167 ( .A1(n7385), .A2(n7384), .ZN(n4503) );
  NOR2_X1 U6168 ( .A1(n6478), .A2(n4713), .ZN(n4504) );
  AND2_X1 U6169 ( .A1(n4808), .A2(n4807), .ZN(n4505) );
  INV_X1 U6170 ( .A(n10225), .ZN(n10207) );
  INV_X1 U6171 ( .A(n8076), .ZN(n6939) );
  INV_X1 U6172 ( .A(n10193), .ZN(n10167) );
  NAND2_X1 U6173 ( .A1(n6606), .A2(n6605), .ZN(n10091) );
  INV_X1 U6174 ( .A(n10091), .ZN(n4591) );
  AND2_X1 U6175 ( .A1(n6096), .A2(n7403), .ZN(n9578) );
  AND2_X1 U6176 ( .A1(n4812), .A2(n4811), .ZN(n4506) );
  AND2_X1 U6177 ( .A1(n4797), .A2(n6857), .ZN(n4507) );
  AND2_X1 U6178 ( .A1(n4840), .A2(n4445), .ZN(n4508) );
  INV_X1 U6179 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4603) );
  INV_X1 U6180 ( .A(n5704), .ZN(n6351) );
  NAND2_X1 U6181 ( .A1(n5704), .A2(n5703), .ZN(n5706) );
  OAI21_X1 U6182 ( .B1(n5716), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4836) );
  OAI21_X1 U6183 ( .B1(n5716), .B2(n4922), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5717) );
  OR2_X1 U6184 ( .A1(n5716), .A2(n4924), .ZN(n9857) );
  NAND2_X1 U6185 ( .A1(n5704), .A2(n5693), .ZN(n5749) );
  XNOR2_X1 U6186 ( .A(n8359), .B(n8373), .ZN(n8340) );
  MUX2_X1 U6187 ( .A(n7625), .B(n7621), .S(n9487), .Z(n7622) );
  AOI21_X1 U6188 ( .B1(n7678), .B2(n7625), .A(n7454), .ZN(n7455) );
  OAI22_X1 U6189 ( .A1(n4686), .A2(n4683), .B1(n7625), .B2(n7473), .ZN(n4682)
         );
  NOR2_X1 U6190 ( .A1(n4685), .A2(n7625), .ZN(n4684) );
  INV_X1 U6191 ( .A(n7625), .ZN(n4677) );
  NAND2_X1 U6192 ( .A1(n9245), .A2(n9246), .ZN(n9244) );
  NAND2_X1 U6193 ( .A1(n4666), .A2(n9347), .ZN(n4665) );
  XNOR2_X2 U6194 ( .A(n7813), .B(n7830), .ZN(n7845) );
  AOI21_X2 U6195 ( .B1(n4877), .B2(n4876), .A(n4490), .ZN(n7159) );
  INV_X1 U6196 ( .A(n7800), .ZN(n4518) );
  NAND2_X2 U6197 ( .A1(n5721), .A2(n9865), .ZN(n7440) );
  XNOR2_X2 U6198 ( .A(n5719), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U6199 ( .A1(n4709), .A2(n4708), .ZN(n7962) );
  NAND2_X1 U6200 ( .A1(n7874), .A2(n7873), .ZN(n4710) );
  NAND2_X1 U6201 ( .A1(n4725), .A2(n7953), .ZN(n7955) );
  INV_X1 U6202 ( .A(n4714), .ZN(n4712) );
  NAND2_X1 U6203 ( .A1(n7914), .A2(n4728), .ZN(n4727) );
  XNOR2_X1 U6204 ( .A(n7308), .B(n7334), .ZN(n7363) );
  AOI21_X1 U6205 ( .B1(n8435), .B2(n9885), .A(n4524), .ZN(n4523) );
  AND2_X1 U6206 ( .A1(n4525), .A2(n4523), .ZN(n8436) );
  NAND2_X1 U6207 ( .A1(n5616), .A2(n8199), .ZN(n8513) );
  NOR2_X1 U6208 ( .A1(n7865), .A2(n8444), .ZN(n7870) );
  OAI21_X1 U6209 ( .B1(n8465), .B2(n8228), .A(n8230), .ZN(n8453) );
  XNOR2_X1 U6210 ( .A(n9061), .B(n9062), .ZN(n9170) );
  AOI21_X2 U6211 ( .B1(n4518), .B2(n4517), .A(n4516), .ZN(n9688) );
  INV_X1 U6212 ( .A(n4635), .ZN(n4634) );
  AOI21_X1 U6213 ( .B1(n6358), .B2(n10116), .A(n10118), .ZN(n10136) );
  NAND2_X1 U6214 ( .A1(n4521), .A2(n4843), .ZN(n8386) );
  NOR2_X1 U6215 ( .A1(n7363), .A2(n7055), .ZN(n7362) );
  NOR2_X1 U6216 ( .A1(n7336), .A2(n7364), .ZN(n7340) );
  NOR2_X1 U6217 ( .A1(n10133), .A2(n10305), .ZN(n10132) );
  INV_X1 U6218 ( .A(n6367), .ZN(n4795) );
  AOI21_X2 U6219 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n10155), .A(n10147), .ZN(
        n6995) );
  INV_X1 U6220 ( .A(n7090), .ZN(n4877) );
  NAND2_X1 U6221 ( .A1(n7159), .A2(n4494), .ZN(n7161) );
  NAND2_X1 U6222 ( .A1(n4881), .A2(n4879), .ZN(n7813) );
  NAND2_X1 U6223 ( .A1(n4637), .A2(n4634), .ZN(P1_U3519) );
  OAI21_X1 U6224 ( .B1(n7845), .B2(n9842), .A(n4636), .ZN(n4635) );
  NAND3_X1 U6225 ( .A1(n8245), .A2(n4538), .A3(n4419), .ZN(n4529) );
  NAND3_X1 U6226 ( .A1(n4535), .A2(n4533), .A3(n4531), .ZN(n4540) );
  NAND2_X1 U6227 ( .A1(n4540), .A2(n4539), .ZN(n8257) );
  NAND2_X1 U6228 ( .A1(n8255), .A2(n8244), .ZN(n4541) );
  NAND2_X1 U6229 ( .A1(n5425), .A2(n4422), .ZN(n4542) );
  NAND2_X1 U6230 ( .A1(n5425), .A2(n5136), .ZN(n5441) );
  NAND2_X1 U6231 ( .A1(n5287), .A2(n4553), .ZN(n4550) );
  NAND3_X1 U6232 ( .A1(n4565), .A2(n4567), .A3(n4482), .ZN(n4563) );
  NAND3_X1 U6233 ( .A1(n8222), .A2(n5528), .A3(n4573), .ZN(n8227) );
  NAND4_X1 U6234 ( .A1(n4577), .A2(n8212), .A3(n4575), .A4(n4574), .ZN(n4573)
         );
  NAND2_X1 U6235 ( .A1(n6277), .A2(n6260), .ZN(n6259) );
  AND2_X1 U6236 ( .A1(n9514), .A2(n4583), .ZN(n9488) );
  OR2_X1 U6237 ( .A1(n9514), .A2(n9793), .ZN(n4581) );
  NAND2_X1 U6238 ( .A1(n9514), .A2(n9505), .ZN(n9498) );
  NAND3_X1 U6239 ( .A1(n4581), .A2(n4580), .A3(n4578), .ZN(n9481) );
  NAND3_X1 U6240 ( .A1(n9514), .A2(n4582), .A3(n9793), .ZN(n4580) );
  NAND2_X1 U6241 ( .A1(n4595), .A2(n5188), .ZN(n5069) );
  XNOR2_X1 U6242 ( .A(n4595), .B(n5188), .ZN(n5992) );
  NAND2_X1 U6243 ( .A1(n5223), .A2(n5222), .ZN(n4596) );
  NAND2_X1 U6244 ( .A1(n5206), .A2(n5205), .ZN(n4597) );
  INV_X1 U6245 ( .A(n9674), .ZN(n4819) );
  NAND2_X2 U6246 ( .A1(n5091), .A2(n5090), .ZN(n5287) );
  NAND2_X1 U6247 ( .A1(n4607), .A2(n4606), .ZN(n7147) );
  NAND4_X1 U6248 ( .A1(n6703), .A2(n7706), .A3(n7650), .A4(n7654), .ZN(n4607)
         );
  NAND3_X1 U6249 ( .A1(n6703), .A2(n7706), .A3(n7650), .ZN(n4608) );
  NAND2_X1 U6250 ( .A1(n9635), .A2(n4614), .ZN(n4612) );
  AOI21_X1 U6251 ( .B1(n9511), .B2(n9508), .A(n4633), .ZN(n9494) );
  NAND2_X2 U6252 ( .A1(n4641), .A2(n9284), .ZN(n9288) );
  AOI21_X2 U6253 ( .B1(n6081), .B2(n4645), .A(n4644), .ZN(n6113) );
  NAND2_X1 U6254 ( .A1(n9256), .A2(n4651), .ZN(n4649) );
  NAND3_X1 U6255 ( .A1(n4665), .A2(n9160), .A3(n9931), .ZN(n9361) );
  OAI21_X2 U6256 ( .B1(n9323), .B2(n4873), .A(n4668), .ZN(n9061) );
  NAND2_X1 U6257 ( .A1(n9223), .A2(n9111), .ZN(n9116) );
  INV_X1 U6258 ( .A(n5729), .ZN(n5734) );
  INV_X1 U6259 ( .A(n7722), .ZN(n7699) );
  INV_X1 U6260 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4675) );
  INV_X1 U6261 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U6262 ( .A1(n7459), .A2(n7625), .ZN(n4676) );
  NAND4_X2 U6263 ( .A1(n4681), .A2(n5930), .A3(n5929), .A4(n5928), .ZN(n9399)
         );
  OAI21_X1 U6264 ( .B1(n4687), .B2(n4682), .A(n7476), .ZN(n7490) );
  NOR2_X1 U6265 ( .A1(n4688), .A2(n4677), .ZN(n4687) );
  OR2_X1 U6266 ( .A1(n7504), .A2(n4693), .ZN(n4692) );
  OR2_X1 U6267 ( .A1(n7503), .A2(n4694), .ZN(n4691) );
  NAND3_X1 U6268 ( .A1(n4691), .A2(n4692), .A3(n4689), .ZN(n7541) );
  AND3_X1 U6269 ( .A1(n4692), .A2(n4691), .A3(n4478), .ZN(n7538) );
  INV_X1 U6270 ( .A(n7512), .ZN(n4695) );
  NAND2_X1 U6271 ( .A1(n7603), .A2(n4700), .ZN(n4699) );
  NAND3_X1 U6272 ( .A1(n5048), .A2(n4716), .A3(n5045), .ZN(n5411) );
  NAND2_X1 U6273 ( .A1(n7987), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U6274 ( .A1(n4737), .A2(n4476), .ZN(n6956) );
  AND2_X4 U6275 ( .A1(n5649), .A2(n4741), .ZN(n7896) );
  XNOR2_X1 U6276 ( .A(n7896), .B(n10219), .ZN(n6220) );
  XNOR2_X1 U6277 ( .A(n5154), .B(n5051), .ZN(n5595) );
  NAND2_X1 U6278 ( .A1(n8454), .A2(n4744), .ZN(n4743) );
  OAI21_X1 U6279 ( .B1(n8454), .B2(n5569), .A(n5568), .ZN(n7847) );
  OAI21_X1 U6280 ( .B1(n8586), .B2(n4762), .A(n4760), .ZN(n8562) );
  INV_X1 U6281 ( .A(n8562), .ZN(n5437) );
  OAI22_X1 U6282 ( .A1(n8508), .A2(n4764), .B1(n4765), .B2(n5491), .ZN(n8484)
         );
  INV_X1 U6283 ( .A(n8508), .ZN(n4769) );
  NAND2_X1 U6284 ( .A1(n8484), .A2(n5021), .ZN(n5510) );
  NAND2_X1 U6285 ( .A1(n4772), .A2(n4480), .ZN(n5548) );
  NAND2_X1 U6286 ( .A1(n5265), .A2(n4434), .ZN(n6822) );
  NAND3_X1 U6287 ( .A1(n5215), .A2(n4774), .A3(n4773), .ZN(n6544) );
  NAND2_X1 U6288 ( .A1(n4775), .A2(n5214), .ZN(n4773) );
  NAND3_X1 U6289 ( .A1(n5197), .A2(n5214), .A3(n8036), .ZN(n4774) );
  NAND2_X1 U6290 ( .A1(n7256), .A2(n4776), .ZN(n5395) );
  NAND2_X1 U6291 ( .A1(n5439), .A2(n4779), .ZN(n4781) );
  INV_X1 U6292 ( .A(n4781), .ZN(n8550) );
  NAND2_X1 U6293 ( .A1(n5049), .A2(n4786), .ZN(n5153) );
  NAND2_X1 U6294 ( .A1(n5049), .A2(n5013), .ZN(n5587) );
  NAND2_X1 U6295 ( .A1(n6858), .A2(n4801), .ZN(n4796) );
  NAND2_X1 U6296 ( .A1(n4796), .A2(n4798), .ZN(n10147) );
  NAND3_X1 U6297 ( .A1(n4800), .A2(n6857), .A3(n4799), .ZN(n4798) );
  NAND2_X1 U6298 ( .A1(n4800), .A2(n6857), .ZN(n6659) );
  NAND2_X1 U6299 ( .A1(n4802), .A2(n6648), .ZN(n4800) );
  INV_X1 U6300 ( .A(n4808), .ZN(n7331) );
  INV_X1 U6301 ( .A(n7332), .ZN(n4807) );
  NAND2_X1 U6302 ( .A1(n6292), .A2(n4822), .ZN(n4821) );
  NAND3_X1 U6303 ( .A1(n4821), .A2(n6243), .A3(n4820), .ZN(n6261) );
  INV_X2 U6304 ( .A(n10106), .ZN(n4826) );
  INV_X1 U6305 ( .A(n4840), .ZN(n6842) );
  NAND3_X1 U6306 ( .A1(n5166), .A2(n4842), .A3(n4475), .ZN(n4841) );
  NOR2_X1 U6307 ( .A1(n5895), .A2(n5896), .ZN(n6373) );
  NAND2_X1 U6308 ( .A1(n8416), .A2(n4851), .ZN(n4850) );
  NOR2_X1 U6309 ( .A1(n8387), .A2(n8580), .ZN(n8415) );
  INV_X1 U6310 ( .A(n8387), .ZN(n4849) );
  INV_X1 U6311 ( .A(n9879), .ZN(n4851) );
  NAND2_X1 U6312 ( .A1(n4860), .A2(n4861), .ZN(n10139) );
  INV_X1 U6313 ( .A(n6378), .ZN(n4860) );
  NAND2_X1 U6314 ( .A1(n6377), .A2(n6376), .ZN(n4861) );
  NAND2_X1 U6315 ( .A1(n4866), .A2(n4865), .ZN(n6317) );
  INV_X1 U6316 ( .A(n6250), .ZN(n4869) );
  NAND2_X1 U6317 ( .A1(n6251), .A2(n6250), .ZN(n6257) );
  OAI21_X1 U6318 ( .B1(n9521), .B2(n4420), .A(n4882), .ZN(n9492) );
  NAND2_X1 U6319 ( .A1(n9521), .A2(n4426), .ZN(n4881) );
  INV_X1 U6320 ( .A(n9688), .ZN(n4893) );
  NAND2_X1 U6321 ( .A1(n9688), .A2(n4890), .ZN(n4885) );
  NAND2_X1 U6322 ( .A1(n9288), .A2(n9132), .ZN(n9245) );
  NAND2_X1 U6323 ( .A1(n9031), .A2(n9030), .ZN(n4913) );
  NAND2_X1 U6324 ( .A1(n4913), .A2(n9033), .ZN(n4914) );
  NAND3_X1 U6325 ( .A1(n4914), .A2(n4915), .A3(n9922), .ZN(n9920) );
  NAND2_X1 U6326 ( .A1(n9031), .A2(n4916), .ZN(n4915) );
  NOR2_X1 U6327 ( .A1(n9033), .A2(n4917), .ZN(n4916) );
  NAND2_X1 U6328 ( .A1(n6503), .A2(n5015), .ZN(n4919) );
  NAND3_X1 U6329 ( .A1(n4921), .A2(n6122), .A3(n6121), .ZN(n4920) );
  NOR2_X1 U6330 ( .A1(n5716), .A2(n4926), .ZN(n5741) );
  NAND2_X1 U6331 ( .A1(n5571), .A2(n5570), .ZN(n4952) );
  NAND2_X1 U6332 ( .A1(n5504), .A2(n5503), .ZN(n5512) );
  NAND2_X1 U6333 ( .A1(n5504), .A2(n4957), .ZN(n4956) );
  OAI21_X2 U6334 ( .B1(n8480), .B2(n4970), .A(n8225), .ZN(n8465) );
  NAND2_X1 U6335 ( .A1(n5605), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U6336 ( .A1(n6942), .A2(n4979), .ZN(n4978) );
  NAND2_X1 U6337 ( .A1(n5052), .A2(n5051), .ZN(n5054) );
  NAND2_X1 U6338 ( .A1(n5052), .A2(n4984), .ZN(n8724) );
  NAND2_X1 U6339 ( .A1(n4986), .A2(n4985), .ZN(n5612) );
  NAND3_X1 U6340 ( .A1(n4988), .A2(n4987), .A3(n10238), .ZN(n8090) );
  OAI21_X1 U6341 ( .B1(n8513), .B2(n4991), .A(n4435), .ZN(n5619) );
  NAND2_X1 U6342 ( .A1(n8561), .A2(n4994), .ZN(n5615) );
  OAI21_X1 U6343 ( .B1(n8258), .B2(n8259), .A(n4999), .ZN(n8261) );
  NAND2_X1 U6344 ( .A1(n5001), .A2(n5000), .ZN(n4999) );
  AOI21_X1 U6345 ( .B1(n8072), .B2(n6939), .A(n8260), .ZN(n5000) );
  NAND2_X1 U6346 ( .A1(n5003), .A2(n5002), .ZN(n5001) );
  NAND2_X1 U6347 ( .A1(n5005), .A2(n5004), .ZN(n5003) );
  NOR2_X1 U6348 ( .A1(n8070), .A2(n8252), .ZN(n5004) );
  NAND2_X1 U6349 ( .A1(n8071), .A2(n8244), .ZN(n5005) );
  OAI21_X1 U6350 ( .B1(n9161), .B2(n9211), .A(n9931), .ZN(n9168) );
  NAND2_X1 U6351 ( .A1(n5548), .A2(n5547), .ZN(n8454) );
  NAND2_X1 U6352 ( .A1(n5187), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5170) );
  XNOR2_X1 U6353 ( .A(n9492), .B(n9493), .ZN(n9797) );
  NAND2_X1 U6354 ( .A1(n5680), .A2(n10300), .ZN(n5665) );
  AOI21_X1 U6355 ( .B1(n5599), .B2(n10207), .A(n5598), .ZN(n7775) );
  OR2_X1 U6356 ( .A1(n5741), .A2(n5864), .ZN(n5743) );
  CLKBUF_X1 U6357 ( .A(n9256), .Z(n9257) );
  NOR2_X2 U6358 ( .A1(n9529), .A2(n9724), .ZN(n9514) );
  AOI21_X2 U6359 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10184), .A(n10189), .ZN(
        n7308) );
  OAI21_X2 U6360 ( .B1(n9554), .B2(n7807), .A(n7806), .ZN(n9543) );
  AND2_X1 U6361 ( .A1(n8561), .A2(n8560), .ZN(n8638) );
  AOI21_X2 U6362 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8351), .A(n8339), .ZN(
        n8359) );
  INV_X1 U6363 ( .A(n8559), .ZN(n5614) );
  CLKBUF_X1 U6364 ( .A(n7264), .Z(n7265) );
  CLKBUF_X1 U6365 ( .A(n8594), .Z(n8595) );
  CLKBUF_X1 U6366 ( .A(n7203), .Z(n7204) );
  OR2_X2 U6367 ( .A1(n5600), .A2(n8078), .ZN(n6193) );
  XOR2_X1 U6368 ( .A(n9523), .B(n9521), .Z(n9805) );
  NAND2_X1 U6369 ( .A1(n6061), .A2(n5183), .ZN(n10223) );
  AOI22_X1 U6370 ( .A1(n5990), .A2(n5989), .B1(n5988), .B2(n5987), .ZN(n6081)
         );
  INV_X1 U6371 ( .A(n8283), .ZN(n10222) );
  CLKBUF_X1 U6372 ( .A(n5595), .Z(n5877) );
  INV_X2 U6373 ( .A(n10302), .ZN(n10300) );
  INV_X1 U6374 ( .A(n8702), .ZN(n5662) );
  NAND2_X2 U6375 ( .A1(n6170), .A2(n10217), .ZN(n8601) );
  AND2_X2 U6376 ( .A1(n6164), .A2(n5679), .ZN(n10325) );
  OR2_X1 U6377 ( .A1(n9828), .A2(n9227), .ZN(n5008) );
  AND2_X1 U6378 ( .A1(n5664), .A2(n5663), .ZN(n5010) );
  AND2_X1 U6379 ( .A1(n5936), .A2(n9204), .ZN(n5011) );
  AND2_X1 U6380 ( .A1(n5442), .A2(n5445), .ZN(n5013) );
  OR2_X1 U6381 ( .A1(n6669), .A2(n9396), .ZN(n5014) );
  OR2_X1 U6382 ( .A1(n6416), .A2(n6415), .ZN(n5015) );
  OR2_X1 U6383 ( .A1(n6428), .A2(n9394), .ZN(n5016) );
  OR3_X1 U6384 ( .A1(n6499), .A2(n6628), .A3(n6500), .ZN(n5017) );
  OR2_X1 U6385 ( .A1(n9669), .A2(n9272), .ZN(n5018) );
  AND2_X1 U6386 ( .A1(n5101), .A2(n5100), .ZN(n5019) );
  XNOR2_X1 U6387 ( .A(n5698), .B(n5700), .ZN(n5902) );
  OR2_X1 U6388 ( .A1(n6253), .A2(n9411), .ZN(n5020) );
  INV_X1 U6389 ( .A(n7946), .ZN(n8551) );
  AND4_X1 U6390 ( .A1(n5465), .A2(n5464), .A3(n5463), .A4(n5462), .ZN(n7946)
         );
  AOI21_X1 U6391 ( .B1(n8524), .B2(n8523), .A(n5480), .ZN(n8508) );
  INV_X1 U6392 ( .A(n8632), .ZN(n5466) );
  OR2_X1 U6393 ( .A1(n8501), .A2(n8672), .ZN(n5021) );
  INV_X1 U6394 ( .A(n6752), .ZN(n6076) );
  OR2_X1 U6395 ( .A1(n7181), .A2(n8277), .ZN(n5022) );
  INV_X1 U6396 ( .A(n7755), .ZN(n6098) );
  OR2_X1 U6397 ( .A1(n6432), .A2(n6322), .ZN(n10098) );
  INV_X1 U6398 ( .A(n8165), .ZN(n5379) );
  OR2_X1 U6399 ( .A1(n8012), .A2(n8475), .ZN(n5023) );
  INV_X1 U6400 ( .A(n7912), .ZN(n8658) );
  INV_X1 U6401 ( .A(n8472), .ZN(n5528) );
  NAND2_X1 U6402 ( .A1(n6824), .A2(n6690), .ZN(n5263) );
  INV_X1 U6403 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5043) );
  INV_X1 U6404 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5688) );
  INV_X1 U6405 ( .A(n9028), .ZN(n9029) );
  INV_X1 U6406 ( .A(n5779), .ZN(n5686) );
  NAND2_X1 U6407 ( .A1(n9027), .A2(n9029), .ZN(n9030) );
  INV_X1 U6408 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5694) );
  INV_X1 U6409 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U6410 ( .A1(n8672), .A2(n8501), .ZN(n5509) );
  NAND2_X1 U6411 ( .A1(n5153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5154) );
  AND2_X1 U6412 ( .A1(n9286), .A2(n9124), .ZN(n9187) );
  INV_X1 U6413 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6444) );
  INV_X1 U6414 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6709) );
  AND2_X1 U6415 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n7439), .ZN(n7428) );
  INV_X1 U6416 ( .A(SI_19_), .ZN(n8922) );
  INV_X1 U6417 ( .A(n5349), .ZN(n5114) );
  INV_X1 U6418 ( .A(SI_8_), .ZN(n5092) );
  INV_X1 U6419 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5030) );
  AND2_X1 U6420 ( .A1(n6144), .A2(n6143), .ZN(n8018) );
  NAND2_X1 U6421 ( .A1(n7912), .A2(n8463), .ZN(n5568) );
  INV_X1 U6422 ( .A(n8563), .ZN(n5613) );
  INV_X1 U6423 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5025) );
  OR2_X1 U6424 ( .A1(n8256), .A2(n5621), .ZN(n6141) );
  AND2_X1 U6425 ( .A1(n7586), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7588) );
  NOR2_X1 U6426 ( .A1(n6802), .A2(n6801), .ZN(n6925) );
  INV_X1 U6427 ( .A(n6076), .ZN(n9137) );
  INV_X1 U6428 ( .A(n7407), .ZN(n7430) );
  OR2_X1 U6429 ( .A1(n7592), .A2(n5720), .ZN(n5723) );
  INV_X1 U6430 ( .A(n9793), .ZN(n9480) );
  INV_X1 U6431 ( .A(n6205), .ZN(n7439) );
  AND2_X1 U6432 ( .A1(n7573), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7586) );
  AND2_X1 U6433 ( .A1(n6925), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7080) );
  OR2_X1 U6434 ( .A1(n9395), .A2(n10046), .ZN(n6250) );
  NAND2_X1 U6435 ( .A1(n6240), .A2(n7646), .ZN(n6234) );
  NAND2_X1 U6436 ( .A1(n5729), .A2(n5730), .ZN(n5709) );
  NOR2_X1 U6437 ( .A1(n5129), .A2(SI_17_), .ZN(n5130) );
  OR2_X1 U6438 ( .A1(n6040), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6138) );
  AND2_X1 U6439 ( .A1(n5250), .A2(n5080), .ZN(n5079) );
  INV_X1 U6440 ( .A(n8578), .ZN(n7967) );
  INV_X1 U6441 ( .A(n8422), .ZN(n8419) );
  OR2_X1 U6442 ( .A1(n5575), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8440) );
  INV_X1 U6443 ( .A(n8223), .ZN(n8464) );
  NOR2_X1 U6444 ( .A1(n8202), .A2(n8206), .ZN(n8512) );
  INV_X1 U6445 ( .A(n8239), .ZN(n8242) );
  AND3_X1 U6446 ( .A1(n5669), .A2(P2_STATE_REG_SCAN_IN), .A3(n6046), .ZN(n5670) );
  INV_X1 U6447 ( .A(n8274), .ZN(n7290) );
  AND2_X1 U6448 ( .A1(n5654), .A2(n6147), .ZN(n10225) );
  NOR2_X1 U6449 ( .A1(n6044), .A2(n5656), .ZN(n6057) );
  NAND2_X1 U6450 ( .A1(n9170), .A2(n9171), .ZN(n9169) );
  OR2_X1 U6451 ( .A1(n5923), .A2(n5922), .ZN(n5925) );
  INV_X1 U6452 ( .A(n9184), .ZN(n9582) );
  NAND2_X1 U6453 ( .A1(n7516), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7532) );
  AND2_X1 U6454 ( .A1(n10019), .A2(n6881), .ZN(n6882) );
  AND2_X1 U6455 ( .A1(n7783), .A2(n7782), .ZN(n10027) );
  OR2_X1 U6456 ( .A1(n9525), .A2(n9578), .ZN(n9527) );
  INV_X1 U6457 ( .A(n9813), .ZN(n9558) );
  INV_X1 U6458 ( .A(n7665), .ZN(n7731) );
  INV_X1 U6459 ( .A(n7539), .ZN(n7732) );
  OR2_X1 U6460 ( .A1(n9172), .A2(n9385), .ZN(n7209) );
  NAND2_X1 U6461 ( .A1(n6610), .A2(n6609), .ZN(n6612) );
  OR2_X1 U6462 ( .A1(n7625), .A2(n6098), .ZN(n6283) );
  AND2_X1 U6463 ( .A1(n5572), .A2(n5557), .ZN(n5570) );
  AND2_X1 U6464 ( .A1(n5503), .A2(n5152), .ZN(n5501) );
  OR2_X1 U6465 ( .A1(n5084), .A2(n5083), .ZN(n5085) );
  INV_X1 U6466 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n8964) );
  NAND2_X1 U6467 ( .A1(n6060), .A2(n10217), .ZN(n7969) );
  AND2_X1 U6468 ( .A1(n5527), .A2(n5526), .ZN(n8486) );
  AND4_X1 U6469 ( .A1(n5408), .A2(n5407), .A3(n5406), .A4(n5405), .ZN(n7875)
         );
  OR2_X1 U6470 ( .A1(P2_U3150), .A2(n5897), .ZN(n10183) );
  NOR2_X1 U6471 ( .A1(n8290), .A2(n8289), .ZN(n8311) );
  XNOR2_X1 U6472 ( .A(n7847), .B(n5583), .ZN(n5599) );
  INV_X1 U6473 ( .A(n8677), .ZN(n8505) );
  INV_X1 U6474 ( .A(n10218), .ZN(n7262) );
  INV_X1 U6475 ( .A(n6573), .ZN(n10254) );
  AND2_X1 U6476 ( .A1(n6142), .A2(n8249), .ZN(n10202) );
  INV_X1 U6477 ( .A(n8516), .ZN(n10210) );
  AND2_X1 U6478 ( .A1(n10325), .A2(n10299), .ZN(n8646) );
  AND2_X1 U6479 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  INV_X1 U6480 ( .A(n10299), .ZN(n10282) );
  AND2_X1 U6481 ( .A1(n8177), .A2(n8179), .ZN(n8585) );
  INV_X1 U6482 ( .A(n10294), .ZN(n10275) );
  INV_X1 U6483 ( .A(n7280), .ZN(n5856) );
  AND2_X1 U6484 ( .A1(n5879), .A2(n5853), .ZN(n6059) );
  INV_X1 U6485 ( .A(n9357), .ZN(n9926) );
  INV_X1 U6486 ( .A(n9935), .ZN(n9359) );
  AND4_X1 U6487 ( .A1(n7434), .A2(n7433), .A3(n7432), .A4(n7431), .ZN(n9248)
         );
  AND3_X1 U6488 ( .A1(n7520), .A2(n7519), .A3(n7518), .ZN(n9340) );
  INV_X1 U6489 ( .A(n10028), .ZN(n9474) );
  OR2_X1 U6490 ( .A1(n10012), .A2(n10011), .ZN(n10019) );
  AND2_X1 U6491 ( .A1(n7692), .A2(n7691), .ZN(n9604) );
  INV_X1 U6492 ( .A(n9578), .ZN(n9697) );
  INV_X1 U6493 ( .A(n6260), .ZN(n10046) );
  INV_X1 U6494 ( .A(n9789), .ZN(n9773) );
  AND2_X1 U6495 ( .A1(n7688), .A2(n7825), .ZN(n9523) );
  NAND2_X1 U6496 ( .A1(n6290), .A2(n6283), .ZN(n10096) );
  AND3_X1 U6497 ( .A1(n5918), .A2(P1_STATE_REG_SCAN_IN), .A3(n5774), .ZN(n9853) );
  AND2_X1 U6498 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7016), .ZN(n10350) );
  NOR2_X1 U6499 ( .A1(n10345), .A2(n10344), .ZN(n7034) );
  NOR2_X1 U6500 ( .A1(n7045), .A2(n7044), .ZN(n10331) );
  INV_X1 U6501 ( .A(n7062), .ZN(n10277) );
  AND2_X1 U6502 ( .A1(n6056), .A2(n6055), .ZN(n7972) );
  INV_X1 U6503 ( .A(n7969), .ZN(n8025) );
  INV_X1 U6504 ( .A(n8565), .ZN(n8588) );
  INV_X1 U6505 ( .A(n9885), .ZN(n10191) );
  INV_X1 U6506 ( .A(n10213), .ZN(n8605) );
  INV_X1 U6507 ( .A(n8601), .ZN(n10235) );
  NAND2_X1 U6508 ( .A1(n8239), .A2(n8646), .ZN(n5684) );
  INV_X1 U6509 ( .A(n8646), .ZN(n8640) );
  NAND2_X1 U6510 ( .A1(n10325), .A2(n10275), .ZN(n8649) );
  INV_X1 U6511 ( .A(n10325), .ZN(n10323) );
  XNOR2_X1 U6512 ( .A(n8453), .B(n4438), .ZN(n8661) );
  OR2_X1 U6513 ( .A1(n10302), .A2(n10282), .ZN(n8702) );
  OR2_X1 U6514 ( .A1(n10302), .A2(n10294), .ZN(n8721) );
  AND2_X1 U6515 ( .A1(n5661), .A2(n5660), .ZN(n10302) );
  INV_X1 U6516 ( .A(n5862), .ZN(n5863) );
  INV_X1 U6517 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8871) );
  INV_X1 U6518 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8840) );
  INV_X1 U6519 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8880) );
  XNOR2_X1 U6520 ( .A(n5711), .B(n5710), .ZN(n5774) );
  INV_X1 U6521 ( .A(n9752), .ZN(n9614) );
  AND2_X1 U6522 ( .A1(n5921), .A2(n7768), .ZN(n9935) );
  AOI21_X1 U6523 ( .B1(n5932), .B2(n6332), .A(n10065), .ZN(n9928) );
  AND4_X1 U6524 ( .A1(n6209), .A2(n6208), .A3(n6207), .A4(n6206), .ZN(n9353)
         );
  AOI21_X1 U6525 ( .B1(n9556), .B2(n7594), .A(n6019), .ZN(n9247) );
  INV_X1 U6526 ( .A(n9050), .ZN(n9386) );
  INV_X1 U6527 ( .A(n9948), .ZN(n10039) );
  INV_X1 U6528 ( .A(n9487), .ZN(n9937) );
  AND2_X1 U6529 ( .A1(n6412), .A2(n6328), .ZN(n9701) );
  INV_X1 U6530 ( .A(n10067), .ZN(n9712) );
  INV_X1 U6531 ( .A(n9846), .ZN(n9783) );
  NAND2_X1 U6532 ( .A1(n10100), .A2(n9767), .ZN(n9852) );
  INV_X2 U6533 ( .A(n10098), .ZN(n10100) );
  INV_X1 U6534 ( .A(n10077), .ZN(n10078) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7599) );
  INV_X1 U6536 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6014) );
  NOR2_X1 U6537 ( .A1(n7035), .A2(n7034), .ZN(n10343) );
  NAND2_X1 U6538 ( .A1(n5665), .A2(n5010), .ZN(P2_U3455) );
  AND2_X1 U6539 ( .A1(n5712), .A2(n5774), .ZN(P1_U3973) );
  INV_X4 U6540 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10212) );
  NAND2_X1 U6541 ( .A1(n10212), .A2(n5025), .ZN(n5231) );
  INV_X1 U6542 ( .A(n5231), .ZN(n5027) );
  OR2_X2 U6543 ( .A1(n5244), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5266) );
  INV_X1 U6544 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5033) );
  INV_X1 U6545 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5035) );
  INV_X1 U6546 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5037) );
  INV_X1 U6547 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8977) );
  INV_X1 U6548 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5040) );
  OR2_X2 U6549 ( .A1(n5485), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6550 ( .A1(n5487), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5042) );
  NAND2_X1 U6551 ( .A1(n5494), .A2(n5042), .ZN(n8504) );
  INV_X1 U6552 ( .A(n5153), .ZN(n5052) );
  INV_X1 U6553 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U6554 ( .A1(n8504), .A2(n5432), .ZN(n5059) );
  NOR2_X2 U6555 ( .A1(n8729), .A2(n5159), .ZN(n5187) );
  AOI22_X1 U6556 ( .A1(n4414), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n7854), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n5058) );
  INV_X1 U6557 ( .A(n8729), .ZN(n5161) );
  AND2_X2 U6558 ( .A1(n5161), .A2(n5159), .ZN(n5184) );
  BUF_X1 U6559 ( .A(n5184), .Z(n5216) );
  NAND2_X1 U6560 ( .A1(n5184), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5057) );
  AND2_X1 U6561 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5060) );
  NAND2_X1 U6562 ( .A1(n5179), .A2(n5060), .ZN(n5739) );
  NAND3_X1 U6563 ( .A1(n5939), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5061) );
  NAND2_X1 U6564 ( .A1(n5739), .A2(n5061), .ZN(n5162) );
  INV_X1 U6565 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5816) );
  INV_X1 U6566 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U6567 ( .A1(n5162), .A2(n5163), .ZN(n5065) );
  INV_X1 U6568 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6569 ( .A1(n5063), .A2(SI_1_), .ZN(n5064) );
  INV_X1 U6570 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5815) );
  MUX2_X1 U6571 ( .A(n5815), .B(n5991), .S(n5179), .Z(n5066) );
  XNOR2_X1 U6572 ( .A(n5066), .B(SI_2_), .ZN(n5188) );
  INV_X1 U6573 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6574 ( .A1(n5067), .A2(SI_2_), .ZN(n5068) );
  NAND2_X1 U6575 ( .A1(n5069), .A2(n5068), .ZN(n5206) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5817) );
  INV_X1 U6577 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6069) );
  MUX2_X1 U6578 ( .A(n5817), .B(n6069), .S(n5179), .Z(n5070) );
  XNOR2_X1 U6579 ( .A(n5070), .B(SI_3_), .ZN(n5205) );
  INV_X1 U6580 ( .A(n5070), .ZN(n5071) );
  NAND2_X1 U6581 ( .A1(n5071), .A2(SI_3_), .ZN(n5072) );
  MUX2_X1 U6582 ( .A(n5818), .B(n6116), .S(n5179), .Z(n5073) );
  XNOR2_X1 U6583 ( .A(n5073), .B(SI_4_), .ZN(n5222) );
  INV_X1 U6584 ( .A(n5073), .ZN(n5074) );
  NAND2_X1 U6585 ( .A1(n5074), .A2(SI_4_), .ZN(n5075) );
  MUX2_X1 U6586 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5179), .Z(n5081) );
  XNOR2_X1 U6587 ( .A(n5081), .B(SI_5_), .ZN(n5237) );
  INV_X1 U6588 ( .A(n5237), .ZN(n5250) );
  MUX2_X1 U6589 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5179), .Z(n5076) );
  NAND2_X1 U6590 ( .A1(n5076), .A2(SI_6_), .ZN(n5082) );
  INV_X1 U6591 ( .A(n5082), .ZN(n5078) );
  XNOR2_X1 U6592 ( .A(n5076), .B(SI_6_), .ZN(n5254) );
  INV_X1 U6593 ( .A(n5254), .ZN(n5077) );
  NAND2_X1 U6594 ( .A1(n5251), .A2(n5079), .ZN(n5086) );
  INV_X1 U6595 ( .A(n5080), .ZN(n5084) );
  NAND2_X1 U6596 ( .A1(n5081), .A2(SI_5_), .ZN(n5252) );
  AND2_X1 U6597 ( .A1(n5252), .A2(n5082), .ZN(n5083) );
  NAND2_X1 U6598 ( .A1(n5086), .A2(n5085), .ZN(n5273) );
  MUX2_X1 U6599 ( .A(n5831), .B(n5087), .S(n5179), .Z(n5088) );
  XNOR2_X1 U6600 ( .A(n5088), .B(SI_7_), .ZN(n5272) );
  NAND2_X1 U6601 ( .A1(n5273), .A2(n5272), .ZN(n5091) );
  INV_X1 U6602 ( .A(n5088), .ZN(n5089) );
  NAND2_X1 U6603 ( .A1(n5089), .A2(SI_7_), .ZN(n5090) );
  MUX2_X1 U6604 ( .A(n5849), .B(n8825), .S(n5179), .Z(n5093) );
  NAND2_X1 U6605 ( .A1(n5093), .A2(n5092), .ZN(n5096) );
  INV_X1 U6606 ( .A(n5093), .ZN(n5094) );
  NAND2_X1 U6607 ( .A1(n5094), .A2(SI_8_), .ZN(n5095) );
  NAND2_X1 U6608 ( .A1(n5096), .A2(n5095), .ZN(n5286) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5097) );
  MUX2_X1 U6610 ( .A(n5097), .B(n8980), .S(n5179), .Z(n5098) );
  NAND2_X1 U6611 ( .A1(n5098), .A2(n8798), .ZN(n5101) );
  INV_X1 U6612 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6613 ( .A1(n5099), .A2(SI_9_), .ZN(n5100) );
  MUX2_X1 U6614 ( .A(n5867), .B(n5865), .S(n5179), .Z(n5102) );
  XNOR2_X1 U6615 ( .A(n5102), .B(SI_10_), .ZN(n5306) );
  INV_X1 U6616 ( .A(n5306), .ZN(n5105) );
  INV_X1 U6617 ( .A(n5102), .ZN(n5103) );
  NAND2_X1 U6618 ( .A1(n5103), .A2(SI_10_), .ZN(n5104) );
  MUX2_X1 U6619 ( .A(n8800), .B(n5106), .S(n5534), .Z(n5107) );
  INV_X1 U6620 ( .A(n5107), .ZN(n5108) );
  NAND2_X1 U6621 ( .A1(n5108), .A2(SI_11_), .ZN(n5109) );
  NAND2_X1 U6622 ( .A1(n5110), .A2(n5109), .ZN(n5318) );
  MUX2_X1 U6623 ( .A(n8880), .B(n6014), .S(n5534), .Z(n5111) );
  INV_X1 U6624 ( .A(n5111), .ZN(n5112) );
  MUX2_X1 U6625 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5534), .Z(n5115) );
  NAND2_X1 U6626 ( .A1(n5350), .A2(n5114), .ZN(n5117) );
  NAND2_X1 U6627 ( .A1(n5115), .A2(SI_13_), .ZN(n5116) );
  MUX2_X1 U6628 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5534), .Z(n5362) );
  NAND2_X1 U6629 ( .A1(n5119), .A2(n5118), .ZN(n5120) );
  MUX2_X1 U6630 ( .A(n5121), .B(n6180), .S(n5534), .Z(n5382) );
  NOR2_X1 U6631 ( .A1(n5122), .A2(SI_15_), .ZN(n5123) );
  MUX2_X1 U6632 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5534), .Z(n5396) );
  NAND2_X1 U6633 ( .A1(n5125), .A2(n5124), .ZN(n5126) );
  INV_X1 U6634 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5127) );
  MUX2_X1 U6635 ( .A(n8967), .B(n5127), .S(n5534), .Z(n5128) );
  INV_X1 U6636 ( .A(n5128), .ZN(n5129) );
  AOI21_X1 U6637 ( .B1(n5410), .B2(n5409), .A(n5130), .ZN(n5421) );
  MUX2_X1 U6638 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5534), .Z(n5131) );
  NAND2_X1 U6639 ( .A1(n5131), .A2(SI_18_), .ZN(n5136) );
  INV_X1 U6640 ( .A(n5131), .ZN(n5133) );
  INV_X1 U6641 ( .A(SI_18_), .ZN(n5132) );
  NAND2_X1 U6642 ( .A1(n5133), .A2(n5132), .ZN(n5134) );
  NAND2_X1 U6643 ( .A1(n5136), .A2(n5134), .ZN(n5422) );
  INV_X1 U6644 ( .A(n5422), .ZN(n5135) );
  NAND2_X1 U6645 ( .A1(n5421), .A2(n5135), .ZN(n5425) );
  MUX2_X1 U6646 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n5534), .Z(n5137) );
  XNOR2_X1 U6647 ( .A(n5137), .B(SI_19_), .ZN(n5440) );
  INV_X1 U6648 ( .A(n5137), .ZN(n5138) );
  NAND2_X1 U6649 ( .A1(n5138), .A2(n8922), .ZN(n5139) );
  MUX2_X1 U6650 ( .A(n6869), .B(n7543), .S(n5534), .Z(n5141) );
  INV_X1 U6651 ( .A(SI_20_), .ZN(n5140) );
  MUX2_X1 U6652 ( .A(n8840), .B(n8932), .S(n5534), .Z(n5468) );
  INV_X1 U6653 ( .A(SI_21_), .ZN(n5142) );
  INV_X1 U6654 ( .A(n5468), .ZN(n5143) );
  MUX2_X1 U6655 ( .A(n6941), .B(n7781), .S(n5534), .Z(n5145) );
  INV_X1 U6656 ( .A(SI_22_), .ZN(n5144) );
  NAND2_X1 U6657 ( .A1(n5145), .A2(n5144), .ZN(n5148) );
  INV_X1 U6658 ( .A(n5145), .ZN(n5146) );
  NAND2_X1 U6659 ( .A1(n5146), .A2(SI_22_), .ZN(n5147) );
  NAND2_X1 U6660 ( .A1(n5148), .A2(n5147), .ZN(n5481) );
  INV_X1 U6661 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5149) );
  MUX2_X1 U6662 ( .A(n5149), .B(n8814), .S(n5534), .Z(n5150) );
  INV_X1 U6663 ( .A(SI_23_), .ZN(n8946) );
  NAND2_X1 U6664 ( .A1(n5150), .A2(n8946), .ZN(n5503) );
  INV_X1 U6665 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6666 ( .A1(n5151), .A2(SI_23_), .ZN(n5152) );
  NAND2_X1 U6667 ( .A1(n7583), .A2(n8060), .ZN(n5158) );
  AND2_X2 U6668 ( .A1(n5181), .A2(n5179), .ZN(n5288) );
  NAND2_X1 U6669 ( .A1(n8061), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6670 ( .A1(n5185), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6671 ( .A1(n5186), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5172) );
  AND2_X1 U6672 ( .A1(n5159), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6673 ( .A1(n5161), .A2(n5160), .ZN(n5171) );
  NAND2_X1 U6674 ( .A1(n5288), .A2(n5816), .ZN(n5169) );
  XNOR2_X1 U6675 ( .A(n5163), .B(n5162), .ZN(n5938) );
  INV_X1 U6676 ( .A(n5938), .ZN(n5164) );
  NAND2_X1 U6677 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5165) );
  MUX2_X1 U6678 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5165), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5166) );
  NAND2_X1 U6679 ( .A1(n5256), .A2(n6356), .ZN(n5167) );
  NAND4_X1 U6680 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n5174)
         );
  NAND2_X1 U6681 ( .A1(n5601), .A2(n8080), .ZN(n5600) );
  NAND2_X1 U6682 ( .A1(n5184), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6683 ( .A1(n5185), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6684 ( .A1(n5187), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U6685 ( .A1(n5186), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5175) );
  NAND4_X2 U6686 ( .A1(n5178), .A2(n5177), .A3(n5176), .A4(n5175), .ZN(n8286)
         );
  NAND2_X1 U6687 ( .A1(n5939), .A2(SI_0_), .ZN(n5180) );
  XNOR2_X1 U6688 ( .A(n5180), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9026) );
  MUX2_X1 U6689 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9026), .S(n5181), .Z(n6172) );
  NAND2_X1 U6690 ( .A1(n8286), .A2(n6172), .ZN(n6196) );
  NAND2_X1 U6691 ( .A1(n5600), .A2(n6196), .ZN(n6195) );
  INV_X1 U6692 ( .A(n5182), .ZN(n8284) );
  INV_X1 U6693 ( .A(n8284), .ZN(n6061) );
  NAND2_X1 U6694 ( .A1(n6195), .A2(n10223), .ZN(n5197) );
  NAND2_X1 U6695 ( .A1(n5185), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5195) );
  NAND2_X1 U6696 ( .A1(n5186), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6697 ( .A1(n5187), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6698 ( .A1(n5288), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6699 ( .A1(n5256), .A2(n6375), .ZN(n5191) );
  OAI211_X1 U6700 ( .C1(n5426), .C2(n5992), .A(n5192), .B(n5191), .ZN(n10238)
         );
  INV_X1 U6701 ( .A(n10238), .ZN(n10219) );
  NAND2_X1 U6702 ( .A1(n5198), .A2(n10219), .ZN(n5199) );
  NAND2_X1 U6703 ( .A1(n5432), .A2(n10212), .ZN(n5204) );
  NAND2_X1 U6704 ( .A1(n5186), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5203) );
  NAND2_X1 U6705 ( .A1(n5216), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U6706 ( .A1(n4414), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5201) );
  XNOR2_X1 U6707 ( .A(n5206), .B(n5205), .ZN(n6068) );
  NAND2_X1 U6708 ( .A1(n5288), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5213) );
  NOR2_X1 U6709 ( .A1(n5209), .A2(n8725), .ZN(n5207) );
  MUX2_X1 U6710 ( .A(n8725), .B(n5207), .S(P2_IR_REG_3__SCAN_IN), .Z(n5211) );
  NAND2_X1 U6711 ( .A1(n5209), .A2(n5208), .ZN(n5238) );
  INV_X1 U6712 ( .A(n5238), .ZN(n5210) );
  NOR2_X2 U6713 ( .A1(n5211), .A2(n5210), .ZN(n6376) );
  NAND2_X1 U6714 ( .A1(n5256), .A2(n6376), .ZN(n5212) );
  OAI211_X1 U6715 ( .C1(n5426), .C2(n6068), .A(n5213), .B(n5212), .ZN(n10243)
         );
  NAND2_X1 U6716 ( .A1(n8283), .A2(n10243), .ZN(n5214) );
  INV_X1 U6717 ( .A(n10243), .ZN(n8088) );
  NAND2_X1 U6718 ( .A1(n10222), .A2(n8088), .ZN(n5215) );
  NAND2_X1 U6719 ( .A1(n5186), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6720 ( .A1(n5216), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5220) );
  NAND2_X1 U6721 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5217) );
  NAND2_X1 U6722 ( .A1(n5231), .A2(n5217), .ZN(n6550) );
  NAND2_X1 U6723 ( .A1(n5432), .A2(n6550), .ZN(n5219) );
  NAND2_X1 U6724 ( .A1(n4414), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5218) );
  XNOR2_X1 U6725 ( .A(n5223), .B(n5222), .ZN(n6114) );
  NAND2_X1 U6726 ( .A1(n5288), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6727 ( .A1(n5238), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5225) );
  INV_X1 U6728 ( .A(n6655), .ZN(n5226) );
  NAND2_X1 U6729 ( .A1(n5256), .A2(n5226), .ZN(n5227) );
  OAI211_X1 U6730 ( .C1(n5426), .C2(n6114), .A(n5228), .B(n5227), .ZN(n10249)
         );
  NOR2_X1 U6731 ( .A1(n10203), .A2(n10249), .ZN(n5230) );
  NAND2_X1 U6732 ( .A1(n10203), .A2(n10249), .ZN(n5229) );
  NAND2_X1 U6733 ( .A1(n4414), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5236) );
  NAND2_X1 U6734 ( .A1(n5186), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U6735 ( .A1(n5231), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5232) );
  NAND2_X1 U6736 ( .A1(n5244), .A2(n5232), .ZN(n6682) );
  NAND2_X1 U6737 ( .A1(n5432), .A2(n6682), .ZN(n5234) );
  NAND2_X1 U6738 ( .A1(n5216), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5233) );
  XNOR2_X1 U6739 ( .A(n5251), .B(n5237), .ZN(n6252) );
  NAND2_X1 U6740 ( .A1(n8060), .A2(n6252), .ZN(n5242) );
  NAND2_X1 U6741 ( .A1(n5288), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5241) );
  NOR2_X1 U6742 ( .A1(n5238), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5258) );
  OR2_X1 U6743 ( .A1(n5258), .A2(n8725), .ZN(n5239) );
  XNOR2_X1 U6744 ( .A(n5239), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6648) );
  NAND2_X1 U6745 ( .A1(n5256), .A2(n6648), .ZN(n5240) );
  NAND2_X1 U6746 ( .A1(n6575), .A2(n6573), .ZN(n6676) );
  NAND2_X1 U6747 ( .A1(n6678), .A2(n6676), .ZN(n5243) );
  NAND2_X1 U6748 ( .A1(n8282), .A2(n10254), .ZN(n6675) );
  NAND2_X1 U6749 ( .A1(n5243), .A2(n6675), .ZN(n6686) );
  NAND2_X1 U6750 ( .A1(n4414), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6751 ( .A1(n5186), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6752 ( .A1(n5244), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5245) );
  NAND2_X1 U6753 ( .A1(n5266), .A2(n5245), .ZN(n6582) );
  NAND2_X1 U6754 ( .A1(n5432), .A2(n6582), .ZN(n5247) );
  NAND2_X1 U6755 ( .A1(n5184), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U6756 ( .A1(n5251), .A2(n5250), .ZN(n5253) );
  NAND2_X1 U6757 ( .A1(n5253), .A2(n5252), .ZN(n5255) );
  XNOR2_X1 U6758 ( .A(n5255), .B(n5254), .ZN(n6301) );
  NAND2_X1 U6759 ( .A1(n8060), .A2(n6301), .ZN(n5262) );
  NAND2_X1 U6760 ( .A1(n5288), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U6761 ( .A1(n5258), .A2(n5257), .ZN(n5274) );
  NAND2_X1 U6762 ( .A1(n5274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5259) );
  XNOR2_X1 U6763 ( .A(n5259), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U6764 ( .A1(n5447), .A2(n6860), .ZN(n5260) );
  NAND2_X1 U6765 ( .A1(n6686), .A2(n5263), .ZN(n5265) );
  INV_X1 U6766 ( .A(n6690), .ZN(n10260) );
  NAND2_X1 U6767 ( .A1(n8281), .A2(n10260), .ZN(n5264) );
  NAND2_X1 U6768 ( .A1(n4414), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6769 ( .A1(n7854), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5270) );
  NAND2_X1 U6770 ( .A1(n5266), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5267) );
  NAND2_X1 U6771 ( .A1(n5278), .A2(n5267), .ZN(n6829) );
  NAND2_X1 U6772 ( .A1(n5432), .A2(n6829), .ZN(n5269) );
  NAND2_X1 U6773 ( .A1(n5216), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6774 ( .A(n5273), .B(n5272), .ZN(n6437) );
  NAND2_X1 U6775 ( .A1(n5288), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n5277) );
  OAI21_X1 U6776 ( .B1(n5274), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5275) );
  XNOR2_X1 U6777 ( .A(n5275), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U6778 ( .A1(n5447), .A2(n6996), .ZN(n5276) );
  OAI211_X1 U6779 ( .C1(n5426), .C2(n6437), .A(n5277), .B(n5276), .ZN(n6832)
         );
  NAND2_X1 U6780 ( .A1(n6962), .A2(n6832), .ZN(n8125) );
  INV_X1 U6781 ( .A(n6962), .ZN(n8280) );
  INV_X1 U6782 ( .A(n6832), .ZN(n10265) );
  NAND2_X1 U6783 ( .A1(n8280), .A2(n10265), .ZN(n6901) );
  NAND2_X1 U6784 ( .A1(n4414), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6785 ( .A1(n7854), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6786 ( .A1(n5278), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5279) );
  NAND2_X1 U6787 ( .A1(n5293), .A2(n5279), .ZN(n6964) );
  NAND2_X1 U6788 ( .A1(n5432), .A2(n6964), .ZN(n5281) );
  NAND2_X1 U6789 ( .A1(n5216), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5280) );
  OR2_X1 U6790 ( .A1(n5284), .A2(n8725), .ZN(n5285) );
  XNOR2_X1 U6791 ( .A(n5285), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6999) );
  XNOR2_X1 U6792 ( .A(n5287), .B(n5286), .ZN(n6441) );
  NAND2_X1 U6793 ( .A1(n6441), .A2(n8060), .ZN(n5290) );
  NAND2_X1 U6794 ( .A1(n5288), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n5289) );
  OAI211_X1 U6795 ( .C1(n5181), .C2(n10171), .A(n5290), .B(n5289), .ZN(n6957)
         );
  NAND2_X1 U6796 ( .A1(n6959), .A2(n6957), .ZN(n8126) );
  NAND2_X1 U6797 ( .A1(n8279), .A2(n10272), .ZN(n8118) );
  NAND2_X1 U6798 ( .A1(n8126), .A2(n8118), .ZN(n8041) );
  NAND2_X1 U6799 ( .A1(n6962), .A2(n10265), .ZN(n6905) );
  AND2_X1 U6800 ( .A1(n8041), .A2(n6905), .ZN(n5291) );
  NAND2_X1 U6801 ( .A1(n8279), .A2(n6957), .ZN(n5292) );
  NAND2_X1 U6802 ( .A1(n6904), .A2(n5292), .ZN(n6893) );
  NAND2_X1 U6803 ( .A1(n4414), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U6804 ( .A1(n7854), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6805 ( .A1(n5293), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5294) );
  NAND2_X1 U6806 ( .A1(n5312), .A2(n5294), .ZN(n7071) );
  NAND2_X1 U6807 ( .A1(n5432), .A2(n7071), .ZN(n5296) );
  NAND2_X1 U6808 ( .A1(n5216), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5295) );
  NAND4_X1 U6809 ( .A1(n5298), .A2(n5297), .A3(n5296), .A4(n5295), .ZN(n8278)
         );
  NAND2_X1 U6810 ( .A1(n9023), .A2(n8060), .ZN(n5303) );
  INV_X1 U6811 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6812 ( .A1(n5284), .A2(n5300), .ZN(n5308) );
  NAND2_X1 U6813 ( .A1(n5308), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5301) );
  XNOR2_X1 U6814 ( .A(n5301), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9021) );
  AOI22_X1 U6815 ( .A1(n8061), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5447), .B2(
        n9021), .ZN(n5302) );
  NAND2_X1 U6816 ( .A1(n5303), .A2(n5302), .ZN(n7062) );
  AND2_X1 U6817 ( .A1(n8278), .A2(n7062), .ZN(n5304) );
  INV_X1 U6818 ( .A(n8278), .ZN(n7179) );
  NAND2_X1 U6819 ( .A1(n7179), .A2(n10277), .ZN(n5305) );
  XNOR2_X1 U6820 ( .A(n5307), .B(n5306), .ZN(n6704) );
  NAND2_X1 U6821 ( .A1(n6704), .A2(n8060), .ZN(n5311) );
  NAND2_X1 U6822 ( .A1(n5320), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6823 ( .A(n5309), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7333) );
  AOI22_X1 U6824 ( .A1(n8061), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5447), .B2(
        n7333), .ZN(n5310) );
  NAND2_X1 U6825 ( .A1(n4414), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6826 ( .A1(n7854), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6827 ( .A1(n5312), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6828 ( .A1(n5328), .A2(n5313), .ZN(n7176) );
  NAND2_X1 U6829 ( .A1(n5432), .A2(n7176), .ZN(n5315) );
  NAND2_X1 U6830 ( .A1(n5216), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5314) );
  NAND4_X1 U6831 ( .A1(n5317), .A2(n5316), .A3(n5315), .A4(n5314), .ZN(n8277)
         );
  NAND2_X1 U6832 ( .A1(n7181), .A2(n8277), .ZN(n7050) );
  XNOR2_X1 U6833 ( .A(n5319), .B(n5318), .ZN(n6794) );
  NAND2_X1 U6834 ( .A1(n6794), .A2(n8060), .ZN(n5327) );
  NOR2_X1 U6835 ( .A1(n5320), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5324) );
  NOR2_X1 U6836 ( .A1(n5324), .A2(n8725), .ZN(n5321) );
  MUX2_X1 U6837 ( .A(n8725), .B(n5321), .S(P2_IR_REG_11__SCAN_IN), .Z(n5322)
         );
  INV_X1 U6838 ( .A(n5322), .ZN(n5325) );
  INV_X1 U6839 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6840 ( .A1(n5324), .A2(n5323), .ZN(n5351) );
  AOI22_X1 U6841 ( .A1(n8061), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5447), .B2(
        n7334), .ZN(n5326) );
  NAND2_X1 U6842 ( .A1(n4414), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5333) );
  NAND2_X1 U6843 ( .A1(n7854), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U6844 ( .A1(n5328), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6845 ( .A1(n5342), .A2(n5329), .ZN(n7236) );
  NAND2_X1 U6846 ( .A1(n5432), .A2(n7236), .ZN(n5331) );
  NAND2_X1 U6847 ( .A1(n5184), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5330) );
  INV_X1 U6848 ( .A(n7124), .ZN(n8276) );
  NAND2_X1 U6849 ( .A1(n10292), .A2(n8276), .ZN(n5334) );
  AND2_X1 U6850 ( .A1(n7050), .A2(n5334), .ZN(n5336) );
  INV_X1 U6851 ( .A(n5334), .ZN(n5335) );
  OR2_X1 U6852 ( .A1(n10292), .A2(n7124), .ZN(n8140) );
  NAND2_X1 U6853 ( .A1(n10292), .A2(n7124), .ZN(n8141) );
  XNOR2_X1 U6854 ( .A(n5338), .B(n5337), .ZN(n6912) );
  NAND2_X1 U6855 ( .A1(n6912), .A2(n8060), .ZN(n5341) );
  NAND2_X1 U6856 ( .A1(n5351), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5339) );
  XNOR2_X1 U6857 ( .A(n5339), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7344) );
  AOI22_X1 U6858 ( .A1(n8061), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5447), .B2(
        n7344), .ZN(n5340) );
  NAND2_X1 U6859 ( .A1(n4414), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U6860 ( .A1(n7854), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6861 ( .A1(n5342), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6862 ( .A1(n5355), .A2(n5343), .ZN(n7287) );
  NAND2_X1 U6863 ( .A1(n5432), .A2(n7287), .ZN(n5345) );
  NAND2_X1 U6864 ( .A1(n5184), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5344) );
  NAND4_X1 U6865 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n8275)
         );
  AND2_X1 U6866 ( .A1(n10298), .A2(n8275), .ZN(n5348) );
  OAI22_X1 U6867 ( .A1(n7101), .A2(n5348), .B1(n8275), .B2(n10298), .ZN(n7200)
         );
  XNOR2_X1 U6868 ( .A(n5350), .B(n5349), .ZN(n7074) );
  NAND2_X1 U6869 ( .A1(n7074), .A2(n8060), .ZN(n5354) );
  NAND2_X1 U6870 ( .A1(n5352), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5366) );
  XNOR2_X1 U6871 ( .A(n5366), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8327) );
  AOI22_X1 U6872 ( .A1(n8061), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5447), .B2(
        n8327), .ZN(n5353) );
  NAND2_X1 U6873 ( .A1(n7854), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6874 ( .A1(n4414), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5359) );
  NAND2_X1 U6875 ( .A1(n5355), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6876 ( .A1(n5373), .A2(n5356), .ZN(n7202) );
  NAND2_X1 U6877 ( .A1(n5432), .A2(n7202), .ZN(n5358) );
  NAND2_X1 U6878 ( .A1(n5184), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5357) );
  NAND4_X1 U6879 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n8274)
         );
  NAND2_X1 U6880 ( .A1(n8154), .A2(n8274), .ZN(n8155) );
  NAND2_X1 U6881 ( .A1(n7200), .A2(n8047), .ZN(n5361) );
  NAND2_X1 U6882 ( .A1(n5361), .A2(n8158), .ZN(n7257) );
  INV_X1 U6883 ( .A(n7257), .ZN(n5380) );
  XNOR2_X1 U6884 ( .A(n5362), .B(SI_14_), .ZN(n5363) );
  XNOR2_X1 U6885 ( .A(n5364), .B(n5363), .ZN(n7144) );
  NAND2_X1 U6886 ( .A1(n7144), .A2(n8060), .ZN(n5372) );
  INV_X1 U6887 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6888 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  NAND2_X1 U6889 ( .A1(n5367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5369) );
  INV_X1 U6890 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5368) );
  NAND2_X1 U6891 ( .A1(n5369), .A2(n5368), .ZN(n5385) );
  OR2_X1 U6892 ( .A1(n5369), .A2(n5368), .ZN(n5370) );
  NAND2_X1 U6893 ( .A1(n5385), .A2(n5370), .ZN(n8351) );
  INV_X1 U6894 ( .A(n8351), .ZN(n8322) );
  AOI22_X1 U6895 ( .A1(n8061), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5447), .B2(
        n8322), .ZN(n5371) );
  NAND2_X1 U6896 ( .A1(n7854), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6897 ( .A1(n5184), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6898 ( .A1(n5373), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6899 ( .A1(n5389), .A2(n5374), .ZN(n7261) );
  NAND2_X1 U6900 ( .A1(n5432), .A2(n7261), .ZN(n5376) );
  NAND2_X1 U6901 ( .A1(n4414), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6902 ( .A1(n7274), .A2(n7243), .ZN(n8163) );
  INV_X1 U6903 ( .A(n7243), .ZN(n8598) );
  NAND2_X1 U6904 ( .A1(n7274), .A2(n8598), .ZN(n5381) );
  XNOR2_X1 U6905 ( .A(n5382), .B(SI_15_), .ZN(n5383) );
  XNOR2_X1 U6906 ( .A(n5384), .B(n5383), .ZN(n7211) );
  NAND2_X1 U6907 ( .A1(n7211), .A2(n8060), .ZN(n5388) );
  NAND2_X1 U6908 ( .A1(n5385), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5386) );
  XNOR2_X1 U6909 ( .A(n5386), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8373) );
  AOI22_X1 U6910 ( .A1(n8061), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5447), .B2(
        n8373), .ZN(n5387) );
  NAND2_X1 U6911 ( .A1(n4414), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6912 ( .A1(n7854), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U6913 ( .A1(n5389), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6914 ( .A1(n5403), .A2(n5390), .ZN(n8602) );
  NAND2_X1 U6915 ( .A1(n5432), .A2(n8602), .ZN(n5392) );
  NAND2_X1 U6916 ( .A1(n5184), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5391) );
  NAND4_X1 U6917 ( .A1(n5394), .A2(n5393), .A3(n5392), .A4(n5391), .ZN(n8587)
         );
  AND2_X1 U6918 ( .A1(n8718), .A2(n8587), .ZN(n8050) );
  OR2_X1 U6919 ( .A1(n8718), .A2(n8587), .ZN(n8049) );
  NAND2_X1 U6920 ( .A1(n5395), .A2(n8049), .ZN(n8586) );
  XNOR2_X1 U6921 ( .A(n5396), .B(SI_16_), .ZN(n5397) );
  XNOR2_X1 U6922 ( .A(n5398), .B(n5397), .ZN(n7496) );
  NAND2_X1 U6923 ( .A1(n7496), .A2(n8060), .ZN(n5402) );
  NAND2_X1 U6924 ( .A1(n5399), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5400) );
  XNOR2_X1 U6925 ( .A(n5400), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8376) );
  AOI22_X1 U6926 ( .A1(n8061), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5447), .B2(
        n8376), .ZN(n5401) );
  NAND2_X1 U6927 ( .A1(n4414), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5408) );
  NAND2_X1 U6928 ( .A1(n7854), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6929 ( .A1(n5403), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6930 ( .A1(n5415), .A2(n5404), .ZN(n8591) );
  NAND2_X1 U6931 ( .A1(n5432), .A2(n8591), .ZN(n5406) );
  NAND2_X1 U6932 ( .A1(n5184), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6933 ( .A1(n8712), .A2(n7875), .ZN(n8179) );
  INV_X1 U6934 ( .A(n8712), .ZN(n7300) );
  XNOR2_X1 U6935 ( .A(n5410), .B(n5409), .ZN(n7513) );
  NAND2_X1 U6936 ( .A1(n7513), .A2(n8060), .ZN(n5414) );
  NAND2_X1 U6937 ( .A1(n5411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5412) );
  XNOR2_X1 U6938 ( .A(n5412), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8414) );
  AOI22_X1 U6939 ( .A1(n8061), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5447), .B2(
        n8414), .ZN(n5413) );
  NAND2_X1 U6940 ( .A1(n4414), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6941 ( .A1(n7854), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U6942 ( .A1(n5415), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6943 ( .A1(n5430), .A2(n5416), .ZN(n8581) );
  NAND2_X1 U6944 ( .A1(n5432), .A2(n8581), .ZN(n5418) );
  NAND2_X1 U6945 ( .A1(n5184), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5417) );
  NAND2_X1 U6946 ( .A1(n8706), .A2(n8565), .ZN(n8185) );
  NAND2_X1 U6947 ( .A1(n8180), .A2(n8185), .ZN(n8175) );
  INV_X1 U6948 ( .A(n5421), .ZN(n5423) );
  NAND2_X1 U6949 ( .A1(n5423), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6950 ( .A1(n5425), .A2(n5424), .ZN(n7522) );
  NAND2_X1 U6951 ( .A1(n5427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  XNOR2_X1 U6952 ( .A(n5443), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8408) );
  AOI22_X1 U6953 ( .A1(n8061), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5447), .B2(
        n8408), .ZN(n5428) );
  NAND2_X1 U6954 ( .A1(n4414), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U6955 ( .A1(n7854), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6956 ( .A1(n5430), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6957 ( .A1(n5450), .A2(n5431), .ZN(n8567) );
  NAND2_X1 U6958 ( .A1(n5432), .A2(n8567), .ZN(n5434) );
  NAND2_X1 U6959 ( .A1(n5184), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5433) );
  NAND4_X1 U6960 ( .A1(n5436), .A2(n5435), .A3(n5434), .A4(n5433), .ZN(n8578)
         );
  NAND2_X1 U6961 ( .A1(n5437), .A2(n4486), .ZN(n5439) );
  OR2_X1 U6962 ( .A1(n8571), .A2(n8578), .ZN(n5438) );
  XNOR2_X1 U6963 ( .A(n5441), .B(n5440), .ZN(n7525) );
  NAND2_X1 U6964 ( .A1(n7525), .A2(n8060), .ZN(n5449) );
  NAND2_X1 U6965 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  NAND2_X1 U6966 ( .A1(n5444), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5446) );
  AOI22_X1 U6967 ( .A1(n8061), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8409), .B2(
        n5447), .ZN(n5448) );
  NAND2_X1 U6968 ( .A1(n7854), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U6969 ( .A1(n5184), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U6970 ( .A1(n5450), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U6971 ( .A1(n5460), .A2(n5451), .ZN(n8555) );
  NAND2_X1 U6972 ( .A1(n5432), .A2(n8555), .ZN(n5453) );
  NAND2_X1 U6973 ( .A1(n4414), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6974 ( .A1(n8556), .A2(n8566), .ZN(n8192) );
  INV_X1 U6975 ( .A(n8566), .ZN(n8535) );
  XNOR2_X1 U6976 ( .A(n5457), .B(n5456), .ZN(n7542) );
  NAND2_X1 U6977 ( .A1(n7542), .A2(n8060), .ZN(n5459) );
  NAND2_X1 U6978 ( .A1(n8061), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6979 ( .A1(n7854), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U6980 ( .A1(n4414), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6981 ( .A1(n5460), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6982 ( .A1(n5475), .A2(n5461), .ZN(n8539) );
  NAND2_X1 U6983 ( .A1(n5432), .A2(n8539), .ZN(n5463) );
  NAND2_X1 U6984 ( .A1(n5184), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U6985 ( .A1(n8632), .A2(n7946), .ZN(n8520) );
  NAND2_X1 U6986 ( .A1(n8196), .A2(n8520), .ZN(n8533) );
  NAND2_X1 U6987 ( .A1(n8532), .A2(n5467), .ZN(n8524) );
  XNOR2_X1 U6988 ( .A(n5468), .B(SI_21_), .ZN(n5469) );
  XNOR2_X1 U6989 ( .A(n5470), .B(n5469), .ZN(n7558) );
  NAND2_X1 U6990 ( .A1(n7558), .A2(n8060), .ZN(n5472) );
  NAND2_X1 U6991 ( .A1(n8061), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6992 ( .A1(n7854), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6993 ( .A1(n5184), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5473) );
  AND2_X1 U6994 ( .A1(n5474), .A2(n5473), .ZN(n5479) );
  NAND2_X1 U6995 ( .A1(n5475), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6996 ( .A1(n5485), .A2(n5476), .ZN(n8528) );
  NAND2_X1 U6997 ( .A1(n8528), .A2(n5432), .ZN(n5478) );
  NAND2_X1 U6998 ( .A1(n4414), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6999 ( .A1(n8687), .A2(n8510), .ZN(n8197) );
  NAND2_X1 U7000 ( .A1(n8199), .A2(n8197), .ZN(n8523) );
  INV_X1 U7001 ( .A(n8687), .ZN(n7950) );
  XNOR2_X1 U7002 ( .A(n5482), .B(n5481), .ZN(n7570) );
  NAND2_X1 U7003 ( .A1(n7570), .A2(n8060), .ZN(n5484) );
  NAND2_X1 U7004 ( .A1(n8061), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5483) );
  INV_X1 U7005 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U7006 ( .A1(n5485), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U7007 ( .A1(n5487), .A2(n5486), .ZN(n8514) );
  NAND2_X1 U7008 ( .A1(n8514), .A2(n5432), .ZN(n5489) );
  AOI22_X1 U7009 ( .A1(n4414), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n7854), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5488) );
  INV_X1 U7010 ( .A(n8525), .ZN(n8500) );
  INV_X1 U7011 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7012 ( .A1(n5494), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7013 ( .A1(n5521), .A2(n5495), .ZN(n8488) );
  NAND2_X1 U7014 ( .A1(n8488), .A2(n5432), .ZN(n5500) );
  INV_X1 U7015 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8828) );
  NAND2_X1 U7016 ( .A1(n4414), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7017 ( .A1(n7854), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5496) );
  OAI211_X1 U7018 ( .C1(n8828), .C2(n7857), .A(n5497), .B(n5496), .ZN(n5498)
         );
  INV_X1 U7019 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7020 ( .A1(n5502), .A2(n5501), .ZN(n5504) );
  MUX2_X1 U7021 ( .A(n8865), .B(n7599), .S(n5534), .Z(n5505) );
  INV_X1 U7022 ( .A(SI_24_), .ZN(n8953) );
  NAND2_X1 U7023 ( .A1(n5505), .A2(n8953), .ZN(n5513) );
  INV_X1 U7024 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U7025 ( .A1(n5506), .A2(SI_24_), .ZN(n5507) );
  NAND2_X1 U7026 ( .A1(n8061), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7027 ( .A1(n5510), .A2(n5509), .ZN(n8473) );
  INV_X1 U7028 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7185) );
  INV_X1 U7029 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8981) );
  MUX2_X1 U7030 ( .A(n7185), .B(n8981), .S(n5534), .Z(n5515) );
  INV_X1 U7031 ( .A(SI_25_), .ZN(n5514) );
  NAND2_X1 U7032 ( .A1(n5515), .A2(n5514), .ZN(n5532) );
  INV_X1 U7033 ( .A(n5515), .ZN(n5516) );
  NAND2_X1 U7034 ( .A1(n5516), .A2(SI_25_), .ZN(n5517) );
  NAND2_X1 U7035 ( .A1(n7435), .A2(n8060), .ZN(n5519) );
  NAND2_X1 U7036 ( .A1(n8061), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5518) );
  INV_X1 U7037 ( .A(n5521), .ZN(n5520) );
  INV_X1 U7038 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U7039 ( .A1(n5521), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7040 ( .A1(n5540), .A2(n5522), .ZN(n8479) );
  NAND2_X1 U7041 ( .A1(n8479), .A2(n5432), .ZN(n5527) );
  INV_X1 U7042 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8803) );
  NAND2_X1 U7043 ( .A1(n4414), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5524) );
  NAND2_X1 U7044 ( .A1(n7854), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5523) );
  OAI211_X1 U7045 ( .C1(n8803), .C2(n7857), .A(n5524), .B(n5523), .ZN(n5525)
         );
  INV_X1 U7046 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7047 ( .A1(n8667), .A2(n8486), .ZN(n8225) );
  INV_X1 U7048 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7425) );
  MUX2_X1 U7049 ( .A(n8871), .B(n7425), .S(n5534), .Z(n5535) );
  INV_X1 U7050 ( .A(SI_26_), .ZN(n8944) );
  NAND2_X1 U7051 ( .A1(n5535), .A2(n8944), .ZN(n5551) );
  INV_X1 U7052 ( .A(n5535), .ZN(n5536) );
  NAND2_X1 U7053 ( .A1(n5536), .A2(SI_26_), .ZN(n5537) );
  NAND2_X1 U7054 ( .A1(n7424), .A2(n8060), .ZN(n5539) );
  NAND2_X1 U7055 ( .A1(n8061), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5538) );
  OR2_X2 U7056 ( .A1(n5540), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7057 ( .A1(n5540), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7058 ( .A1(n5561), .A2(n5541), .ZN(n8466) );
  NAND2_X1 U7059 ( .A1(n8466), .A2(n5432), .ZN(n5546) );
  INV_X1 U7060 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U7061 ( .A1(n4414), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U7062 ( .A1(n7854), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5542) );
  OAI211_X1 U7063 ( .C1(n8663), .C2(n7857), .A(n5543), .B(n5542), .ZN(n5544)
         );
  INV_X1 U7064 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U7065 ( .A1(n8012), .A2(n8475), .ZN(n5547) );
  INV_X1 U7066 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5553) );
  INV_X1 U7067 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U7068 ( .A(n5553), .B(n7776), .S(n5534), .Z(n5555) );
  INV_X1 U7069 ( .A(SI_27_), .ZN(n5554) );
  NAND2_X1 U7070 ( .A1(n5555), .A2(n5554), .ZN(n5572) );
  INV_X1 U7071 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7072 ( .A1(n5556), .A2(SI_27_), .ZN(n5557) );
  NAND2_X1 U7073 ( .A1(n7421), .A2(n8060), .ZN(n5559) );
  NAND2_X1 U7074 ( .A1(n8061), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5558) );
  INV_X1 U7075 ( .A(n5561), .ZN(n5560) );
  INV_X1 U7076 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U7077 ( .A1(n5560), .A2(n8853), .ZN(n5575) );
  NAND2_X1 U7078 ( .A1(n5561), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U7079 ( .A1(n5575), .A2(n5562), .ZN(n8458) );
  NAND2_X1 U7080 ( .A1(n8458), .A2(n5432), .ZN(n5567) );
  INV_X1 U7081 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U7082 ( .A1(n4414), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7083 ( .A1(n7854), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5563) );
  OAI211_X1 U7084 ( .C1(n8657), .C2(n7857), .A(n5564), .B(n5563), .ZN(n5565)
         );
  INV_X1 U7085 ( .A(n5565), .ZN(n5566) );
  NOR2_X1 U7086 ( .A1(n7912), .A2(n8463), .ZN(n5569) );
  MUX2_X1 U7087 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n5534), .Z(n7383) );
  INV_X1 U7088 ( .A(SI_28_), .ZN(n7384) );
  XNOR2_X1 U7089 ( .A(n7383), .B(n7384), .ZN(n7381) );
  NAND2_X1 U7090 ( .A1(n7412), .A2(n8060), .ZN(n5574) );
  NAND2_X1 U7091 ( .A1(n8061), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7092 ( .A1(n5575), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7093 ( .A1(n8440), .A2(n5576), .ZN(n7935) );
  NAND2_X1 U7094 ( .A1(n7935), .A2(n5432), .ZN(n5582) );
  INV_X1 U7095 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7096 ( .A1(n4414), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7097 ( .A1(n7854), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5577) );
  OAI211_X1 U7098 ( .C1(n5579), .C2(n7857), .A(n5578), .B(n5577), .ZN(n5580)
         );
  INV_X1 U7099 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7100 ( .A1(n4430), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7101 ( .A1(n8264), .A2(n8409), .ZN(n5654) );
  NAND2_X1 U7102 ( .A1(n4447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5585) );
  MUX2_X1 U7103 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5585), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5586) );
  NAND2_X1 U7104 ( .A1(n5587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5589) );
  INV_X1 U7105 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5588) );
  INV_X1 U7106 ( .A(n8260), .ZN(n5672) );
  NAND2_X1 U7107 ( .A1(n8076), .A2(n5672), .ZN(n6147) );
  INV_X1 U7108 ( .A(n8440), .ZN(n5590) );
  NAND2_X1 U7109 ( .A1(n5590), .A2(n5432), .ZN(n8032) );
  INV_X1 U7110 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7866) );
  NAND2_X1 U7111 ( .A1(n4414), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7112 ( .A1(n7854), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7113 ( .C1(n7866), .C2(n7857), .A(n5592), .B(n5591), .ZN(n5593)
         );
  INV_X1 U7114 ( .A(n5593), .ZN(n5594) );
  OR2_X1 U7115 ( .A1(n7938), .A2(n8256), .ZN(n8074) );
  INV_X1 U7116 ( .A(n5877), .ZN(n5891) );
  INV_X4 U7117 ( .A(n7294), .ZN(n8426) );
  NAND2_X1 U7118 ( .A1(n5891), .A2(n8426), .ZN(n8262) );
  NAND2_X1 U7119 ( .A1(n5877), .A2(n7294), .ZN(n5882) );
  INV_X1 U7120 ( .A(n6142), .ZN(n5597) );
  OAI22_X1 U7121 ( .A1(n8074), .A2(n5597), .B1(n8463), .B2(n10220), .ZN(n5598)
         );
  INV_X1 U7122 ( .A(n8286), .ZN(n6145) );
  NAND2_X1 U7123 ( .A1(n6145), .A2(n6172), .ZN(n8078) );
  NAND2_X1 U7124 ( .A1(n6193), .A2(n5601), .ZN(n10216) );
  INV_X1 U7125 ( .A(n8036), .ZN(n10224) );
  NAND2_X1 U7126 ( .A1(n10216), .A2(n10224), .ZN(n5602) );
  NAND2_X1 U7127 ( .A1(n5602), .A2(n8090), .ZN(n10209) );
  XNOR2_X1 U7128 ( .A(n8283), .B(n10243), .ZN(n10208) );
  NAND2_X1 U7129 ( .A1(n10209), .A2(n10208), .ZN(n5603) );
  NAND2_X1 U7130 ( .A1(n10222), .A2(n10243), .ZN(n8098) );
  NAND2_X1 U7131 ( .A1(n5603), .A2(n8098), .ZN(n6541) );
  XNOR2_X1 U7132 ( .A(n10203), .B(n10249), .ZN(n8096) );
  NAND2_X1 U7133 ( .A1(n6541), .A2(n8096), .ZN(n5604) );
  INV_X1 U7134 ( .A(n10203), .ZN(n6474) );
  NAND2_X1 U7135 ( .A1(n6474), .A2(n10249), .ZN(n8105) );
  NAND2_X1 U7136 ( .A1(n5604), .A2(n8105), .ZN(n6677) );
  NAND2_X1 U7137 ( .A1(n8282), .A2(n6573), .ZN(n8108) );
  NAND2_X1 U7138 ( .A1(n6677), .A2(n8108), .ZN(n6688) );
  NAND2_X1 U7139 ( .A1(n6824), .A2(n10260), .ZN(n8112) );
  NAND2_X1 U7140 ( .A1(n6575), .A2(n10254), .ZN(n8110) );
  AND2_X1 U7141 ( .A1(n8112), .A2(n8110), .ZN(n8102) );
  NAND2_X1 U7142 ( .A1(n6688), .A2(n8102), .ZN(n5605) );
  NAND2_X1 U7143 ( .A1(n8281), .A2(n6690), .ZN(n8114) );
  AND2_X1 U7144 ( .A1(n8118), .A2(n6901), .ZN(n8130) );
  NAND2_X1 U7145 ( .A1(n7179), .A2(n7062), .ZN(n8127) );
  NAND2_X1 U7146 ( .A1(n8278), .A2(n10277), .ZN(n8119) );
  NAND2_X1 U7147 ( .A1(n8127), .A2(n8119), .ZN(n6892) );
  OR2_X2 U7148 ( .A1(n6890), .A2(n6892), .ZN(n6942) );
  OR2_X1 U7149 ( .A1(n7114), .A2(n7181), .ZN(n8139) );
  AND2_X1 U7150 ( .A1(n8139), .A2(n8119), .ZN(n8129) );
  NAND2_X1 U7151 ( .A1(n7181), .A2(n7114), .ZN(n8136) );
  INV_X1 U7152 ( .A(n8134), .ZN(n8045) );
  XNOR2_X1 U7153 ( .A(n10298), .B(n8148), .ZN(n8152) );
  OR2_X1 U7154 ( .A1(n10298), .A2(n8148), .ZN(n8150) );
  NAND2_X1 U7155 ( .A1(n7100), .A2(n8150), .ZN(n7203) );
  NAND2_X1 U7156 ( .A1(n8154), .A2(n7290), .ZN(n5607) );
  NAND2_X1 U7157 ( .A1(n7203), .A2(n5607), .ZN(n5609) );
  OR2_X1 U7158 ( .A1(n8154), .A2(n7290), .ZN(n5608) );
  NAND2_X1 U7159 ( .A1(n5609), .A2(n5608), .ZN(n7264) );
  NAND2_X1 U7160 ( .A1(n7264), .A2(n8163), .ZN(n5610) );
  NAND2_X1 U7161 ( .A1(n5610), .A2(n8171), .ZN(n8594) );
  INV_X1 U7162 ( .A(n8587), .ZN(n7245) );
  NAND2_X1 U7163 ( .A1(n8718), .A2(n7245), .ZN(n8170) );
  NAND2_X1 U7164 ( .A1(n8594), .A2(n8170), .ZN(n5611) );
  OR2_X1 U7165 ( .A1(n8718), .A2(n7245), .ZN(n8167) );
  NAND2_X1 U7166 ( .A1(n5611), .A2(n8167), .ZN(n8584) );
  NAND2_X1 U7167 ( .A1(n5612), .A2(n8185), .ZN(n8559) );
  NAND2_X1 U7168 ( .A1(n8571), .A2(n7967), .ZN(n8191) );
  NAND2_X1 U7169 ( .A1(n8186), .A2(n8191), .ZN(n8563) );
  NAND2_X1 U7170 ( .A1(n8531), .A2(n8196), .ZN(n8521) );
  AND2_X1 U7171 ( .A1(n8197), .A2(n8520), .ZN(n8200) );
  NAND2_X1 U7172 ( .A1(n8521), .A2(n8200), .ZN(n5616) );
  INV_X1 U7173 ( .A(n8206), .ZN(n8207) );
  INV_X1 U7174 ( .A(n8202), .ZN(n5617) );
  NAND2_X1 U7175 ( .A1(n5618), .A2(n8501), .ZN(n8215) );
  NAND2_X1 U7176 ( .A1(n8505), .A2(n8511), .ZN(n8489) );
  AND2_X1 U7177 ( .A1(n8215), .A2(n8489), .ZN(n8219) );
  NAND2_X1 U7178 ( .A1(n5619), .A2(n8217), .ZN(n8480) );
  NAND2_X1 U7179 ( .A1(n8658), .A2(n8463), .ZN(n8033) );
  NAND2_X1 U7180 ( .A1(n5620), .A2(n8058), .ZN(n7852) );
  OAI21_X1 U7181 ( .B1(n5620), .B2(n8058), .A(n7852), .ZN(n7773) );
  INV_X1 U7182 ( .A(n7773), .ZN(n5623) );
  AND2_X1 U7183 ( .A1(n8431), .A2(n8260), .ZN(n5666) );
  INV_X1 U7184 ( .A(n5666), .ZN(n5621) );
  INV_X1 U7185 ( .A(n8264), .ZN(n6940) );
  AOI21_X1 U7186 ( .B1(n6940), .B2(n5672), .A(n8409), .ZN(n5622) );
  NAND2_X1 U7187 ( .A1(n6940), .A2(n6194), .ZN(n10284) );
  INV_X1 U7188 ( .A(n10284), .ZN(n10255) );
  NAND2_X1 U7189 ( .A1(n7775), .A2(n5009), .ZN(n5680) );
  NAND2_X1 U7190 ( .A1(n5653), .A2(n5652), .ZN(n5624) );
  XNOR2_X1 U7191 ( .A(n7143), .B(P2_B_REG_SCAN_IN), .ZN(n5631) );
  NAND2_X1 U7192 ( .A1(n7187), .A2(n5631), .ZN(n5635) );
  NAND2_X1 U7193 ( .A1(n4467), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5632) );
  MUX2_X1 U7194 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5632), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5633) );
  NAND2_X1 U7195 ( .A1(n7187), .A2(n7280), .ZN(n5636) );
  NOR2_X1 U7196 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n5641) );
  NOR4_X1 U7197 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5640) );
  NOR4_X1 U7198 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_16__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5639) );
  NOR4_X1 U7199 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n5638) );
  NAND4_X1 U7200 ( .A1(n5641), .A2(n5640), .A3(n5639), .A4(n5638), .ZN(n5647)
         );
  NOR4_X1 U7201 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5645) );
  NOR4_X1 U7202 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n5644) );
  NOR4_X1 U7203 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5643) );
  NOR4_X1 U7204 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5642) );
  NAND4_X1 U7205 ( .A1(n5645), .A2(n5644), .A3(n5643), .A4(n5642), .ZN(n5646)
         );
  NOR2_X1 U7206 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  INV_X1 U7207 ( .A(n5669), .ZN(n5655) );
  NOR2_X1 U7208 ( .A1(n6162), .A2(n5655), .ZN(n5650) );
  NAND2_X1 U7209 ( .A1(n7143), .A2(n7280), .ZN(n5851) );
  INV_X1 U7210 ( .A(n4497), .ZN(n5674) );
  NOR2_X1 U7211 ( .A1(n7143), .A2(n7280), .ZN(n5651) );
  OR2_X1 U7212 ( .A1(n5654), .A2(n8260), .ZN(n5657) );
  NAND3_X1 U7213 ( .A1(n10282), .A2(n8256), .A3(n5657), .ZN(n6053) );
  INV_X1 U7214 ( .A(n6194), .ZN(n6148) );
  NAND2_X1 U7215 ( .A1(n10299), .A2(n6148), .ZN(n10218) );
  NAND2_X1 U7216 ( .A1(n6053), .A2(n10218), .ZN(n6043) );
  NAND2_X1 U7217 ( .A1(n6144), .A2(n6043), .ZN(n5661) );
  NAND2_X1 U7218 ( .A1(n6162), .A2(n4497), .ZN(n5671) );
  OR2_X1 U7219 ( .A1(n5671), .A2(n5655), .ZN(n6044) );
  INV_X1 U7220 ( .A(n6059), .ZN(n5656) );
  INV_X1 U7221 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7222 ( .A1(n5658), .A2(n6939), .ZN(n6051) );
  NAND2_X1 U7223 ( .A1(n6051), .A2(n6141), .ZN(n5659) );
  NAND2_X1 U7224 ( .A1(n6057), .A2(n5659), .ZN(n5660) );
  NAND2_X1 U7225 ( .A1(n8239), .A2(n5662), .ZN(n5664) );
  NAND2_X1 U7226 ( .A1(n10302), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5663) );
  OAI21_X1 U7227 ( .B1(n8256), .B2(n5666), .A(n5880), .ZN(n5667) );
  INV_X1 U7228 ( .A(n5667), .ZN(n5668) );
  AND2_X1 U7229 ( .A1(n5879), .A2(n5668), .ZN(n6046) );
  AND2_X1 U7230 ( .A1(n10299), .A2(n6194), .ZN(n6058) );
  NAND3_X1 U7231 ( .A1(n8264), .A2(n5672), .A3(n8431), .ZN(n5673) );
  AND2_X1 U7232 ( .A1(n8256), .A2(n5673), .ZN(n6161) );
  OAI21_X1 U7233 ( .B1(n5674), .B2(n6058), .A(n6161), .ZN(n5678) );
  INV_X1 U7234 ( .A(n6162), .ZN(n5676) );
  INV_X1 U7235 ( .A(n6161), .ZN(n5675) );
  NAND2_X1 U7236 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  NAND2_X1 U7237 ( .A1(n5680), .A2(n10325), .ZN(n5683) );
  INV_X1 U7238 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5681) );
  OR2_X1 U7239 ( .A1(n10325), .A2(n5681), .ZN(n5682) );
  NAND2_X1 U7240 ( .A1(n5024), .A2(n5684), .ZN(P2_U3487) );
  NAND2_X1 U7241 ( .A1(n5687), .A2(n5686), .ZN(n5859) );
  NOR2_X1 U7242 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5691) );
  NAND4_X1 U7243 ( .A1(n5691), .A2(n5690), .A3(n5689), .A4(n5688), .ZN(n5692)
         );
  INV_X1 U7244 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5693) );
  NAND3_X1 U7245 ( .A1(n5750), .A2(n5752), .A3(n5694), .ZN(n5695) );
  NAND2_X1 U7246 ( .A1(n5745), .A2(n5710), .ZN(n5697) );
  NAND4_X1 U7247 ( .A1(n5699), .A2(n5745), .A3(n5693), .A4(n5750), .ZN(n5702)
         );
  NAND4_X1 U7248 ( .A1(n5710), .A2(n5730), .A3(n5752), .A4(n5700), .ZN(n5701)
         );
  NAND2_X1 U7249 ( .A1(n5716), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7250 ( .A1(n5706), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5707) );
  MUX2_X1 U7251 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5707), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5708) );
  NAND2_X1 U7252 ( .A1(n5708), .A2(n5716), .ZN(n7184) );
  OR3_X2 U7253 ( .A1(n5902), .A2(n7255), .A3(n7184), .ZN(n5918) );
  NOR2_X1 U7254 ( .A1(n5918), .A2(P1_U3086), .ZN(n5712) );
  NAND2_X1 U7255 ( .A1(n5709), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7256 ( .A1(n5746), .A2(n5745), .ZN(n5748) );
  NAND2_X1 U7257 ( .A1(n5748), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7258 ( .A1(n5879), .A2(n8256), .ZN(n5713) );
  NAND2_X1 U7259 ( .A1(n5713), .A2(n5880), .ZN(n5714) );
  NAND2_X1 U7260 ( .A1(n5714), .A2(n5181), .ZN(n5715) );
  NAND2_X1 U7261 ( .A1(n5715), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7262 ( .A(n5853), .ZN(n5855) );
  INV_X1 U7263 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9945) );
  OR2_X1 U7264 ( .A1(n7440), .A2(n9945), .ZN(n5724) );
  INV_X1 U7265 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5720) );
  INV_X1 U7266 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5935) );
  OR2_X1 U7267 ( .A1(n7534), .A2(n5935), .ZN(n5722) );
  INV_X1 U7268 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5726) );
  INV_X1 U7269 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7270 ( .A1(n5732), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  MUX2_X1 U7271 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5733), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5735) );
  INV_X1 U7272 ( .A(n6326), .ZN(n5736) );
  AND2_X2 U7273 ( .A1(n5918), .A2(n5736), .ZN(n6752) );
  NAND2_X1 U7274 ( .A1(n6231), .A2(n6752), .ZN(n5761) );
  NAND2_X1 U7275 ( .A1(n5534), .A2(SI_0_), .ZN(n5738) );
  INV_X1 U7276 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7277 ( .A1(n5738), .A2(n5737), .ZN(n5740) );
  NAND2_X1 U7278 ( .A1(n5740), .A2(n5739), .ZN(n9873) );
  MUX2_X1 U7279 ( .A(n4675), .B(n9873), .S(n6253), .Z(n10061) );
  INV_X1 U7280 ( .A(n10061), .ZN(n6230) );
  NAND2_X1 U7281 ( .A1(n6485), .A2(n5750), .ZN(n5751) );
  NAND2_X1 U7282 ( .A1(n6642), .A2(n5752), .ZN(n5753) );
  AND2_X1 U7283 ( .A1(n5756), .A2(n6326), .ZN(n5755) );
  INV_X1 U7284 ( .A(n7835), .ZN(n5757) );
  NAND2_X1 U7285 ( .A1(n7684), .A2(n6326), .ZN(n5758) );
  NAND2_X1 U7286 ( .A1(n6230), .A2(n4417), .ZN(n5760) );
  OR2_X1 U7287 ( .A1(n5918), .A2(n9945), .ZN(n5762) );
  NAND2_X1 U7288 ( .A1(n5936), .A2(n5762), .ZN(n5767) );
  INV_X2 U7289 ( .A(n9201), .ZN(n9081) );
  NAND2_X1 U7290 ( .A1(n6231), .A2(n9081), .ZN(n5765) );
  OAI22_X1 U7291 ( .A1(n10061), .A2(n6076), .B1(n5918), .B2(n4675), .ZN(n5763)
         );
  INV_X1 U7292 ( .A(n5763), .ZN(n5764) );
  NAND2_X1 U7293 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NOR2_X1 U7294 ( .A1(n5767), .A2(n5766), .ZN(n5768) );
  NOR2_X1 U7295 ( .A1(n5937), .A2(n5768), .ZN(n5931) );
  INV_X1 U7296 ( .A(n7769), .ZN(n5946) );
  NAND2_X1 U7297 ( .A1(n5946), .A2(n4416), .ZN(n5771) );
  OAI21_X1 U7298 ( .B1(n4416), .B2(P1_REG2_REG_0__SCAN_IN), .A(n5946), .ZN(
        n9944) );
  INV_X1 U7299 ( .A(n4416), .ZN(n5769) );
  AND2_X1 U7300 ( .A1(n5946), .A2(n5769), .ZN(n7763) );
  AND2_X1 U7301 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9405) );
  AOI22_X1 U7302 ( .A1(n9944), .A2(n4675), .B1(n7763), .B2(n9405), .ZN(n5770)
         );
  OAI211_X1 U7303 ( .C1(n5931), .C2(n5771), .A(P1_U3973), .B(n5770), .ZN(n9425) );
  INV_X1 U7304 ( .A(n9425), .ZN(n5814) );
  INV_X1 U7305 ( .A(n5774), .ZN(n5772) );
  NAND2_X1 U7306 ( .A1(n5772), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7768) );
  INV_X1 U7307 ( .A(n7768), .ZN(n5773) );
  OR2_X1 U7308 ( .A1(n9853), .A2(n5773), .ZN(n5778) );
  NAND2_X1 U7309 ( .A1(n5774), .A2(n7752), .ZN(n5775) );
  AND2_X1 U7310 ( .A1(n5775), .A2(n6253), .ZN(n5777) );
  INV_X1 U7311 ( .A(n5777), .ZN(n5776) );
  AND2_X1 U7312 ( .A1(n5778), .A2(n5776), .ZN(n9948) );
  INV_X1 U7313 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7314 ( .A1(n5778), .A2(n5777), .ZN(n9950) );
  NOR2_X2 U7315 ( .A1(n9950), .A2(n5946), .ZN(n10031) );
  OR2_X1 U7316 ( .A1(n5797), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n5780) );
  NOR2_X1 U7317 ( .A1(n5780), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5822) );
  INV_X1 U7318 ( .A(n5822), .ZN(n5783) );
  NAND2_X1 U7319 ( .A1(n5780), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5781) );
  MUX2_X1 U7320 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5781), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5782) );
  NAND2_X1 U7321 ( .A1(n5783), .A2(n5782), .ZN(n6115) );
  INV_X1 U7322 ( .A(n6115), .ZN(n5968) );
  NAND2_X1 U7323 ( .A1(n10031), .A2(n5968), .ZN(n5784) );
  NAND2_X1 U7324 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n6132) );
  OAI211_X1 U7325 ( .C1(n10039), .C2(n5785), .A(n5784), .B(n6132), .ZN(n5813)
         );
  INV_X1 U7326 ( .A(n9950), .ZN(n5786) );
  NAND2_X1 U7327 ( .A1(n5786), .A2(n4416), .ZN(n10028) );
  INV_X1 U7328 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5787) );
  MUX2_X1 U7329 ( .A(n5787), .B(P1_REG1_REG_4__SCAN_IN), .S(n6115), .Z(n5802)
         );
  INV_X1 U7330 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5792) );
  NOR2_X1 U7331 ( .A1(n5788), .A2(n5864), .ZN(n5789) );
  MUX2_X1 U7332 ( .A(n5864), .B(n5789), .S(P1_IR_REG_2__SCAN_IN), .Z(n5790) );
  INV_X1 U7333 ( .A(n5790), .ZN(n5791) );
  NAND2_X1 U7334 ( .A1(n5791), .A2(n5797), .ZN(n9411) );
  MUX2_X1 U7335 ( .A(n5792), .B(P1_REG1_REG_2__SCAN_IN), .S(n9411), .Z(n9418)
         );
  NAND2_X1 U7336 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5793) );
  MUX2_X1 U7337 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5793), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5795) );
  INV_X1 U7338 ( .A(n5788), .ZN(n5794) );
  NAND2_X1 U7339 ( .A1(n5795), .A2(n5794), .ZN(n5941) );
  INV_X1 U7340 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10101) );
  MUX2_X1 U7341 ( .A(n10101), .B(P1_REG1_REG_1__SCAN_IN), .S(n5941), .Z(n9402)
         );
  AND2_X1 U7342 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9401) );
  NAND2_X1 U7343 ( .A1(n9402), .A2(n9401), .ZN(n9400) );
  OAI21_X1 U7344 ( .B1(n10101), .B2(n5941), .A(n9400), .ZN(n9417) );
  NAND2_X1 U7345 ( .A1(n9418), .A2(n9417), .ZN(n9416) );
  OR2_X1 U7346 ( .A1(n9411), .A2(n5792), .ZN(n5796) );
  NAND2_X1 U7347 ( .A1(n9416), .A2(n5796), .ZN(n9432) );
  NAND2_X1 U7348 ( .A1(n5797), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  INV_X1 U7349 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U7350 ( .A(n5799), .B(n5798), .ZN(n9426) );
  XNOR2_X1 U7351 ( .A(n9426), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U7352 ( .A1(n9432), .A2(n9433), .ZN(n9431) );
  INV_X1 U7353 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6000) );
  OR2_X1 U7354 ( .A1(n9426), .A2(n6000), .ZN(n5800) );
  NAND2_X1 U7355 ( .A1(n9431), .A2(n5800), .ZN(n5801) );
  NAND2_X1 U7356 ( .A1(n5801), .A2(n5802), .ZN(n5970) );
  OAI21_X1 U7357 ( .B1(n5802), .B2(n5801), .A(n5970), .ZN(n5811) );
  MUX2_X1 U7358 ( .A(n10044), .B(P1_REG2_REG_4__SCAN_IN), .S(n6115), .Z(n5809)
         );
  INV_X1 U7359 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5803) );
  MUX2_X1 U7360 ( .A(n5803), .B(P1_REG2_REG_2__SCAN_IN), .S(n9411), .Z(n9421)
         );
  INV_X1 U7361 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U7362 ( .A(n8866), .B(P1_REG2_REG_1__SCAN_IN), .S(n5941), .Z(n9406)
         );
  NAND2_X1 U7363 ( .A1(n9406), .A2(n9405), .ZN(n9404) );
  INV_X1 U7364 ( .A(n5941), .ZN(n9403) );
  NAND2_X1 U7365 ( .A1(n9403), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7366 ( .A1(n9404), .A2(n5804), .ZN(n9420) );
  NAND2_X1 U7367 ( .A1(n9421), .A2(n9420), .ZN(n9419) );
  OR2_X1 U7368 ( .A1(n9411), .A2(n5803), .ZN(n5805) );
  NAND2_X1 U7369 ( .A1(n9419), .A2(n5805), .ZN(n9435) );
  XNOR2_X1 U7370 ( .A(n9426), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U7371 ( .A1(n9435), .A2(n9436), .ZN(n9434) );
  INV_X1 U7372 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6341) );
  OR2_X1 U7373 ( .A1(n9426), .A2(n6341), .ZN(n5806) );
  NAND2_X1 U7374 ( .A1(n9434), .A2(n5806), .ZN(n5808) );
  INV_X1 U7375 ( .A(n7763), .ZN(n5807) );
  NOR2_X2 U7376 ( .A1(n9950), .A2(n5807), .ZN(n10024) );
  NAND2_X1 U7377 ( .A1(n5808), .A2(n5809), .ZN(n5958) );
  OAI211_X1 U7378 ( .C1(n5809), .C2(n5808), .A(n10024), .B(n5958), .ZN(n5810)
         );
  OAI21_X1 U7379 ( .B1(n10028), .B2(n5811), .A(n5810), .ZN(n5812) );
  OR3_X1 U7380 ( .A1(n5814), .A2(n5813), .A3(n5812), .ZN(P1_U3247) );
  AND2_X1 U7381 ( .A1(n5534), .A2(P2_U3151), .ZN(n9020) );
  INV_X1 U7382 ( .A(n9020), .ZN(n7278) );
  AND2_X1 U7383 ( .A1(n5939), .A2(P2_U3151), .ZN(n9022) );
  INV_X2 U7384 ( .A(n9022), .ZN(n8733) );
  INV_X1 U7385 ( .A(n6375), .ZN(n10116) );
  OAI222_X1 U7386 ( .A1(n7278), .A2(n5815), .B1(n8733), .B2(n5992), .C1(
        P2_U3151), .C2(n10116), .ZN(P2_U3293) );
  AND2_X1 U7387 ( .A1(n5534), .A2(P1_U3086), .ZN(n6978) );
  INV_X2 U7388 ( .A(n6978), .ZN(n9872) );
  OAI222_X1 U7389 ( .A1(n9868), .A2(n5940), .B1(n9872), .B2(n5938), .C1(
        P1_U3086), .C2(n5941), .ZN(P1_U3354) );
  OAI222_X1 U7390 ( .A1(n6356), .A2(P2_U3151), .B1(n8733), .B2(n5938), .C1(
        n5816), .C2(n7278), .ZN(P2_U3294) );
  INV_X1 U7391 ( .A(n6376), .ZN(n10140) );
  OAI222_X1 U7392 ( .A1(n7278), .A2(n5817), .B1(n8733), .B2(n6068), .C1(
        P2_U3151), .C2(n10140), .ZN(P2_U3292) );
  OAI222_X1 U7393 ( .A1(n7278), .A2(n5818), .B1(n8733), .B2(n6114), .C1(
        P2_U3151), .C2(n6655), .ZN(P2_U3291) );
  OAI222_X1 U7394 ( .A1(n9868), .A2(n6116), .B1(n9872), .B2(n6114), .C1(
        P1_U3086), .C2(n6115), .ZN(P1_U3351) );
  OAI222_X1 U7395 ( .A1(n9868), .A2(n6069), .B1(n9872), .B2(n6068), .C1(
        P1_U3086), .C2(n9426), .ZN(P1_U3352) );
  OAI222_X1 U7396 ( .A1(n9868), .A2(n5991), .B1(n9872), .B2(n5992), .C1(
        P1_U3086), .C2(n9411), .ZN(P1_U3353) );
  INV_X1 U7397 ( .A(n6252), .ZN(n5827) );
  OR2_X1 U7398 ( .A1(n5822), .A2(n5864), .ZN(n5819) );
  XNOR2_X1 U7399 ( .A(n5819), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9443) );
  INV_X1 U7400 ( .A(n9868), .ZN(n6486) );
  AOI22_X1 U7401 ( .A1(n9443), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n6486), .ZN(n5820) );
  OAI21_X1 U7402 ( .B1(n5827), .B2(n9872), .A(n5820), .ZN(P1_U3350) );
  NOR2_X1 U7403 ( .A1(n9948), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U7404 ( .A1(n5822), .A2(n5821), .ZN(n5844) );
  NAND2_X1 U7405 ( .A1(n5844), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U7406 ( .A1(n5829), .A2(n5823), .ZN(n5824) );
  NAND2_X1 U7407 ( .A1(n5824), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5825) );
  XNOR2_X1 U7408 ( .A(n5825), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U7409 ( .A1(n9469), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n6486), .ZN(n5826) );
  OAI21_X1 U7410 ( .B1(n6437), .B2(n9872), .A(n5826), .ZN(P1_U3348) );
  INV_X1 U7411 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5828) );
  OAI222_X1 U7412 ( .A1(n7278), .A2(n5828), .B1(n8733), .B2(n5827), .C1(
        P2_U3151), .C2(n6847), .ZN(P2_U3290) );
  INV_X1 U7413 ( .A(n6301), .ZN(n5832) );
  XNOR2_X1 U7414 ( .A(n5829), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9456) );
  AOI22_X1 U7415 ( .A1(n9456), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n6486), .ZN(n5830) );
  OAI21_X1 U7416 ( .B1(n5832), .B2(n9872), .A(n5830), .ZN(P1_U3349) );
  INV_X1 U7417 ( .A(n6996), .ZN(n6988) );
  OAI222_X1 U7418 ( .A1(n7278), .A2(n5831), .B1(n8733), .B2(n6437), .C1(
        P2_U3151), .C2(n6988), .ZN(P2_U3288) );
  INV_X1 U7419 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5833) );
  OAI222_X1 U7420 ( .A1(n7278), .A2(n5833), .B1(n8733), .B2(n5832), .C1(
        P2_U3151), .C2(n10155), .ZN(P2_U3289) );
  INV_X1 U7421 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U7422 ( .A1(n6231), .A2(P1_U3973), .ZN(n5834) );
  OAI21_X1 U7423 ( .B1(P1_U3973), .B2(n5835), .A(n5834), .ZN(P1_U3554) );
  INV_X1 U7424 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8952) );
  INV_X1 U7425 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U7426 ( .A1(n7616), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5838) );
  INV_X1 U7427 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8934) );
  OR2_X1 U7428 ( .A1(n5836), .A2(n8934), .ZN(n5837) );
  OAI211_X1 U7429 ( .C1(n7592), .C2(n9791), .A(n5838), .B(n5837), .ZN(n9484)
         );
  NAND2_X1 U7430 ( .A1(n9484), .A2(P1_U3973), .ZN(n5839) );
  OAI21_X1 U7431 ( .B1(P1_U3973), .B2(n8952), .A(n5839), .ZN(P1_U3585) );
  NAND2_X1 U7432 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6123) );
  NAND2_X1 U7433 ( .A1(n6264), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7434 ( .A1(n6615), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6710) );
  INV_X1 U7435 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n7150) );
  INV_X1 U7436 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7217) );
  XNOR2_X1 U7437 ( .A(n7532), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n9666) );
  INV_X1 U7438 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9835) );
  NAND2_X1 U7439 ( .A1(n7589), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7440 ( .A1(n7616), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5840) );
  OAI211_X1 U7441 ( .C1(n9835), .C2(n7592), .A(n5841), .B(n5840), .ZN(n5842)
         );
  AOI21_X1 U7442 ( .B1(n9666), .B2(n7594), .A(n5842), .ZN(n9272) );
  NAND2_X1 U7443 ( .A1(n9398), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n5843) );
  OAI21_X1 U7444 ( .B1(n9272), .B2(n9398), .A(n5843), .ZN(P1_U3572) );
  INV_X1 U7445 ( .A(n6441), .ZN(n5848) );
  NAND2_X1 U7446 ( .A1(n5845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  XNOR2_X1 U7447 ( .A(n5846), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9916) );
  INV_X1 U7448 ( .A(n9916), .ZN(n5847) );
  OAI222_X1 U7449 ( .A1(n9868), .A2(n8825), .B1(n9872), .B2(n5848), .C1(
        P1_U3086), .C2(n5847), .ZN(P1_U3347) );
  OAI222_X1 U7450 ( .A1(n7278), .A2(n5849), .B1(n8733), .B2(n5848), .C1(
        P2_U3151), .C2(n10171), .ZN(P2_U3287) );
  INV_X1 U7451 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5854) );
  INV_X1 U7452 ( .A(n5851), .ZN(n5852) );
  AOI22_X1 U7453 ( .A1(n5862), .A2(n5854), .B1(n5853), .B2(n5852), .ZN(
        P2_U3376) );
  INV_X1 U7454 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8990) );
  NOR3_X1 U7455 ( .A1(n5857), .A2(n5856), .A3(n5855), .ZN(n5858) );
  AOI21_X1 U7456 ( .B1(n8990), .B2(n5862), .A(n5858), .ZN(P2_U3377) );
  AND2_X1 U7457 ( .A1(n5862), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U7458 ( .A1(n5862), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7459 ( .A1(n5862), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7460 ( .A1(n5862), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7461 ( .A1(n5862), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7462 ( .A1(n5862), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7463 ( .A1(n5862), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7464 ( .A1(n5862), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7465 ( .A1(n5862), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7466 ( .A1(n5862), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7467 ( .A1(n5862), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7468 ( .A1(n5862), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7469 ( .A1(n5862), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7470 ( .A1(n5862), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7471 ( .A1(n5862), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7472 ( .A1(n5862), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7473 ( .A1(n5862), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7474 ( .A1(n5862), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7475 ( .A1(n5862), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7476 ( .A1(n5862), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7477 ( .A1(n5862), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7478 ( .A1(n5862), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7479 ( .A1(n5862), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7480 ( .A1(n5862), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  INV_X1 U7481 ( .A(n9023), .ZN(n5861) );
  NAND2_X1 U7482 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5860) );
  XNOR2_X1 U7483 ( .A(n5860), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6604) );
  INV_X1 U7484 ( .A(n6604), .ZN(n5982) );
  OAI222_X1 U7485 ( .A1(n9872), .A2(n5861), .B1(n5982), .B2(P1_U3086), .C1(
        n8980), .C2(n9868), .ZN(P1_U3346) );
  INV_X1 U7486 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8920) );
  NOR2_X1 U7487 ( .A1(n5863), .A2(n8920), .ZN(P2_U3251) );
  INV_X1 U7488 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n8937) );
  NOR2_X1 U7489 ( .A1(n5863), .A2(n8937), .ZN(P2_U3248) );
  INV_X1 U7490 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n8999) );
  NOR2_X1 U7491 ( .A1(n5863), .A2(n8999), .ZN(P2_U3238) );
  INV_X1 U7492 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n8882) );
  NOR2_X1 U7493 ( .A1(n5863), .A2(n8882), .ZN(P2_U3259) );
  INV_X1 U7494 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n8883) );
  NOR2_X1 U7495 ( .A1(n5863), .A2(n8883), .ZN(P2_U3241) );
  INV_X1 U7496 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n8910) );
  NOR2_X1 U7497 ( .A1(n5863), .A2(n8910), .ZN(P2_U3246) );
  INV_X1 U7498 ( .A(n6704), .ZN(n5866) );
  NOR2_X1 U7499 ( .A1(n5859), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6012) );
  OR2_X1 U7500 ( .A1(n6012), .A2(n5864), .ZN(n5869) );
  XNOR2_X1 U7501 ( .A(n5869), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9902) );
  INV_X1 U7502 ( .A(n9902), .ZN(n6024) );
  OAI222_X1 U7503 ( .A1(n9872), .A2(n5866), .B1(n6024), .B2(P1_U3086), .C1(
        n5865), .C2(n9868), .ZN(P1_U3345) );
  OAI222_X1 U7504 ( .A1(n7278), .A2(n5867), .B1(n8733), .B2(n5866), .C1(n10184), .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U7505 ( .A(n6794), .ZN(n5873) );
  INV_X1 U7506 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U7507 ( .A1(n5869), .A2(n5868), .ZN(n5870) );
  NAND2_X1 U7508 ( .A1(n5870), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5871) );
  XNOR2_X1 U7509 ( .A(n5871), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9960) );
  AOI22_X1 U7510 ( .A1(n9960), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n6486), .ZN(n5872) );
  OAI21_X1 U7511 ( .B1(n5873), .B2(n9872), .A(n5872), .ZN(P1_U3344) );
  OAI222_X1 U7512 ( .A1(n7278), .A2(n8800), .B1(n8733), .B2(n5873), .C1(
        P2_U3151), .C2(n7368), .ZN(P2_U3284) );
  MUX2_X1 U7513 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5596), .Z(n6357) );
  XNOR2_X1 U7514 ( .A(n6357), .B(n6356), .ZN(n5875) );
  INV_X1 U7515 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6105) );
  MUX2_X1 U7516 ( .A(n5893), .B(n6105), .S(n8426), .Z(n10107) );
  AND2_X1 U7517 ( .A1(n10107), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5874) );
  NAND2_X1 U7518 ( .A1(P2_U3893), .A2(n5877), .ZN(n10193) );
  AOI211_X1 U7519 ( .C1(n5875), .C2(n5874), .A(n10193), .B(n6355), .ZN(n5901)
         );
  INV_X1 U7520 ( .A(n5880), .ZN(n5876) );
  NOR2_X1 U7521 ( .A1(n5879), .A2(n5876), .ZN(n5897) );
  NOR2_X1 U7522 ( .A1(n5877), .A2(P2_U3151), .ZN(n7379) );
  NAND2_X1 U7523 ( .A1(n5897), .A2(n7379), .ZN(n5885) );
  AND2_X1 U7524 ( .A1(n8256), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7525 ( .A1(n5879), .A2(n5878), .ZN(n5881) );
  OR2_X1 U7526 ( .A1(n5880), .A2(P2_U3151), .ZN(n8267) );
  NAND2_X1 U7527 ( .A1(n5881), .A2(n8267), .ZN(n5892) );
  INV_X1 U7528 ( .A(n5882), .ZN(n5883) );
  NAND2_X1 U7529 ( .A1(n5892), .A2(n5883), .ZN(n5884) );
  INV_X1 U7530 ( .A(n8262), .ZN(n5886) );
  INV_X1 U7531 ( .A(n10199), .ZN(n10127) );
  INV_X1 U7532 ( .A(n6356), .ZN(n5888) );
  INV_X1 U7533 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10112) );
  NAND2_X1 U7534 ( .A1(n10112), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5887) );
  AND2_X1 U7535 ( .A1(n5894), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6363) );
  XNOR2_X1 U7536 ( .A(n6362), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n5889) );
  AOI22_X1 U7537 ( .A1(n10127), .A2(n5889), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        P2_U3151), .ZN(n5890) );
  OAI21_X1 U7538 ( .B1(n10185), .B2(n6356), .A(n5890), .ZN(n5900) );
  AND2_X1 U7539 ( .A1(n5892), .A2(n5891), .ZN(n10109) );
  AND2_X1 U7540 ( .A1(n10109), .A2(n7294), .ZN(n9885) );
  INV_X1 U7541 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5896) );
  INV_X1 U7542 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U7543 ( .A1(n5894), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6371) );
  AOI21_X1 U7544 ( .B1(n5896), .B2(n5895), .A(n6373), .ZN(n5898) );
  INV_X1 U7545 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10328) );
  OAI22_X1 U7546 ( .A1(n10191), .A2(n5898), .B1(n10328), .B2(n10183), .ZN(
        n5899) );
  OR3_X1 U7547 ( .A1(n5901), .A2(n5900), .A3(n5899), .ZN(P2_U3183) );
  NAND2_X1 U7548 ( .A1(n7779), .A2(n7699), .ZN(n6095) );
  NOR2_X1 U7549 ( .A1(n6095), .A2(n7755), .ZN(n6332) );
  INV_X1 U7550 ( .A(n7684), .ZN(n5926) );
  NAND2_X1 U7551 ( .A1(n7184), .A2(P1_B_REG_SCAN_IN), .ZN(n5903) );
  MUX2_X1 U7552 ( .A(P1_B_REG_SCAN_IN), .B(n5903), .S(n5902), .Z(n5905) );
  INV_X1 U7553 ( .A(n7255), .ZN(n5904) );
  OR2_X1 U7554 ( .A1(n9854), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7555 ( .A1(n5902), .A2(n7255), .ZN(n9856) );
  OR2_X1 U7556 ( .A1(n9854), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5907) );
  NAND2_X1 U7557 ( .A1(n7255), .A2(n7184), .ZN(n9855) );
  NOR4_X1 U7558 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5916) );
  NOR4_X1 U7559 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5915) );
  INV_X1 U7560 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10074) );
  INV_X1 U7561 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10073) );
  INV_X1 U7562 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10076) );
  INV_X1 U7563 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10070) );
  NAND4_X1 U7564 ( .A1(n10074), .A2(n10073), .A3(n10076), .A4(n10070), .ZN(
        n5913) );
  NOR4_X1 U7565 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5911) );
  NOR4_X1 U7566 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5910) );
  NOR4_X1 U7567 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5909) );
  NOR4_X1 U7568 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5908) );
  NAND4_X1 U7569 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n5912)
         );
  NOR4_X1 U7570 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5913), .A4(n5912), .ZN(n5914) );
  AND3_X1 U7571 ( .A1(n5916), .A2(n5915), .A3(n5914), .ZN(n5917) );
  OR2_X1 U7572 ( .A1(n9854), .A2(n5917), .ZN(n6093) );
  NAND3_X1 U7573 ( .A1(n6322), .A2(n6325), .A3(n6093), .ZN(n5923) );
  OAI21_X1 U7574 ( .B1(n6332), .B2(n10094), .A(n5923), .ZN(n5919) );
  NAND2_X1 U7575 ( .A1(n7752), .A2(n7684), .ZN(n6091) );
  NAND3_X1 U7576 ( .A1(n5919), .A2(n5918), .A3(n6091), .ZN(n5920) );
  NAND2_X1 U7577 ( .A1(n5920), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5921) );
  NOR2_X1 U7578 ( .A1(n9359), .A2(P1_U3086), .ZN(n6010) );
  INV_X1 U7579 ( .A(n9853), .ZN(n5922) );
  INV_X1 U7580 ( .A(n7752), .ZN(n7753) );
  NAND2_X1 U7581 ( .A1(n7753), .A2(n10094), .ZN(n5924) );
  INV_X1 U7582 ( .A(n5925), .ZN(n5932) );
  NAND2_X1 U7583 ( .A1(n5932), .A2(n5926), .ZN(n9357) );
  INV_X1 U7584 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6399) );
  INV_X1 U7585 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5927) );
  OR2_X1 U7586 ( .A1(n7592), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7587 ( .A1(n7589), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5928) );
  INV_X1 U7588 ( .A(n9399), .ZN(n7643) );
  NAND2_X1 U7589 ( .A1(n7752), .A2(n7769), .ZN(n9352) );
  NOR2_X1 U7590 ( .A1(n7643), .A2(n9352), .ZN(n10057) );
  AOI22_X1 U7591 ( .A1(n5931), .A2(n9931), .B1(n9926), .B2(n10057), .ZN(n5934)
         );
  NAND2_X1 U7592 ( .A1(n9368), .A2(n6230), .ZN(n5933) );
  OAI211_X1 U7593 ( .C1(n6010), .C2(n5935), .A(n5934), .B(n5933), .ZN(P1_U3232) );
  INV_X2 U7594 ( .A(n6074), .ZN(n9204) );
  NAND2_X1 U7595 ( .A1(n9399), .A2(n6752), .ZN(n5943) );
  NAND2_X1 U7596 ( .A1(n4417), .A2(n7642), .ZN(n5942) );
  NAND2_X1 U7597 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  XNOR2_X1 U7598 ( .A(n5944), .B(n6074), .ZN(n5986) );
  AOI22_X1 U7599 ( .A1(n9399), .A2(n9081), .B1(n9082), .B2(n7642), .ZN(n5988)
         );
  XNOR2_X1 U7600 ( .A(n5986), .B(n5988), .ZN(n5989) );
  XNOR2_X1 U7601 ( .A(n5990), .B(n5989), .ZN(n5945) );
  NAND2_X1 U7602 ( .A1(n5945), .A2(n9931), .ZN(n5955) );
  NAND2_X1 U7603 ( .A1(n7752), .A2(n5946), .ZN(n9350) );
  INV_X1 U7604 ( .A(n9350), .ZN(n9296) );
  NAND2_X1 U7605 ( .A1(n6231), .A2(n9296), .ZN(n5953) );
  NAND2_X1 U7606 ( .A1(n7589), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5951) );
  INV_X1 U7607 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9413) );
  OR2_X1 U7608 ( .A1(n7534), .A2(n9413), .ZN(n5950) );
  OR2_X1 U7609 ( .A1(n7440), .A2(n5792), .ZN(n5949) );
  INV_X1 U7610 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7611 ( .A1(n7592), .A2(n5947), .ZN(n5948) );
  INV_X1 U7612 ( .A(n9352), .ZN(n9229) );
  NAND2_X1 U7613 ( .A1(n9397), .A2(n9229), .ZN(n5952) );
  NAND2_X1 U7614 ( .A1(n5953), .A2(n5952), .ZN(n6394) );
  AOI22_X1 U7615 ( .A1(n9368), .A2(n7642), .B1(n9926), .B2(n6394), .ZN(n5954)
         );
  OAI211_X1 U7616 ( .C1(n6010), .C2(n6399), .A(n5955), .B(n5954), .ZN(P1_U3222) );
  NOR2_X1 U7617 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n6604), .ZN(n5956) );
  AOI21_X1 U7618 ( .B1(n6604), .B2(P1_REG2_REG_9__SCAN_IN), .A(n5956), .ZN(
        n5967) );
  NAND2_X1 U7619 ( .A1(n5968), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7620 ( .A1(n5958), .A2(n5957), .ZN(n9448) );
  INV_X1 U7621 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6333) );
  XNOR2_X1 U7622 ( .A(n9443), .B(n6333), .ZN(n9449) );
  NAND2_X1 U7623 ( .A1(n9448), .A2(n9449), .ZN(n9447) );
  NAND2_X1 U7624 ( .A1(n9443), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U7625 ( .A1(n9447), .A2(n5959), .ZN(n9461) );
  INV_X1 U7626 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5960) );
  XNOR2_X1 U7627 ( .A(n9456), .B(n5960), .ZN(n9462) );
  NAND2_X1 U7628 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
  NAND2_X1 U7629 ( .A1(n9456), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5961) );
  NAND2_X1 U7630 ( .A1(n9460), .A2(n5961), .ZN(n9471) );
  INV_X1 U7631 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U7632 ( .A(n9469), .B(n6530), .ZN(n9472) );
  NAND2_X1 U7633 ( .A1(n9471), .A2(n9472), .ZN(n9470) );
  NAND2_X1 U7634 ( .A1(n9469), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5962) );
  NAND2_X1 U7635 ( .A1(n9470), .A2(n5962), .ZN(n9910) );
  OR2_X1 U7636 ( .A1(n9916), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U7637 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n9916), .ZN(n5963) );
  NAND2_X1 U7638 ( .A1(n5964), .A2(n5963), .ZN(n9912) );
  INV_X1 U7639 ( .A(n9912), .ZN(n5965) );
  AND2_X1 U7640 ( .A1(n9910), .A2(n5965), .ZN(n9911) );
  AOI21_X1 U7641 ( .B1(n9916), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9911), .ZN(
        n5966) );
  NAND2_X1 U7642 ( .A1(n5967), .A2(n5966), .ZN(n6029) );
  OAI21_X1 U7643 ( .B1(n5967), .B2(n5966), .A(n6029), .ZN(n5984) );
  INV_X1 U7644 ( .A(n10031), .ZN(n10015) );
  INV_X1 U7645 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U7646 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n6604), .B1(n5982), .B2(
        n10104), .ZN(n5978) );
  NAND2_X1 U7647 ( .A1(n5968), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7648 ( .A1(n5970), .A2(n5969), .ZN(n9445) );
  INV_X1 U7649 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6125) );
  XNOR2_X1 U7650 ( .A(n9443), .B(n6125), .ZN(n9446) );
  NAND2_X1 U7651 ( .A1(n9445), .A2(n9446), .ZN(n9444) );
  NAND2_X1 U7652 ( .A1(n9443), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7653 ( .A1(n9444), .A2(n5971), .ZN(n9458) );
  INV_X1 U7654 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6266) );
  XNOR2_X1 U7655 ( .A(n9456), .B(n6266), .ZN(n9459) );
  NAND2_X1 U7656 ( .A1(n9458), .A2(n9459), .ZN(n9457) );
  NAND2_X1 U7657 ( .A1(n9456), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7658 ( .A1(n9457), .A2(n5972), .ZN(n9475) );
  INV_X1 U7659 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6308) );
  XNOR2_X1 U7660 ( .A(n9469), .B(n6308), .ZN(n9476) );
  NAND2_X1 U7661 ( .A1(n9475), .A2(n9476), .ZN(n9473) );
  NAND2_X1 U7662 ( .A1(n9469), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7663 ( .A1(n9473), .A2(n5973), .ZN(n9906) );
  OR2_X1 U7664 ( .A1(n9916), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7665 ( .A1(P1_REG1_REG_8__SCAN_IN), .A2(n9916), .ZN(n5974) );
  NAND2_X1 U7666 ( .A1(n5975), .A2(n5974), .ZN(n9908) );
  INV_X1 U7667 ( .A(n9908), .ZN(n5976) );
  AND2_X1 U7668 ( .A1(n9906), .A2(n5976), .ZN(n9907) );
  AOI21_X1 U7669 ( .B1(n9916), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9907), .ZN(
        n5977) );
  NAND2_X1 U7670 ( .A1(n5978), .A2(n5977), .ZN(n6025) );
  OAI21_X1 U7671 ( .B1(n5978), .B2(n5977), .A(n6025), .ZN(n5979) );
  NAND2_X1 U7672 ( .A1(n5979), .A2(n9474), .ZN(n5981) );
  NOR2_X1 U7673 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6453), .ZN(n6773) );
  AOI21_X1 U7674 ( .B1(n9948), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n6773), .ZN(
        n5980) );
  OAI211_X1 U7675 ( .C1(n10015), .C2(n5982), .A(n5981), .B(n5980), .ZN(n5983)
         );
  AOI21_X1 U7676 ( .B1(n10024), .B2(n5984), .A(n5983), .ZN(n5985) );
  INV_X1 U7677 ( .A(n5985), .ZN(P1_U3252) );
  INV_X1 U7678 ( .A(n5986), .ZN(n5987) );
  NAND2_X1 U7679 ( .A1(n9397), .A2(n6752), .ZN(n5997) );
  OR2_X1 U7680 ( .A1(n7613), .A2(n5991), .ZN(n5995) );
  OR2_X1 U7681 ( .A1(n7521), .A2(n5992), .ZN(n5993) );
  NAND2_X1 U7682 ( .A1(n4514), .A2(n6672), .ZN(n5996) );
  NAND2_X1 U7683 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  INV_X1 U7684 ( .A(n9397), .ZN(n6240) );
  INV_X1 U7685 ( .A(n6672), .ZN(n7646) );
  OAI22_X1 U7686 ( .A1(n6240), .A2(n9201), .B1(n7646), .B2(n9207), .ZN(n6079)
         );
  XNOR2_X1 U7687 ( .A(n6081), .B(n6080), .ZN(n5999) );
  NAND2_X1 U7688 ( .A1(n5999), .A2(n9931), .ZN(n6009) );
  NAND2_X1 U7689 ( .A1(n9399), .A2(n9296), .ZN(n6007) );
  NAND2_X1 U7690 ( .A1(n7589), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6005) );
  OR2_X1 U7691 ( .A1(n7440), .A2(n6000), .ZN(n6004) );
  INV_X1 U7692 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7693 ( .A1(n7592), .A2(n6001), .ZN(n6003) );
  OR2_X1 U7694 ( .A1(n7534), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6002) );
  NAND4_X1 U7695 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n9396)
         );
  NAND2_X1 U7696 ( .A1(n9396), .A2(n9229), .ZN(n6006) );
  NAND2_X1 U7697 ( .A1(n6007), .A2(n6006), .ZN(n6293) );
  AOI22_X1 U7698 ( .A1(n9368), .A2(n6672), .B1(n9926), .B2(n6293), .ZN(n6008)
         );
  OAI211_X1 U7699 ( .C1(n6010), .C2(n9413), .A(n6009), .B(n6008), .ZN(P1_U3237) );
  INV_X1 U7700 ( .A(n6912), .ZN(n6039) );
  NOR2_X1 U7701 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6011) );
  NAND2_X1 U7702 ( .A1(n6012), .A2(n6011), .ZN(n6040) );
  NAND2_X1 U7703 ( .A1(n6040), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6013) );
  XNOR2_X1 U7704 ( .A(n6013), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6913) );
  INV_X1 U7705 ( .A(n6913), .ZN(n6038) );
  OAI222_X1 U7706 ( .A1(n9872), .A2(n6039), .B1(n6038), .B2(P1_U3086), .C1(
        n6014), .C2(n9868), .ZN(P1_U3343) );
  NAND2_X1 U7707 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n6015) );
  INV_X1 U7708 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9299) );
  INV_X1 U7709 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9230) );
  OR2_X1 U7710 ( .A1(n7588), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7711 ( .A1(n6016), .A2(n6205), .ZN(n9283) );
  INV_X1 U7712 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n8992) );
  NAND2_X1 U7713 ( .A1(n7589), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7714 ( .A1(n6082), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6017) );
  OAI211_X1 U7715 ( .C1(n8992), .C2(n7440), .A(n6018), .B(n6017), .ZN(n6019)
         );
  NAND2_X1 U7716 ( .A1(n9398), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6020) );
  OAI21_X1 U7717 ( .B1(n9247), .B2(n9398), .A(n6020), .ZN(P1_U3578) );
  INV_X1 U7718 ( .A(n9960), .ZN(n6022) );
  NOR2_X1 U7719 ( .A1(n6022), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6021) );
  AOI21_X1 U7720 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6022), .A(n6021), .ZN(
        n9954) );
  NOR2_X1 U7721 ( .A1(n6024), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6023) );
  AOI21_X1 U7722 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6024), .A(n6023), .ZN(
        n9895) );
  OAI21_X1 U7723 ( .B1(n6604), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6025), .ZN(
        n9896) );
  NOR2_X1 U7724 ( .A1(n9895), .A2(n9896), .ZN(n9894) );
  AOI21_X1 U7725 ( .B1(n9902), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9894), .ZN(
        n9953) );
  NOR2_X1 U7726 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  AOI21_X1 U7727 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9960), .A(n9952), .ZN(
        n6027) );
  INV_X1 U7728 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6975) );
  AOI22_X1 U7729 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n6913), .B1(n6038), .B2(
        n6975), .ZN(n6026) );
  NAND2_X1 U7730 ( .A1(n6027), .A2(n6026), .ZN(n6870) );
  OAI21_X1 U7731 ( .B1(n6027), .B2(n6026), .A(n6870), .ZN(n6034) );
  XNOR2_X1 U7732 ( .A(n9960), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9956) );
  NAND2_X1 U7733 ( .A1(n9902), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6028) );
  OAI21_X1 U7734 ( .B1(n9902), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6028), .ZN(
        n9898) );
  OAI21_X1 U7735 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6604), .A(n6029), .ZN(
        n9899) );
  NOR2_X1 U7736 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  AOI21_X1 U7737 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9902), .A(n9897), .ZN(
        n9957) );
  NOR2_X1 U7738 ( .A1(n9956), .A2(n9957), .ZN(n9955) );
  AOI21_X1 U7739 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9960), .A(n9955), .ZN(
        n6032) );
  NOR2_X1 U7740 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6913), .ZN(n6030) );
  AOI21_X1 U7741 ( .B1(n6913), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6030), .ZN(
        n6031) );
  NAND2_X1 U7742 ( .A1(n6031), .A2(n6032), .ZN(n6876) );
  OAI21_X1 U7743 ( .B1(n6032), .B2(n6031), .A(n6876), .ZN(n6033) );
  AOI22_X1 U7744 ( .A1(n9474), .A2(n6034), .B1(n10024), .B2(n6033), .ZN(n6037)
         );
  NAND2_X1 U7745 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9238) );
  INV_X1 U7746 ( .A(n9238), .ZN(n6035) );
  AOI21_X1 U7747 ( .B1(n9948), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n6035), .ZN(
        n6036) );
  OAI211_X1 U7748 ( .C1(n6038), .C2(n10015), .A(n6037), .B(n6036), .ZN(
        P1_U3255) );
  INV_X1 U7749 ( .A(n7344), .ZN(n7324) );
  OAI222_X1 U7750 ( .A1(n7278), .A2(n8880), .B1(n8733), .B2(n6039), .C1(n7324), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U7751 ( .A(n7074), .ZN(n6066) );
  NAND2_X1 U7752 ( .A1(n6138), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6041) );
  XNOR2_X1 U7753 ( .A(n6041), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9969) );
  AOI22_X1 U7754 ( .A1(n9969), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n6486), .ZN(n6042) );
  OAI21_X1 U7755 ( .B1(n6066), .B2(n9872), .A(n6042), .ZN(P1_U3342) );
  NAND2_X1 U7756 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  OAI211_X1 U7757 ( .C1(n6048), .C2(n6051), .A(n6046), .B(n6045), .ZN(n6047)
         );
  NAND2_X1 U7758 ( .A1(n6047), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6050) );
  INV_X1 U7759 ( .A(n6141), .ZN(n6165) );
  NAND2_X1 U7760 ( .A1(n6059), .A2(n6165), .ZN(n8263) );
  OR2_X1 U7761 ( .A1(n6048), .A2(n8263), .ZN(n6049) );
  NAND2_X2 U7762 ( .A1(n6050), .A2(n6049), .ZN(n8022) );
  NOR2_X1 U7763 ( .A1(n8022), .A2(P2_U3151), .ZN(n6191) );
  INV_X1 U7764 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6065) );
  INV_X1 U7765 ( .A(n6172), .ZN(n6153) );
  NAND2_X1 U7766 ( .A1(n8286), .A2(n6153), .ZN(n8084) );
  NAND2_X1 U7767 ( .A1(n8078), .A2(n8084), .ZN(n8037) );
  INV_X1 U7768 ( .A(n6051), .ZN(n6052) );
  NAND2_X1 U7769 ( .A1(n6144), .A2(n6052), .ZN(n6056) );
  INV_X1 U7770 ( .A(n6053), .ZN(n6054) );
  NAND2_X1 U7771 ( .A1(n6057), .A2(n6054), .ZN(n6055) );
  NAND2_X1 U7772 ( .A1(n6057), .A2(n7262), .ZN(n6060) );
  AND2_X1 U7773 ( .A1(n6142), .A2(n6165), .ZN(n6062) );
  OAI22_X1 U7774 ( .A1(n8025), .A2(n6153), .B1(n6061), .B2(n8020), .ZN(n6063)
         );
  AOI21_X1 U7775 ( .B1(n8037), .B2(n8016), .A(n6063), .ZN(n6064) );
  OAI21_X1 U7776 ( .B1(n6191), .B2(n6065), .A(n6064), .ZN(P2_U3172) );
  INV_X1 U7777 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6067) );
  INV_X1 U7778 ( .A(n8327), .ZN(n8316) );
  OAI222_X1 U7779 ( .A1(n7278), .A2(n6067), .B1(n8733), .B2(n6066), .C1(
        P2_U3151), .C2(n8316), .ZN(P2_U3282) );
  OR2_X1 U7780 ( .A1(n7521), .A2(n6068), .ZN(n6072) );
  OR2_X1 U7781 ( .A1(n7613), .A2(n6069), .ZN(n6071) );
  OR2_X1 U7782 ( .A1(n6253), .A2(n9426), .ZN(n6070) );
  AOI22_X1 U7783 ( .A1(n9396), .A2(n9137), .B1(n6669), .B2(n4417), .ZN(n6075)
         );
  XNOR2_X1 U7784 ( .A(n6075), .B(n6074), .ZN(n6111) );
  NAND2_X1 U7785 ( .A1(n9396), .A2(n9081), .ZN(n6078) );
  NAND2_X1 U7786 ( .A1(n6669), .A2(n9082), .ZN(n6077) );
  NAND2_X1 U7787 ( .A1(n6078), .A2(n6077), .ZN(n6109) );
  XNOR2_X1 U7788 ( .A(n6111), .B(n6109), .ZN(n6112) );
  XOR2_X1 U7789 ( .A(n6112), .B(n6113), .Z(n6090) );
  NAND2_X1 U7790 ( .A1(n6082), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6086) );
  INV_X1 U7791 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10044) );
  OR2_X1 U7792 ( .A1(n5836), .A2(n10044), .ZN(n6085) );
  OAI21_X1 U7793 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6123), .ZN(n10043) );
  OR2_X1 U7794 ( .A1(n7534), .A2(n10043), .ZN(n6084) );
  OR2_X1 U7795 ( .A1(n7440), .A2(n5787), .ZN(n6083) );
  AOI22_X1 U7796 ( .A1(n9296), .A2(n9397), .B1(n9395), .B2(n9229), .ZN(n6279)
         );
  INV_X1 U7797 ( .A(n6279), .ZN(n6087) );
  AOI22_X1 U7798 ( .A1(n9368), .A2(n6669), .B1(n9926), .B2(n6087), .ZN(n6089)
         );
  MUX2_X1 U7799 ( .A(n9935), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6088) );
  OAI211_X1 U7800 ( .C1(n6090), .C2(n9370), .A(n6089), .B(n6088), .ZN(P1_U3218) );
  AND2_X1 U7801 ( .A1(n9853), .A2(n6091), .ZN(n6092) );
  NAND2_X1 U7802 ( .A1(n6093), .A2(n6092), .ZN(n6323) );
  INV_X1 U7803 ( .A(n6095), .ZN(n6101) );
  OR2_X1 U7804 ( .A1(n7779), .A2(n5757), .ZN(n6096) );
  NAND2_X1 U7805 ( .A1(n7722), .A2(n6098), .ZN(n7403) );
  NOR2_X1 U7806 ( .A1(n5756), .A2(n6326), .ZN(n7764) );
  NOR2_X1 U7807 ( .A1(n7764), .A2(n6101), .ZN(n10058) );
  NAND2_X1 U7808 ( .A1(n5756), .A2(n7684), .ZN(n6097) );
  NAND2_X1 U7809 ( .A1(n10058), .A2(n6097), .ZN(n6290) );
  NAND2_X1 U7810 ( .A1(n7779), .A2(n4418), .ZN(n7625) );
  INV_X1 U7811 ( .A(n10096), .ZN(n9778) );
  NOR2_X1 U7812 ( .A1(n6231), .A2(n10061), .ZN(n6393) );
  INV_X1 U7813 ( .A(n6393), .ZN(n6099) );
  NAND2_X1 U7814 ( .A1(n6231), .A2(n10061), .ZN(n7641) );
  AND2_X1 U7815 ( .A1(n6099), .A2(n7641), .ZN(n10056) );
  AOI21_X1 U7816 ( .B1(n9578), .B2(n9778), .A(n10056), .ZN(n6100) );
  AOI211_X1 U7817 ( .C1(n6101), .C2(n6230), .A(n10057), .B(n6100), .ZN(n6435)
         );
  OR2_X1 U7818 ( .A1(n6435), .A2(n10098), .ZN(n6102) );
  OAI21_X1 U7819 ( .B1(n10100), .B2(n5720), .A(n6102), .ZN(P1_U3453) );
  OAI21_X1 U7820 ( .B1(n10207), .B2(n10275), .A(n8037), .ZN(n6103) );
  NAND2_X1 U7821 ( .A1(n8284), .A2(n10202), .ZN(n6167) );
  OAI211_X1 U7822 ( .C1(n10282), .C2(n6153), .A(n6103), .B(n6167), .ZN(n6106)
         );
  NAND2_X1 U7823 ( .A1(n6106), .A2(n10325), .ZN(n6104) );
  OAI21_X1 U7824 ( .B1(n10325), .B2(n6105), .A(n6104), .ZN(P2_U3459) );
  INV_X1 U7825 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7826 ( .A1(n6106), .A2(n10300), .ZN(n6107) );
  OAI21_X1 U7827 ( .B1(n6108), .B2(n10300), .A(n6107), .ZN(P2_U3390) );
  INV_X1 U7828 ( .A(n6109), .ZN(n6110) );
  AOI22_X2 U7829 ( .A1(n6113), .A2(n6112), .B1(n6111), .B2(n6110), .ZN(n6122)
         );
  OR2_X1 U7830 ( .A1(n6114), .A2(n7521), .ZN(n6119) );
  OR2_X1 U7831 ( .A1(n6253), .A2(n6115), .ZN(n6118) );
  OR2_X1 U7832 ( .A1(n7613), .A2(n6116), .ZN(n6117) );
  AOI22_X1 U7833 ( .A1(n9137), .A2(n9395), .B1(n10046), .B2(n4514), .ZN(n6120)
         );
  XNOR2_X1 U7834 ( .A(n6120), .B(n9140), .ZN(n6416) );
  INV_X1 U7835 ( .A(n9395), .ZN(n6262) );
  OAI22_X1 U7836 ( .A1(n6262), .A2(n9201), .B1(n6260), .B2(n9207), .ZN(n6414)
         );
  XNOR2_X1 U7837 ( .A(n6416), .B(n6414), .ZN(n6121) );
  OAI211_X1 U7838 ( .C1(n6122), .C2(n6121), .A(n6417), .B(n9931), .ZN(n6136)
         );
  NAND2_X1 U7839 ( .A1(n9396), .A2(n9296), .ZN(n6131) );
  NAND2_X1 U7840 ( .A1(n7589), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6129) );
  OR2_X1 U7841 ( .A1(n7592), .A2(n6272), .ZN(n6128) );
  AND2_X1 U7842 ( .A1(n6123), .A2(n6425), .ZN(n6124) );
  OR2_X1 U7843 ( .A1(n6124), .A2(n6264), .ZN(n6431) );
  OR2_X1 U7844 ( .A1(n7534), .A2(n6431), .ZN(n6127) );
  OR2_X1 U7845 ( .A1(n7440), .A2(n6125), .ZN(n6126) );
  NAND4_X1 U7846 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(n9394)
         );
  NAND2_X1 U7847 ( .A1(n9394), .A2(n9229), .ZN(n6130) );
  NAND2_X1 U7848 ( .A1(n6131), .A2(n6130), .ZN(n6244) );
  INV_X1 U7849 ( .A(n6244), .ZN(n6133) );
  OAI21_X1 U7850 ( .B1(n9357), .B2(n6133), .A(n6132), .ZN(n6134) );
  AOI21_X1 U7851 ( .B1(n9368), .B2(n10046), .A(n6134), .ZN(n6135) );
  OAI211_X1 U7852 ( .C1(n9935), .C2(n10043), .A(n6136), .B(n6135), .ZN(
        P1_U3230) );
  INV_X1 U7853 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6137) );
  INV_X1 U7854 ( .A(n7144), .ZN(n6140) );
  OAI222_X1 U7855 ( .A1(n7278), .A2(n6137), .B1(n8733), .B2(n6140), .C1(
        P2_U3151), .C2(n8351), .ZN(P2_U3281) );
  INV_X1 U7856 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8988) );
  OAI21_X1 U7857 ( .B1(n6138), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6177) );
  XNOR2_X1 U7858 ( .A(n6177), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9986) );
  INV_X1 U7859 ( .A(n9986), .ZN(n6139) );
  OAI222_X1 U7860 ( .A1(n9868), .A2(n8988), .B1(n9872), .B2(n6140), .C1(
        P1_U3086), .C2(n6139), .ZN(P1_U3341) );
  INV_X1 U7861 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6160) );
  NOR2_X1 U7862 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  INV_X1 U7863 ( .A(n8018), .ZN(n7999) );
  OAI22_X1 U7864 ( .A1(n7999), .A2(n6145), .B1(n5198), .B2(n8020), .ZN(n6146)
         );
  AOI21_X1 U7865 ( .B1(n6211), .B2(n7969), .A(n6146), .ZN(n6159) );
  OAI21_X1 U7866 ( .B1(n6148), .B2(n8076), .A(n6147), .ZN(n6149) );
  INV_X1 U7867 ( .A(n6149), .ZN(n6150) );
  XNOR2_X1 U7868 ( .A(n7896), .B(n6211), .ZN(n6151) );
  OR2_X1 U7869 ( .A1(n6151), .A2(n6061), .ZN(n6152) );
  NAND2_X1 U7870 ( .A1(n6151), .A2(n6061), .ZN(n6182) );
  AND2_X1 U7871 ( .A1(n6152), .A2(n6182), .ZN(n6156) );
  NAND2_X1 U7872 ( .A1(n6153), .A2(n7932), .ZN(n6154) );
  NAND2_X1 U7873 ( .A1(n8078), .A2(n6154), .ZN(n6155) );
  NAND2_X1 U7874 ( .A1(n6156), .A2(n6155), .ZN(n6183) );
  OAI21_X1 U7875 ( .B1(n6156), .B2(n6155), .A(n6183), .ZN(n6157) );
  NAND2_X1 U7876 ( .A1(n6157), .A2(n8016), .ZN(n6158) );
  OAI211_X1 U7877 ( .C1(n6191), .C2(n6160), .A(n6159), .B(n6158), .ZN(P2_U3162) );
  MUX2_X1 U7878 ( .A(n4497), .B(n6162), .S(n6161), .Z(n6163) );
  INV_X1 U7879 ( .A(n8037), .ZN(n6166) );
  NOR3_X1 U7880 ( .A1(n6166), .A2(n6165), .A3(n10299), .ZN(n6169) );
  INV_X1 U7881 ( .A(n6167), .ZN(n6168) );
  OAI21_X1 U7882 ( .B1(n6169), .B2(n6168), .A(n8601), .ZN(n6174) );
  INV_X1 U7883 ( .A(n6170), .ZN(n6171) );
  AOI22_X1 U7884 ( .A1(n10210), .A2(n6172), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10211), .ZN(n6173) );
  OAI211_X1 U7885 ( .C1(n5893), .C2(n8601), .A(n6174), .B(n6173), .ZN(P2_U3233) );
  INV_X1 U7886 ( .A(n7211), .ZN(n6181) );
  AOI22_X1 U7887 ( .A1(n8373), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9020), .ZN(n6175) );
  OAI21_X1 U7888 ( .B1(n6181), .B2(n8733), .A(n6175), .ZN(P2_U3280) );
  INV_X1 U7889 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7890 ( .A1(n6177), .A2(n6176), .ZN(n6178) );
  NAND2_X1 U7891 ( .A1(n6178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6179) );
  XNOR2_X1 U7892 ( .A(n6179), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10006) );
  INV_X1 U7893 ( .A(n10006), .ZN(n6878) );
  OAI222_X1 U7894 ( .A1(n9872), .A2(n6181), .B1(n6878), .B2(P1_U3086), .C1(
        n6180), .C2(n9868), .ZN(P1_U3340) );
  INV_X1 U7895 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6190) );
  XNOR2_X1 U7896 ( .A(n5198), .B(n6220), .ZN(n6185) );
  NAND2_X1 U7897 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  NAND2_X1 U7898 ( .A1(n6184), .A2(n6185), .ZN(n6226) );
  OAI21_X1 U7899 ( .B1(n6185), .B2(n6184), .A(n6226), .ZN(n6186) );
  NAND2_X1 U7900 ( .A1(n6186), .A2(n8016), .ZN(n6189) );
  OAI22_X1 U7901 ( .A1(n7999), .A2(n6061), .B1(n10222), .B2(n8020), .ZN(n6187)
         );
  AOI21_X1 U7902 ( .B1(n10238), .B2(n7969), .A(n6187), .ZN(n6188) );
  OAI211_X1 U7903 ( .C1(n6191), .C2(n6190), .A(n6189), .B(n6188), .ZN(P2_U3177) );
  NAND2_X1 U7904 ( .A1(n5600), .A2(n8078), .ZN(n6192) );
  NAND2_X1 U7905 ( .A1(n6193), .A2(n6192), .ZN(n6212) );
  INV_X1 U7906 ( .A(n6212), .ZN(n6203) );
  AND2_X1 U7907 ( .A1(n8076), .A2(n6194), .ZN(n10233) );
  NAND2_X1 U7908 ( .A1(n8601), .A2(n10233), .ZN(n8451) );
  NAND2_X1 U7909 ( .A1(n6212), .A2(n10230), .ZN(n6200) );
  OAI21_X1 U7910 ( .B1(n6196), .B2(n5600), .A(n6195), .ZN(n6197) );
  NAND2_X1 U7911 ( .A1(n6197), .A2(n10207), .ZN(n6199) );
  AOI22_X1 U7912 ( .A1(n10205), .A2(n10202), .B1(n10204), .B2(n8286), .ZN(
        n6198) );
  AND3_X1 U7913 ( .A1(n6200), .A2(n6199), .A3(n6198), .ZN(n6214) );
  MUX2_X1 U7914 ( .A(n6214), .B(n5896), .S(n10235), .Z(n6202) );
  AOI22_X1 U7915 ( .A1(n10210), .A2(n6211), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10211), .ZN(n6201) );
  OAI211_X1 U7916 ( .C1(n6203), .C2(n8451), .A(n6202), .B(n6201), .ZN(P2_U3232) );
  NAND2_X1 U7917 ( .A1(n7616), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6209) );
  INV_X1 U7918 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6204) );
  OR2_X1 U7919 ( .A1(n5836), .A2(n6204), .ZN(n6208) );
  INV_X1 U7920 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9799) );
  OR2_X1 U7921 ( .A1(n7592), .A2(n9799), .ZN(n6207) );
  INV_X1 U7922 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9165) );
  XNOR2_X1 U7923 ( .A(n7430), .B(n9165), .ZN(n9162) );
  OR2_X1 U7924 ( .A1(n7534), .A2(n9162), .ZN(n6206) );
  NAND2_X1 U7925 ( .A1(n9398), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6210) );
  OAI21_X1 U7926 ( .B1(n9353), .B2(n9398), .A(n6210), .ZN(P1_U3581) );
  AOI22_X1 U7927 ( .A1(n6212), .A2(n10255), .B1(n6211), .B2(n10299), .ZN(n6213) );
  AND2_X1 U7928 ( .A1(n6214), .A2(n6213), .ZN(n10236) );
  INV_X1 U7929 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6215) );
  MUX2_X1 U7930 ( .A(n10236), .B(n6215), .S(n10323), .Z(n6216) );
  INV_X1 U7931 ( .A(n6216), .ZN(P2_U3460) );
  NAND2_X1 U7932 ( .A1(n8018), .A2(n10205), .ZN(n6217) );
  OR2_X1 U7933 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10212), .ZN(n10144) );
  OAI211_X1 U7934 ( .C1(n6474), .C2(n8020), .A(n6217), .B(n10144), .ZN(n6219)
         );
  INV_X1 U7935 ( .A(n8022), .ZN(n6583) );
  NOR2_X1 U7936 ( .A1(n6583), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6218) );
  AOI211_X1 U7937 ( .C1(n10243), .C2(n7969), .A(n6219), .B(n6218), .ZN(n6229)
         );
  INV_X1 U7938 ( .A(n6226), .ZN(n6222) );
  INV_X1 U7939 ( .A(n6220), .ZN(n6221) );
  AND2_X1 U7940 ( .A1(n6221), .A2(n5198), .ZN(n6223) );
  XNOR2_X1 U7941 ( .A(n7932), .B(n10243), .ZN(n6471) );
  XNOR2_X1 U7942 ( .A(n6471), .B(n8283), .ZN(n6224) );
  OAI21_X1 U7943 ( .B1(n6222), .B2(n6223), .A(n6224), .ZN(n6227) );
  NOR2_X1 U7944 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NAND2_X1 U7945 ( .A1(n6226), .A2(n6225), .ZN(n6473) );
  NAND3_X1 U7946 ( .A1(n6227), .A2(n8016), .A3(n6473), .ZN(n6228) );
  NAND2_X1 U7947 ( .A1(n6229), .A2(n6228), .ZN(P2_U3158) );
  INV_X1 U7948 ( .A(n6238), .ZN(n6232) );
  NAND2_X1 U7949 ( .A1(n6231), .A2(n6230), .ZN(n6387) );
  NAND2_X1 U7950 ( .A1(n6232), .A2(n6387), .ZN(n6390) );
  NAND2_X1 U7951 ( .A1(n7643), .A2(n10080), .ZN(n6233) );
  NAND2_X1 U7952 ( .A1(n6390), .A2(n6233), .ZN(n6285) );
  INV_X1 U7953 ( .A(n7698), .ZN(n6284) );
  NAND2_X1 U7954 ( .A1(n6285), .A2(n6284), .ZN(n6287) );
  NAND2_X1 U7955 ( .A1(n6287), .A2(n6234), .ZN(n6276) );
  XNOR2_X1 U7956 ( .A(n9396), .B(n6342), .ZN(n7702) );
  NAND2_X1 U7957 ( .A1(n6276), .A2(n7702), .ZN(n6275) );
  XNOR2_X1 U7958 ( .A(n9395), .B(n6260), .ZN(n7703) );
  OAI21_X1 U7959 ( .B1(n6235), .B2(n7703), .A(n6251), .ZN(n10052) );
  INV_X1 U7960 ( .A(n6277), .ZN(n6237) );
  INV_X1 U7961 ( .A(n6259), .ZN(n6236) );
  AOI211_X1 U7962 ( .C1(n10046), .C2(n6237), .A(n9664), .B(n6236), .ZN(n10041)
         );
  NAND2_X1 U7963 ( .A1(n6238), .A2(n6393), .ZN(n6392) );
  NAND2_X1 U7964 ( .A1(n7643), .A2(n7642), .ZN(n6239) );
  NAND2_X1 U7965 ( .A1(n6392), .A2(n6239), .ZN(n6292) );
  NAND2_X1 U7966 ( .A1(n6240), .A2(n6672), .ZN(n6241) );
  NAND2_X1 U7967 ( .A1(n9396), .A2(n6342), .ZN(n7640) );
  INV_X1 U7968 ( .A(n9396), .ZN(n6242) );
  NAND2_X1 U7969 ( .A1(n6242), .A2(n6669), .ZN(n6243) );
  XOR2_X1 U7970 ( .A(n7703), .B(n6261), .Z(n6245) );
  AOI21_X1 U7971 ( .B1(n6245), .B2(n9697), .A(n6244), .ZN(n10055) );
  INV_X1 U7972 ( .A(n10055), .ZN(n6246) );
  AOI211_X1 U7973 ( .C1(n10096), .C2(n10052), .A(n10041), .B(n6246), .ZN(n6668) );
  INV_X1 U7974 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6247) );
  OAI22_X1 U7975 ( .A1(n9852), .A2(n6260), .B1(n10100), .B2(n6247), .ZN(n6248)
         );
  INV_X1 U7976 ( .A(n6248), .ZN(n6249) );
  OAI21_X1 U7977 ( .B1(n6668), .B2(n10098), .A(n6249), .ZN(P1_U3465) );
  NAND2_X1 U7978 ( .A1(n6252), .A2(n7612), .ZN(n6255) );
  AOI22_X1 U7979 ( .A1(n7527), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n7526), .B2(
        n9443), .ZN(n6254) );
  INV_X1 U7980 ( .A(n7465), .ZN(n6256) );
  NAND2_X1 U7981 ( .A1(n6488), .A2(n9394), .ZN(n7648) );
  OAI21_X1 U7982 ( .B1(n6257), .B2(n7700), .A(n6317), .ZN(n6329) );
  INV_X1 U7983 ( .A(n6316), .ZN(n6258) );
  AOI211_X1 U7984 ( .C1(n6428), .C2(n6259), .A(n9664), .B(n6258), .ZN(n6336)
         );
  NAND2_X1 U7985 ( .A1(n9395), .A2(n6260), .ZN(n7647) );
  NAND2_X1 U7986 ( .A1(n6262), .A2(n10046), .ZN(n7463) );
  XNOR2_X1 U7987 ( .A(n6300), .B(n7700), .ZN(n6271) );
  NAND2_X1 U7988 ( .A1(n7589), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6270) );
  INV_X1 U7989 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6263) );
  OR2_X1 U7990 ( .A1(n7592), .A2(n6263), .ZN(n6269) );
  OR2_X1 U7991 ( .A1(n6264), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7992 ( .A1(n6306), .A2(n6265), .ZN(n6554) );
  OR2_X1 U7993 ( .A1(n7534), .A2(n6554), .ZN(n6268) );
  OR2_X1 U7994 ( .A1(n7440), .A2(n6266), .ZN(n6267) );
  INV_X1 U7995 ( .A(n6510), .ZN(n9393) );
  AOI22_X1 U7996 ( .A1(n9393), .A2(n9229), .B1(n9296), .B2(n9395), .ZN(n6426)
         );
  OAI21_X1 U7997 ( .B1(n6271), .B2(n9578), .A(n6426), .ZN(n6330) );
  AOI211_X1 U7998 ( .C1(n10096), .C2(n6329), .A(n6336), .B(n6330), .ZN(n6491)
         );
  INV_X1 U7999 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6272) );
  OAI22_X1 U8000 ( .A1(n9852), .A2(n6488), .B1(n10100), .B2(n6272), .ZN(n6273)
         );
  INV_X1 U8001 ( .A(n6273), .ZN(n6274) );
  OAI21_X1 U8002 ( .B1(n6491), .B2(n10098), .A(n6274), .ZN(P1_U3468) );
  OAI21_X1 U8003 ( .B1(n6276), .B2(n7702), .A(n6275), .ZN(n6340) );
  AOI211_X1 U8004 ( .C1(n6669), .C2(n6288), .A(n9664), .B(n6277), .ZN(n6345)
         );
  XNOR2_X1 U8005 ( .A(n6278), .B(n7702), .ZN(n6280) );
  OAI21_X1 U8006 ( .B1(n6280), .B2(n9578), .A(n6279), .ZN(n6346) );
  AOI211_X1 U8007 ( .C1(n10096), .C2(n6340), .A(n6345), .B(n6346), .ZN(n6671)
         );
  OAI22_X1 U8008 ( .A1(n9852), .A2(n6342), .B1(n10100), .B2(n6001), .ZN(n6281)
         );
  INV_X1 U8009 ( .A(n6281), .ZN(n6282) );
  OAI21_X1 U8010 ( .B1(n6671), .B2(n10098), .A(n6282), .ZN(P1_U3462) );
  INV_X1 U8011 ( .A(n6283), .ZN(n10082) );
  OR2_X1 U8012 ( .A1(n6285), .A2(n6284), .ZN(n6286) );
  NAND2_X1 U8013 ( .A1(n6287), .A2(n6286), .ZN(n6405) );
  INV_X1 U8014 ( .A(n6398), .ZN(n6289) );
  INV_X1 U8015 ( .A(n9664), .ZN(n9939) );
  OAI211_X1 U8016 ( .C1(n6289), .C2(n7646), .A(n9939), .B(n6288), .ZN(n6408)
         );
  INV_X1 U8017 ( .A(n6408), .ZN(n6297) );
  INV_X1 U8018 ( .A(n6290), .ZN(n6391) );
  NAND2_X1 U8019 ( .A1(n6405), .A2(n6391), .ZN(n6296) );
  OAI21_X1 U8020 ( .B1(n6292), .B2(n7698), .A(n6291), .ZN(n6294) );
  AOI21_X1 U8021 ( .B1(n6294), .B2(n9697), .A(n6293), .ZN(n6295) );
  NAND2_X1 U8022 ( .A1(n6296), .A2(n6295), .ZN(n6406) );
  AOI211_X1 U8023 ( .C1(n10082), .C2(n6405), .A(n6297), .B(n6406), .ZN(n6674)
         );
  OAI22_X1 U8024 ( .A1(n9852), .A2(n7646), .B1(n10100), .B2(n5947), .ZN(n6298)
         );
  INV_X1 U8025 ( .A(n6298), .ZN(n6299) );
  OAI21_X1 U8026 ( .B1(n6674), .B2(n10098), .A(n6299), .ZN(P1_U3459) );
  NAND2_X1 U8027 ( .A1(n6301), .A2(n7612), .ZN(n6303) );
  AOI22_X1 U8028 ( .A1(n7527), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7526), .B2(
        n9456), .ZN(n6302) );
  NAND2_X1 U8029 ( .A1(n6303), .A2(n6302), .ZN(n6498) );
  OR2_X1 U8030 ( .A1(n6510), .A2(n6498), .ZN(n7461) );
  NAND2_X1 U8031 ( .A1(n6498), .A2(n6510), .ZN(n7467) );
  NAND2_X1 U8032 ( .A1(n7461), .A2(n7467), .ZN(n6318) );
  INV_X1 U8033 ( .A(n6318), .ZN(n6436) );
  XNOR2_X1 U8034 ( .A(n6697), .B(n6436), .ZN(n6315) );
  NAND2_X1 U8035 ( .A1(n7589), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6312) );
  INV_X1 U8036 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6304) );
  OR2_X1 U8037 ( .A1(n7592), .A2(n6304), .ZN(n6311) );
  NAND2_X1 U8038 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  NAND2_X1 U8039 ( .A1(n6445), .A2(n6307), .ZN(n6529) );
  OR2_X1 U8040 ( .A1(n7534), .A2(n6529), .ZN(n6310) );
  OR2_X1 U8041 ( .A1(n7440), .A2(n6308), .ZN(n6309) );
  OR2_X1 U8042 ( .A1(n6504), .A2(n9352), .ZN(n6314) );
  NAND2_X1 U8043 ( .A1(n9394), .A2(n9296), .ZN(n6313) );
  AND2_X1 U8044 ( .A1(n6314), .A2(n6313), .ZN(n6636) );
  OAI21_X1 U8045 ( .B1(n6315), .B2(n9578), .A(n6636), .ZN(n6558) );
  AOI211_X1 U8046 ( .C1(n6498), .C2(n6316), .A(n9664), .B(n6526), .ZN(n6557)
         );
  NOR2_X1 U8047 ( .A1(n6558), .A2(n6557), .ZN(n6494) );
  NAND2_X1 U8048 ( .A1(n6317), .A2(n5016), .ZN(n6319) );
  NAND2_X1 U8049 ( .A1(n6319), .A2(n6318), .ZN(n6464) );
  OAI21_X1 U8050 ( .B1(n6319), .B2(n6318), .A(n6464), .ZN(n6553) );
  INV_X1 U8051 ( .A(n9842), .ZN(n6469) );
  INV_X1 U8052 ( .A(n6498), .ZN(n6641) );
  OAI22_X1 U8053 ( .A1(n9852), .A2(n6641), .B1(n10100), .B2(n6263), .ZN(n6320)
         );
  AOI21_X1 U8054 ( .B1(n6553), .B2(n6469), .A(n6320), .ZN(n6321) );
  OAI21_X1 U8055 ( .B1(n6494), .B2(n10098), .A(n6321), .ZN(P1_U3471) );
  INV_X1 U8056 ( .A(n6322), .ZN(n6433) );
  INV_X1 U8057 ( .A(n6323), .ZN(n6324) );
  NAND3_X1 U8058 ( .A1(n6433), .A2(n6325), .A3(n6324), .ZN(n6331) );
  NOR2_X1 U8059 ( .A1(n5757), .A2(n6326), .ZN(n6327) );
  NAND2_X1 U8060 ( .A1(n10067), .A2(n6327), .ZN(n6412) );
  NAND2_X1 U8061 ( .A1(n10067), .A2(n6391), .ZN(n6328) );
  INV_X1 U8062 ( .A(n6329), .ZN(n6339) );
  NAND2_X1 U8063 ( .A1(n6330), .A2(n10067), .ZN(n6338) );
  NOR2_X1 U8064 ( .A1(n10062), .A2(n6488), .ZN(n6335) );
  OAI22_X1 U8065 ( .A1(n10067), .A2(n6333), .B1(n6431), .B2(n10042), .ZN(n6334) );
  AOI211_X1 U8066 ( .C1(n6336), .C2(n9665), .A(n6335), .B(n6334), .ZN(n6337)
         );
  OAI211_X1 U8067 ( .C1(n9701), .C2(n6339), .A(n6338), .B(n6337), .ZN(P1_U3288) );
  INV_X1 U8068 ( .A(n6340), .ZN(n6349) );
  OAI22_X1 U8069 ( .A1(n10067), .A2(n6341), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10042), .ZN(n6344) );
  NOR2_X1 U8070 ( .A1(n10062), .A2(n6342), .ZN(n6343) );
  AOI211_X1 U8071 ( .C1(n6345), .C2(n9665), .A(n6344), .B(n6343), .ZN(n6348)
         );
  NAND2_X1 U8072 ( .A1(n6346), .A2(n10067), .ZN(n6347) );
  OAI211_X1 U8073 ( .C1(n6349), .C2(n9701), .A(n6348), .B(n6347), .ZN(P1_U3290) );
  INV_X1 U8074 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6350) );
  INV_X1 U8075 ( .A(n7496), .ZN(n6353) );
  INV_X1 U8076 ( .A(n8376), .ZN(n8397) );
  OAI222_X1 U8077 ( .A1(n7278), .A2(n6350), .B1(n8733), .B2(n6353), .C1(
        P2_U3151), .C2(n8397), .ZN(P2_U3279) );
  INV_X1 U8078 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8079 ( .A1(n6351), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U8080 ( .A(n6352), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7497) );
  INV_X1 U8081 ( .A(n7497), .ZN(n10016) );
  OAI222_X1 U8082 ( .A1(n9868), .A2(n6354), .B1(n9872), .B2(n6353), .C1(
        P1_U3086), .C2(n10016), .ZN(P1_U3339) );
  MUX2_X1 U8083 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8426), .Z(n6650) );
  XNOR2_X1 U8084 ( .A(n6650), .B(n6655), .ZN(n6361) );
  MUX2_X1 U8085 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8426), .Z(n6359) );
  MUX2_X1 U8086 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8426), .Z(n6358) );
  AOI21_X1 U8087 ( .B1(n6357), .B2(n6356), .A(n6355), .ZN(n10119) );
  XOR2_X1 U8088 ( .A(n6375), .B(n6358), .Z(n10120) );
  NOR2_X1 U8089 ( .A1(n10119), .A2(n10120), .ZN(n10118) );
  XNOR2_X1 U8090 ( .A(n6359), .B(n6376), .ZN(n10135) );
  NAND2_X1 U8091 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U8092 ( .B1(n6359), .B2(n10140), .A(n10134), .ZN(n6360) );
  AOI211_X1 U8093 ( .C1(n6361), .C2(n6360), .A(n10193), .B(n6649), .ZN(n6386)
         );
  XNOR2_X1 U8094 ( .A(n6375), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U8095 ( .A1(n6362), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6365) );
  INV_X1 U8096 ( .A(n6363), .ZN(n6364) );
  NAND2_X1 U8097 ( .A1(n6365), .A2(n6364), .ZN(n10124) );
  AOI21_X1 U8098 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n10116), .A(n10129), .ZN(
        n6366) );
  INV_X1 U8099 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U8100 ( .A1(n6367), .A2(n10132), .ZN(n6657) );
  NAND2_X1 U8101 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6655), .ZN(n6368) );
  OAI21_X1 U8102 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6655), .A(n6368), .ZN(
        n6656) );
  XNOR2_X1 U8103 ( .A(n6657), .B(n6656), .ZN(n6369) );
  AND2_X1 U8104 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6481) );
  AOI21_X1 U8105 ( .B1(n10127), .B2(n6369), .A(n6481), .ZN(n6370) );
  OAI21_X1 U8106 ( .B1(n10185), .B2(n6655), .A(n6370), .ZN(n6385) );
  INV_X1 U8107 ( .A(n6371), .ZN(n6372) );
  NOR2_X1 U8108 ( .A1(n6373), .A2(n6372), .ZN(n10114) );
  NOR2_X1 U8109 ( .A1(n10114), .A2(n10115), .ZN(n10113) );
  NOR2_X1 U8110 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  INV_X1 U8111 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10215) );
  NAND2_X1 U8112 ( .A1(P2_REG2_REG_4__SCAN_IN), .A2(n6655), .ZN(n6379) );
  OAI21_X1 U8113 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6655), .A(n6379), .ZN(
        n6380) );
  NOR2_X1 U8114 ( .A1(n6381), .A2(n6380), .ZN(n6645) );
  AOI21_X1 U8115 ( .B1(n6381), .B2(n6380), .A(n6645), .ZN(n6383) );
  INV_X1 U8116 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6382) );
  OAI22_X1 U8117 ( .A1(n10191), .A2(n6383), .B1(n10183), .B2(n6382), .ZN(n6384) );
  OR3_X1 U8118 ( .A1(n6386), .A2(n6385), .A3(n6384), .ZN(P2_U3186) );
  INV_X1 U8119 ( .A(n6387), .ZN(n6388) );
  NAND2_X1 U8120 ( .A1(n6238), .A2(n6388), .ZN(n6389) );
  NAND2_X1 U8121 ( .A1(n6390), .A2(n6389), .ZN(n10083) );
  NAND2_X1 U8122 ( .A1(n10083), .A2(n6391), .ZN(n6397) );
  OAI21_X1 U8123 ( .B1(n6393), .B2(n6238), .A(n6392), .ZN(n6395) );
  AOI21_X1 U8124 ( .B1(n6395), .B2(n9697), .A(n6394), .ZN(n6396) );
  AND2_X1 U8125 ( .A1(n6397), .A2(n6396), .ZN(n10085) );
  NOR2_X1 U8126 ( .A1(n10067), .A2(n8866), .ZN(n6401) );
  OAI211_X1 U8127 ( .C1(n10080), .C2(n10061), .A(n9939), .B(n6398), .ZN(n10079) );
  OAI22_X1 U8128 ( .A1(n10049), .A2(n10079), .B1(n6399), .B2(n10042), .ZN(
        n6400) );
  AOI211_X1 U8129 ( .C1(n10047), .C2(n7642), .A(n6401), .B(n6400), .ZN(n6404)
         );
  INV_X1 U8130 ( .A(n6412), .ZN(n6402) );
  NAND2_X1 U8131 ( .A1(n6402), .A2(n10083), .ZN(n6403) );
  OAI211_X1 U8132 ( .C1(n9712), .C2(n10085), .A(n6404), .B(n6403), .ZN(
        P1_U3292) );
  INV_X1 U8133 ( .A(n6405), .ZN(n6413) );
  MUX2_X1 U8134 ( .A(n6406), .B(P1_REG2_REG_2__SCAN_IN), .S(n9712), .Z(n6407)
         );
  INV_X1 U8135 ( .A(n6407), .ZN(n6411) );
  OAI22_X1 U8136 ( .A1(n10049), .A2(n6408), .B1(n9413), .B2(n10042), .ZN(n6409) );
  AOI21_X1 U8137 ( .B1(n10047), .B2(n6672), .A(n6409), .ZN(n6410) );
  OAI211_X1 U8138 ( .C1(n6413), .C2(n6412), .A(n6411), .B(n6410), .ZN(P1_U3291) );
  INV_X1 U8139 ( .A(n6414), .ZN(n6415) );
  INV_X1 U8140 ( .A(n6073), .ZN(n9112) );
  NAND2_X1 U8141 ( .A1(n9394), .A2(n9082), .ZN(n6418) );
  OAI21_X1 U8142 ( .B1(n6488), .B2(n9112), .A(n6418), .ZN(n6419) );
  XNOR2_X1 U8143 ( .A(n6419), .B(n9140), .ZN(n6628) );
  XOR2_X1 U8144 ( .A(n6627), .B(n6628), .Z(n6423) );
  OR2_X1 U8145 ( .A1(n6488), .A2(n9207), .ZN(n6421) );
  NAND2_X1 U8146 ( .A1(n9394), .A2(n9081), .ZN(n6420) );
  NAND2_X1 U8147 ( .A1(n6421), .A2(n6420), .ZN(n6500) );
  INV_X1 U8148 ( .A(n6500), .ZN(n6422) );
  NAND2_X1 U8149 ( .A1(n6423), .A2(n6422), .ZN(n6626) );
  OAI21_X1 U8150 ( .B1(n6423), .B2(n6422), .A(n6626), .ZN(n6424) );
  NAND2_X1 U8151 ( .A1(n6424), .A2(n9931), .ZN(n6430) );
  OAI22_X1 U8152 ( .A1(n9357), .A2(n6426), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6425), .ZN(n6427) );
  AOI21_X1 U8153 ( .B1(n9368), .B2(n6428), .A(n6427), .ZN(n6429) );
  OAI211_X1 U8154 ( .C1(n9935), .C2(n6431), .A(n6430), .B(n6429), .ZN(P1_U3227) );
  NOR2_X4 U8155 ( .A1(n6433), .A2(n6432), .ZN(n10106) );
  NAND2_X1 U8156 ( .A1(n4826), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6434) );
  OAI21_X1 U8157 ( .B1(n6435), .B2(n4826), .A(n6434), .ZN(P1_U3522) );
  NAND2_X1 U8158 ( .A1(n6697), .A2(n6436), .ZN(n6517) );
  OR2_X1 U8159 ( .A1(n6437), .A2(n7521), .ZN(n6439) );
  AOI22_X1 U8160 ( .A1(n7527), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7526), .B2(
        n9469), .ZN(n6438) );
  NAND2_X1 U8161 ( .A1(n6439), .A2(n6438), .ZN(n6532) );
  OR2_X1 U8162 ( .A1(n6532), .A2(n6504), .ZN(n6699) );
  NAND2_X1 U8163 ( .A1(n6532), .A2(n6504), .ZN(n6695) );
  AND2_X1 U8164 ( .A1(n7471), .A2(n7461), .ZN(n6440) );
  NAND2_X1 U8165 ( .A1(n6517), .A2(n6440), .ZN(n6602) );
  NAND2_X1 U8166 ( .A1(n6602), .A2(n6695), .ZN(n6452) );
  NAND2_X1 U8167 ( .A1(n6441), .A2(n7612), .ZN(n6443) );
  AOI22_X1 U8168 ( .A1(n7527), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7526), .B2(
        n9916), .ZN(n6442) );
  NAND2_X1 U8169 ( .A1(n6443), .A2(n6442), .ZN(n6757) );
  NAND2_X1 U8170 ( .A1(n6082), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6451) );
  INV_X1 U8171 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6563) );
  OR2_X1 U8172 ( .A1(n5836), .A2(n6563), .ZN(n6450) );
  NAND2_X1 U8173 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  NAND2_X1 U8174 ( .A1(n6454), .A2(n6446), .ZN(n6787) );
  OR2_X1 U8175 ( .A1(n7534), .A2(n6787), .ZN(n6449) );
  INV_X1 U8176 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6447) );
  OR2_X1 U8177 ( .A1(n7440), .A2(n6447), .ZN(n6448) );
  OR2_X1 U8178 ( .A1(n6757), .A2(n6753), .ZN(n6700) );
  NAND2_X1 U8179 ( .A1(n6757), .A2(n6753), .ZN(n7475) );
  NAND2_X1 U8180 ( .A1(n6700), .A2(n7475), .ZN(n6465) );
  INV_X1 U8181 ( .A(n6465), .ZN(n6601) );
  XNOR2_X1 U8182 ( .A(n6452), .B(n6601), .ZN(n6463) );
  OR2_X1 U8183 ( .A1(n6504), .A2(n9350), .ZN(n6462) );
  NAND2_X1 U8184 ( .A1(n6082), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6460) );
  INV_X1 U8185 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6613) );
  OR2_X1 U8186 ( .A1(n5836), .A2(n6613), .ZN(n6459) );
  OR2_X1 U8187 ( .A1(n7440), .A2(n10104), .ZN(n6458) );
  INV_X1 U8188 ( .A(n6615), .ZN(n6456) );
  NAND2_X1 U8189 ( .A1(n6454), .A2(n6453), .ZN(n6455) );
  NAND2_X1 U8190 ( .A1(n6456), .A2(n6455), .ZN(n6776) );
  OR2_X1 U8191 ( .A1(n7534), .A2(n6776), .ZN(n6457) );
  OR2_X1 U8192 ( .A1(n6763), .A2(n9352), .ZN(n6461) );
  NAND2_X1 U8193 ( .A1(n6462), .A2(n6461), .ZN(n6785) );
  AOI21_X1 U8194 ( .B1(n6463), .B2(n9697), .A(n6785), .ZN(n6570) );
  INV_X1 U8195 ( .A(n6532), .ZN(n10087) );
  INV_X1 U8196 ( .A(n6757), .ZN(n6783) );
  OAI211_X1 U8197 ( .C1(n6527), .C2(n6783), .A(n9939), .B(n6614), .ZN(n6566)
         );
  AND2_X1 U8198 ( .A1(n6570), .A2(n6566), .ZN(n6540) );
  INV_X1 U8199 ( .A(n6504), .ZN(n9392) );
  INV_X1 U8200 ( .A(n7471), .ZN(n6524) );
  NAND2_X1 U8201 ( .A1(n6525), .A2(n6524), .ZN(n6523) );
  OAI21_X1 U8202 ( .B1(n6532), .B2(n9392), .A(n6523), .ZN(n6466) );
  NAND2_X1 U8203 ( .A1(n6466), .A2(n6465), .ZN(n6610) );
  OAI21_X1 U8204 ( .B1(n6466), .B2(n6465), .A(n6610), .ZN(n6568) );
  INV_X1 U8205 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n6467) );
  OAI22_X1 U8206 ( .A1(n6783), .A2(n9852), .B1(n10100), .B2(n6467), .ZN(n6468)
         );
  AOI21_X1 U8207 ( .B1(n6568), .B2(n6469), .A(n6468), .ZN(n6470) );
  OAI21_X1 U8208 ( .B1(n6540), .B2(n10098), .A(n6470), .ZN(P1_U3477) );
  NAND2_X1 U8209 ( .A1(n6471), .A2(n8283), .ZN(n6472) );
  XNOR2_X1 U8210 ( .A(n7896), .B(n10249), .ZN(n6475) );
  NAND2_X1 U8211 ( .A1(n6475), .A2(n6474), .ZN(n6571) );
  INV_X1 U8212 ( .A(n6475), .ZN(n6476) );
  NAND2_X1 U8213 ( .A1(n6476), .A2(n10203), .ZN(n6477) );
  NAND2_X1 U8214 ( .A1(n6571), .A2(n6477), .ZN(n6479) );
  INV_X1 U8215 ( .A(n6572), .ZN(n6478) );
  INV_X1 U8216 ( .A(n10249), .ZN(n8099) );
  NOR2_X1 U8217 ( .A1(n8020), .A2(n6575), .ZN(n6480) );
  AOI211_X1 U8218 ( .C1(n8018), .C2(n8283), .A(n6481), .B(n6480), .ZN(n6482)
         );
  OAI21_X1 U8219 ( .B1(n8099), .B2(n8025), .A(n6482), .ZN(n6483) );
  AOI21_X1 U8220 ( .B1(n6550), .B2(n8022), .A(n6483), .ZN(n6484) );
  OAI21_X1 U8221 ( .B1(n4504), .B2(n7972), .A(n6484), .ZN(P2_U3170) );
  INV_X1 U8222 ( .A(n7513), .ZN(n6562) );
  XNOR2_X1 U8223 ( .A(n6485), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7787) );
  AOI22_X1 U8224 ( .A1(n7787), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6486), .ZN(n6487) );
  OAI21_X1 U8225 ( .B1(n6562), .B2(n9872), .A(n6487), .ZN(P1_U3338) );
  NAND2_X1 U8226 ( .A1(n10106), .A2(n9767), .ZN(n9789) );
  OAI22_X1 U8227 ( .A1(n9789), .A2(n6488), .B1(n10106), .B2(n6125), .ZN(n6489)
         );
  INV_X1 U8228 ( .A(n6489), .ZN(n6490) );
  OAI21_X1 U8229 ( .B1(n6491), .B2(n4826), .A(n6490), .ZN(P1_U3527) );
  NAND2_X1 U8230 ( .A1(n10106), .A2(n10096), .ZN(n9775) );
  INV_X1 U8231 ( .A(n9775), .ZN(n6538) );
  OAI22_X1 U8232 ( .A1(n9789), .A2(n6641), .B1(n10106), .B2(n6266), .ZN(n6492)
         );
  AOI21_X1 U8233 ( .B1(n6553), .B2(n6538), .A(n6492), .ZN(n6493) );
  OAI21_X1 U8234 ( .B1(n6494), .B2(n4826), .A(n6493), .ZN(P1_U3528) );
  NAND2_X1 U8235 ( .A1(n6498), .A2(n4514), .ZN(n6496) );
  OR2_X1 U8236 ( .A1(n6510), .A2(n9207), .ZN(n6495) );
  NAND2_X1 U8237 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  XNOR2_X1 U8238 ( .A(n6497), .B(n9204), .ZN(n6631) );
  AOI22_X1 U8239 ( .A1(n9393), .A2(n9081), .B1(n6498), .B2(n9137), .ZN(n6630)
         );
  NOR2_X1 U8240 ( .A1(n6631), .A2(n6630), .ZN(n6629) );
  INV_X1 U8241 ( .A(n6630), .ZN(n6499) );
  OAI21_X1 U8242 ( .B1(n6628), .B2(n6500), .A(n6499), .ZN(n6501) );
  OAI22_X1 U8243 ( .A1(n10087), .A2(n9112), .B1(n6504), .B2(n9207), .ZN(n6505)
         );
  XOR2_X1 U8244 ( .A(n9140), .B(n6505), .Z(n6507) );
  AOI22_X1 U8245 ( .A1(n6532), .A2(n9082), .B1(n9081), .B2(n9392), .ZN(n6506)
         );
  NAND2_X1 U8246 ( .A1(n6507), .A2(n6506), .ZN(n6750) );
  OAI21_X1 U8247 ( .B1(n6507), .B2(n6506), .A(n6750), .ZN(n6508) );
  AOI21_X1 U8248 ( .B1(n6509), .B2(n6508), .A(n6751), .ZN(n6516) );
  OR2_X1 U8249 ( .A1(n6753), .A2(n9352), .ZN(n6512) );
  OR2_X1 U8250 ( .A1(n6510), .A2(n9350), .ZN(n6511) );
  AND2_X1 U8251 ( .A1(n6512), .A2(n6511), .ZN(n6521) );
  NAND2_X1 U8252 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9466) );
  OAI21_X1 U8253 ( .B1(n9357), .B2(n6521), .A(n9466), .ZN(n6514) );
  NOR2_X1 U8254 ( .A1(n9935), .A2(n6529), .ZN(n6513) );
  AOI211_X1 U8255 ( .C1(n6532), .C2(n9368), .A(n6514), .B(n6513), .ZN(n6515)
         );
  OAI21_X1 U8256 ( .B1(n6516), .B2(n9370), .A(n6515), .ZN(P1_U3213) );
  NAND2_X1 U8257 ( .A1(n6517), .A2(n7461), .ZN(n6518) );
  NAND2_X1 U8258 ( .A1(n6518), .A2(n6524), .ZN(n6519) );
  NAND2_X1 U8259 ( .A1(n6519), .A2(n6602), .ZN(n6520) );
  NAND2_X1 U8260 ( .A1(n6520), .A2(n9697), .ZN(n6522) );
  NAND2_X1 U8261 ( .A1(n6522), .A2(n6521), .ZN(n10089) );
  INV_X1 U8262 ( .A(n10089), .ZN(n6536) );
  OAI21_X1 U8263 ( .B1(n6525), .B2(n6524), .A(n6523), .ZN(n10090) );
  OAI21_X1 U8264 ( .B1(n6526), .B2(n10087), .A(n9939), .ZN(n6528) );
  OR2_X1 U8265 ( .A1(n6528), .A2(n6527), .ZN(n10086) );
  OAI22_X1 U8266 ( .A1(n10067), .A2(n6530), .B1(n6529), .B2(n10042), .ZN(n6531) );
  AOI21_X1 U8267 ( .B1(n10047), .B2(n6532), .A(n6531), .ZN(n6533) );
  OAI21_X1 U8268 ( .B1(n10086), .B2(n10049), .A(n6533), .ZN(n6534) );
  AOI21_X1 U8269 ( .B1(n10090), .B2(n10053), .A(n6534), .ZN(n6535) );
  OAI21_X1 U8270 ( .B1(n9712), .B2(n6536), .A(n6535), .ZN(P1_U3286) );
  OAI22_X1 U8271 ( .A1(n6783), .A2(n9789), .B1(n10106), .B2(n6447), .ZN(n6537)
         );
  AOI21_X1 U8272 ( .B1(n6568), .B2(n6538), .A(n6537), .ZN(n6539) );
  OAI21_X1 U8273 ( .B1(n6540), .B2(n4826), .A(n6539), .ZN(P1_U3530) );
  INV_X1 U8274 ( .A(n8096), .ZN(n6545) );
  XNOR2_X1 U8275 ( .A(n6541), .B(n6545), .ZN(n10248) );
  INV_X1 U8276 ( .A(n10230), .ZN(n6948) );
  INV_X1 U8277 ( .A(n10233), .ZN(n6542) );
  NAND2_X1 U8278 ( .A1(n6948), .A2(n6542), .ZN(n6543) );
  INV_X1 U8279 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6549) );
  XNOR2_X1 U8280 ( .A(n6544), .B(n6545), .ZN(n6548) );
  NAND2_X1 U8281 ( .A1(n8283), .A2(n10204), .ZN(n6546) );
  OAI21_X1 U8282 ( .B1(n6575), .B2(n10221), .A(n6546), .ZN(n6547) );
  AOI21_X1 U8283 ( .B1(n6548), .B2(n10207), .A(n6547), .ZN(n10252) );
  MUX2_X1 U8284 ( .A(n6549), .B(n10252), .S(n8601), .Z(n6552) );
  AOI22_X1 U8285 ( .A1(n10210), .A2(n10249), .B1(n10211), .B2(n6550), .ZN(
        n6551) );
  OAI211_X1 U8286 ( .C1(n10248), .C2(n8605), .A(n6552), .B(n6551), .ZN(
        P2_U3229) );
  INV_X1 U8287 ( .A(n6553), .ZN(n6561) );
  INV_X1 U8288 ( .A(n6554), .ZN(n6638) );
  AOI22_X1 U8289 ( .A1(n9712), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n6638), .B2(
        n10065), .ZN(n6555) );
  OAI21_X1 U8290 ( .B1(n6641), .B2(n10062), .A(n6555), .ZN(n6556) );
  AOI21_X1 U8291 ( .B1(n6557), .B2(n9665), .A(n6556), .ZN(n6560) );
  NAND2_X1 U8292 ( .A1(n6558), .A2(n10067), .ZN(n6559) );
  OAI211_X1 U8293 ( .C1(n6561), .C2(n9701), .A(n6560), .B(n6559), .ZN(P1_U3287) );
  INV_X1 U8294 ( .A(n8414), .ZN(n8424) );
  OAI222_X1 U8295 ( .A1(n7278), .A2(n8967), .B1(n8733), .B2(n6562), .C1(n8424), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OAI22_X1 U8296 ( .A1(n10067), .A2(n6563), .B1(n6787), .B2(n10042), .ZN(n6564) );
  AOI21_X1 U8297 ( .B1(n10047), .B2(n6757), .A(n6564), .ZN(n6565) );
  OAI21_X1 U8298 ( .B1(n6566), .B2(n10049), .A(n6565), .ZN(n6567) );
  AOI21_X1 U8299 ( .B1(n6568), .B2(n10053), .A(n6567), .ZN(n6569) );
  OAI21_X1 U8300 ( .B1(n9712), .B2(n6570), .A(n6569), .ZN(P1_U3285) );
  NAND2_X1 U8301 ( .A1(n6572), .A2(n6571), .ZN(n6590) );
  XNOR2_X1 U8302 ( .A(n7896), .B(n6573), .ZN(n6574) );
  XNOR2_X1 U8303 ( .A(n6574), .B(n6575), .ZN(n6591) );
  XNOR2_X1 U8304 ( .A(n7896), .B(n6690), .ZN(n6739) );
  XNOR2_X1 U8305 ( .A(n6739), .B(n6824), .ZN(n6578) );
  INV_X1 U8306 ( .A(n6574), .ZN(n6576) );
  NAND2_X1 U8307 ( .A1(n6576), .A2(n6575), .ZN(n6579) );
  AND2_X1 U8308 ( .A1(n6578), .A2(n6579), .ZN(n6577) );
  NAND2_X1 U8309 ( .A1(n6741), .A2(n8016), .ZN(n6588) );
  AOI21_X1 U8310 ( .B1(n6589), .B2(n6579), .A(n6578), .ZN(n6587) );
  NAND2_X1 U8311 ( .A1(n8018), .A2(n8282), .ZN(n6581) );
  INV_X1 U8312 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6580) );
  OR2_X1 U8313 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6580), .ZN(n10159) );
  OAI211_X1 U8314 ( .C1(n6962), .C2(n8020), .A(n6581), .B(n10159), .ZN(n6585)
         );
  INV_X1 U8315 ( .A(n6582), .ZN(n6691) );
  NOR2_X1 U8316 ( .A1(n6583), .A2(n6691), .ZN(n6584) );
  AOI211_X1 U8317 ( .C1(n10260), .C2(n7969), .A(n6585), .B(n6584), .ZN(n6586)
         );
  OAI21_X1 U8318 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(P2_U3179) );
  OAI21_X1 U8319 ( .B1(n6591), .B2(n6590), .A(n6589), .ZN(n6597) );
  AND2_X1 U8320 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6654) );
  AOI21_X1 U8321 ( .B1(n8018), .B2(n10203), .A(n6654), .ZN(n6595) );
  NAND2_X1 U8322 ( .A1(n8022), .A2(n6682), .ZN(n6594) );
  NAND2_X1 U8323 ( .A1(n7969), .A2(n10254), .ZN(n6593) );
  OR2_X1 U8324 ( .A1(n8020), .A2(n6824), .ZN(n6592) );
  NAND4_X1 U8325 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6596)
         );
  AOI21_X1 U8326 ( .B1(n6597), .B2(n8016), .A(n6596), .ZN(n6598) );
  INV_X1 U8327 ( .A(n6598), .ZN(P2_U3167) );
  NAND2_X1 U8328 ( .A1(n8285), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6599) );
  OAI21_X1 U8329 ( .B1(n7938), .B2(n8285), .A(n6599), .ZN(P2_U3520) );
  INV_X1 U8330 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6600) );
  INV_X1 U8331 ( .A(n8408), .ZN(n9888) );
  OAI222_X1 U8332 ( .A1(n7278), .A2(n6600), .B1(n8733), .B2(n7522), .C1(n9888), 
        .C2(P2_U3151), .ZN(P2_U3277) );
  NAND3_X1 U8333 ( .A1(n6602), .A2(n6601), .A3(n6695), .ZN(n6603) );
  NAND2_X1 U8334 ( .A1(n6603), .A2(n6700), .ZN(n6607) );
  AOI22_X1 U8335 ( .A1(n7527), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7526), .B2(
        n6604), .ZN(n6605) );
  NAND2_X1 U8336 ( .A1(n10091), .A2(n6763), .ZN(n7489) );
  NAND2_X1 U8337 ( .A1(n7477), .A2(n7489), .ZN(n6611) );
  XNOR2_X1 U8338 ( .A(n6607), .B(n6611), .ZN(n6608) );
  NOR2_X1 U8339 ( .A1(n6753), .A2(n9350), .ZN(n6771) );
  AOI21_X1 U8340 ( .B1(n6608), .B2(n9697), .A(n6771), .ZN(n10093) );
  INV_X1 U8341 ( .A(n6753), .ZN(n9391) );
  NAND2_X1 U8342 ( .A1(n6612), .A2(n6611), .ZN(n6723) );
  OAI21_X1 U8343 ( .B1(n6612), .B2(n6611), .A(n6723), .ZN(n10097) );
  NAND2_X1 U8344 ( .A1(n10097), .A2(n10053), .ZN(n6625) );
  OAI22_X1 U8345 ( .A1(n10067), .A2(n6613), .B1(n6776), .B2(n10042), .ZN(n6623) );
  AOI21_X1 U8346 ( .B1(n6614), .B2(n10091), .A(n9664), .ZN(n6621) );
  NAND2_X1 U8347 ( .A1(n6082), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6620) );
  NAND2_X1 U8348 ( .A1(n7616), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6619) );
  INV_X1 U8349 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6727) );
  OR2_X1 U8350 ( .A1(n5836), .A2(n6727), .ZN(n6618) );
  OR2_X1 U8351 ( .A1(n6615), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6616) );
  NAND2_X1 U8352 ( .A1(n6710), .A2(n6616), .ZN(n9934) );
  OR2_X1 U8353 ( .A1(n7534), .A2(n9934), .ZN(n6617) );
  NAND4_X1 U8354 ( .A1(n6620), .A2(n6619), .A3(n6618), .A4(n6617), .ZN(n9389)
         );
  AND2_X1 U8355 ( .A1(n9389), .A2(n9229), .ZN(n6772) );
  AOI21_X1 U8356 ( .B1(n6621), .B2(n6726), .A(n6772), .ZN(n10092) );
  NOR2_X1 U8357 ( .A1(n10092), .A2(n10049), .ZN(n6622) );
  AOI211_X1 U8358 ( .C1(n10047), .C2(n10091), .A(n6623), .B(n6622), .ZN(n6624)
         );
  OAI211_X1 U8359 ( .C1(n9712), .C2(n10093), .A(n6625), .B(n6624), .ZN(
        P1_U3284) );
  OAI21_X1 U8360 ( .B1(n6628), .B2(n6627), .A(n6626), .ZN(n6633) );
  AOI21_X1 U8361 ( .B1(n6631), .B2(n6630), .A(n6629), .ZN(n6632) );
  XNOR2_X1 U8362 ( .A(n6633), .B(n6632), .ZN(n6634) );
  NAND2_X1 U8363 ( .A1(n6634), .A2(n9931), .ZN(n6640) );
  INV_X1 U8364 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6635) );
  OAI22_X1 U8365 ( .A1(n9357), .A2(n6636), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6635), .ZN(n6637) );
  AOI21_X1 U8366 ( .B1(n9359), .B2(n6638), .A(n6637), .ZN(n6639) );
  OAI211_X1 U8367 ( .C1(n6641), .C2(n9928), .A(n6640), .B(n6639), .ZN(P1_U3239) );
  INV_X1 U8368 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8947) );
  XNOR2_X1 U8369 ( .A(n6642), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10032) );
  INV_X1 U8370 ( .A(n10032), .ZN(n6643) );
  OAI222_X1 U8371 ( .A1(n9868), .A2(n8947), .B1(n6643), .B2(P1_U3086), .C1(
        n9872), .C2(n7522), .ZN(P1_U3337) );
  INV_X1 U8372 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6647) );
  AND2_X1 U8373 ( .A1(n6655), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6644) );
  AOI21_X1 U8374 ( .B1(n6647), .B2(n6646), .A(n6842), .ZN(n6666) );
  MUX2_X1 U8375 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8426), .Z(n6848) );
  XOR2_X1 U8376 ( .A(n6648), .B(n6848), .Z(n6652) );
  AOI211_X1 U8377 ( .C1(n6652), .C2(n6651), .A(n10193), .B(n6846), .ZN(n6653)
         );
  INV_X1 U8378 ( .A(n6653), .ZN(n6665) );
  INV_X1 U8379 ( .A(n10183), .ZN(n10175) );
  INV_X1 U8380 ( .A(n6654), .ZN(n6662) );
  NAND2_X1 U8381 ( .A1(n6658), .A2(n6847), .ZN(n6857) );
  INV_X1 U8382 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10309) );
  AND2_X1 U8383 ( .A1(n6659), .A2(n10309), .ZN(n6660) );
  OAI21_X1 U8384 ( .B1(n6859), .B2(n6660), .A(n10127), .ZN(n6661) );
  OAI211_X1 U8385 ( .C1(n10185), .C2(n6847), .A(n6662), .B(n6661), .ZN(n6663)
         );
  AOI21_X1 U8386 ( .B1(n10175), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6663), .ZN(
        n6664) );
  OAI211_X1 U8387 ( .C1(n6666), .C2(n10191), .A(n6665), .B(n6664), .ZN(
        P2_U3187) );
  AOI22_X1 U8388 ( .A1(n9773), .A2(n10046), .B1(n4826), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U8389 ( .B1(n6668), .B2(n4826), .A(n6667), .ZN(P1_U3526) );
  AOI22_X1 U8390 ( .A1(n9773), .A2(n6669), .B1(n4826), .B2(
        P1_REG1_REG_3__SCAN_IN), .ZN(n6670) );
  OAI21_X1 U8391 ( .B1(n6671), .B2(n4826), .A(n6670), .ZN(P1_U3525) );
  AOI22_X1 U8392 ( .A1(n9773), .A2(n6672), .B1(n4826), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6673) );
  OAI21_X1 U8393 ( .B1(n6674), .B2(n4826), .A(n6673), .ZN(P1_U3524) );
  NAND2_X1 U8394 ( .A1(n6676), .A2(n6675), .ZN(n8038) );
  XNOR2_X1 U8395 ( .A(n6677), .B(n8038), .ZN(n10256) );
  INV_X1 U8396 ( .A(n10256), .ZN(n6685) );
  XOR2_X1 U8397 ( .A(n6678), .B(n8038), .Z(n6680) );
  AOI22_X1 U8398 ( .A1(n8281), .A2(n10202), .B1(n10204), .B2(n10203), .ZN(
        n6679) );
  OAI21_X1 U8399 ( .B1(n6680), .B2(n10225), .A(n6679), .ZN(n6681) );
  AOI21_X1 U8400 ( .B1(n10230), .B2(n10256), .A(n6681), .ZN(n10258) );
  MUX2_X1 U8401 ( .A(n6647), .B(n10258), .S(n8601), .Z(n6684) );
  AOI22_X1 U8402 ( .A1(n10210), .A2(n10254), .B1(n10211), .B2(n6682), .ZN(
        n6683) );
  OAI211_X1 U8403 ( .C1(n6685), .C2(n8451), .A(n6684), .B(n6683), .ZN(P2_U3228) );
  NAND2_X1 U8404 ( .A1(n8112), .A2(n8114), .ZN(n8040) );
  XOR2_X1 U8405 ( .A(n6686), .B(n8040), .Z(n6687) );
  AOI222_X1 U8406 ( .A1(n10207), .A2(n6687), .B1(n8280), .B2(n10202), .C1(
        n8282), .C2(n10204), .ZN(n10263) );
  NAND2_X1 U8407 ( .A1(n6688), .A2(n8110), .ZN(n6689) );
  XOR2_X1 U8408 ( .A(n8040), .B(n6689), .Z(n10261) );
  NOR2_X1 U8409 ( .A1(n8516), .A2(n6690), .ZN(n6693) );
  INV_X1 U8410 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6843) );
  OAI22_X1 U8411 ( .A1(n8601), .A2(n6843), .B1(n6691), .B2(n10217), .ZN(n6692)
         );
  AOI211_X1 U8412 ( .C1(n10261), .C2(n10213), .A(n6693), .B(n6692), .ZN(n6694)
         );
  OAI21_X1 U8413 ( .B1(n10263), .B2(n10235), .A(n6694), .ZN(P2_U3227) );
  NAND2_X1 U8414 ( .A1(n7475), .A2(n6695), .ZN(n7470) );
  NAND2_X1 U8415 ( .A1(n6696), .A2(n7489), .ZN(n6698) );
  NOR2_X1 U8416 ( .A1(n6698), .A2(n4685), .ZN(n7707) );
  NAND2_X1 U8417 ( .A1(n7707), .A2(n6697), .ZN(n6703) );
  INV_X1 U8418 ( .A(n6698), .ZN(n6702) );
  AND2_X1 U8419 ( .A1(n6700), .A2(n6699), .ZN(n7473) );
  AND3_X1 U8420 ( .A1(n7477), .A2(n7473), .A3(n7461), .ZN(n7705) );
  INV_X1 U8421 ( .A(n7705), .ZN(n6701) );
  NAND2_X1 U8422 ( .A1(n6702), .A2(n6701), .ZN(n7650) );
  NAND2_X1 U8423 ( .A1(n6704), .A2(n7612), .ZN(n6706) );
  AOI22_X1 U8424 ( .A1(n7527), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7526), .B2(
        n9902), .ZN(n6705) );
  AND2_X1 U8425 ( .A1(n9929), .A2(n9389), .ZN(n7651) );
  INV_X1 U8426 ( .A(n7651), .ZN(n6708) );
  INV_X1 U8427 ( .A(n9389), .ZN(n6707) );
  XNOR2_X1 U8428 ( .A(n7653), .B(n7706), .ZN(n6721) );
  OR2_X1 U8429 ( .A1(n6763), .A2(n9350), .ZN(n6719) );
  NAND2_X1 U8430 ( .A1(n7589), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8431 ( .A1(n6710), .A2(n6709), .ZN(n6711) );
  NAND2_X1 U8432 ( .A1(n6802), .A2(n6711), .ZN(n9331) );
  OR2_X1 U8433 ( .A1(n7534), .A2(n9331), .ZN(n6716) );
  INV_X1 U8434 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6712) );
  OR2_X1 U8435 ( .A1(n7440), .A2(n6712), .ZN(n6715) );
  INV_X1 U8436 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6713) );
  OR2_X1 U8437 ( .A1(n7592), .A2(n6713), .ZN(n6714) );
  OR2_X1 U8438 ( .A1(n9038), .A2(n9352), .ZN(n6718) );
  NAND2_X1 U8439 ( .A1(n6719), .A2(n6718), .ZN(n9925) );
  INV_X1 U8440 ( .A(n9925), .ZN(n6720) );
  OAI21_X1 U8441 ( .B1(n6721), .B2(n9578), .A(n6720), .ZN(n6733) );
  INV_X1 U8442 ( .A(n6733), .ZN(n6732) );
  INV_X1 U8443 ( .A(n6763), .ZN(n9390) );
  NAND2_X1 U8444 ( .A1(n6724), .A2(n6797), .ZN(n6793) );
  OAI21_X1 U8445 ( .B1(n6724), .B2(n6797), .A(n6793), .ZN(n6735) );
  NAND2_X1 U8446 ( .A1(n6735), .A2(n10053), .ZN(n6731) );
  INV_X1 U8447 ( .A(n6812), .ZN(n6725) );
  AOI211_X1 U8448 ( .C1(n9034), .C2(n6726), .A(n9664), .B(n6725), .ZN(n6734)
         );
  NOR2_X1 U8449 ( .A1(n9929), .A2(n10062), .ZN(n6729) );
  OAI22_X1 U8450 ( .A1(n10067), .A2(n6727), .B1(n9934), .B2(n10042), .ZN(n6728) );
  AOI211_X1 U8451 ( .C1(n6734), .C2(n9665), .A(n6729), .B(n6728), .ZN(n6730)
         );
  OAI211_X1 U8452 ( .C1(n9712), .C2(n6732), .A(n6731), .B(n6730), .ZN(P1_U3283) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8891) );
  INV_X1 U8454 ( .A(n7525), .ZN(n7778) );
  OAI222_X1 U8455 ( .A1(n7278), .A2(n8891), .B1(n8733), .B2(n7778), .C1(
        P2_U3151), .C2(n8431), .ZN(P2_U3276) );
  AOI211_X1 U8456 ( .C1(n6735), .C2(n10096), .A(n6734), .B(n6733), .ZN(n6738)
         );
  AOI22_X1 U8457 ( .A1(n9034), .A2(n9847), .B1(n10098), .B2(
        P1_REG0_REG_10__SCAN_IN), .ZN(n6736) );
  OAI21_X1 U8458 ( .B1(n6738), .B2(n10098), .A(n6736), .ZN(P1_U3483) );
  AOI22_X1 U8459 ( .A1(n9034), .A2(n9773), .B1(n4826), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n6737) );
  OAI21_X1 U8460 ( .B1(n6738), .B2(n4826), .A(n6737), .ZN(P1_U3532) );
  XNOR2_X1 U8461 ( .A(n7896), .B(n6832), .ZN(n6954) );
  XNOR2_X1 U8462 ( .A(n6954), .B(n6962), .ZN(n6744) );
  INV_X1 U8463 ( .A(n6739), .ZN(n6740) );
  INV_X1 U8464 ( .A(n6956), .ZN(n6742) );
  AOI21_X1 U8465 ( .B1(n6744), .B2(n6743), .A(n6742), .ZN(n6749) );
  AND2_X1 U8466 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6853) );
  AOI21_X1 U8467 ( .B1(n8018), .B2(n8281), .A(n6853), .ZN(n6746) );
  NAND2_X1 U8468 ( .A1(n8022), .A2(n6829), .ZN(n6745) );
  OAI211_X1 U8469 ( .C1(n6959), .C2(n8020), .A(n6746), .B(n6745), .ZN(n6747)
         );
  AOI21_X1 U8470 ( .B1(n6832), .B2(n7969), .A(n6747), .ZN(n6748) );
  OAI21_X1 U8471 ( .B1(n6749), .B2(n7972), .A(n6748), .ZN(P2_U3153) );
  NAND2_X1 U8472 ( .A1(n6757), .A2(n4514), .ZN(n6755) );
  OR2_X1 U8473 ( .A1(n6753), .A2(n9207), .ZN(n6754) );
  NAND2_X1 U8474 ( .A1(n6755), .A2(n6754), .ZN(n6756) );
  XNOR2_X1 U8475 ( .A(n6756), .B(n9204), .ZN(n6758) );
  AOI22_X1 U8476 ( .A1(n6757), .A2(n9082), .B1(n9081), .B2(n9391), .ZN(n6782)
         );
  NAND2_X1 U8477 ( .A1(n6781), .A2(n6782), .ZN(n6768) );
  NAND2_X1 U8478 ( .A1(n6759), .A2(n6758), .ZN(n6770) );
  INV_X1 U8479 ( .A(n6770), .ZN(n6766) );
  NAND2_X1 U8480 ( .A1(n10091), .A2(n4514), .ZN(n6761) );
  OR2_X1 U8481 ( .A1(n6763), .A2(n9207), .ZN(n6760) );
  NAND2_X1 U8482 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  XNOR2_X1 U8483 ( .A(n6762), .B(n9140), .ZN(n9027) );
  NOR2_X1 U8484 ( .A1(n6763), .A2(n9201), .ZN(n6764) );
  AOI21_X1 U8485 ( .B1(n10091), .B2(n9137), .A(n6764), .ZN(n9028) );
  XNOR2_X1 U8486 ( .A(n9027), .B(n9028), .ZN(n6769) );
  INV_X1 U8487 ( .A(n6769), .ZN(n6765) );
  NOR2_X1 U8488 ( .A1(n6766), .A2(n6765), .ZN(n6767) );
  NAND2_X1 U8489 ( .A1(n6768), .A2(n6767), .ZN(n9031) );
  NAND2_X1 U8490 ( .A1(n9031), .A2(n9931), .ZN(n6780) );
  AOI21_X1 U8491 ( .B1(n6768), .B2(n6770), .A(n6769), .ZN(n6779) );
  OAI21_X1 U8492 ( .B1(n6772), .B2(n6771), .A(n9926), .ZN(n6775) );
  INV_X1 U8493 ( .A(n6773), .ZN(n6774) );
  OAI211_X1 U8494 ( .C1(n9935), .C2(n6776), .A(n6775), .B(n6774), .ZN(n6777)
         );
  AOI21_X1 U8495 ( .B1(n10091), .B2(n9368), .A(n6777), .ZN(n6778) );
  OAI21_X1 U8496 ( .B1(n6780), .B2(n6779), .A(n6778), .ZN(P1_U3231) );
  OAI21_X1 U8497 ( .B1(n6782), .B2(n6781), .A(n6768), .ZN(n6790) );
  NOR2_X1 U8498 ( .A1(n9928), .A2(n6783), .ZN(n6789) );
  NAND2_X1 U8499 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9917) );
  INV_X1 U8500 ( .A(n9917), .ZN(n6784) );
  AOI21_X1 U8501 ( .B1(n9926), .B2(n6785), .A(n6784), .ZN(n6786) );
  OAI21_X1 U8502 ( .B1(n9935), .B2(n6787), .A(n6786), .ZN(n6788) );
  AOI211_X1 U8503 ( .C1(n6790), .C2(n9931), .A(n6789), .B(n6788), .ZN(n6791)
         );
  INV_X1 U8504 ( .A(n6791), .ZN(P1_U3221) );
  NAND2_X1 U8505 ( .A1(n6794), .A2(n7612), .ZN(n6796) );
  AOI22_X1 U8506 ( .A1(n7527), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7526), .B2(
        n9960), .ZN(n6795) );
  OR2_X1 U8507 ( .A1(n9333), .A2(n9038), .ZN(n7077) );
  AND2_X1 U8508 ( .A1(n9333), .A2(n9038), .ZN(n7078) );
  INV_X1 U8509 ( .A(n7078), .ZN(n7485) );
  NAND2_X1 U8510 ( .A1(n7077), .A2(n7485), .ZN(n7709) );
  XNOR2_X1 U8511 ( .A(n6917), .B(n7709), .ZN(n6837) );
  INV_X1 U8512 ( .A(n6837), .ZN(n6818) );
  INV_X1 U8513 ( .A(n7709), .ZN(n6798) );
  XNOR2_X1 U8514 ( .A(n7079), .B(n6798), .ZN(n6799) );
  NAND2_X1 U8515 ( .A1(n6799), .A2(n9697), .ZN(n6811) );
  NAND2_X1 U8516 ( .A1(n6082), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6807) );
  INV_X1 U8517 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6800) );
  OR2_X1 U8518 ( .A1(n5836), .A2(n6800), .ZN(n6806) );
  AND2_X1 U8519 ( .A1(n6802), .A2(n6801), .ZN(n6803) );
  OR2_X1 U8520 ( .A1(n6803), .A2(n6925), .ZN(n9239) );
  OR2_X1 U8521 ( .A1(n7534), .A2(n9239), .ZN(n6805) );
  OR2_X1 U8522 ( .A1(n7440), .A2(n6975), .ZN(n6804) );
  OR2_X1 U8523 ( .A1(n9042), .A2(n9352), .ZN(n6809) );
  NAND2_X1 U8524 ( .A1(n9389), .A2(n9296), .ZN(n6808) );
  NAND2_X1 U8525 ( .A1(n6809), .A2(n6808), .ZN(n9329) );
  INV_X1 U8526 ( .A(n9329), .ZN(n6810) );
  NAND2_X1 U8527 ( .A1(n6811), .A2(n6810), .ZN(n6835) );
  INV_X1 U8528 ( .A(n9333), .ZN(n6916) );
  AOI211_X1 U8529 ( .C1(n9333), .C2(n6812), .A(n9664), .B(n6919), .ZN(n6836)
         );
  NAND2_X1 U8530 ( .A1(n6836), .A2(n9665), .ZN(n6815) );
  INV_X1 U8531 ( .A(n9331), .ZN(n6813) );
  AOI22_X1 U8532 ( .A1(n9712), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n6813), .B2(
        n10065), .ZN(n6814) );
  OAI211_X1 U8533 ( .C1(n6916), .C2(n10062), .A(n6815), .B(n6814), .ZN(n6816)
         );
  AOI21_X1 U8534 ( .B1(n10067), .B2(n6835), .A(n6816), .ZN(n6817) );
  OAI21_X1 U8535 ( .B1(n6818), .B2(n9701), .A(n6817), .ZN(P1_U3282) );
  INV_X1 U8536 ( .A(n7542), .ZN(n6868) );
  OAI222_X1 U8537 ( .A1(n9872), .A2(n6868), .B1(n7755), .B2(P1_U3086), .C1(
        n7543), .C2(n9868), .ZN(P1_U3335) );
  OR2_X1 U8538 ( .A1(n6819), .A2(n8122), .ZN(n6820) );
  AND2_X1 U8539 ( .A1(n6902), .A2(n6820), .ZN(n6826) );
  INV_X1 U8540 ( .A(n6826), .ZN(n10266) );
  INV_X1 U8541 ( .A(n6822), .ZN(n6823) );
  AOI21_X1 U8542 ( .B1(n8122), .B2(n6821), .A(n6823), .ZN(n6828) );
  OAI22_X1 U8543 ( .A1(n6824), .A2(n10220), .B1(n6959), .B2(n10221), .ZN(n6825) );
  AOI21_X1 U8544 ( .B1(n6826), .B2(n10230), .A(n6825), .ZN(n6827) );
  OAI21_X1 U8545 ( .B1(n6828), .B2(n10225), .A(n6827), .ZN(n10268) );
  NAND2_X1 U8546 ( .A1(n10268), .A2(n8601), .ZN(n6834) );
  INV_X1 U8547 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6845) );
  INV_X1 U8548 ( .A(n6829), .ZN(n6830) );
  OAI22_X1 U8549 ( .A1(n8601), .A2(n6845), .B1(n6830), .B2(n10217), .ZN(n6831)
         );
  AOI21_X1 U8550 ( .B1(n10210), .B2(n6832), .A(n6831), .ZN(n6833) );
  OAI211_X1 U8551 ( .C1(n10266), .C2(n8451), .A(n6834), .B(n6833), .ZN(
        P2_U3226) );
  AOI211_X1 U8552 ( .C1(n6837), .C2(n10096), .A(n6836), .B(n6835), .ZN(n6840)
         );
  AOI22_X1 U8553 ( .A1(n9333), .A2(n9773), .B1(n4826), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n6838) );
  OAI21_X1 U8554 ( .B1(n6840), .B2(n4826), .A(n6838), .ZN(P1_U3533) );
  AOI22_X1 U8555 ( .A1(n9333), .A2(n9847), .B1(n10098), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n6839) );
  OAI21_X1 U8556 ( .B1(n6840), .B2(n10098), .A(n6839), .ZN(P1_U3486) );
  AOI22_X1 U8557 ( .A1(n6860), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n6843), .B2(
        n10155), .ZN(n10154) );
  AOI21_X1 U8558 ( .B1(n6845), .B2(n6844), .A(n6981), .ZN(n6867) );
  MUX2_X1 U8559 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8426), .Z(n6989) );
  XNOR2_X1 U8560 ( .A(n6989), .B(n6996), .ZN(n6852) );
  MUX2_X1 U8561 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8426), .Z(n6849) );
  OR2_X1 U8562 ( .A1(n6849), .A2(n10155), .ZN(n6850) );
  XNOR2_X1 U8563 ( .A(n6849), .B(n6860), .ZN(n10150) );
  NAND2_X1 U8564 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  NAND2_X1 U8565 ( .A1(n6850), .A2(n10149), .ZN(n6851) );
  NAND2_X1 U8566 ( .A1(n6852), .A2(n6851), .ZN(n6987) );
  OAI21_X1 U8567 ( .B1(n6852), .B2(n6851), .A(n6987), .ZN(n6865) );
  INV_X1 U8568 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n6856) );
  OR2_X1 U8569 ( .A1(n10185), .A2(n6988), .ZN(n6855) );
  INV_X1 U8570 ( .A(n6853), .ZN(n6854) );
  OAI211_X1 U8571 ( .C1(n10183), .C2(n6856), .A(n6855), .B(n6854), .ZN(n6864)
         );
  INV_X1 U8572 ( .A(n6857), .ZN(n6858) );
  INV_X1 U8573 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U8574 ( .A1(n6860), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10311), .B2(
        n10155), .ZN(n10148) );
  INV_X1 U8575 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10313) );
  AOI21_X1 U8576 ( .B1(n6861), .B2(n10313), .A(n6997), .ZN(n6862) );
  NOR2_X1 U8577 ( .A1(n6862), .A2(n10199), .ZN(n6863) );
  AOI211_X1 U8578 ( .C1(n10167), .C2(n6865), .A(n6864), .B(n6863), .ZN(n6866)
         );
  OAI21_X1 U8579 ( .B1(n6867), .B2(n10191), .A(n6866), .ZN(P2_U3189) );
  OAI222_X1 U8580 ( .A1(n7278), .A2(n6869), .B1(n8733), .B2(n6868), .C1(n8260), 
        .C2(P2_U3151), .ZN(P2_U3275) );
  XNOR2_X1 U8581 ( .A(n7787), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n7788) );
  XNOR2_X1 U8582 ( .A(n9969), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n9965) );
  OR2_X1 U8583 ( .A1(n6913), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U8584 ( .A1(n6871), .A2(n6870), .ZN(n9964) );
  NOR2_X1 U8585 ( .A1(n9965), .A2(n9964), .ZN(n9966) );
  AOI21_X1 U8586 ( .B1(n9969), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9966), .ZN(
        n9981) );
  XNOR2_X1 U8587 ( .A(n9986), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U8588 ( .A1(n9981), .A2(n9982), .ZN(n9983) );
  AOI21_X1 U8589 ( .B1(n9986), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9983), .ZN(
        n6872) );
  NOR2_X1 U8590 ( .A1(n6872), .A2(n6878), .ZN(n6873) );
  INV_X1 U8591 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9999) );
  XNOR2_X1 U8592 ( .A(n6878), .B(n6872), .ZN(n10000) );
  NOR2_X1 U8593 ( .A1(n9999), .A2(n10000), .ZN(n9998) );
  NOR2_X1 U8594 ( .A1(n6873), .A2(n9998), .ZN(n10013) );
  INV_X1 U8595 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9781) );
  XNOR2_X1 U8596 ( .A(n7497), .B(n9781), .ZN(n10014) );
  AOI22_X1 U8597 ( .A1(n10013), .A2(n10014), .B1(n10016), .B2(n9781), .ZN(
        n7789) );
  XOR2_X1 U8598 ( .A(n7788), .B(n7789), .Z(n6889) );
  INV_X1 U8599 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6874) );
  XNOR2_X1 U8600 ( .A(n7787), .B(n6874), .ZN(n6883) );
  NAND2_X1 U8601 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n9969), .ZN(n6875) );
  OAI21_X1 U8602 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9969), .A(n6875), .ZN(
        n9972) );
  OAI21_X1 U8603 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6913), .A(n6876), .ZN(
        n9971) );
  NOR2_X1 U8604 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  AOI21_X1 U8605 ( .B1(n9969), .B2(P1_REG2_REG_13__SCAN_IN), .A(n9970), .ZN(
        n9988) );
  NAND2_X1 U8606 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9986), .ZN(n6877) );
  OAI21_X1 U8607 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9986), .A(n6877), .ZN(
        n9989) );
  NOR2_X1 U8608 ( .A1(n9988), .A2(n9989), .ZN(n9987) );
  AOI21_X1 U8609 ( .B1(n9986), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9987), .ZN(
        n6879) );
  NOR2_X1 U8610 ( .A1(n6879), .A2(n6878), .ZN(n6880) );
  INV_X1 U8611 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10002) );
  XOR2_X1 U8612 ( .A(n10006), .B(n6879), .Z(n10003) );
  NOR2_X1 U8613 ( .A1(n10002), .A2(n10003), .ZN(n10001) );
  NOR2_X1 U8614 ( .A1(n6880), .A2(n10001), .ZN(n10012) );
  XNOR2_X1 U8615 ( .A(n7497), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n10011) );
  NAND2_X1 U8616 ( .A1(n7497), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6881) );
  NAND2_X1 U8617 ( .A1(n6882), .A2(n6883), .ZN(n7783) );
  OAI21_X1 U8618 ( .B1(n6883), .B2(n6882), .A(n7783), .ZN(n6884) );
  NAND2_X1 U8619 ( .A1(n6884), .A2(n10024), .ZN(n6888) );
  INV_X1 U8620 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U8621 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9275) );
  OAI21_X1 U8622 ( .B1(n10039), .B2(n6885), .A(n9275), .ZN(n6886) );
  AOI21_X1 U8623 ( .B1(n7787), .B2(n10031), .A(n6886), .ZN(n6887) );
  OAI211_X1 U8624 ( .C1(n10028), .C2(n6889), .A(n6888), .B(n6887), .ZN(
        P1_U3260) );
  NAND2_X1 U8625 ( .A1(n6890), .A2(n6892), .ZN(n6891) );
  NAND2_X1 U8626 ( .A1(n6942), .A2(n6891), .ZN(n10278) );
  INV_X1 U8627 ( .A(n6892), .ZN(n8043) );
  XNOR2_X1 U8628 ( .A(n6893), .B(n8043), .ZN(n6894) );
  NAND2_X1 U8629 ( .A1(n6894), .A2(n10207), .ZN(n6896) );
  AOI22_X1 U8630 ( .A1(n8279), .A2(n10204), .B1(n10202), .B2(n8277), .ZN(n6895) );
  OAI211_X1 U8631 ( .C1(n6948), .C2(n10278), .A(n6896), .B(n6895), .ZN(n10280)
         );
  NAND2_X1 U8632 ( .A1(n10280), .A2(n8601), .ZN(n6900) );
  INV_X1 U8633 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6984) );
  INV_X1 U8634 ( .A(n7071), .ZN(n6897) );
  OAI22_X1 U8635 ( .A1(n8601), .A2(n6984), .B1(n6897), .B2(n10217), .ZN(n6898)
         );
  AOI21_X1 U8636 ( .B1(n10210), .B2(n7062), .A(n6898), .ZN(n6899) );
  OAI211_X1 U8637 ( .C1(n10278), .C2(n8451), .A(n6900), .B(n6899), .ZN(
        P2_U3224) );
  INV_X1 U8638 ( .A(n7558), .ZN(n6938) );
  OAI222_X1 U8639 ( .A1(n9872), .A2(n6938), .B1(n7699), .B2(P1_U3086), .C1(
        n8932), .C2(n9868), .ZN(P1_U3334) );
  NAND2_X1 U8640 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  XOR2_X1 U8641 ( .A(n8041), .B(n6903), .Z(n10270) );
  NOR2_X1 U8642 ( .A1(n6962), .A2(n10220), .ZN(n6909) );
  INV_X1 U8643 ( .A(n6904), .ZN(n6907) );
  AOI21_X1 U8644 ( .B1(n6822), .B2(n6905), .A(n8041), .ZN(n6906) );
  NOR3_X1 U8645 ( .A1(n6907), .A2(n6906), .A3(n10225), .ZN(n6908) );
  AOI211_X1 U8646 ( .C1(n10202), .C2(n8278), .A(n6909), .B(n6908), .ZN(n10271)
         );
  MUX2_X1 U8647 ( .A(n8810), .B(n10271), .S(n8601), .Z(n6911) );
  AOI22_X1 U8648 ( .A1(n10210), .A2(n6957), .B1(n10211), .B2(n6964), .ZN(n6910) );
  OAI211_X1 U8649 ( .C1(n10270), .C2(n8605), .A(n6911), .B(n6910), .ZN(
        P2_U3225) );
  NAND2_X1 U8650 ( .A1(n6912), .A2(n7612), .ZN(n6915) );
  AOI22_X1 U8651 ( .A1(n7527), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7526), .B2(
        n6913), .ZN(n6914) );
  XOR2_X1 U8652 ( .A(n9241), .B(n9387), .Z(n7710) );
  INV_X1 U8653 ( .A(n9038), .ZN(n9388) );
  NAND2_X1 U8654 ( .A1(n6917), .A2(n5006), .ZN(n6918) );
  XOR2_X1 U8655 ( .A(n7090), .B(n7710), .Z(n6970) );
  INV_X1 U8656 ( .A(n6919), .ZN(n6921) );
  INV_X1 U8657 ( .A(n9241), .ZN(n7091) );
  INV_X1 U8658 ( .A(n7093), .ZN(n6920) );
  AOI21_X1 U8659 ( .B1(n9241), .B2(n6921), .A(n6920), .ZN(n6967) );
  NOR2_X1 U8660 ( .A1(n10049), .A2(n9664), .ZN(n10060) );
  INV_X1 U8661 ( .A(n9239), .ZN(n6922) );
  AOI22_X1 U8662 ( .A1(n9712), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6922), .B2(
        n10065), .ZN(n6923) );
  OAI21_X1 U8663 ( .B1(n7091), .B2(n10062), .A(n6923), .ZN(n6936) );
  OAI21_X1 U8664 ( .B1(n7079), .B2(n7078), .A(n7077), .ZN(n6924) );
  XNOR2_X1 U8665 ( .A(n6924), .B(n7710), .ZN(n6934) );
  NAND2_X1 U8666 ( .A1(n6082), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6931) );
  INV_X1 U8667 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7094) );
  OR2_X1 U8668 ( .A1(n5836), .A2(n7094), .ZN(n6930) );
  NOR2_X1 U8669 ( .A1(n6925), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6926) );
  OR2_X1 U8670 ( .A1(n7080), .A2(n6926), .ZN(n9307) );
  OR2_X1 U8671 ( .A1(n7534), .A2(n9307), .ZN(n6929) );
  INV_X1 U8672 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6927) );
  OR2_X1 U8673 ( .A1(n7440), .A2(n6927), .ZN(n6928) );
  OR2_X1 U8674 ( .A1(n9050), .A2(n9352), .ZN(n6933) );
  OR2_X1 U8675 ( .A1(n9038), .A2(n9350), .ZN(n6932) );
  NAND2_X1 U8676 ( .A1(n6933), .A2(n6932), .ZN(n9236) );
  AOI21_X1 U8677 ( .B1(n6934), .B2(n9697), .A(n9236), .ZN(n6969) );
  INV_X1 U8678 ( .A(n10067), .ZN(n9581) );
  NOR2_X1 U8679 ( .A1(n6969), .A2(n9581), .ZN(n6935) );
  AOI211_X1 U8680 ( .C1(n6967), .C2(n10060), .A(n6936), .B(n6935), .ZN(n6937)
         );
  OAI21_X1 U8681 ( .B1(n6970), .B2(n9701), .A(n6937), .ZN(P1_U3281) );
  OAI222_X1 U8682 ( .A1(P2_U3151), .A2(n6939), .B1(n8733), .B2(n6938), .C1(
        n8840), .C2(n7278), .ZN(P2_U3274) );
  INV_X1 U8683 ( .A(n7570), .ZN(n7780) );
  OAI222_X1 U8684 ( .A1(n7278), .A2(n6941), .B1(n8733), .B2(n7780), .C1(
        P2_U3151), .C2(n6940), .ZN(P2_U3273) );
  NAND2_X1 U8685 ( .A1(n6942), .A2(n8119), .ZN(n6943) );
  XNOR2_X1 U8686 ( .A(n6943), .B(n8044), .ZN(n10285) );
  XOR2_X1 U8687 ( .A(n6944), .B(n8044), .Z(n6945) );
  NAND2_X1 U8688 ( .A1(n6945), .A2(n10207), .ZN(n6947) );
  AOI22_X1 U8689 ( .A1(n8276), .A2(n10202), .B1(n10204), .B2(n8278), .ZN(n6946) );
  OAI211_X1 U8690 ( .C1(n10285), .C2(n6948), .A(n6947), .B(n6946), .ZN(n10287)
         );
  NAND2_X1 U8691 ( .A1(n10287), .A2(n8601), .ZN(n6953) );
  INV_X1 U8692 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6950) );
  INV_X1 U8693 ( .A(n7176), .ZN(n6949) );
  OAI22_X1 U8694 ( .A1(n8601), .A2(n6950), .B1(n6949), .B2(n10217), .ZN(n6951)
         );
  AOI21_X1 U8695 ( .B1(n10210), .B2(n7181), .A(n6951), .ZN(n6952) );
  OAI211_X1 U8696 ( .C1(n10285), .C2(n8451), .A(n6953), .B(n6952), .ZN(
        P2_U3223) );
  NAND2_X1 U8697 ( .A1(n6954), .A2(n6962), .ZN(n6955) );
  NAND2_X1 U8698 ( .A1(n6956), .A2(n6955), .ZN(n7061) );
  XNOR2_X1 U8699 ( .A(n6957), .B(n4415), .ZN(n7059) );
  NAND2_X1 U8700 ( .A1(n6958), .A2(n6959), .ZN(n7066) );
  OAI21_X1 U8701 ( .B1(n6959), .B2(n6958), .A(n7066), .ZN(n6960) );
  NAND2_X1 U8702 ( .A1(n6960), .A2(n8016), .ZN(n6966) );
  INV_X1 U8703 ( .A(n8020), .ZN(n7997) );
  INV_X1 U8704 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8935) );
  NOR2_X1 U8705 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8935), .ZN(n10176) );
  AOI21_X1 U8706 ( .B1(n7997), .B2(n8278), .A(n10176), .ZN(n6961) );
  OAI21_X1 U8707 ( .B1(n6962), .B2(n7999), .A(n6961), .ZN(n6963) );
  AOI21_X1 U8708 ( .B1(n6964), .B2(n8022), .A(n6963), .ZN(n6965) );
  OAI211_X1 U8709 ( .C1(n10272), .C2(n8025), .A(n6966), .B(n6965), .ZN(
        P2_U3161) );
  INV_X1 U8710 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6972) );
  AOI22_X1 U8711 ( .A1(n6967), .A2(n9939), .B1(n9767), .B2(n9241), .ZN(n6968)
         );
  OAI211_X1 U8712 ( .C1(n6970), .C2(n9778), .A(n6969), .B(n6968), .ZN(n6973)
         );
  NAND2_X1 U8713 ( .A1(n6973), .A2(n10100), .ZN(n6971) );
  OAI21_X1 U8714 ( .B1(n10100), .B2(n6972), .A(n6971), .ZN(P1_U3489) );
  NAND2_X1 U8715 ( .A1(n6973), .A2(n10106), .ZN(n6974) );
  OAI21_X1 U8716 ( .B1(n10106), .B2(n6975), .A(n6974), .ZN(P1_U3534) );
  INV_X1 U8717 ( .A(n7583), .ZN(n6977) );
  NAND2_X1 U8718 ( .A1(n9020), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6976) );
  OAI211_X1 U8719 ( .C1(n6977), .C2(n8733), .A(n8267), .B(n6976), .ZN(P2_U3272) );
  NAND2_X1 U8720 ( .A1(n7583), .A2(n6978), .ZN(n6979) );
  OAI211_X1 U8721 ( .C1(n8814), .C2(n9868), .A(n6979), .B(n7768), .ZN(P1_U3332) );
  NOR2_X1 U8722 ( .A1(n6996), .A2(n6980), .ZN(n6982) );
  INV_X1 U8723 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8810) );
  AOI22_X1 U8724 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6999), .B1(n10171), .B2(
        n8810), .ZN(n10170) );
  AOI21_X1 U8725 ( .B1(n6984), .B2(n6983), .A(n7306), .ZN(n7006) );
  MUX2_X1 U8726 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8426), .Z(n6985) );
  INV_X1 U8727 ( .A(n9021), .ZN(n6994) );
  NOR2_X1 U8728 ( .A1(n6985), .A2(n6994), .ZN(n7315) );
  AND2_X1 U8729 ( .A1(n6985), .A2(n6994), .ZN(n7314) );
  NOR2_X1 U8730 ( .A1(n7315), .A2(n7314), .ZN(n6991) );
  MUX2_X1 U8731 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8426), .Z(n6986) );
  OR2_X1 U8732 ( .A1(n6986), .A2(n10171), .ZN(n6990) );
  XNOR2_X1 U8733 ( .A(n6986), .B(n6999), .ZN(n10165) );
  OAI21_X1 U8734 ( .B1(n6989), .B2(n6988), .A(n6987), .ZN(n10166) );
  NAND2_X1 U8735 ( .A1(n10165), .A2(n10166), .ZN(n10164) );
  NAND2_X1 U8736 ( .A1(n6990), .A2(n10164), .ZN(n7316) );
  XNOR2_X1 U8737 ( .A(n6991), .B(n7316), .ZN(n6992) );
  NAND2_X1 U8738 ( .A1(n6992), .A2(n10167), .ZN(n7005) );
  AND2_X1 U8739 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7068) );
  INV_X1 U8740 ( .A(n7068), .ZN(n6993) );
  OAI21_X1 U8741 ( .B1(n10185), .B2(n6994), .A(n6993), .ZN(n7003) );
  NOR2_X1 U8742 ( .A1(n6996), .A2(n6995), .ZN(n6998) );
  INV_X1 U8743 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10315) );
  AOI22_X1 U8744 ( .A1(P2_REG1_REG_8__SCAN_IN), .A2(n6999), .B1(n10171), .B2(
        n10315), .ZN(n10163) );
  INV_X1 U8745 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10317) );
  AOI21_X1 U8746 ( .B1(n7000), .B2(n10317), .A(n7331), .ZN(n7001) );
  NOR2_X1 U8747 ( .A1(n7001), .A2(n10199), .ZN(n7002) );
  AOI211_X1 U8748 ( .C1(n10175), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7003), .B(
        n7002), .ZN(n7004) );
  OAI211_X1 U8749 ( .C1(n7006), .C2(n10191), .A(n7005), .B(n7004), .ZN(
        P2_U3191) );
  INV_X1 U8750 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U8751 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7045) );
  NOR2_X1 U8752 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7043) );
  NOR2_X1 U8753 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7041) );
  NOR2_X1 U8754 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7039) );
  NOR2_X1 U8755 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7037) );
  NOR2_X1 U8756 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7035) );
  INV_X1 U8757 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7007) );
  INV_X1 U8758 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7346) );
  AOI22_X1 U8759 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n7007), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n7346), .ZN(n10345) );
  NAND2_X1 U8760 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7033) );
  INV_X1 U8761 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9963) );
  INV_X1 U8762 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7367) );
  AOI22_X1 U8763 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .B1(n9963), .B2(n7367), .ZN(n10347) );
  NAND2_X1 U8764 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7031) );
  XOR2_X1 U8765 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P2_ADDR_REG_10__SCAN_IN), 
        .Z(n10349) );
  NOR2_X1 U8766 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7015) );
  XNOR2_X1 U8767 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10362) );
  NAND2_X1 U8768 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7013) );
  XOR2_X1 U8769 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10360) );
  NAND2_X1 U8770 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7011) );
  AOI21_X1 U8771 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10326) );
  NAND2_X1 U8772 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7008) );
  NOR2_X1 U8773 ( .A1(n8964), .A2(n7008), .ZN(n10327) );
  NOR2_X1 U8774 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10327), .ZN(n7009) );
  NOR2_X1 U8775 ( .A1(n10326), .A2(n7009), .ZN(n10358) );
  XOR2_X1 U8776 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10357) );
  NAND2_X1 U8777 ( .A1(n10358), .A2(n10357), .ZN(n7010) );
  NAND2_X1 U8778 ( .A1(n7011), .A2(n7010), .ZN(n10359) );
  NAND2_X1 U8779 ( .A1(n10360), .A2(n10359), .ZN(n7012) );
  NAND2_X1 U8780 ( .A1(n7013), .A2(n7012), .ZN(n10361) );
  NOR2_X1 U8781 ( .A1(n10362), .A2(n10361), .ZN(n7014) );
  NOR2_X1 U8782 ( .A1(n7015), .A2(n7014), .ZN(n7016) );
  NOR2_X1 U8783 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n7016), .ZN(n10351) );
  NAND2_X1 U8784 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n7018), .ZN(n7020) );
  XOR2_X1 U8785 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n7018), .Z(n10356) );
  NAND2_X1 U8786 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10356), .ZN(n7019) );
  NAND2_X1 U8787 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  NAND2_X1 U8788 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7021), .ZN(n7023) );
  XOR2_X1 U8789 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7021), .Z(n10354) );
  NAND2_X1 U8790 ( .A1(n10354), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8791 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8792 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7024), .ZN(n7026) );
  XOR2_X1 U8793 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7024), .Z(n10355) );
  NAND2_X1 U8794 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10355), .ZN(n7025) );
  NAND2_X1 U8795 ( .A1(n7026), .A2(n7025), .ZN(n7027) );
  NAND2_X1 U8796 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7027), .ZN(n7029) );
  XOR2_X1 U8797 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7027), .Z(n10353) );
  NAND2_X1 U8798 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10353), .ZN(n7028) );
  NAND2_X1 U8799 ( .A1(n7029), .A2(n7028), .ZN(n10348) );
  NAND2_X1 U8800 ( .A1(n10349), .A2(n10348), .ZN(n7030) );
  NAND2_X1 U8801 ( .A1(n7031), .A2(n7030), .ZN(n10346) );
  NAND2_X1 U8802 ( .A1(n10347), .A2(n10346), .ZN(n7032) );
  NAND2_X1 U8803 ( .A1(n7033), .A2(n7032), .ZN(n10344) );
  INV_X1 U8804 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9980) );
  INV_X1 U8805 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8304) );
  AOI22_X1 U8806 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(n9980), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n8304), .ZN(n10342) );
  INV_X1 U8807 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9997) );
  INV_X1 U8808 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8325) );
  AOI22_X1 U8809 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9997), .B1(
        P1_ADDR_REG_14__SCAN_IN), .B2(n8325), .ZN(n10340) );
  INV_X1 U8810 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10009) );
  INV_X1 U8811 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8349) );
  AOI22_X1 U8812 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n10009), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n8349), .ZN(n10338) );
  NOR2_X1 U8813 ( .A1(n10339), .A2(n10338), .ZN(n7040) );
  NOR2_X1 U8814 ( .A1(n7041), .A2(n7040), .ZN(n10337) );
  INV_X1 U8815 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10023) );
  INV_X1 U8816 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8371) );
  AOI22_X1 U8817 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n10023), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n8371), .ZN(n10336) );
  NOR2_X1 U8818 ( .A1(n10337), .A2(n10336), .ZN(n7042) );
  NOR2_X1 U8819 ( .A1(n7043), .A2(n7042), .ZN(n10335) );
  INV_X1 U8820 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9002) );
  AOI22_X1 U8821 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n6885), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9002), .ZN(n10334) );
  NOR2_X1 U8822 ( .A1(n10335), .A2(n10334), .ZN(n7044) );
  NAND2_X1 U8823 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10331), .ZN(n7046) );
  NOR2_X1 U8824 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10331), .ZN(n10330) );
  AOI21_X1 U8825 ( .B1(n10332), .B2(n7046), .A(n10330), .ZN(n7048) );
  XNOR2_X1 U8826 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7047) );
  XNOR2_X1 U8827 ( .A(n7048), .B(n7047), .ZN(ADD_1068_U4) );
  XNOR2_X1 U8828 ( .A(n7049), .B(n8134), .ZN(n10289) );
  NAND2_X1 U8829 ( .A1(n7051), .A2(n7050), .ZN(n7052) );
  XNOR2_X1 U8830 ( .A(n7052), .B(n8134), .ZN(n7053) );
  OAI222_X1 U8831 ( .A1(n10221), .A2(n8148), .B1(n10220), .B2(n7114), .C1(
        n7053), .C2(n10225), .ZN(n10290) );
  NAND2_X1 U8832 ( .A1(n10290), .A2(n8601), .ZN(n7058) );
  INV_X1 U8833 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7055) );
  INV_X1 U8834 ( .A(n7236), .ZN(n7054) );
  OAI22_X1 U8835 ( .A1(n8601), .A2(n7055), .B1(n7054), .B2(n10217), .ZN(n7056)
         );
  AOI21_X1 U8836 ( .B1(n10210), .B2(n10292), .A(n7056), .ZN(n7057) );
  OAI211_X1 U8837 ( .C1(n8605), .C2(n10289), .A(n7058), .B(n7057), .ZN(
        P2_U3222) );
  INV_X1 U8838 ( .A(n7059), .ZN(n7060) );
  NAND2_X1 U8839 ( .A1(n7061), .A2(n7060), .ZN(n7065) );
  XNOR2_X1 U8840 ( .A(n7062), .B(n4415), .ZN(n7113) );
  XNOR2_X1 U8841 ( .A(n7113), .B(n7179), .ZN(n7064) );
  AND2_X1 U8842 ( .A1(n7065), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U8843 ( .A1(n7066), .A2(n7063), .ZN(n7121) );
  INV_X1 U8844 ( .A(n7121), .ZN(n7172) );
  AOI21_X1 U8845 ( .B1(n7066), .B2(n7065), .A(n7064), .ZN(n7067) );
  OR3_X1 U8846 ( .A1(n7172), .A2(n7067), .A3(n7972), .ZN(n7073) );
  AOI21_X1 U8847 ( .B1(n8018), .B2(n8279), .A(n7068), .ZN(n7069) );
  OAI21_X1 U8848 ( .B1(n7114), .B2(n8020), .A(n7069), .ZN(n7070) );
  AOI21_X1 U8849 ( .B1(n7071), .B2(n8022), .A(n7070), .ZN(n7072) );
  OAI211_X1 U8850 ( .C1(n10277), .C2(n8025), .A(n7073), .B(n7072), .ZN(
        P2_U3171) );
  NAND2_X1 U8851 ( .A1(n7074), .A2(n7612), .ZN(n7076) );
  AOI22_X1 U8852 ( .A1(n7527), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7526), .B2(
        n9969), .ZN(n7075) );
  XNOR2_X1 U8853 ( .A(n9309), .B(n9386), .ZN(n7712) );
  OR2_X1 U8854 ( .A1(n9241), .A2(n9042), .ZN(n7482) );
  AND2_X1 U8855 ( .A1(n7482), .A2(n7077), .ZN(n7654) );
  AND2_X1 U8856 ( .A1(n9241), .A2(n9042), .ZN(n7481) );
  AOI21_X1 U8857 ( .B1(n7654), .B2(n7078), .A(n7481), .ZN(n7637) );
  XOR2_X1 U8858 ( .A(n7712), .B(n7147), .Z(n7089) );
  OR2_X1 U8859 ( .A1(n9042), .A2(n9350), .ZN(n7087) );
  INV_X1 U8860 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7163) );
  OR2_X1 U8861 ( .A1(n5836), .A2(n7163), .ZN(n7085) );
  INV_X1 U8862 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9850) );
  OR2_X1 U8863 ( .A1(n7592), .A2(n9850), .ZN(n7084) );
  OR2_X1 U8864 ( .A1(n7080), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7081) );
  NAND2_X1 U8865 ( .A1(n7151), .A2(n7081), .ZN(n9176) );
  OR2_X1 U8866 ( .A1(n7534), .A2(n9176), .ZN(n7083) );
  INV_X1 U8867 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9787) );
  OR2_X1 U8868 ( .A1(n7440), .A2(n9787), .ZN(n7082) );
  OR2_X1 U8869 ( .A1(n9057), .A2(n9352), .ZN(n7086) );
  NAND2_X1 U8870 ( .A1(n7087), .A2(n7086), .ZN(n9305) );
  INV_X1 U8871 ( .A(n9305), .ZN(n7088) );
  OAI21_X1 U8872 ( .B1(n7089), .B2(n9578), .A(n7088), .ZN(n7107) );
  INV_X1 U8873 ( .A(n7107), .ZN(n7099) );
  XOR2_X1 U8874 ( .A(n7712), .B(n7159), .Z(n7109) );
  NAND2_X1 U8875 ( .A1(n7109), .A2(n10053), .ZN(n7098) );
  INV_X1 U8876 ( .A(n7162), .ZN(n7092) );
  AOI211_X1 U8877 ( .C1(n9309), .C2(n7093), .A(n9664), .B(n7092), .ZN(n7108)
         );
  INV_X1 U8878 ( .A(n9309), .ZN(n7160) );
  NOR2_X1 U8879 ( .A1(n7160), .A2(n10062), .ZN(n7096) );
  OAI22_X1 U8880 ( .A1(n10067), .A2(n7094), .B1(n9307), .B2(n10042), .ZN(n7095) );
  AOI211_X1 U8881 ( .C1(n7108), .C2(n9665), .A(n7096), .B(n7095), .ZN(n7097)
         );
  OAI211_X1 U8882 ( .C1(n9712), .C2(n7099), .A(n7098), .B(n7097), .ZN(P1_U3280) );
  OAI21_X1 U8883 ( .B1(n4437), .B2(n5606), .A(n7100), .ZN(n10295) );
  XNOR2_X1 U8884 ( .A(n7101), .B(n8152), .ZN(n7102) );
  OAI222_X1 U8885 ( .A1(n10221), .A2(n7290), .B1(n10220), .B2(n7124), .C1(
        n10225), .C2(n7102), .ZN(n10296) );
  NAND2_X1 U8886 ( .A1(n10296), .A2(n8601), .ZN(n7106) );
  INV_X1 U8887 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8993) );
  INV_X1 U8888 ( .A(n7287), .ZN(n7103) );
  OAI22_X1 U8889 ( .A1(n8601), .A2(n8993), .B1(n7103), .B2(n10217), .ZN(n7104)
         );
  AOI21_X1 U8890 ( .B1(n10298), .B2(n10210), .A(n7104), .ZN(n7105) );
  OAI211_X1 U8891 ( .C1(n8605), .C2(n10295), .A(n7106), .B(n7105), .ZN(
        P2_U3221) );
  AOI211_X1 U8892 ( .C1(n7109), .C2(n10096), .A(n7108), .B(n7107), .ZN(n7112)
         );
  AOI22_X1 U8893 ( .A1(n9309), .A2(n9773), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n4826), .ZN(n7110) );
  OAI21_X1 U8894 ( .B1(n7112), .B2(n4826), .A(n7110), .ZN(P1_U3535) );
  AOI22_X1 U8895 ( .A1(n9309), .A2(n9847), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10098), .ZN(n7111) );
  OAI21_X1 U8896 ( .B1(n7112), .B2(n10098), .A(n7111), .ZN(P1_U3492) );
  INV_X1 U8897 ( .A(n7598), .ZN(n7142) );
  OAI222_X1 U8898 ( .A1(n9872), .A2(n7142), .B1(n5902), .B2(P1_U3086), .C1(
        n7599), .C2(n9868), .ZN(P1_U3331) );
  INV_X1 U8899 ( .A(n8154), .ZN(n7141) );
  XNOR2_X1 U8900 ( .A(n10298), .B(n4415), .ZN(n7131) );
  XNOR2_X1 U8901 ( .A(n7131), .B(n8148), .ZN(n7122) );
  XNOR2_X1 U8902 ( .A(n8134), .B(n7896), .ZN(n7281) );
  NAND2_X1 U8903 ( .A1(n7113), .A2(n8278), .ZN(n7170) );
  NAND2_X1 U8904 ( .A1(n7170), .A2(n7114), .ZN(n7169) );
  NAND2_X1 U8905 ( .A1(n7181), .A2(n7896), .ZN(n7116) );
  INV_X1 U8906 ( .A(n7181), .ZN(n10283) );
  NAND3_X1 U8907 ( .A1(n8134), .A2(n10283), .A3(n4415), .ZN(n7115) );
  OAI21_X1 U8908 ( .B1(n8134), .B2(n7116), .A(n7115), .ZN(n7117) );
  NAND2_X1 U8909 ( .A1(n7117), .A2(n7170), .ZN(n7118) );
  OAI21_X1 U8910 ( .B1(n7281), .B2(n7169), .A(n7118), .ZN(n7119) );
  AND2_X1 U8911 ( .A1(n7122), .A2(n7119), .ZN(n7120) );
  NAND2_X1 U8912 ( .A1(n7121), .A2(n7120), .ZN(n7130) );
  INV_X1 U8913 ( .A(n7122), .ZN(n7284) );
  NOR2_X1 U8914 ( .A1(n8277), .A2(n4415), .ZN(n7123) );
  AOI22_X1 U8915 ( .A1(n7123), .A2(n7181), .B1(n7124), .B2(n4415), .ZN(n7127)
         );
  NOR2_X1 U8916 ( .A1(n8277), .A2(n7896), .ZN(n7125) );
  AOI22_X1 U8917 ( .A1(n10283), .A2(n7125), .B1(n7124), .B2(n7896), .ZN(n7126)
         );
  MUX2_X1 U8918 ( .A(n7127), .B(n7126), .S(n8134), .Z(n7128) );
  OR2_X1 U8919 ( .A1(n7284), .A2(n7128), .ZN(n7129) );
  INV_X1 U8920 ( .A(n7131), .ZN(n7132) );
  NAND2_X1 U8921 ( .A1(n7132), .A2(n8148), .ZN(n7134) );
  INV_X1 U8922 ( .A(n7134), .ZN(n7133) );
  NOR2_X1 U8923 ( .A1(n7283), .A2(n7133), .ZN(n7136) );
  XNOR2_X1 U8924 ( .A(n8154), .B(n4415), .ZN(n7188) );
  XNOR2_X1 U8925 ( .A(n7188), .B(n7290), .ZN(n7135) );
  OAI211_X1 U8926 ( .C1(n7136), .C2(n7135), .A(n8016), .B(n7192), .ZN(n7140)
         );
  AND2_X1 U8927 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8301) );
  AOI21_X1 U8928 ( .B1(n7997), .B2(n8598), .A(n8301), .ZN(n7137) );
  OAI21_X1 U8929 ( .B1(n8148), .B2(n7999), .A(n7137), .ZN(n7138) );
  AOI21_X1 U8930 ( .B1(n7202), .B2(n8022), .A(n7138), .ZN(n7139) );
  OAI211_X1 U8931 ( .C1(n7141), .C2(n8025), .A(n7140), .B(n7139), .ZN(P2_U3174) );
  OAI222_X1 U8932 ( .A1(n7143), .A2(P2_U3151), .B1(n8733), .B2(n7142), .C1(
        n8865), .C2(n7278), .ZN(P2_U3271) );
  NAND2_X1 U8933 ( .A1(n7144), .A2(n7612), .ZN(n7146) );
  AOI22_X1 U8934 ( .A1(n7527), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7526), .B2(
        n9986), .ZN(n7145) );
  OR2_X1 U8935 ( .A1(n9172), .A2(n9057), .ZN(n7457) );
  NAND2_X1 U8936 ( .A1(n9172), .A2(n9057), .ZN(n7505) );
  NAND2_X1 U8937 ( .A1(n7457), .A2(n7505), .ZN(n7711) );
  NAND2_X1 U8938 ( .A1(n7147), .A2(n7712), .ZN(n7148) );
  AND2_X1 U8939 ( .A1(n9309), .A2(n9050), .ZN(n7638) );
  INV_X1 U8940 ( .A(n7638), .ZN(n7501) );
  NAND2_X1 U8941 ( .A1(n7148), .A2(n7501), .ZN(n7149) );
  OR2_X1 U8942 ( .A1(n7149), .A2(n7711), .ZN(n7215) );
  INV_X1 U8943 ( .A(n7215), .ZN(n7214) );
  AOI211_X1 U8944 ( .C1(n7711), .C2(n7149), .A(n9578), .B(n7214), .ZN(n7158)
         );
  NAND2_X1 U8945 ( .A1(n6082), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7156) );
  OR2_X1 U8946 ( .A1(n5836), .A2(n10002), .ZN(n7155) );
  NAND2_X1 U8947 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NAND2_X1 U8948 ( .A1(n7218), .A2(n7152), .ZN(n9704) );
  OR2_X1 U8949 ( .A1(n7534), .A2(n9704), .ZN(n7154) );
  OR2_X1 U8950 ( .A1(n7440), .A2(n9999), .ZN(n7153) );
  OR2_X1 U8951 ( .A1(n9050), .A2(n9350), .ZN(n7157) );
  OAI21_X1 U8952 ( .B1(n9068), .B2(n9352), .A(n7157), .ZN(n9173) );
  OR2_X1 U8953 ( .A1(n7158), .A2(n9173), .ZN(n9784) );
  INV_X1 U8954 ( .A(n9784), .ZN(n7168) );
  XNOR2_X1 U8955 ( .A(n7208), .B(n7711), .ZN(n9786) );
  NAND2_X1 U8956 ( .A1(n9786), .A2(n10053), .ZN(n7167) );
  AOI211_X1 U8957 ( .C1(n9172), .C2(n7162), .A(n9664), .B(n4496), .ZN(n9785)
         );
  NOR2_X1 U8958 ( .A1(n4588), .A2(n10062), .ZN(n7165) );
  OAI22_X1 U8959 ( .A1(n10067), .A2(n7163), .B1(n9176), .B2(n10042), .ZN(n7164) );
  AOI211_X1 U8960 ( .C1(n9785), .C2(n9665), .A(n7165), .B(n7164), .ZN(n7166)
         );
  OAI211_X1 U8961 ( .C1(n9712), .C2(n7168), .A(n7167), .B(n7166), .ZN(P1_U3279) );
  NOR2_X1 U8962 ( .A1(n7172), .A2(n7169), .ZN(n7235) );
  INV_X1 U8963 ( .A(n7235), .ZN(n7173) );
  INV_X1 U8964 ( .A(n7170), .ZN(n7171) );
  OAI21_X1 U8965 ( .B1(n7172), .B2(n7171), .A(n8277), .ZN(n7233) );
  NAND2_X1 U8966 ( .A1(n7173), .A2(n7233), .ZN(n7174) );
  XNOR2_X1 U8967 ( .A(n7181), .B(n7896), .ZN(n7234) );
  XNOR2_X1 U8968 ( .A(n7174), .B(n7234), .ZN(n7183) );
  INV_X1 U8969 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7175) );
  NOR2_X1 U8970 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7175), .ZN(n10197) );
  AOI21_X1 U8971 ( .B1(n7997), .B2(n8276), .A(n10197), .ZN(n7178) );
  NAND2_X1 U8972 ( .A1(n8022), .A2(n7176), .ZN(n7177) );
  OAI211_X1 U8973 ( .C1(n7179), .C2(n7999), .A(n7178), .B(n7177), .ZN(n7180)
         );
  AOI21_X1 U8974 ( .B1(n7181), .B2(n7969), .A(n7180), .ZN(n7182) );
  OAI21_X1 U8975 ( .B1(n7183), .B2(n7972), .A(n7182), .ZN(P2_U3157) );
  INV_X1 U8976 ( .A(n7435), .ZN(n7186) );
  OAI222_X1 U8977 ( .A1(n9872), .A2(n7186), .B1(n7184), .B2(P1_U3086), .C1(
        n8981), .C2(n9868), .ZN(P1_U3330) );
  OAI222_X1 U8978 ( .A1(n7187), .A2(P2_U3151), .B1(n8733), .B2(n7186), .C1(
        n7185), .C2(n7278), .ZN(P2_U3270) );
  INV_X1 U8979 ( .A(n7274), .ZN(n7199) );
  XNOR2_X1 U8980 ( .A(n7274), .B(n4415), .ZN(n7242) );
  XNOR2_X1 U8981 ( .A(n7242), .B(n7243), .ZN(n7190) );
  NAND2_X1 U8982 ( .A1(n7188), .A2(n8274), .ZN(n7191) );
  AND2_X1 U8983 ( .A1(n7190), .A2(n7191), .ZN(n7189) );
  INV_X1 U8984 ( .A(n7247), .ZN(n7194) );
  AOI21_X1 U8985 ( .B1(n7192), .B2(n7191), .A(n7190), .ZN(n7193) );
  OAI21_X1 U8986 ( .B1(n7194), .B2(n7193), .A(n8016), .ZN(n7198) );
  NAND2_X1 U8987 ( .A1(n8018), .A2(n8274), .ZN(n7195) );
  NAND2_X1 U8988 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8323) );
  OAI211_X1 U8989 ( .C1(n7245), .C2(n8020), .A(n7195), .B(n8323), .ZN(n7196)
         );
  AOI21_X1 U8990 ( .B1(n7261), .B2(n8022), .A(n7196), .ZN(n7197) );
  OAI211_X1 U8991 ( .C1(n7199), .C2(n8025), .A(n7198), .B(n7197), .ZN(P2_U3155) );
  XOR2_X1 U8992 ( .A(n7200), .B(n8047), .Z(n7201) );
  OAI222_X1 U8993 ( .A1(n10221), .A2(n7243), .B1(n10220), .B2(n8148), .C1(
        n7201), .C2(n10225), .ZN(n7352) );
  AOI21_X1 U8994 ( .B1(n7262), .B2(n8154), .A(n7352), .ZN(n7207) );
  AOI22_X1 U8995 ( .A1(n10235), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10211), 
        .B2(n7202), .ZN(n7206) );
  XNOR2_X1 U8996 ( .A(n7204), .B(n8047), .ZN(n7359) );
  NAND2_X1 U8997 ( .A1(n7359), .A2(n10213), .ZN(n7205) );
  OAI211_X1 U8998 ( .C1(n7207), .C2(n10235), .A(n7206), .B(n7205), .ZN(
        P2_U3220) );
  NAND2_X1 U8999 ( .A1(n7208), .A2(n5007), .ZN(n7210) );
  INV_X1 U9000 ( .A(n9057), .ZN(n9385) );
  NAND2_X1 U9001 ( .A1(n7210), .A2(n7209), .ZN(n7800) );
  NAND2_X1 U9002 ( .A1(n7211), .A2(n7612), .ZN(n7213) );
  AOI22_X1 U9003 ( .A1(n7527), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7526), .B2(
        n10006), .ZN(n7212) );
  OR2_X1 U9004 ( .A1(n9708), .A2(n9068), .ZN(n7508) );
  NAND2_X1 U9005 ( .A1(n9708), .A2(n9068), .ZN(n7729) );
  XNOR2_X1 U9006 ( .A(n7800), .B(n7714), .ZN(n9702) );
  AOI22_X1 U9007 ( .A1(n9708), .A2(n9773), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n4826), .ZN(n7229) );
  INV_X1 U9008 ( .A(n7457), .ZN(n7657) );
  NOR2_X1 U9009 ( .A1(n7214), .A2(n7657), .ZN(n7216) );
  NAND3_X1 U9010 ( .A1(n7215), .A2(n7714), .A3(n7457), .ZN(n7730) );
  OAI21_X1 U9011 ( .B1(n7216), .B2(n7714), .A(n7730), .ZN(n7226) );
  OR2_X1 U9012 ( .A1(n9057), .A2(n9350), .ZN(n7225) );
  AND2_X1 U9013 ( .A1(n7218), .A2(n7217), .ZN(n7219) );
  OR2_X1 U9014 ( .A1(n7219), .A2(n7516), .ZN(n9689) );
  NAND2_X1 U9015 ( .A1(n7589), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7221) );
  NAND2_X1 U9016 ( .A1(n6082), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n7220) );
  AND2_X1 U9017 ( .A1(n7221), .A2(n7220), .ZN(n7223) );
  OR2_X1 U9018 ( .A1(n7440), .A2(n9781), .ZN(n7222) );
  OAI211_X1 U9019 ( .C1(n9689), .C2(n7534), .A(n7223), .B(n7222), .ZN(n9383)
         );
  NAND2_X1 U9020 ( .A1(n9383), .A2(n9229), .ZN(n7224) );
  NAND2_X1 U9021 ( .A1(n7225), .A2(n7224), .ZN(n9365) );
  AOI21_X1 U9022 ( .B1(n7226), .B2(n9697), .A(n9365), .ZN(n9711) );
  INV_X1 U9023 ( .A(n9708), .ZN(n7801) );
  OAI21_X1 U9024 ( .B1(n4496), .B2(n7801), .A(n9939), .ZN(n7227) );
  OR2_X1 U9025 ( .A1(n7227), .A2(n9691), .ZN(n9705) );
  NAND2_X1 U9026 ( .A1(n9711), .A2(n9705), .ZN(n7230) );
  NAND2_X1 U9027 ( .A1(n7230), .A2(n10106), .ZN(n7228) );
  OAI211_X1 U9028 ( .C1(n9702), .C2(n9775), .A(n7229), .B(n7228), .ZN(P1_U3537) );
  AOI22_X1 U9029 ( .A1(n9708), .A2(n9847), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n10098), .ZN(n7232) );
  NAND2_X1 U9030 ( .A1(n7230), .A2(n10100), .ZN(n7231) );
  OAI211_X1 U9031 ( .C1(n9702), .C2(n9842), .A(n7232), .B(n7231), .ZN(P1_U3498) );
  OAI21_X1 U9032 ( .B1(n7235), .B2(n7234), .A(n7233), .ZN(n7282) );
  XOR2_X1 U9033 ( .A(n7281), .B(n7282), .Z(n7241) );
  AND2_X1 U9034 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7375) );
  AOI21_X1 U9035 ( .B1(n8018), .B2(n8277), .A(n7375), .ZN(n7238) );
  NAND2_X1 U9036 ( .A1(n8022), .A2(n7236), .ZN(n7237) );
  OAI211_X1 U9037 ( .C1(n8148), .C2(n8020), .A(n7238), .B(n7237), .ZN(n7239)
         );
  AOI21_X1 U9038 ( .B1(n10292), .B2(n7969), .A(n7239), .ZN(n7240) );
  OAI21_X1 U9039 ( .B1(n7241), .B2(n7972), .A(n7240), .ZN(P2_U3176) );
  INV_X1 U9040 ( .A(n8718), .ZN(n7254) );
  INV_X1 U9041 ( .A(n7242), .ZN(n7244) );
  NAND2_X1 U9042 ( .A1(n7244), .A2(n7243), .ZN(n7246) );
  AND2_X1 U9043 ( .A1(n7247), .A2(n7246), .ZN(n7249) );
  XNOR2_X1 U9044 ( .A(n8718), .B(n4415), .ZN(n7296) );
  XNOR2_X1 U9045 ( .A(n7296), .B(n7245), .ZN(n7248) );
  OAI211_X1 U9046 ( .C1(n7249), .C2(n7248), .A(n8016), .B(n7298), .ZN(n7253)
         );
  NAND2_X1 U9047 ( .A1(n8018), .A2(n8598), .ZN(n7250) );
  NAND2_X1 U9048 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U9049 ( .C1(n7875), .C2(n8020), .A(n7250), .B(n8347), .ZN(n7251)
         );
  AOI21_X1 U9050 ( .B1(n8602), .B2(n8022), .A(n7251), .ZN(n7252) );
  OAI211_X1 U9051 ( .C1(n7254), .C2(n8025), .A(n7253), .B(n7252), .ZN(P2_U3181) );
  INV_X1 U9052 ( .A(n7424), .ZN(n7279) );
  OAI222_X1 U9053 ( .A1(n9872), .A2(n7279), .B1(n7255), .B2(P1_U3086), .C1(
        n7425), .C2(n9868), .ZN(P1_U3329) );
  NAND2_X1 U9054 ( .A1(n7257), .A2(n8165), .ZN(n7258) );
  NAND3_X1 U9055 ( .A1(n7256), .A2(n10207), .A3(n7258), .ZN(n7260) );
  AOI22_X1 U9056 ( .A1(n10204), .A2(n8274), .B1(n8587), .B2(n10202), .ZN(n7259) );
  AOI22_X1 U9057 ( .A1(n7274), .A2(n7262), .B1(n10211), .B2(n7261), .ZN(n7263)
         );
  AOI21_X1 U9058 ( .B1(n7272), .B2(n7263), .A(n10235), .ZN(n7268) );
  XNOR2_X1 U9059 ( .A(n7265), .B(n8165), .ZN(n7277) );
  INV_X1 U9060 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7266) );
  OAI22_X1 U9061 ( .A1(n7277), .A2(n8605), .B1(n7266), .B2(n8601), .ZN(n7267)
         );
  OR2_X1 U9062 ( .A1(n7268), .A2(n7267), .ZN(P2_U3219) );
  INV_X1 U9063 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7269) );
  MUX2_X1 U9064 ( .A(n7269), .B(n7272), .S(n10325), .Z(n7271) );
  NAND2_X1 U9065 ( .A1(n7274), .A2(n8646), .ZN(n7270) );
  OAI211_X1 U9066 ( .C1(n7277), .C2(n8649), .A(n7271), .B(n7270), .ZN(P2_U3473) );
  INV_X1 U9067 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7273) );
  MUX2_X1 U9068 ( .A(n7273), .B(n7272), .S(n10300), .Z(n7276) );
  NAND2_X1 U9069 ( .A1(n7274), .A2(n5662), .ZN(n7275) );
  OAI211_X1 U9070 ( .C1(n7277), .C2(n8721), .A(n7276), .B(n7275), .ZN(P2_U3432) );
  OAI222_X1 U9071 ( .A1(n7280), .A2(P2_U3151), .B1(n8733), .B2(n7279), .C1(
        n8871), .C2(n7278), .ZN(P2_U3269) );
  MUX2_X1 U9072 ( .A(n7282), .B(n8276), .S(n7281), .Z(n7285) );
  AOI21_X1 U9073 ( .B1(n7285), .B2(n7284), .A(n7283), .ZN(n7293) );
  NOR2_X1 U9074 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7286), .ZN(n7343) );
  AOI21_X1 U9075 ( .B1(n8018), .B2(n8276), .A(n7343), .ZN(n7289) );
  NAND2_X1 U9076 ( .A1(n8022), .A2(n7287), .ZN(n7288) );
  OAI211_X1 U9077 ( .C1(n7290), .C2(n8020), .A(n7289), .B(n7288), .ZN(n7291)
         );
  AOI21_X1 U9078 ( .B1(n10298), .B2(n7969), .A(n7291), .ZN(n7292) );
  OAI21_X1 U9079 ( .B1(n7293), .B2(n7972), .A(n7292), .ZN(P2_U3164) );
  INV_X1 U9080 ( .A(n7421), .ZN(n7777) );
  AOI22_X1 U9081 ( .A1(n7294), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9020), .ZN(n7295) );
  OAI21_X1 U9082 ( .B1(n7777), .B2(n8733), .A(n7295), .ZN(P2_U3268) );
  NAND2_X1 U9083 ( .A1(n7296), .A2(n8587), .ZN(n7297) );
  NAND2_X1 U9084 ( .A1(n7298), .A2(n7297), .ZN(n7874) );
  XNOR2_X1 U9085 ( .A(n8712), .B(n4415), .ZN(n7876) );
  XNOR2_X1 U9086 ( .A(n7876), .B(n7875), .ZN(n7873) );
  XNOR2_X1 U9087 ( .A(n7874), .B(n7873), .ZN(n7304) );
  NAND2_X1 U9088 ( .A1(n8018), .A2(n8587), .ZN(n7299) );
  NAND2_X1 U9089 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8369) );
  OAI211_X1 U9090 ( .C1(n8565), .C2(n8020), .A(n7299), .B(n8369), .ZN(n7302)
         );
  NOR2_X1 U9091 ( .A1(n7300), .A2(n8025), .ZN(n7301) );
  AOI211_X1 U9092 ( .C1(n8591), .C2(n8022), .A(n7302), .B(n7301), .ZN(n7303)
         );
  OAI21_X1 U9093 ( .B1(n7304), .B2(n7972), .A(n7303), .ZN(P2_U3166) );
  NOR2_X1 U9094 ( .A1(n9021), .A2(n7305), .ZN(n7307) );
  AOI22_X1 U9095 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7333), .B1(n10184), .B2(
        n6950), .ZN(n10190) );
  NOR2_X1 U9096 ( .A1(n7334), .A2(n7308), .ZN(n7309) );
  OR2_X1 U9097 ( .A1(n7344), .A2(n8993), .ZN(n8287) );
  NAND2_X1 U9098 ( .A1(n7344), .A2(n8993), .ZN(n7310) );
  NAND2_X1 U9099 ( .A1(n8287), .A2(n7310), .ZN(n7312) );
  INV_X1 U9100 ( .A(n8288), .ZN(n7311) );
  AOI21_X1 U9101 ( .B1(n7313), .B2(n7312), .A(n7311), .ZN(n7351) );
  MUX2_X1 U9102 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8426), .Z(n7321) );
  NOR2_X1 U9103 ( .A1(n7321), .A2(n7368), .ZN(n7323) );
  MUX2_X1 U9104 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8426), .Z(n7318) );
  NOR2_X1 U9105 ( .A1(n7318), .A2(n10184), .ZN(n7320) );
  INV_X1 U9106 ( .A(n7314), .ZN(n7317) );
  AOI21_X1 U9107 ( .B1(n7318), .B2(n10184), .A(n7320), .ZN(n7319) );
  INV_X1 U9108 ( .A(n7319), .ZN(n10187) );
  AOI21_X1 U9109 ( .B1(n7321), .B2(n7368), .A(n7323), .ZN(n7322) );
  INV_X1 U9110 ( .A(n7322), .ZN(n7371) );
  MUX2_X1 U9111 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8426), .Z(n7325) );
  AND2_X1 U9112 ( .A1(n7325), .A2(n7324), .ZN(n8291) );
  INV_X1 U9113 ( .A(n8291), .ZN(n7327) );
  INV_X1 U9114 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7337) );
  MUX2_X1 U9115 ( .A(n8993), .B(n7337), .S(n8426), .Z(n7326) );
  NAND2_X1 U9116 ( .A1(n7326), .A2(n7344), .ZN(n8292) );
  NAND2_X1 U9117 ( .A1(n7327), .A2(n8292), .ZN(n7328) );
  XNOR2_X1 U9118 ( .A(n8293), .B(n7328), .ZN(n7329) );
  NAND2_X1 U9119 ( .A1(n7329), .A2(n10167), .ZN(n7350) );
  NOR2_X1 U9120 ( .A1(n9021), .A2(n7330), .ZN(n7332) );
  INV_X1 U9121 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10319) );
  AOI22_X1 U9122 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7333), .B1(n10184), .B2(
        n10319), .ZN(n10181) );
  NOR2_X1 U9123 ( .A1(n7334), .A2(n7335), .ZN(n7336) );
  INV_X1 U9124 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10321) );
  NOR2_X1 U9125 ( .A1(n10321), .A2(n7365), .ZN(n7364) );
  INV_X1 U9126 ( .A(n7340), .ZN(n7342) );
  OR2_X1 U9127 ( .A1(n7344), .A2(n7337), .ZN(n8297) );
  NAND2_X1 U9128 ( .A1(n7344), .A2(n7337), .ZN(n7338) );
  NAND2_X1 U9129 ( .A1(n8297), .A2(n7338), .ZN(n7339) );
  INV_X1 U9130 ( .A(n7339), .ZN(n7341) );
  OAI21_X1 U9131 ( .B1(n7342), .B2(n7341), .A(n8298), .ZN(n7348) );
  INV_X1 U9132 ( .A(n10185), .ZN(n8393) );
  AOI21_X1 U9133 ( .B1(n8393), .B2(n7344), .A(n7343), .ZN(n7345) );
  OAI21_X1 U9134 ( .B1(n7346), .B2(n10183), .A(n7345), .ZN(n7347) );
  AOI21_X1 U9135 ( .B1(n7348), .B2(n10127), .A(n7347), .ZN(n7349) );
  OAI211_X1 U9136 ( .C1(n7351), .C2(n10191), .A(n7350), .B(n7349), .ZN(
        P2_U3194) );
  INV_X1 U9137 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7353) );
  INV_X1 U9138 ( .A(n7352), .ZN(n7357) );
  MUX2_X1 U9139 ( .A(n7353), .B(n7357), .S(n10300), .Z(n7356) );
  INV_X1 U9140 ( .A(n8721), .ZN(n7354) );
  AOI22_X1 U9141 ( .A1(n7359), .A2(n7354), .B1(n5662), .B2(n8154), .ZN(n7355)
         );
  NAND2_X1 U9142 ( .A1(n7356), .A2(n7355), .ZN(P2_U3429) );
  INV_X1 U9143 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8300) );
  MUX2_X1 U9144 ( .A(n8300), .B(n7357), .S(n10325), .Z(n7361) );
  INV_X1 U9145 ( .A(n8649), .ZN(n7358) );
  AOI22_X1 U9146 ( .A1(n7359), .A2(n7358), .B1(n8646), .B2(n8154), .ZN(n7360)
         );
  NAND2_X1 U9147 ( .A1(n7361), .A2(n7360), .ZN(P2_U3472) );
  AOI21_X1 U9148 ( .B1(n7055), .B2(n7363), .A(n7362), .ZN(n7378) );
  AOI21_X1 U9149 ( .B1(n10321), .B2(n7365), .A(n7364), .ZN(n7366) );
  NOR2_X1 U9150 ( .A1(n7366), .A2(n10199), .ZN(n7376) );
  OAI22_X1 U9151 ( .A1(n10185), .A2(n7368), .B1(n10183), .B2(n7367), .ZN(n7374) );
  AOI21_X1 U9152 ( .B1(n7371), .B2(n7370), .A(n7369), .ZN(n7372) );
  NOR2_X1 U9153 ( .A1(n7372), .A2(n10193), .ZN(n7373) );
  NOR4_X1 U9154 ( .A1(n7376), .A2(n7375), .A3(n7374), .A4(n7373), .ZN(n7377)
         );
  OAI21_X1 U9155 ( .B1(n7378), .B2(n10191), .A(n7377), .ZN(P2_U3193) );
  INV_X1 U9156 ( .A(n7412), .ZN(n7770) );
  AOI21_X1 U9157 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n9020), .A(n7379), .ZN(
        n7380) );
  OAI21_X1 U9158 ( .B1(n7770), .B2(n8733), .A(n7380), .ZN(P2_U3267) );
  INV_X1 U9159 ( .A(n7383), .ZN(n7385) );
  INV_X1 U9160 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7386) );
  INV_X1 U9161 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9869) );
  MUX2_X1 U9162 ( .A(n7386), .B(n9869), .S(n5534), .Z(n7388) );
  INV_X1 U9163 ( .A(SI_29_), .ZN(n7387) );
  INV_X1 U9164 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7392) );
  INV_X1 U9165 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9867) );
  MUX2_X1 U9166 ( .A(n7392), .B(n9867), .S(n5534), .Z(n7394) );
  INV_X1 U9167 ( .A(SI_30_), .ZN(n7393) );
  NAND2_X1 U9168 ( .A1(n7394), .A2(n7393), .ZN(n7397) );
  INV_X1 U9169 ( .A(n7394), .ZN(n7395) );
  NAND2_X1 U9170 ( .A1(n7395), .A2(SI_30_), .ZN(n7396) );
  NAND2_X1 U9171 ( .A1(n7397), .A2(n7396), .ZN(n7610) );
  INV_X1 U9172 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9859) );
  MUX2_X1 U9173 ( .A(n8952), .B(n9859), .S(n5534), .Z(n7398) );
  XNOR2_X1 U9174 ( .A(n7398), .B(SI_31_), .ZN(n7399) );
  NAND2_X1 U9175 ( .A1(n8723), .A2(n7612), .ZN(n7402) );
  OR2_X1 U9176 ( .A1(n7613), .A2(n9859), .ZN(n7401) );
  NAND2_X1 U9177 ( .A1(n9793), .A2(n9484), .ZN(n7754) );
  AOI211_X1 U9178 ( .C1(n7721), .C2(n4418), .A(n7766), .B(n7403), .ZN(n7762)
         );
  INV_X1 U9179 ( .A(n9484), .ZN(n7404) );
  NAND2_X1 U9180 ( .A1(n9480), .A2(n7404), .ZN(n7757) );
  NAND2_X1 U9181 ( .A1(n7589), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7411) );
  INV_X1 U9182 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7832) );
  OR2_X1 U9183 ( .A1(n7592), .A2(n7832), .ZN(n7410) );
  AND2_X1 U9184 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n7406) );
  NAND2_X1 U9185 ( .A1(n7407), .A2(n7406), .ZN(n7837) );
  OR2_X1 U9186 ( .A1(n7534), .A2(n7837), .ZN(n7409) );
  INV_X1 U9187 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7833) );
  OR2_X1 U9188 ( .A1(n7440), .A2(n7833), .ZN(n7408) );
  INV_X1 U9189 ( .A(n7687), .ZN(n7681) );
  NAND2_X1 U9190 ( .A1(n7412), .A2(n7612), .ZN(n7414) );
  INV_X1 U9191 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8870) );
  OR2_X1 U9192 ( .A1(n7613), .A2(n8870), .ZN(n7413) );
  NAND2_X1 U9193 ( .A1(n7589), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n7420) );
  INV_X1 U9194 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9795) );
  OR2_X1 U9195 ( .A1(n7592), .A2(n9795), .ZN(n7419) );
  INV_X1 U9196 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U9197 ( .B1(n7430), .B2(n9165), .A(n7415), .ZN(n7416) );
  NAND2_X1 U9198 ( .A1(n7416), .A2(n7837), .ZN(n9501) );
  OR2_X1 U9199 ( .A1(n7534), .A2(n9501), .ZN(n7418) );
  INV_X1 U9200 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9720) );
  OR2_X1 U9201 ( .A1(n7440), .A2(n9720), .ZN(n7417) );
  AND4_X2 U9202 ( .A1(n7420), .A2(n7419), .A3(n7418), .A4(n7417), .ZN(n9208)
         );
  NAND2_X1 U9203 ( .A1(n9719), .A2(n9208), .ZN(n7828) );
  NAND2_X1 U9204 ( .A1(n7421), .A2(n7612), .ZN(n7423) );
  OR2_X1 U9205 ( .A1(n7613), .A2(n7776), .ZN(n7422) );
  NAND2_X1 U9206 ( .A1(n9724), .A2(n9353), .ZN(n7827) );
  NAND2_X2 U9207 ( .A1(n7675), .A2(n7827), .ZN(n9510) );
  NAND2_X1 U9208 ( .A1(n7424), .A2(n7612), .ZN(n7427) );
  OR2_X1 U9209 ( .A1(n7613), .A2(n7425), .ZN(n7426) );
  NAND2_X1 U9210 ( .A1(n7589), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n7434) );
  INV_X1 U9211 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9730) );
  OR2_X1 U9212 ( .A1(n7440), .A2(n9730), .ZN(n7433) );
  INV_X1 U9213 ( .A(n7428), .ZN(n7438) );
  INV_X1 U9214 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U9215 ( .A1(n7438), .A2(n9356), .ZN(n7429) );
  NAND2_X1 U9216 ( .A1(n7430), .A2(n7429), .ZN(n9349) );
  OR2_X1 U9217 ( .A1(n7534), .A2(n9349), .ZN(n7432) );
  INV_X1 U9218 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9803) );
  OR2_X1 U9219 ( .A1(n7592), .A2(n9803), .ZN(n7431) );
  INV_X1 U9220 ( .A(n9248), .ZN(n9375) );
  NAND2_X1 U9221 ( .A1(n9729), .A2(n9248), .ZN(n7825) );
  NAND2_X1 U9222 ( .A1(n7435), .A2(n7612), .ZN(n7437) );
  OR2_X1 U9223 ( .A1(n7613), .A2(n8981), .ZN(n7436) );
  NAND2_X1 U9224 ( .A1(n6082), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n7444) );
  INV_X1 U9225 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9546) );
  OR2_X1 U9226 ( .A1(n5836), .A2(n9546), .ZN(n7443) );
  OAI21_X1 U9227 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n7439), .A(n7438), .ZN(
        n9545) );
  OR2_X1 U9228 ( .A1(n7534), .A2(n9545), .ZN(n7442) );
  INV_X1 U9229 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8854) );
  OR2_X1 U9230 ( .A1(n7440), .A2(n8854), .ZN(n7441) );
  NAND2_X1 U9231 ( .A1(n9808), .A2(n9351), .ZN(n7689) );
  NAND2_X1 U9232 ( .A1(n7825), .A2(n7689), .ZN(n7604) );
  NAND2_X1 U9233 ( .A1(n7688), .A2(n7604), .ZN(n7448) );
  NOR4_X1 U9234 ( .A1(n7829), .A2(n9510), .A3(n7625), .A4(n7448), .ZN(n7446)
         );
  NAND2_X1 U9235 ( .A1(n7828), .A2(n7827), .ZN(n7680) );
  INV_X1 U9236 ( .A(n7680), .ZN(n7740) );
  INV_X1 U9237 ( .A(n7450), .ZN(n7677) );
  NOR3_X1 U9238 ( .A1(n7740), .A2(n7677), .A3(n7625), .ZN(n7445) );
  AOI211_X1 U9239 ( .C1(n7681), .C2(n4677), .A(n7446), .B(n7445), .ZN(n7456)
         );
  INV_X1 U9240 ( .A(n7814), .ZN(n7841) );
  INV_X1 U9241 ( .A(n9212), .ZN(n9373) );
  NAND2_X1 U9242 ( .A1(n7841), .A2(n9373), .ZN(n7686) );
  INV_X1 U9243 ( .A(n7686), .ZN(n7678) );
  INV_X1 U9244 ( .A(n7604), .ZN(n7447) );
  AOI21_X1 U9245 ( .B1(n7447), .B2(n9522), .A(n4677), .ZN(n7449) );
  NAND4_X1 U9246 ( .A1(n9493), .A2(n9508), .A3(n7449), .A4(n7448), .ZN(n7453)
         );
  NAND2_X1 U9247 ( .A1(n7680), .A2(n7450), .ZN(n7451) );
  OAI211_X1 U9248 ( .C1(n7829), .C2(n9510), .A(n7625), .B(n7451), .ZN(n7452)
         );
  AOI21_X1 U9249 ( .B1(n7453), .B2(n7452), .A(n7681), .ZN(n7454) );
  NAND2_X1 U9250 ( .A1(n7457), .A2(n7625), .ZN(n7506) );
  INV_X1 U9251 ( .A(n7458), .ZN(n7459) );
  INV_X1 U9252 ( .A(n7466), .ZN(n7460) );
  NOR2_X1 U9253 ( .A1(n7460), .A2(n7465), .ZN(n7462) );
  NAND2_X1 U9254 ( .A1(n7461), .A2(n7648), .ZN(n7468) );
  INV_X1 U9255 ( .A(n7463), .ZN(n7464) );
  NOR3_X1 U9256 ( .A1(n7466), .A2(n7465), .A3(n7464), .ZN(n7469) );
  OAI21_X1 U9257 ( .B1(n7469), .B2(n7468), .A(n7467), .ZN(n7472) );
  MUX2_X1 U9258 ( .A(n7475), .B(n7474), .S(n7625), .Z(n7476) );
  INV_X1 U9259 ( .A(n7490), .ZN(n7480) );
  INV_X1 U9260 ( .A(n7477), .ZN(n7479) );
  OAI211_X1 U9261 ( .C1(n7480), .C2(n7479), .A(n7489), .B(n7478), .ZN(n7488)
         );
  INV_X1 U9262 ( .A(n7654), .ZN(n7492) );
  NOR2_X1 U9263 ( .A1(n7492), .A2(n7651), .ZN(n7487) );
  INV_X1 U9264 ( .A(n7481), .ZN(n7484) );
  INV_X1 U9265 ( .A(n7482), .ZN(n7483) );
  AOI21_X1 U9266 ( .B1(n7485), .B2(n7484), .A(n7483), .ZN(n7486) );
  AOI21_X1 U9267 ( .B1(n7488), .B2(n7487), .A(n7486), .ZN(n7495) );
  AOI21_X1 U9268 ( .B1(n7490), .B2(n7489), .A(n7651), .ZN(n7491) );
  NOR2_X1 U9269 ( .A1(n7491), .A2(n7655), .ZN(n7493) );
  OAI21_X1 U9270 ( .B1(n7493), .B2(n7492), .A(n7637), .ZN(n7494) );
  MUX2_X1 U9271 ( .A(n7495), .B(n7494), .S(n7625), .Z(n7502) );
  OR2_X1 U9272 ( .A1(n9309), .A2(n9050), .ZN(n7500) );
  AOI211_X1 U9273 ( .C1(n7502), .C2(n7500), .A(n7638), .B(n7711), .ZN(n7504)
         );
  NAND2_X1 U9274 ( .A1(n7496), .A2(n7612), .ZN(n7499) );
  AOI22_X1 U9275 ( .A1(n7527), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7526), .B2(
        n7497), .ZN(n7498) );
  INV_X1 U9276 ( .A(n9383), .ZN(n7802) );
  OR2_X1 U9277 ( .A1(n9846), .A2(n7802), .ZN(n7697) );
  NAND2_X1 U9278 ( .A1(n7697), .A2(n7508), .ZN(n7661) );
  INV_X1 U9279 ( .A(n7500), .ZN(n7658) );
  AOI211_X1 U9280 ( .C1(n7502), .C2(n7501), .A(n7658), .B(n7711), .ZN(n7503)
         );
  NAND2_X1 U9281 ( .A1(n7729), .A2(n7505), .ZN(n7663) );
  NAND2_X1 U9282 ( .A1(n7663), .A2(n7506), .ZN(n7512) );
  INV_X1 U9283 ( .A(n7697), .ZN(n7507) );
  NOR3_X1 U9284 ( .A1(n7507), .A2(n4677), .A3(n7729), .ZN(n7511) );
  OAI21_X1 U9285 ( .B1(n7665), .B2(n7508), .A(n7697), .ZN(n7509) );
  MUX2_X1 U9286 ( .A(n7509), .B(n7665), .S(n7625), .Z(n7510) );
  NAND2_X1 U9287 ( .A1(n7513), .A2(n7612), .ZN(n7515) );
  AOI22_X1 U9288 ( .A1(n7527), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7526), .B2(
        n7787), .ZN(n7514) );
  OR2_X1 U9289 ( .A1(n7516), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n7517) );
  AND2_X1 U9290 ( .A1(n7532), .A2(n7517), .ZN(n9682) );
  NAND2_X1 U9291 ( .A1(n9682), .A2(n7594), .ZN(n7520) );
  AOI22_X1 U9292 ( .A1(n7589), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n7616), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n7519) );
  INV_X1 U9293 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n8829) );
  OR2_X1 U9294 ( .A1(n7592), .A2(n8829), .ZN(n7518) );
  OR2_X1 U9295 ( .A1(n9840), .A2(n9340), .ZN(n9653) );
  NAND2_X1 U9296 ( .A1(n9840), .A2(n9340), .ZN(n7540) );
  NAND2_X1 U9297 ( .A1(n9653), .A2(n7540), .ZN(n9673) );
  INV_X1 U9298 ( .A(n9653), .ZN(n7666) );
  OR2_X1 U9299 ( .A1(n7522), .A2(n7521), .ZN(n7524) );
  AOI22_X1 U9300 ( .A1(n7527), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n7526), .B2(
        n10032), .ZN(n7523) );
  NOR2_X1 U9301 ( .A1(n9766), .A2(n9272), .ZN(n7693) );
  NAND2_X1 U9302 ( .A1(n7525), .A2(n7612), .ZN(n7529) );
  AOI22_X1 U9303 ( .A1(n7527), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4418), .B2(
        n7526), .ZN(n7528) );
  INV_X1 U9304 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7531) );
  INV_X1 U9305 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7530) );
  OAI21_X1 U9306 ( .B1(n7532), .B2(n7531), .A(n7530), .ZN(n7533) );
  NAND2_X1 U9307 ( .A1(n7533), .A2(n7546), .ZN(n9642) );
  OR2_X1 U9308 ( .A1(n9642), .A2(n7534), .ZN(n7537) );
  AOI22_X1 U9309 ( .A1(n6082), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n7589), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n7536) );
  NAND2_X1 U9310 ( .A1(n7616), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n7535) );
  AND2_X1 U9311 ( .A1(n9648), .A2(n9341), .ZN(n7733) );
  AND2_X1 U9312 ( .A1(n9766), .A2(n9272), .ZN(n7539) );
  NOR3_X1 U9313 ( .A1(n7538), .A2(n7733), .A3(n7539), .ZN(n7556) );
  NAND2_X1 U9314 ( .A1(n7732), .A2(n7540), .ZN(n7669) );
  NOR2_X1 U9315 ( .A1(n9648), .A2(n9341), .ZN(n7557) );
  NOR2_X1 U9316 ( .A1(n7557), .A2(n7693), .ZN(n7668) );
  OAI21_X1 U9317 ( .B1(n7541), .B2(n7669), .A(n7668), .ZN(n7554) );
  INV_X1 U9318 ( .A(n7733), .ZN(n7695) );
  NAND2_X1 U9319 ( .A1(n7542), .A2(n7612), .ZN(n7545) );
  OR2_X1 U9320 ( .A1(n7613), .A2(n7543), .ZN(n7544) );
  NAND2_X1 U9321 ( .A1(n7546), .A2(n9299), .ZN(n7547) );
  AND2_X1 U9322 ( .A1(n7561), .A2(n7547), .ZN(n9629) );
  NAND2_X1 U9323 ( .A1(n9629), .A2(n7594), .ZN(n7553) );
  INV_X1 U9324 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n7550) );
  NAND2_X1 U9325 ( .A1(n6082), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n7549) );
  NAND2_X1 U9326 ( .A1(n7616), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n7548) );
  OAI211_X1 U9327 ( .C1(n5836), .C2(n7550), .A(n7549), .B(n7548), .ZN(n7551)
         );
  INV_X1 U9328 ( .A(n7551), .ZN(n7552) );
  NAND2_X1 U9329 ( .A1(n9627), .A2(n9227), .ZN(n7817) );
  NAND3_X1 U9330 ( .A1(n7554), .A2(n7695), .A3(n7817), .ZN(n7555) );
  MUX2_X1 U9331 ( .A(n7556), .B(n7555), .S(n7625), .Z(n7569) );
  OR2_X1 U9332 ( .A1(n9627), .A2(n9227), .ZN(n9606) );
  INV_X1 U9333 ( .A(n7557), .ZN(n7696) );
  AOI21_X1 U9334 ( .B1(n9606), .B2(n7696), .A(n7625), .ZN(n7568) );
  NAND2_X1 U9335 ( .A1(n7558), .A2(n7612), .ZN(n7560) );
  OR2_X1 U9336 ( .A1(n7613), .A2(n8932), .ZN(n7559) );
  AND2_X1 U9337 ( .A1(n7561), .A2(n9230), .ZN(n7562) );
  NOR2_X1 U9338 ( .A1(n7573), .A2(n7562), .ZN(n9611) );
  INV_X1 U9339 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n7565) );
  NAND2_X1 U9340 ( .A1(n7589), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n7564) );
  NAND2_X1 U9341 ( .A1(n7616), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n7563) );
  OAI211_X1 U9342 ( .C1(n7592), .C2(n7565), .A(n7564), .B(n7563), .ZN(n7566)
         );
  AOI21_X1 U9343 ( .B1(n9611), .B2(n7594), .A(n7566), .ZN(n9316) );
  NAND2_X1 U9344 ( .A1(n9752), .A2(n9316), .ZN(n7691) );
  AND2_X1 U9345 ( .A1(n7691), .A2(n7817), .ZN(n7631) );
  OR2_X1 U9346 ( .A1(n9752), .A2(n9316), .ZN(n7692) );
  AND2_X1 U9347 ( .A1(n7692), .A2(n9606), .ZN(n7734) );
  MUX2_X1 U9348 ( .A(n7631), .B(n7734), .S(n7625), .Z(n7567) );
  OAI21_X1 U9349 ( .B1(n7569), .B2(n7568), .A(n7567), .ZN(n7582) );
  MUX2_X1 U9350 ( .A(n7692), .B(n7691), .S(n7625), .Z(n7581) );
  NAND2_X1 U9351 ( .A1(n7570), .A2(n7612), .ZN(n7572) );
  OR2_X1 U9352 ( .A1(n7613), .A2(n7781), .ZN(n7571) );
  NOR2_X1 U9353 ( .A1(n7573), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n7574) );
  OR2_X1 U9354 ( .A1(n7586), .A2(n7574), .ZN(n9596) );
  INV_X1 U9355 ( .A(n9596), .ZN(n7575) );
  NAND2_X1 U9356 ( .A1(n7575), .A2(n7594), .ZN(n7580) );
  INV_X1 U9357 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U9358 ( .A1(n6082), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9359 ( .A1(n7616), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n7576) );
  OAI211_X1 U9360 ( .C1(n5836), .C2(n9595), .A(n7577), .B(n7576), .ZN(n7578)
         );
  INV_X1 U9361 ( .A(n7578), .ZN(n7579) );
  OR2_X1 U9362 ( .A1(n9600), .A2(n9180), .ZN(n7819) );
  NAND2_X1 U9363 ( .A1(n9600), .A2(n9180), .ZN(n7820) );
  NAND2_X1 U9364 ( .A1(n7819), .A2(n7820), .ZN(n9592) );
  AOI21_X1 U9365 ( .B1(n7582), .B2(n7581), .A(n9592), .ZN(n7595) );
  NAND2_X1 U9366 ( .A1(n7583), .A2(n7612), .ZN(n7585) );
  OR2_X1 U9367 ( .A1(n7613), .A2(n8814), .ZN(n7584) );
  NOR2_X1 U9368 ( .A1(n7586), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7587) );
  OR2_X1 U9369 ( .A1(n7588), .A2(n7587), .ZN(n9184) );
  INV_X1 U9370 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U9371 ( .A1(n7589), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n7591) );
  NAND2_X1 U9372 ( .A1(n7616), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n7590) );
  OAI211_X1 U9373 ( .C1(n7592), .C2(n9817), .A(n7591), .B(n7590), .ZN(n7593)
         );
  AOI21_X1 U9374 ( .B1(n9582), .B2(n7594), .A(n7593), .ZN(n9315) );
  OR2_X1 U9375 ( .A1(n9742), .A2(n9315), .ZN(n7690) );
  NAND2_X1 U9376 ( .A1(n7690), .A2(n7819), .ZN(n7626) );
  NAND2_X1 U9377 ( .A1(n9742), .A2(n9315), .ZN(n7822) );
  OAI21_X1 U9378 ( .B1(n7595), .B2(n7626), .A(n7822), .ZN(n7597) );
  NAND2_X1 U9379 ( .A1(n7822), .A2(n7820), .ZN(n7630) );
  OAI21_X1 U9380 ( .B1(n7595), .B2(n7630), .A(n7690), .ZN(n7596) );
  MUX2_X1 U9381 ( .A(n7597), .B(n7596), .S(n7625), .Z(n7603) );
  NAND2_X1 U9382 ( .A1(n7598), .A2(n7612), .ZN(n7601) );
  OR2_X1 U9383 ( .A1(n7613), .A2(n7599), .ZN(n7600) );
  OR2_X1 U9384 ( .A1(n9813), .A2(n9247), .ZN(n7823) );
  NAND2_X1 U9385 ( .A1(n9813), .A2(n9247), .ZN(n7633) );
  NAND2_X1 U9386 ( .A1(n7823), .A2(n7633), .ZN(n9559) );
  MUX2_X1 U9387 ( .A(n7823), .B(n7633), .S(n7625), .Z(n7602) );
  NOR4_X1 U9388 ( .A1(n7829), .A2(n9510), .A3(n4677), .A4(n7604), .ZN(n7608)
         );
  NAND2_X1 U9389 ( .A1(n9522), .A2(n4677), .ZN(n7605) );
  NOR4_X1 U9390 ( .A1(n7829), .A2(n9510), .A3(n7606), .A4(n7605), .ZN(n7607)
         );
  AOI22_X1 U9391 ( .A1(n7687), .A2(n7608), .B1(n7686), .B2(n7607), .ZN(n7609)
         );
  NAND2_X1 U9392 ( .A1(n8728), .A2(n7612), .ZN(n7615) );
  OR2_X1 U9393 ( .A1(n7613), .A2(n9867), .ZN(n7614) );
  INV_X1 U9394 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U9395 ( .A1(n7616), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7618) );
  NAND2_X1 U9396 ( .A1(n6082), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7617) );
  OAI211_X1 U9397 ( .C1(n5836), .C2(n7619), .A(n7618), .B(n7617), .ZN(n9372)
         );
  NAND2_X1 U9398 ( .A1(n9372), .A2(n9484), .ZN(n7747) );
  NAND3_X1 U9399 ( .A1(n7620), .A2(n7754), .A3(n7747), .ZN(n7624) );
  NAND3_X1 U9400 ( .A1(n7622), .A2(n9480), .A3(n9372), .ZN(n7623) );
  NAND3_X1 U9401 ( .A1(n7624), .A2(n7623), .A3(n7757), .ZN(n7685) );
  OAI21_X1 U9402 ( .B1(n7625), .B2(n7757), .A(n7685), .ZN(n7761) );
  NAND2_X1 U9403 ( .A1(n7626), .A2(n7822), .ZN(n7627) );
  NAND2_X1 U9404 ( .A1(n7823), .A2(n7627), .ZN(n7628) );
  NAND2_X1 U9405 ( .A1(n7628), .A2(n7633), .ZN(n7629) );
  AND2_X1 U9406 ( .A1(n9522), .A2(n7629), .ZN(n7728) );
  INV_X1 U9407 ( .A(n7630), .ZN(n7634) );
  INV_X1 U9408 ( .A(n7631), .ZN(n7632) );
  NAND2_X1 U9409 ( .A1(n7632), .A2(n7692), .ZN(n7818) );
  NAND3_X1 U9410 ( .A1(n7634), .A2(n7633), .A3(n7818), .ZN(n7636) );
  INV_X1 U9411 ( .A(n7689), .ZN(n7635) );
  AOI21_X1 U9412 ( .B1(n7728), .B2(n7636), .A(n7635), .ZN(n7727) );
  INV_X1 U9413 ( .A(n7637), .ZN(n7639) );
  NOR2_X1 U9414 ( .A1(n7639), .A2(n7638), .ZN(n7660) );
  INV_X1 U9415 ( .A(n7640), .ZN(n7645) );
  OAI211_X1 U9416 ( .C1(n7643), .C2(n7642), .A(n7722), .B(n7641), .ZN(n7644)
         );
  AOI211_X1 U9417 ( .C1(n7646), .C2(n9397), .A(n7645), .B(n7644), .ZN(n7649)
         );
  NAND4_X1 U9418 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7647), .ZN(n7652)
         );
  AOI21_X1 U9419 ( .B1(n7653), .B2(n7652), .A(n7651), .ZN(n7656) );
  OAI21_X1 U9420 ( .B1(n7656), .B2(n7655), .A(n7654), .ZN(n7659) );
  AOI211_X1 U9421 ( .C1(n7660), .C2(n7659), .A(n7658), .B(n7657), .ZN(n7664)
         );
  INV_X1 U9422 ( .A(n7661), .ZN(n7662) );
  OAI21_X1 U9423 ( .B1(n7664), .B2(n7663), .A(n7662), .ZN(n7667) );
  AOI21_X1 U9424 ( .B1(n7667), .B2(n7731), .A(n7666), .ZN(n7670) );
  OAI21_X1 U9425 ( .B1(n7670), .B2(n7669), .A(n7668), .ZN(n7673) );
  INV_X1 U9426 ( .A(n9606), .ZN(n7672) );
  INV_X1 U9427 ( .A(n7692), .ZN(n7671) );
  AOI211_X1 U9428 ( .C1(n7695), .C2(n7673), .A(n7672), .B(n7671), .ZN(n7674)
         );
  INV_X1 U9429 ( .A(n7825), .ZN(n7737) );
  AOI21_X1 U9430 ( .B1(n7728), .B2(n7674), .A(n7737), .ZN(n7676) );
  NAND2_X1 U9431 ( .A1(n7675), .A2(n7688), .ZN(n7741) );
  AOI21_X1 U9432 ( .B1(n7727), .B2(n7676), .A(n7741), .ZN(n7679) );
  NOR2_X1 U9433 ( .A1(n7678), .A2(n7677), .ZN(n7746) );
  OAI21_X1 U9434 ( .B1(n7680), .B2(n7679), .A(n7746), .ZN(n7682) );
  INV_X1 U9435 ( .A(n9372), .ZN(n7831) );
  AOI21_X1 U9436 ( .B1(n7831), .B2(n9487), .A(n7681), .ZN(n7743) );
  AOI22_X1 U9437 ( .A1(n7682), .A2(n7743), .B1(n9937), .B2(n9372), .ZN(n7683)
         );
  OAI21_X1 U9438 ( .B1(n7683), .B2(n7721), .A(n7757), .ZN(n7725) );
  NAND2_X1 U9439 ( .A1(n7685), .A2(n7766), .ZN(n7723) );
  XOR2_X1 U9440 ( .A(n9372), .B(n9487), .Z(n7720) );
  NAND2_X1 U9441 ( .A1(n7687), .A2(n7686), .ZN(n7830) );
  NAND2_X1 U9442 ( .A1(n9522), .A2(n7689), .ZN(n7824) );
  NAND2_X1 U9443 ( .A1(n7690), .A2(n7822), .ZN(n9574) );
  INV_X1 U9444 ( .A(n9592), .ZN(n9588) );
  INV_X1 U9445 ( .A(n7693), .ZN(n7694) );
  NAND2_X1 U9446 ( .A1(n7694), .A2(n7732), .ZN(n9654) );
  NAND2_X1 U9447 ( .A1(n7696), .A2(n7695), .ZN(n9639) );
  NAND4_X1 U9448 ( .A1(n10056), .A2(n7699), .A3(n7698), .A4(n6238), .ZN(n7701)
         );
  NOR4_X1 U9449 ( .A1(n7703), .A2(n7702), .A3(n7701), .A4(n7700), .ZN(n7704)
         );
  NAND4_X1 U9450 ( .A1(n7707), .A2(n7706), .A3(n7705), .A4(n7704), .ZN(n7708)
         );
  NOR4_X1 U9451 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n7713)
         );
  NAND4_X1 U9452 ( .A1(n9694), .A2(n7714), .A3(n7713), .A4(n7712), .ZN(n7715)
         );
  NOR4_X1 U9453 ( .A1(n9654), .A2(n9639), .A3(n9673), .A4(n7715), .ZN(n7716)
         );
  XNOR2_X1 U9454 ( .A(n9627), .B(n9380), .ZN(n9618) );
  NAND4_X1 U9455 ( .A1(n9588), .A2(n9604), .A3(n7716), .A4(n9618), .ZN(n7717)
         );
  NOR4_X1 U9456 ( .A1(n7824), .A2(n9559), .A3(n9574), .A4(n7717), .ZN(n7718)
         );
  NAND4_X1 U9457 ( .A1(n9493), .A2(n9508), .A3(n9523), .A4(n7718), .ZN(n7719)
         );
  NOR4_X1 U9458 ( .A1(n7721), .A2(n7720), .A3(n7830), .A4(n7719), .ZN(n7750)
         );
  AOI22_X1 U9459 ( .A1(n7723), .A2(n7722), .B1(n7750), .B2(n7757), .ZN(n7724)
         );
  NOR2_X1 U9460 ( .A1(n7725), .A2(n6098), .ZN(n7726) );
  INV_X1 U9461 ( .A(n7727), .ZN(n7739) );
  INV_X1 U9462 ( .A(n7728), .ZN(n7736) );
  INV_X1 U9463 ( .A(n9639), .ZN(n9636) );
  INV_X1 U9464 ( .A(n7734), .ZN(n7735) );
  NOR3_X1 U9465 ( .A1(n7736), .A2(n9620), .A3(n7735), .ZN(n7738) );
  NOR3_X1 U9466 ( .A1(n7739), .A2(n7738), .A3(n7737), .ZN(n7742) );
  OAI21_X1 U9467 ( .B1(n7742), .B2(n7741), .A(n7740), .ZN(n7745) );
  INV_X1 U9468 ( .A(n7743), .ZN(n7744) );
  AOI21_X1 U9469 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7749) );
  NOR2_X1 U9470 ( .A1(n9487), .A2(n7747), .ZN(n7748) );
  OAI22_X1 U9471 ( .A1(n7749), .A2(n7748), .B1(n9937), .B2(n9484), .ZN(n7751)
         );
  AOI21_X1 U9472 ( .B1(n7752), .B2(n7751), .A(n7750), .ZN(n7756) );
  OAI22_X1 U9473 ( .A1(n7756), .A2(n7755), .B1(n7754), .B2(n7753), .ZN(n7758)
         );
  AND2_X1 U9474 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U9475 ( .A1(n7759), .A2(n5757), .ZN(n7760) );
  NAND3_X1 U9476 ( .A1(n9853), .A2(n7764), .A3(n7763), .ZN(n7765) );
  OAI211_X1 U9477 ( .C1(n7766), .C2(n7768), .A(n7765), .B(P1_B_REG_SCAN_IN), 
        .ZN(n7767) );
  OAI222_X1 U9478 ( .A1(n9872), .A2(n7770), .B1(n7769), .B2(P1_U3086), .C1(
        n8870), .C2(n9868), .ZN(P1_U3327) );
  AOI22_X1 U9479 ( .A1(n7935), .A2(n10211), .B1(n10235), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n7771) );
  OAI21_X1 U9480 ( .B1(n8242), .B2(n8516), .A(n7771), .ZN(n7772) );
  AOI21_X1 U9481 ( .B1(n7773), .B2(n10213), .A(n7772), .ZN(n7774) );
  OAI21_X1 U9482 ( .B1(n7775), .B2(n10235), .A(n7774), .ZN(P2_U3205) );
  OAI222_X1 U9483 ( .A1(n9872), .A2(n7777), .B1(n4416), .B2(P1_U3086), .C1(
        n7776), .C2(n9868), .ZN(P1_U3328) );
  INV_X1 U9484 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8943) );
  OAI222_X1 U9485 ( .A1(n9868), .A2(n8943), .B1(n9872), .B2(n7778), .C1(
        P1_U3086), .C2(n5757), .ZN(P1_U3336) );
  OAI222_X1 U9486 ( .A1(n9868), .A2(n7781), .B1(n9872), .B2(n7780), .C1(
        P1_U3086), .C2(n7779), .ZN(P1_U3333) );
  OR2_X1 U9487 ( .A1(n7787), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7782) );
  NAND2_X1 U9488 ( .A1(n10032), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7785) );
  OR2_X1 U9489 ( .A1(n10032), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7784) );
  AND2_X1 U9490 ( .A1(n7785), .A2(n7784), .ZN(n10026) );
  NAND2_X1 U9491 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  NAND2_X1 U9492 ( .A1(n10025), .A2(n7785), .ZN(n7786) );
  XNOR2_X1 U9493 ( .A(n7786), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n7795) );
  INV_X1 U9494 ( .A(n7795), .ZN(n7792) );
  OAI22_X1 U9495 ( .A1(n7789), .A2(n7788), .B1(P1_REG1_REG_17__SCAN_IN), .B2(
        n7787), .ZN(n10030) );
  NAND2_X1 U9496 ( .A1(n10032), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7790) );
  OAI21_X1 U9497 ( .B1(n10032), .B2(P1_REG1_REG_18__SCAN_IN), .A(n7790), .ZN(
        n10029) );
  OR2_X1 U9498 ( .A1(n10030), .A2(n10029), .ZN(n10033) );
  NAND2_X1 U9499 ( .A1(n10033), .A2(n7790), .ZN(n7791) );
  XOR2_X1 U9500 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n7791), .Z(n7793) );
  AOI22_X1 U9501 ( .A1(n7792), .A2(n10024), .B1(n7793), .B2(n9474), .ZN(n7797)
         );
  NOR2_X1 U9502 ( .A1(n7793), .A2(n10028), .ZN(n7794) );
  AOI211_X1 U9503 ( .C1(n10024), .C2(n7795), .A(n10031), .B(n7794), .ZN(n7796)
         );
  MUX2_X1 U9504 ( .A(n7797), .B(n7796), .S(n4418), .Z(n7799) );
  NAND2_X1 U9505 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n7798) );
  OAI211_X1 U9506 ( .C1(n4603), .C2(n10039), .A(n7799), .B(n7798), .ZN(
        P1_U3262) );
  INV_X1 U9507 ( .A(n9840), .ZN(n9681) );
  INV_X1 U9508 ( .A(n9340), .ZN(n9382) );
  INV_X1 U9509 ( .A(n9068), .ZN(n9384) );
  INV_X1 U9510 ( .A(n9766), .ZN(n9669) );
  INV_X1 U9511 ( .A(n9648), .ZN(n9829) );
  NAND2_X1 U9512 ( .A1(n9829), .A2(n9341), .ZN(n7804) );
  INV_X1 U9513 ( .A(n9341), .ZN(n9381) );
  AOI21_X2 U9514 ( .B1(n9640), .B2(n7804), .A(n7803), .ZN(n9617) );
  NAND2_X1 U9515 ( .A1(n9617), .A2(n5008), .ZN(n7805) );
  INV_X1 U9516 ( .A(n9316), .ZN(n9379) );
  INV_X1 U9517 ( .A(n9315), .ZN(n9377) );
  NOR2_X1 U9518 ( .A1(n9558), .A2(n9247), .ZN(n7807) );
  NAND2_X1 U9519 ( .A1(n9558), .A2(n9247), .ZN(n7806) );
  INV_X1 U9520 ( .A(n9351), .ZN(n9376) );
  NOR2_X1 U9521 ( .A1(n9808), .A2(n9376), .ZN(n7809) );
  NAND2_X1 U9522 ( .A1(n9808), .A2(n9376), .ZN(n7808) );
  NOR2_X1 U9523 ( .A1(n9534), .A2(n9248), .ZN(n7811) );
  INV_X1 U9524 ( .A(n9724), .ZN(n9518) );
  NAND2_X1 U9525 ( .A1(n9518), .A2(n9353), .ZN(n7812) );
  INV_X1 U9526 ( .A(n9208), .ZN(n9374) );
  INV_X1 U9527 ( .A(n9719), .ZN(n9505) );
  NAND2_X1 U9528 ( .A1(n9691), .A2(n9783), .ZN(n9690) );
  NAND2_X1 U9529 ( .A1(n9669), .A2(n9662), .ZN(n9644) );
  NAND2_X1 U9530 ( .A1(n9558), .A2(n9580), .ZN(n9555) );
  NOR2_X1 U9531 ( .A1(n9555), .A2(n9808), .ZN(n9528) );
  NAND2_X1 U9532 ( .A1(n9534), .A2(n9528), .ZN(n9529) );
  AOI211_X1 U9533 ( .C1(n7814), .C2(n9498), .A(n9664), .B(n9488), .ZN(n7836)
         );
  INV_X1 U9534 ( .A(P1_B_REG_SCAN_IN), .ZN(n7815) );
  NOR2_X1 U9535 ( .A1(n4416), .A2(n7815), .ZN(n7816) );
  OR2_X1 U9536 ( .A1(n9352), .A2(n7816), .ZN(n9482) );
  NAND2_X1 U9537 ( .A1(n9589), .A2(n7819), .ZN(n7821) );
  INV_X1 U9538 ( .A(n9574), .ZN(n9570) );
  INV_X1 U9539 ( .A(n7822), .ZN(n9560) );
  INV_X1 U9540 ( .A(n7824), .ZN(n9542) );
  NAND2_X1 U9541 ( .A1(n7826), .A2(n7825), .ZN(n9511) );
  OAI21_X1 U9542 ( .B1(n7845), .B2(n9775), .A(n7834), .ZN(P1_U3551) );
  NOR2_X1 U9543 ( .A1(n9581), .A2(n4418), .ZN(n9628) );
  NAND2_X1 U9544 ( .A1(n7836), .A2(n9628), .ZN(n7840) );
  INV_X1 U9545 ( .A(n7837), .ZN(n7838) );
  AOI22_X1 U9546 ( .A1(n9581), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n7838), .B2(
        n10065), .ZN(n7839) );
  OAI211_X1 U9547 ( .C1(n7841), .C2(n10062), .A(n7840), .B(n7839), .ZN(n7842)
         );
  AOI21_X1 U9548 ( .B1(n7843), .B2(n10067), .A(n7842), .ZN(n7844) );
  OAI21_X1 U9549 ( .B1(n7845), .B2(n9701), .A(n7844), .ZN(P1_U3356) );
  NOR2_X1 U9550 ( .A1(n8239), .A2(n8455), .ZN(n7846) );
  INV_X1 U9551 ( .A(n8455), .ZN(n7908) );
  NAND2_X1 U9552 ( .A1(n7848), .A2(n8060), .ZN(n7850) );
  NAND2_X1 U9553 ( .A1(n8061), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7849) );
  NAND2_X1 U9554 ( .A1(n8445), .A2(n7938), .ZN(n8067) );
  NAND2_X1 U9555 ( .A1(n8244), .A2(n8067), .ZN(n7853) );
  NAND2_X1 U9556 ( .A1(n8239), .A2(n7908), .ZN(n7851) );
  INV_X1 U9557 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U9558 ( .A1(n4414), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7856) );
  NAND2_X1 U9559 ( .A1(n7854), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7855) );
  OAI211_X1 U9560 ( .C1(n7858), .C2(n7857), .A(n7856), .B(n7855), .ZN(n7859)
         );
  INV_X1 U9561 ( .A(n7859), .ZN(n7860) );
  AND2_X1 U9562 ( .A1(n8032), .A2(n7860), .ZN(n8064) );
  NAND2_X1 U9563 ( .A1(n5181), .A2(P2_B_REG_SCAN_IN), .ZN(n7861) );
  NAND2_X1 U9564 ( .A1(n10202), .A2(n7861), .ZN(n8438) );
  OAI22_X1 U9565 ( .A1(n7908), .A2(n10220), .B1(n8064), .B2(n8438), .ZN(n7862)
         );
  AOI21_X1 U9566 ( .B1(n7864), .B2(n10230), .A(n7862), .ZN(n7863) );
  INV_X1 U9567 ( .A(n7864), .ZN(n8452) );
  NOR2_X1 U9568 ( .A1(n8452), .A2(n10284), .ZN(n7865) );
  MUX2_X1 U9569 ( .A(n7866), .B(n7870), .S(n10300), .Z(n7868) );
  NAND2_X1 U9570 ( .A1(n8445), .A2(n5662), .ZN(n7867) );
  NAND2_X1 U9571 ( .A1(n7868), .A2(n7867), .ZN(P2_U3456) );
  INV_X1 U9572 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n7869) );
  MUX2_X1 U9573 ( .A(n7870), .B(n7869), .S(n10323), .Z(n7872) );
  NAND2_X1 U9574 ( .A1(n8445), .A2(n8646), .ZN(n7871) );
  NAND2_X1 U9575 ( .A1(n7872), .A2(n7871), .ZN(P2_U3488) );
  XNOR2_X1 U9576 ( .A(n8667), .B(n4415), .ZN(n7900) );
  XNOR2_X1 U9577 ( .A(n8677), .B(n4415), .ZN(n7913) );
  NAND2_X1 U9578 ( .A1(n7876), .A2(n8599), .ZN(n7877) );
  XNOR2_X1 U9579 ( .A(n8706), .B(n7896), .ZN(n7878) );
  NAND2_X1 U9580 ( .A1(n7878), .A2(n8565), .ZN(n7881) );
  INV_X1 U9581 ( .A(n7878), .ZN(n7879) );
  NAND2_X1 U9582 ( .A1(n7879), .A2(n8588), .ZN(n7880) );
  NAND2_X1 U9583 ( .A1(n7881), .A2(n7880), .ZN(n7965) );
  XNOR2_X1 U9584 ( .A(n8571), .B(n4415), .ZN(n7882) );
  XNOR2_X1 U9585 ( .A(n7882), .B(n7967), .ZN(n8005) );
  NAND2_X1 U9586 ( .A1(n8004), .A2(n8005), .ZN(n8003) );
  XNOR2_X1 U9587 ( .A(n8556), .B(n4415), .ZN(n7888) );
  XNOR2_X1 U9588 ( .A(n7888), .B(n8566), .ZN(n7924) );
  INV_X1 U9589 ( .A(n7882), .ZN(n7883) );
  NAND2_X1 U9590 ( .A1(n7883), .A2(n7967), .ZN(n7923) );
  AND2_X1 U9591 ( .A1(n7924), .A2(n7923), .ZN(n7884) );
  XNOR2_X1 U9592 ( .A(n8632), .B(n7896), .ZN(n7885) );
  NAND2_X1 U9593 ( .A1(n7885), .A2(n7946), .ZN(n7942) );
  INV_X1 U9594 ( .A(n7885), .ZN(n7886) );
  NAND2_X1 U9595 ( .A1(n7886), .A2(n8551), .ZN(n7887) );
  NAND2_X1 U9596 ( .A1(n7942), .A2(n7887), .ZN(n7984) );
  AND2_X1 U9597 ( .A1(n7888), .A2(n8535), .ZN(n7983) );
  NOR2_X1 U9598 ( .A1(n7984), .A2(n7983), .ZN(n7889) );
  XNOR2_X1 U9599 ( .A(n8687), .B(n7896), .ZN(n7890) );
  NAND2_X1 U9600 ( .A1(n7890), .A2(n8510), .ZN(n7893) );
  INV_X1 U9601 ( .A(n7890), .ZN(n7891) );
  INV_X1 U9602 ( .A(n8510), .ZN(n8536) );
  NAND2_X1 U9603 ( .A1(n7891), .A2(n8536), .ZN(n7892) );
  AND2_X1 U9604 ( .A1(n7893), .A2(n7892), .ZN(n7943) );
  XNOR2_X1 U9605 ( .A(n8684), .B(n4415), .ZN(n7894) );
  XNOR2_X1 U9606 ( .A(n7894), .B(n8525), .ZN(n7995) );
  NAND2_X1 U9607 ( .A1(n7994), .A2(n7995), .ZN(n7993) );
  NAND2_X1 U9608 ( .A1(n7894), .A2(n8500), .ZN(n7895) );
  NAND2_X1 U9609 ( .A1(n7993), .A2(n7895), .ZN(n7914) );
  XNOR2_X1 U9610 ( .A(n8672), .B(n7896), .ZN(n7897) );
  NAND2_X1 U9611 ( .A1(n7897), .A2(n8474), .ZN(n7951) );
  INV_X1 U9612 ( .A(n7897), .ZN(n7898) );
  NAND2_X1 U9613 ( .A1(n7898), .A2(n8501), .ZN(n7952) );
  NAND3_X1 U9614 ( .A1(n7951), .A2(n8511), .A3(n7913), .ZN(n7899) );
  XNOR2_X1 U9615 ( .A(n7900), .B(n8486), .ZN(n7953) );
  XNOR2_X1 U9616 ( .A(n8012), .B(n4415), .ZN(n7901) );
  XNOR2_X1 U9617 ( .A(n7903), .B(n7901), .ZN(n8014) );
  NAND2_X1 U9618 ( .A1(n8014), .A2(n8015), .ZN(n8013) );
  INV_X1 U9619 ( .A(n7901), .ZN(n7902) );
  NAND2_X1 U9620 ( .A1(n7903), .A2(n7902), .ZN(n7904) );
  AND2_X1 U9621 ( .A1(n8013), .A2(n7904), .ZN(n7906) );
  XNOR2_X1 U9622 ( .A(n7912), .B(n4415), .ZN(n7931) );
  XNOR2_X1 U9623 ( .A(n7931), .B(n8271), .ZN(n7905) );
  NAND3_X1 U9624 ( .A1(n8013), .A2(n7905), .A3(n7904), .ZN(n7930) );
  OAI211_X1 U9625 ( .C1(n7906), .C2(n7905), .A(n8016), .B(n7930), .ZN(n7911)
         );
  AOI22_X1 U9626 ( .A1(n8475), .A2(n8018), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7907) );
  OAI21_X1 U9627 ( .B1(n7908), .B2(n8020), .A(n7907), .ZN(n7909) );
  AOI21_X1 U9628 ( .B1(n8458), .B2(n8022), .A(n7909), .ZN(n7910) );
  OAI211_X1 U9629 ( .C1(n7912), .C2(n8025), .A(n7911), .B(n7910), .ZN(P2_U3154) );
  OR2_X1 U9630 ( .A1(n7914), .A2(n7913), .ZN(n7916) );
  NAND2_X1 U9631 ( .A1(n7916), .A2(n8511), .ZN(n7976) );
  NAND2_X1 U9632 ( .A1(n7914), .A2(n7913), .ZN(n7975) );
  INV_X1 U9633 ( .A(n7975), .ZN(n7915) );
  NOR2_X1 U9634 ( .A1(n7976), .A2(n7915), .ZN(n7918) );
  AOI21_X1 U9635 ( .B1(n7916), .B2(n7975), .A(n8511), .ZN(n7917) );
  OAI21_X1 U9636 ( .B1(n7918), .B2(n7917), .A(n8016), .ZN(n7922) );
  AOI22_X1 U9637 ( .A1(n8474), .A2(n7997), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7919) );
  OAI21_X1 U9638 ( .B1(n8500), .B2(n7999), .A(n7919), .ZN(n7920) );
  AOI21_X1 U9639 ( .B1(n8504), .B2(n8022), .A(n7920), .ZN(n7921) );
  OAI211_X1 U9640 ( .C1(n8677), .C2(n8025), .A(n7922), .B(n7921), .ZN(P2_U3156) );
  INV_X1 U9641 ( .A(n8556), .ZN(n8695) );
  AND2_X1 U9642 ( .A1(n8003), .A2(n7923), .ZN(n7925) );
  OAI211_X1 U9643 ( .C1(n7925), .C2(n7924), .A(n8016), .B(n7987), .ZN(n7929)
         );
  NOR2_X1 U9644 ( .A1(n8977), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8433) );
  AOI21_X1 U9645 ( .B1(n7997), .B2(n8551), .A(n8433), .ZN(n7926) );
  OAI21_X1 U9646 ( .B1(n7967), .B2(n7999), .A(n7926), .ZN(n7927) );
  AOI21_X1 U9647 ( .B1(n8555), .B2(n8022), .A(n7927), .ZN(n7928) );
  OAI211_X1 U9648 ( .C1(n8695), .C2(n8025), .A(n7929), .B(n7928), .ZN(P2_U3159) );
  OAI21_X1 U9649 ( .B1(n8463), .B2(n7931), .A(n7930), .ZN(n7934) );
  XOR2_X1 U9650 ( .A(n4415), .B(n8058), .Z(n7933) );
  XNOR2_X1 U9651 ( .A(n7934), .B(n7933), .ZN(n7941) );
  AOI22_X1 U9652 ( .A1(n8271), .A2(n8018), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7937) );
  NAND2_X1 U9653 ( .A1(n7935), .A2(n8022), .ZN(n7936) );
  OAI211_X1 U9654 ( .C1(n7938), .C2(n8020), .A(n7937), .B(n7936), .ZN(n7939)
         );
  AOI21_X1 U9655 ( .B1(n8239), .B2(n7969), .A(n7939), .ZN(n7940) );
  OAI21_X1 U9656 ( .B1(n7941), .B2(n7972), .A(n7940), .ZN(P2_U3160) );
  NOR3_X1 U9657 ( .A1(n4439), .A2(n4723), .A3(n7943), .ZN(n7944) );
  OAI21_X1 U9658 ( .B1(n7944), .B2(n4472), .A(n8016), .ZN(n7949) );
  AOI22_X1 U9659 ( .A1(n7997), .A2(n8525), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7945) );
  OAI21_X1 U9660 ( .B1(n7946), .B2(n7999), .A(n7945), .ZN(n7947) );
  AOI21_X1 U9661 ( .B1(n8528), .B2(n8022), .A(n7947), .ZN(n7948) );
  OAI211_X1 U9662 ( .C1(n7950), .C2(n8025), .A(n7949), .B(n7948), .ZN(P2_U3163) );
  INV_X1 U9663 ( .A(n8667), .ZN(n8471) );
  NAND2_X1 U9664 ( .A1(n7951), .A2(n7952), .ZN(n7974) );
  AOI21_X1 U9665 ( .B1(n7976), .B2(n7975), .A(n7974), .ZN(n7978) );
  INV_X1 U9666 ( .A(n7952), .ZN(n7954) );
  NOR3_X1 U9667 ( .A1(n7978), .A2(n7954), .A3(n7953), .ZN(n7957) );
  INV_X1 U9668 ( .A(n7955), .ZN(n7956) );
  OAI21_X1 U9669 ( .B1(n7957), .B2(n7956), .A(n8016), .ZN(n7961) );
  NOR2_X1 U9670 ( .A1(n8501), .A2(n7999), .ZN(n7959) );
  OAI22_X1 U9671 ( .A1(n8015), .A2(n8020), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8831), .ZN(n7958) );
  AOI211_X1 U9672 ( .C1(n8479), .C2(n8022), .A(n7959), .B(n7958), .ZN(n7960)
         );
  OAI211_X1 U9673 ( .C1(n8471), .C2(n8025), .A(n7961), .B(n7960), .ZN(P2_U3165) );
  INV_X1 U9674 ( .A(n7962), .ZN(n7963) );
  AOI21_X1 U9675 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(n7973) );
  NAND2_X1 U9676 ( .A1(n8018), .A2(n8599), .ZN(n7966) );
  NAND2_X1 U9677 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8394) );
  OAI211_X1 U9678 ( .C1(n7967), .C2(n8020), .A(n7966), .B(n8394), .ZN(n7968)
         );
  AOI21_X1 U9679 ( .B1(n8581), .B2(n8022), .A(n7968), .ZN(n7971) );
  NAND2_X1 U9680 ( .A1(n8706), .A2(n7969), .ZN(n7970) );
  OAI211_X1 U9681 ( .C1(n7973), .C2(n7972), .A(n7971), .B(n7970), .ZN(P2_U3168) );
  AND3_X1 U9682 ( .A1(n7976), .A2(n7975), .A3(n7974), .ZN(n7977) );
  OAI21_X1 U9683 ( .B1(n7978), .B2(n7977), .A(n8016), .ZN(n7982) );
  AOI22_X1 U9684 ( .A1(n8272), .A2(n7997), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7979) );
  OAI21_X1 U9685 ( .B1(n8511), .B2(n7999), .A(n7979), .ZN(n7980) );
  AOI21_X1 U9686 ( .B1(n8488), .B2(n8022), .A(n7980), .ZN(n7981) );
  OAI211_X1 U9687 ( .C1(n8672), .C2(n8025), .A(n7982), .B(n7981), .ZN(P2_U3169) );
  INV_X1 U9688 ( .A(n7983), .ZN(n7986) );
  INV_X1 U9689 ( .A(n7984), .ZN(n7985) );
  AOI21_X1 U9690 ( .B1(n7987), .B2(n7986), .A(n7985), .ZN(n7988) );
  OAI21_X1 U9691 ( .B1(n4439), .B2(n7988), .A(n8016), .ZN(n7992) );
  AOI22_X1 U9692 ( .A1(n7997), .A2(n8536), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7989) );
  OAI21_X1 U9693 ( .B1(n8566), .B2(n7999), .A(n7989), .ZN(n7990) );
  AOI21_X1 U9694 ( .B1(n8539), .B2(n8022), .A(n7990), .ZN(n7991) );
  OAI211_X1 U9695 ( .C1(n5466), .C2(n8025), .A(n7992), .B(n7991), .ZN(P2_U3173) );
  OAI21_X1 U9696 ( .B1(n7995), .B2(n7994), .A(n7993), .ZN(n7996) );
  NAND2_X1 U9697 ( .A1(n7996), .A2(n8016), .ZN(n8002) );
  AOI22_X1 U9698 ( .A1(n8273), .A2(n7997), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7998) );
  OAI21_X1 U9699 ( .B1(n8510), .B2(n7999), .A(n7998), .ZN(n8000) );
  AOI21_X1 U9700 ( .B1(n8514), .B2(n8022), .A(n8000), .ZN(n8001) );
  OAI211_X1 U9701 ( .C1(n8684), .C2(n8025), .A(n8002), .B(n8001), .ZN(P2_U3175) );
  INV_X1 U9702 ( .A(n8571), .ZN(n8703) );
  OAI21_X1 U9703 ( .B1(n8005), .B2(n8004), .A(n8003), .ZN(n8006) );
  NAND2_X1 U9704 ( .A1(n8006), .A2(n8016), .ZN(n8011) );
  NAND2_X1 U9705 ( .A1(n8018), .A2(n8588), .ZN(n8008) );
  NAND2_X1 U9706 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9882) );
  OAI211_X1 U9707 ( .C1(n8566), .C2(n8020), .A(n8008), .B(n9882), .ZN(n8009)
         );
  AOI21_X1 U9708 ( .B1(n8567), .B2(n8022), .A(n8009), .ZN(n8010) );
  OAI211_X1 U9709 ( .C1(n8703), .C2(n8025), .A(n8011), .B(n8010), .ZN(P2_U3178) );
  OAI21_X1 U9710 ( .B1(n8015), .B2(n8014), .A(n8013), .ZN(n8017) );
  NAND2_X1 U9711 ( .A1(n8017), .A2(n8016), .ZN(n8024) );
  AOI22_X1 U9712 ( .A1(n8272), .A2(n8018), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8019) );
  OAI21_X1 U9713 ( .B1(n8463), .B2(n8020), .A(n8019), .ZN(n8021) );
  AOI21_X1 U9714 ( .B1(n8466), .B2(n8022), .A(n8021), .ZN(n8023) );
  OAI211_X1 U9715 ( .C1(n8665), .C2(n8025), .A(n8024), .B(n8023), .ZN(P2_U3180) );
  NAND2_X1 U9716 ( .A1(n8723), .A2(n8060), .ZN(n8027) );
  NAND2_X1 U9717 ( .A1(n8061), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8026) );
  NAND2_X1 U9718 ( .A1(n5184), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U9719 ( .A1(n4414), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U9720 ( .A1(n7854), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8028) );
  AND3_X1 U9721 ( .A1(n8030), .A2(n8029), .A3(n8028), .ZN(n8031) );
  NAND2_X1 U9722 ( .A1(n8032), .A2(n8031), .ZN(n8269) );
  NAND2_X1 U9723 ( .A1(n8652), .A2(n8269), .ZN(n8069) );
  INV_X1 U9724 ( .A(n8069), .ZN(n8259) );
  INV_X1 U9725 ( .A(n8033), .ZN(n8234) );
  INV_X1 U9726 ( .A(n8230), .ZN(n8034) );
  NAND2_X1 U9727 ( .A1(n8217), .A2(n8215), .ZN(n8491) );
  INV_X1 U9728 ( .A(n8489), .ZN(n8035) );
  NOR2_X1 U9729 ( .A1(n8213), .A2(n8035), .ZN(n8498) );
  INV_X1 U9730 ( .A(n8523), .ZN(n8056) );
  INV_X1 U9731 ( .A(n8546), .ZN(n8054) );
  NOR3_X1 U9732 ( .A1(n8037), .A2(n5600), .A3(n8036), .ZN(n8039) );
  NAND4_X1 U9733 ( .A1(n8039), .A2(n8038), .A3(n10208), .A4(n8096), .ZN(n8042)
         );
  NOR4_X1 U9734 ( .A1(n8042), .A2(n8041), .A3(n4976), .A4(n8040), .ZN(n8046)
         );
  NAND4_X1 U9735 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(n8048)
         );
  NOR4_X1 U9736 ( .A1(n5379), .A2(n8048), .A3(n8047), .A4(n8152), .ZN(n8052)
         );
  INV_X1 U9737 ( .A(n8049), .ZN(n8051) );
  NAND4_X1 U9738 ( .A1(n5613), .A2(n8585), .A3(n8052), .A4(n8596), .ZN(n8053)
         );
  NOR4_X1 U9739 ( .A1(n8533), .A2(n8054), .A3(n8175), .A4(n8053), .ZN(n8055)
         );
  NAND4_X1 U9740 ( .A1(n8498), .A2(n8512), .A3(n8056), .A4(n8055), .ZN(n8057)
         );
  NOR4_X1 U9741 ( .A1(n8223), .A2(n8472), .A3(n8491), .A4(n8057), .ZN(n8059)
         );
  NAND4_X1 U9742 ( .A1(n4758), .A2(n4438), .A3(n8059), .A4(n8058), .ZN(n8066)
         );
  NAND2_X1 U9743 ( .A1(n8728), .A2(n8060), .ZN(n8063) );
  NAND2_X1 U9744 ( .A1(n8061), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8062) );
  INV_X1 U9745 ( .A(n8064), .ZN(n8270) );
  INV_X1 U9746 ( .A(n8655), .ZN(n8065) );
  NAND2_X1 U9747 ( .A1(n8065), .A2(n8064), .ZN(n8068) );
  INV_X1 U9748 ( .A(n8068), .ZN(n8250) );
  NOR4_X1 U9749 ( .A1(n8259), .A2(n8066), .A3(n8243), .A4(n8250), .ZN(n8072)
         );
  NAND2_X1 U9750 ( .A1(n8068), .A2(n8067), .ZN(n8252) );
  OAI21_X1 U9751 ( .B1(n8655), .B2(n8606), .A(n8069), .ZN(n8070) );
  NAND2_X1 U9752 ( .A1(n8445), .A2(n8249), .ZN(n8073) );
  NAND2_X1 U9753 ( .A1(n8244), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U9754 ( .A1(n8075), .A2(n8074), .ZN(n8240) );
  NAND2_X1 U9755 ( .A1(n8084), .A2(n8076), .ZN(n8077) );
  NAND2_X1 U9756 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  NAND2_X1 U9757 ( .A1(n8079), .A2(n8256), .ZN(n8083) );
  INV_X1 U9758 ( .A(n8080), .ZN(n8081) );
  OAI21_X1 U9759 ( .B1(n8083), .B2(n8081), .A(n8256), .ZN(n8082) );
  MUX2_X1 U9760 ( .A(n8256), .B(n8082), .S(n5601), .Z(n8087) );
  INV_X1 U9761 ( .A(n5600), .ZN(n8085) );
  NAND3_X1 U9762 ( .A1(n8085), .A2(n8084), .A3(n8083), .ZN(n8086) );
  NAND3_X1 U9763 ( .A1(n8087), .A2(n10224), .A3(n8086), .ZN(n8095) );
  NAND2_X1 U9764 ( .A1(n8283), .A2(n8088), .ZN(n8104) );
  NAND2_X1 U9765 ( .A1(n8089), .A2(n8104), .ZN(n8092) );
  NAND2_X1 U9766 ( .A1(n8090), .A2(n8098), .ZN(n8091) );
  MUX2_X1 U9767 ( .A(n8092), .B(n8091), .S(n8256), .Z(n8093) );
  INV_X1 U9768 ( .A(n8093), .ZN(n8094) );
  NAND2_X1 U9769 ( .A1(n8095), .A2(n8094), .ZN(n8097) );
  NAND2_X1 U9770 ( .A1(n8097), .A2(n8096), .ZN(n8107) );
  INV_X1 U9771 ( .A(n8098), .ZN(n8101) );
  NAND2_X1 U9772 ( .A1(n10203), .A2(n8099), .ZN(n8100) );
  OAI211_X1 U9773 ( .C1(n8107), .C2(n8101), .A(n8100), .B(n8108), .ZN(n8103)
         );
  AOI21_X1 U9774 ( .B1(n8103), .B2(n8102), .A(n4973), .ZN(n8117) );
  INV_X1 U9775 ( .A(n8104), .ZN(n8106) );
  OAI21_X1 U9776 ( .B1(n8107), .B2(n8106), .A(n8105), .ZN(n8109) );
  NAND2_X1 U9777 ( .A1(n8109), .A2(n8108), .ZN(n8111) );
  NAND2_X1 U9778 ( .A1(n8111), .A2(n8110), .ZN(n8115) );
  INV_X1 U9779 ( .A(n8112), .ZN(n8113) );
  AOI21_X1 U9780 ( .B1(n8115), .B2(n8114), .A(n8113), .ZN(n8116) );
  MUX2_X1 U9781 ( .A(n8117), .B(n8116), .S(n8256), .Z(n8123) );
  AND2_X1 U9782 ( .A1(n8126), .A2(n8127), .ZN(n8121) );
  AND2_X1 U9783 ( .A1(n8119), .A2(n8118), .ZN(n8120) );
  MUX2_X1 U9784 ( .A(n8121), .B(n8120), .S(n8249), .Z(n8124) );
  NAND3_X1 U9785 ( .A1(n8123), .A2(n8122), .A3(n8124), .ZN(n8147) );
  INV_X1 U9786 ( .A(n8124), .ZN(n8131) );
  AND2_X1 U9787 ( .A1(n8126), .A2(n8125), .ZN(n8128) );
  OAI211_X1 U9788 ( .C1(n8131), .C2(n8128), .A(n8136), .B(n8127), .ZN(n8133)
         );
  OAI21_X1 U9789 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8132) );
  MUX2_X1 U9790 ( .A(n8133), .B(n8132), .S(n8256), .Z(n8135) );
  NOR2_X1 U9791 ( .A1(n8135), .A2(n8134), .ZN(n8146) );
  INV_X1 U9792 ( .A(n8136), .ZN(n8137) );
  NAND2_X1 U9793 ( .A1(n8140), .A2(n8137), .ZN(n8138) );
  NAND2_X1 U9794 ( .A1(n8138), .A2(n8141), .ZN(n8144) );
  NAND2_X1 U9795 ( .A1(n8140), .A2(n8139), .ZN(n8142) );
  AND2_X1 U9796 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  MUX2_X1 U9797 ( .A(n8144), .B(n8143), .S(n8249), .Z(n8145) );
  AOI21_X1 U9798 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8153) );
  NAND2_X1 U9799 ( .A1(n10298), .A2(n8148), .ZN(n8149) );
  MUX2_X1 U9800 ( .A(n8150), .B(n8149), .S(n8256), .Z(n8151) );
  OAI21_X1 U9801 ( .B1(n8153), .B2(n8152), .A(n8151), .ZN(n8157) );
  MUX2_X1 U9802 ( .A(n8274), .B(n8154), .S(n8249), .Z(n8160) );
  NAND2_X1 U9803 ( .A1(n8160), .A2(n8155), .ZN(n8156) );
  NAND2_X1 U9804 ( .A1(n8157), .A2(n8156), .ZN(n8162) );
  INV_X1 U9805 ( .A(n8158), .ZN(n8159) );
  OR2_X1 U9806 ( .A1(n8160), .A2(n8159), .ZN(n8161) );
  NAND2_X1 U9807 ( .A1(n8162), .A2(n8161), .ZN(n8166) );
  NOR2_X1 U9808 ( .A1(n8163), .A2(n8249), .ZN(n8164) );
  AOI21_X1 U9809 ( .B1(n8166), .B2(n8165), .A(n8164), .ZN(n8172) );
  NAND2_X1 U9810 ( .A1(n8177), .A2(n8167), .ZN(n8168) );
  AOI21_X1 U9811 ( .B1(n8172), .B2(n8596), .A(n8168), .ZN(n8169) );
  MUX2_X1 U9812 ( .A(n8170), .B(n8169), .S(n8256), .Z(n8174) );
  NAND3_X1 U9813 ( .A1(n8172), .A2(n8596), .A3(n8171), .ZN(n8173) );
  NAND3_X1 U9814 ( .A1(n8174), .A2(n8179), .A3(n8173), .ZN(n8176) );
  INV_X1 U9815 ( .A(n8175), .ZN(n8576) );
  NAND2_X1 U9816 ( .A1(n8176), .A2(n8576), .ZN(n8182) );
  INV_X1 U9817 ( .A(n8177), .ZN(n8178) );
  NOR2_X1 U9818 ( .A1(n8182), .A2(n8178), .ZN(n8184) );
  INV_X1 U9819 ( .A(n8179), .ZN(n8181) );
  OAI211_X1 U9820 ( .C1(n8182), .C2(n8181), .A(n8180), .B(n8186), .ZN(n8183)
         );
  MUX2_X1 U9821 ( .A(n8184), .B(n8183), .S(n8256), .Z(n8193) );
  NAND2_X1 U9822 ( .A1(n8191), .A2(n8185), .ZN(n8187) );
  OAI211_X1 U9823 ( .C1(n8193), .C2(n8187), .A(n8194), .B(n8186), .ZN(n8190)
         );
  NAND4_X1 U9824 ( .A1(n8197), .A2(n8249), .A3(n8520), .A4(n8192), .ZN(n8188)
         );
  NOR2_X1 U9825 ( .A1(n8206), .A2(n8188), .ZN(n8189) );
  NAND2_X1 U9826 ( .A1(n8190), .A2(n8189), .ZN(n8212) );
  NAND3_X1 U9827 ( .A1(n8193), .A2(n8192), .A3(n8191), .ZN(n8211) );
  NAND4_X1 U9828 ( .A1(n8199), .A2(n8196), .A3(n8194), .A4(n8256), .ZN(n8195)
         );
  NOR2_X1 U9829 ( .A1(n8202), .A2(n8195), .ZN(n8210) );
  NAND2_X1 U9830 ( .A1(n8199), .A2(n8196), .ZN(n8198) );
  NAND3_X1 U9831 ( .A1(n8198), .A2(n8249), .A3(n8197), .ZN(n8205) );
  INV_X1 U9832 ( .A(n8199), .ZN(n8201) );
  OR4_X1 U9833 ( .A1(n8202), .A2(n8201), .A3(n8200), .A4(n8249), .ZN(n8204) );
  NAND2_X1 U9834 ( .A1(n8202), .A2(n8249), .ZN(n8203) );
  OAI211_X1 U9835 ( .C1(n8206), .C2(n8205), .A(n8204), .B(n8203), .ZN(n8209)
         );
  AOI21_X1 U9836 ( .B1(n8489), .B2(n8207), .A(n8249), .ZN(n8208) );
  INV_X1 U9837 ( .A(n8213), .ZN(n8214) );
  NAND2_X1 U9838 ( .A1(n8214), .A2(n8217), .ZN(n8216) );
  NAND2_X1 U9839 ( .A1(n8216), .A2(n8215), .ZN(n8221) );
  INV_X1 U9840 ( .A(n8217), .ZN(n8218) );
  OR2_X1 U9841 ( .A1(n8219), .A2(n8218), .ZN(n8220) );
  MUX2_X1 U9842 ( .A(n8221), .B(n8220), .S(n8249), .Z(n8222) );
  MUX2_X1 U9843 ( .A(n8225), .B(n8224), .S(n8249), .Z(n8226) );
  NAND3_X1 U9844 ( .A1(n8227), .A2(n8464), .A3(n8226), .ZN(n8232) );
  INV_X1 U9845 ( .A(n8228), .ZN(n8229) );
  MUX2_X1 U9846 ( .A(n8230), .B(n8229), .S(n8249), .Z(n8231) );
  NAND3_X1 U9847 ( .A1(n4438), .A2(n8232), .A3(n8231), .ZN(n8237) );
  MUX2_X1 U9848 ( .A(n8234), .B(n8233), .S(n8249), .Z(n8235) );
  INV_X1 U9849 ( .A(n8235), .ZN(n8236) );
  NAND2_X1 U9850 ( .A1(n8237), .A2(n8236), .ZN(n8238) );
  NAND2_X1 U9851 ( .A1(n8240), .A2(n8238), .ZN(n8248) );
  MUX2_X1 U9852 ( .A(n8455), .B(n8239), .S(n8256), .Z(n8246) );
  NAND2_X1 U9853 ( .A1(n8240), .A2(n8246), .ZN(n8241) );
  NAND2_X1 U9854 ( .A1(n8248), .A2(n8241), .ZN(n8251) );
  NAND2_X1 U9855 ( .A1(n8251), .A2(n8242), .ZN(n8245) );
  INV_X1 U9856 ( .A(n8243), .ZN(n8255) );
  INV_X1 U9857 ( .A(n8246), .ZN(n8247) );
  INV_X1 U9858 ( .A(n8251), .ZN(n8254) );
  INV_X1 U9859 ( .A(n8252), .ZN(n8253) );
  INV_X1 U9860 ( .A(n8269), .ZN(n8439) );
  AOI22_X1 U9861 ( .A1(n8257), .A2(n8260), .B1(n8439), .B2(n8606), .ZN(n8258)
         );
  XNOR2_X1 U9862 ( .A(n8261), .B(n8431), .ZN(n8268) );
  NOR2_X1 U9863 ( .A1(n8263), .A2(n8262), .ZN(n8266) );
  OAI21_X1 U9864 ( .B1(n8267), .B2(n8264), .A(P2_B_REG_SCAN_IN), .ZN(n8265) );
  OAI22_X1 U9865 ( .A1(n8268), .A2(n8267), .B1(n8266), .B2(n8265), .ZN(
        P2_U3296) );
  MUX2_X1 U9866 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8269), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9867 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8270), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9868 ( .A(n8455), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8285), .Z(
        P2_U3519) );
  MUX2_X1 U9869 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8271), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9870 ( .A(n8475), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8285), .Z(
        P2_U3517) );
  MUX2_X1 U9871 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8272), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9872 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8474), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9873 ( .A(n8273), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8285), .Z(
        P2_U3514) );
  MUX2_X1 U9874 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8525), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9875 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8536), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9876 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8551), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9877 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8535), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9878 ( .A(n8578), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8285), .Z(
        P2_U3509) );
  MUX2_X1 U9879 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8588), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9880 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8599), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9881 ( .A(n8587), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8285), .Z(
        P2_U3506) );
  MUX2_X1 U9882 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8598), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U9883 ( .A(n8274), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8285), .Z(
        P2_U3504) );
  MUX2_X1 U9884 ( .A(n8275), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8285), .Z(
        P2_U3503) );
  MUX2_X1 U9885 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8276), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U9886 ( .A(n8277), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8285), .Z(
        P2_U3501) );
  MUX2_X1 U9887 ( .A(n8278), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8285), .Z(
        P2_U3500) );
  MUX2_X1 U9888 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8279), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9889 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8280), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9890 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8281), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9891 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8282), .S(P2_U3893), .Z(
        P2_U3496) );
  MUX2_X1 U9892 ( .A(n10203), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8285), .Z(
        P2_U3495) );
  MUX2_X1 U9893 ( .A(n8283), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8285), .Z(
        P2_U3494) );
  MUX2_X1 U9894 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n10205), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9895 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8284), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U9896 ( .A(n8286), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8285), .Z(
        P2_U3491) );
  INV_X1 U9897 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8290) );
  AOI21_X1 U9898 ( .B1(n8290), .B2(n8289), .A(n8311), .ZN(n8309) );
  AOI21_X1 U9899 ( .B1(n8293), .B2(n8292), .A(n8291), .ZN(n8295) );
  MUX2_X1 U9900 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8426), .Z(n8317) );
  XNOR2_X1 U9901 ( .A(n8317), .B(n8327), .ZN(n8294) );
  NAND2_X1 U9902 ( .A1(n8295), .A2(n8294), .ZN(n8318) );
  OAI21_X1 U9903 ( .B1(n8295), .B2(n8294), .A(n8318), .ZN(n8296) );
  NAND2_X1 U9904 ( .A1(n8296), .A2(n10167), .ZN(n8308) );
  AOI21_X1 U9905 ( .B1(n8300), .B2(n8299), .A(n8328), .ZN(n8303) );
  INV_X1 U9906 ( .A(n8301), .ZN(n8302) );
  OAI21_X1 U9907 ( .B1(n10199), .B2(n8303), .A(n8302), .ZN(n8306) );
  NOR2_X1 U9908 ( .A1(n10183), .A2(n8304), .ZN(n8305) );
  AOI211_X1 U9909 ( .C1(n8327), .C2(n8393), .A(n8306), .B(n8305), .ZN(n8307)
         );
  OAI211_X1 U9910 ( .C1(n8309), .C2(n10191), .A(n8308), .B(n8307), .ZN(
        P2_U3195) );
  NOR2_X1 U9911 ( .A1(n8327), .A2(n8310), .ZN(n8312) );
  NAND2_X1 U9912 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8351), .ZN(n8313) );
  OAI21_X1 U9913 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8351), .A(n8313), .ZN(
        n8314) );
  NOR2_X1 U9914 ( .A1(n8315), .A2(n8314), .ZN(n8339) );
  AOI21_X1 U9915 ( .B1(n8315), .B2(n8314), .A(n8339), .ZN(n8338) );
  MUX2_X1 U9916 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8426), .Z(n8342) );
  XNOR2_X1 U9917 ( .A(n8342), .B(n8322), .ZN(n8321) );
  OR2_X1 U9918 ( .A1(n8317), .A2(n8316), .ZN(n8319) );
  NAND2_X1 U9919 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U9920 ( .A1(n8321), .A2(n8320), .ZN(n8343) );
  OAI21_X1 U9921 ( .B1(n8321), .B2(n8320), .A(n8343), .ZN(n8336) );
  NAND2_X1 U9922 ( .A1(n8393), .A2(n8322), .ZN(n8324) );
  OAI211_X1 U9923 ( .C1(n8325), .C2(n10183), .A(n8324), .B(n8323), .ZN(n8335)
         );
  NOR2_X1 U9924 ( .A1(n8327), .A2(n8326), .ZN(n8329) );
  NAND2_X1 U9925 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8351), .ZN(n8330) );
  OAI21_X1 U9926 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n8351), .A(n8330), .ZN(
        n8331) );
  NOR2_X1 U9927 ( .A1(n8332), .A2(n8331), .ZN(n8350) );
  AOI21_X1 U9928 ( .B1(n8332), .B2(n8331), .A(n8350), .ZN(n8333) );
  NOR2_X1 U9929 ( .A1(n8333), .A2(n10199), .ZN(n8334) );
  AOI211_X1 U9930 ( .C1(n10167), .C2(n8336), .A(n8335), .B(n8334), .ZN(n8337)
         );
  OAI21_X1 U9931 ( .B1(n8338), .B2(n10191), .A(n8337), .ZN(P2_U3196) );
  INV_X1 U9932 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8341) );
  AOI21_X1 U9933 ( .B1(n8341), .B2(n8340), .A(n8360), .ZN(n8358) );
  MUX2_X1 U9934 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8426), .Z(n8363) );
  XNOR2_X1 U9935 ( .A(n8363), .B(n8373), .ZN(n8346) );
  OR2_X1 U9936 ( .A1(n8342), .A2(n8351), .ZN(n8344) );
  NAND2_X1 U9937 ( .A1(n8344), .A2(n8343), .ZN(n8345) );
  NAND2_X1 U9938 ( .A1(n8346), .A2(n8345), .ZN(n8365) );
  OAI21_X1 U9939 ( .B1(n8346), .B2(n8345), .A(n8365), .ZN(n8356) );
  NAND2_X1 U9940 ( .A1(n8393), .A2(n8373), .ZN(n8348) );
  OAI211_X1 U9941 ( .C1(n8349), .C2(n10183), .A(n8348), .B(n8347), .ZN(n8355)
         );
  INV_X1 U9942 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8892) );
  AOI21_X1 U9943 ( .B1(n8352), .B2(n8892), .A(n8374), .ZN(n8353) );
  NOR2_X1 U9944 ( .A1(n8353), .A2(n10199), .ZN(n8354) );
  AOI211_X1 U9945 ( .C1(n10167), .C2(n8356), .A(n8355), .B(n8354), .ZN(n8357)
         );
  OAI21_X1 U9946 ( .B1(n8358), .B2(n10191), .A(n8357), .ZN(P2_U3197) );
  NOR2_X1 U9947 ( .A1(n8373), .A2(n8359), .ZN(n8361) );
  NAND2_X1 U9948 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8397), .ZN(n8384) );
  OAI21_X1 U9949 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8397), .A(n8384), .ZN(
        n8362) );
  AOI21_X1 U9950 ( .B1(n4457), .B2(n8362), .A(n8386), .ZN(n8383) );
  MUX2_X1 U9951 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8426), .Z(n8388) );
  XNOR2_X1 U9952 ( .A(n8388), .B(n8376), .ZN(n8368) );
  INV_X1 U9953 ( .A(n8363), .ZN(n8364) );
  NAND2_X1 U9954 ( .A1(n8373), .A2(n8364), .ZN(n8366) );
  NAND2_X1 U9955 ( .A1(n8366), .A2(n8365), .ZN(n8367) );
  NAND2_X1 U9956 ( .A1(n8368), .A2(n8367), .ZN(n8389) );
  OAI21_X1 U9957 ( .B1(n8368), .B2(n8367), .A(n8389), .ZN(n8381) );
  NAND2_X1 U9958 ( .A1(n8393), .A2(n8376), .ZN(n8370) );
  OAI211_X1 U9959 ( .C1(n8371), .C2(n10183), .A(n8370), .B(n8369), .ZN(n8380)
         );
  NOR2_X1 U9960 ( .A1(n8373), .A2(n8372), .ZN(n8375) );
  INV_X1 U9961 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8643) );
  AOI22_X1 U9962 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8376), .B1(n8397), .B2(
        n8643), .ZN(n8377) );
  AOI21_X1 U9963 ( .B1(n4454), .B2(n8377), .A(n8396), .ZN(n8378) );
  NOR2_X1 U9964 ( .A1(n8378), .A2(n10199), .ZN(n8379) );
  AOI211_X1 U9965 ( .C1(n10167), .C2(n8381), .A(n8380), .B(n8379), .ZN(n8382)
         );
  OAI21_X1 U9966 ( .B1(n8383), .B2(n10191), .A(n8382), .ZN(P2_U3198) );
  INV_X1 U9967 ( .A(n8384), .ZN(n8385) );
  OR2_X2 U9968 ( .A1(n8386), .A2(n8385), .ZN(n8412) );
  XNOR2_X2 U9969 ( .A(n8412), .B(n8424), .ZN(n8387) );
  AOI21_X1 U9970 ( .B1(n8580), .B2(n8387), .A(n8415), .ZN(n8404) );
  MUX2_X1 U9971 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8426), .Z(n8425) );
  XNOR2_X1 U9972 ( .A(n8425), .B(n8414), .ZN(n8392) );
  OR2_X1 U9973 ( .A1(n8388), .A2(n8397), .ZN(n8390) );
  NAND2_X1 U9974 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  NAND2_X1 U9975 ( .A1(n8392), .A2(n8391), .ZN(n8423) );
  OAI21_X1 U9976 ( .B1(n8392), .B2(n8391), .A(n8423), .ZN(n8402) );
  NAND2_X1 U9977 ( .A1(n8393), .A2(n8414), .ZN(n8395) );
  OAI211_X1 U9978 ( .C1(n9002), .C2(n10183), .A(n8395), .B(n8394), .ZN(n8401)
         );
  XNOR2_X1 U9979 ( .A(n8414), .B(n8405), .ZN(n8398) );
  INV_X1 U9980 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8857) );
  NOR2_X1 U9981 ( .A1(n8857), .A2(n8398), .ZN(n8406) );
  AOI21_X1 U9982 ( .B1(n8398), .B2(n8857), .A(n8406), .ZN(n8399) );
  NOR2_X1 U9983 ( .A1(n8399), .A2(n10199), .ZN(n8400) );
  AOI211_X1 U9984 ( .C1(n10167), .C2(n8402), .A(n8401), .B(n8400), .ZN(n8403)
         );
  OAI21_X1 U9985 ( .B1(n8404), .B2(n10191), .A(n8403), .ZN(P2_U3199) );
  INV_X1 U9986 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8918) );
  NOR2_X1 U9987 ( .A1(n8414), .A2(n8405), .ZN(n8407) );
  NOR2_X1 U9988 ( .A1(n8407), .A2(n8406), .ZN(n9878) );
  XNOR2_X1 U9989 ( .A(n8408), .B(n8918), .ZN(n9877) );
  OAI21_X1 U9990 ( .B1(n8408), .B2(n8918), .A(n9875), .ZN(n8411) );
  XNOR2_X1 U9991 ( .A(n8409), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8421) );
  INV_X1 U9992 ( .A(n8421), .ZN(n8410) );
  XNOR2_X1 U9993 ( .A(n8411), .B(n8410), .ZN(n8437) );
  NOR2_X1 U9994 ( .A1(n8414), .A2(n8413), .ZN(n8416) );
  NAND2_X1 U9995 ( .A1(n9888), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8417) );
  OAI21_X1 U9996 ( .B1(n9888), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8417), .ZN(
        n9879) );
  INV_X1 U9997 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8418) );
  MUX2_X1 U9998 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8418), .S(n8431), .Z(n8422)
         );
  XNOR2_X1 U9999 ( .A(n8420), .B(n8419), .ZN(n8435) );
  MUX2_X1 U10000 ( .A(n8422), .B(n8421), .S(n8426), .Z(n8430) );
  OAI21_X1 U10001 ( .B1(n8425), .B2(n8424), .A(n8423), .ZN(n8428) );
  INV_X1 U10002 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8569) );
  MUX2_X1 U10003 ( .A(n8569), .B(n8918), .S(n8426), .Z(n8427) );
  NAND2_X1 U10004 ( .A1(n8428), .A2(n8427), .ZN(n9887) );
  NOR2_X1 U10005 ( .A1(n10185), .A2(n8431), .ZN(n8432) );
  AOI211_X1 U10006 ( .C1(n10175), .C2(P2_ADDR_REG_19__SCAN_IN), .A(n8433), .B(
        n8432), .ZN(n8434) );
  OAI21_X1 U10007 ( .B1(n8437), .B2(n10199), .A(n8436), .ZN(P2_U3201) );
  NOR2_X1 U10008 ( .A1(n8439), .A2(n8438), .ZN(n8650) );
  NOR2_X1 U10009 ( .A1(n8440), .A2(n10217), .ZN(n8448) );
  AOI21_X1 U10010 ( .B1(n8650), .B2(n8601), .A(n8448), .ZN(n8443) );
  NAND2_X1 U10011 ( .A1(n10235), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8441) );
  OAI211_X1 U10012 ( .C1(n8652), .C2(n8516), .A(n8443), .B(n8441), .ZN(
        P2_U3202) );
  NAND2_X1 U10013 ( .A1(n10235), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8442) );
  OAI211_X1 U10014 ( .C1(n8655), .C2(n8516), .A(n8443), .B(n8442), .ZN(
        P2_U3203) );
  NAND2_X1 U10015 ( .A1(n8444), .A2(n8601), .ZN(n8450) );
  INV_X1 U10016 ( .A(n8445), .ZN(n8446) );
  NOR2_X1 U10017 ( .A1(n8446), .A2(n8516), .ZN(n8447) );
  AOI211_X1 U10018 ( .C1(n10235), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8448), .B(
        n8447), .ZN(n8449) );
  OAI211_X1 U10019 ( .C1(n8452), .C2(n8451), .A(n8450), .B(n8449), .ZN(
        P2_U3204) );
  INV_X1 U10020 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10021 ( .A(n8454), .B(n4438), .ZN(n8456) );
  AOI222_X1 U10022 ( .A1(n10207), .A2(n8456), .B1(n8455), .B2(n10202), .C1(
        n8475), .C2(n10204), .ZN(n8656) );
  MUX2_X1 U10023 ( .A(n8457), .B(n8656), .S(n8601), .Z(n8460) );
  AOI22_X1 U10024 ( .A1(n8658), .A2(n10210), .B1(n10211), .B2(n8458), .ZN(
        n8459) );
  OAI211_X1 U10025 ( .C1(n8661), .C2(n8605), .A(n8460), .B(n8459), .ZN(
        P2_U3206) );
  XNOR2_X1 U10026 ( .A(n8461), .B(n8464), .ZN(n8462) );
  OAI222_X1 U10027 ( .A1(n10221), .A2(n8463), .B1(n10220), .B2(n8486), .C1(
        n10225), .C2(n8462), .ZN(n8614) );
  INV_X1 U10028 ( .A(n8614), .ZN(n8470) );
  XNOR2_X1 U10029 ( .A(n8465), .B(n8464), .ZN(n8615) );
  AOI22_X1 U10030 ( .A1(n8466), .A2(n10211), .B1(n10235), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8467) );
  OAI21_X1 U10031 ( .B1(n8665), .B2(n8516), .A(n8467), .ZN(n8468) );
  AOI21_X1 U10032 ( .B1(n8615), .B2(n10213), .A(n8468), .ZN(n8469) );
  OAI21_X1 U10033 ( .B1(n8470), .B2(n10235), .A(n8469), .ZN(P2_U3207) );
  NOR2_X1 U10034 ( .A1(n8471), .A2(n10218), .ZN(n8478) );
  XNOR2_X1 U10035 ( .A(n8473), .B(n8472), .ZN(n8476) );
  AOI222_X1 U10036 ( .A1(n10207), .A2(n8476), .B1(n8475), .B2(n10202), .C1(
        n8474), .C2(n10204), .ZN(n8666) );
  INV_X1 U10037 ( .A(n8666), .ZN(n8477) );
  AOI211_X1 U10038 ( .C1(n10211), .C2(n8479), .A(n8478), .B(n8477), .ZN(n8483)
         );
  XNOR2_X1 U10039 ( .A(n8480), .B(n5528), .ZN(n8670) );
  INV_X1 U10040 ( .A(n8670), .ZN(n8481) );
  AOI22_X1 U10041 ( .A1(n8481), .A2(n10213), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10235), .ZN(n8482) );
  OAI21_X1 U10042 ( .B1(n8483), .B2(n10235), .A(n8482), .ZN(P2_U3208) );
  NOR2_X1 U10043 ( .A1(n8672), .A2(n10218), .ZN(n8487) );
  XOR2_X1 U10044 ( .A(n8491), .B(n8484), .Z(n8485) );
  OAI222_X1 U10045 ( .A1(n10221), .A2(n8486), .B1(n10220), .B2(n8511), .C1(
        n8485), .C2(n10225), .ZN(n8671) );
  AOI211_X1 U10046 ( .C1(n10211), .C2(n8488), .A(n8487), .B(n8671), .ZN(n8495)
         );
  NAND2_X1 U10047 ( .A1(n8490), .A2(n8489), .ZN(n8492) );
  XNOR2_X1 U10048 ( .A(n8492), .B(n8491), .ZN(n8673) );
  INV_X1 U10049 ( .A(n8673), .ZN(n8493) );
  AOI22_X1 U10050 ( .A1(n8493), .A2(n10213), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10235), .ZN(n8494) );
  OAI21_X1 U10051 ( .B1(n8495), .B2(n10235), .A(n8494), .ZN(P2_U3209) );
  XNOR2_X1 U10052 ( .A(n8496), .B(n8498), .ZN(n8678) );
  INV_X1 U10053 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8503) );
  XNOR2_X1 U10054 ( .A(n8497), .B(n8498), .ZN(n8499) );
  OAI222_X1 U10055 ( .A1(n10221), .A2(n8501), .B1(n10220), .B2(n8500), .C1(
        n10225), .C2(n8499), .ZN(n8676) );
  INV_X1 U10056 ( .A(n8676), .ZN(n8502) );
  MUX2_X1 U10057 ( .A(n8503), .B(n8502), .S(n8601), .Z(n8507) );
  AOI22_X1 U10058 ( .A1(n8505), .A2(n10210), .B1(n10211), .B2(n8504), .ZN(
        n8506) );
  OAI211_X1 U10059 ( .C1(n8678), .C2(n8605), .A(n8507), .B(n8506), .ZN(
        P2_U3210) );
  XOR2_X1 U10060 ( .A(n8508), .B(n8512), .Z(n8509) );
  OAI222_X1 U10061 ( .A1(n10221), .A2(n8511), .B1(n10220), .B2(n8510), .C1(
        n10225), .C2(n8509), .ZN(n8625) );
  INV_X1 U10062 ( .A(n8625), .ZN(n8519) );
  XOR2_X1 U10063 ( .A(n8513), .B(n8512), .Z(n8626) );
  AOI22_X1 U10064 ( .A1(n10235), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n10211), 
        .B2(n8514), .ZN(n8515) );
  OAI21_X1 U10065 ( .B1(n8684), .B2(n8516), .A(n8515), .ZN(n8517) );
  AOI21_X1 U10066 ( .B1(n8626), .B2(n10213), .A(n8517), .ZN(n8518) );
  OAI21_X1 U10067 ( .B1(n8519), .B2(n10235), .A(n8518), .ZN(P2_U3211) );
  NAND2_X1 U10068 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  XNOR2_X1 U10069 ( .A(n8522), .B(n8523), .ZN(n8690) );
  INV_X1 U10070 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8527) );
  XNOR2_X1 U10071 ( .A(n8524), .B(n8523), .ZN(n8526) );
  AOI222_X1 U10072 ( .A1(n10207), .A2(n8526), .B1(n8525), .B2(n10202), .C1(
        n8551), .C2(n10204), .ZN(n8685) );
  MUX2_X1 U10073 ( .A(n8527), .B(n8685), .S(n8601), .Z(n8530) );
  AOI22_X1 U10074 ( .A1(n8687), .A2(n10210), .B1(n10211), .B2(n8528), .ZN(
        n8529) );
  OAI211_X1 U10075 ( .C1(n8690), .C2(n8605), .A(n8530), .B(n8529), .ZN(
        P2_U3212) );
  XNOR2_X1 U10076 ( .A(n8531), .B(n8533), .ZN(n8693) );
  OAI21_X1 U10077 ( .B1(n8534), .B2(n8533), .A(n8532), .ZN(n8537) );
  AOI222_X1 U10078 ( .A1(n10207), .A2(n8537), .B1(n8536), .B2(n10202), .C1(
        n8535), .C2(n10204), .ZN(n8538) );
  INV_X1 U10079 ( .A(n8538), .ZN(n8631) );
  NAND2_X1 U10080 ( .A1(n8631), .A2(n8601), .ZN(n8544) );
  INV_X1 U10081 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8541) );
  INV_X1 U10082 ( .A(n8539), .ZN(n8540) );
  OAI22_X1 U10083 ( .A1(n8601), .A2(n8541), .B1(n8540), .B2(n10217), .ZN(n8542) );
  AOI21_X1 U10084 ( .B1(n8632), .B2(n10210), .A(n8542), .ZN(n8543) );
  OAI211_X1 U10085 ( .C1(n8693), .C2(n8605), .A(n8544), .B(n8543), .ZN(
        P2_U3213) );
  XNOR2_X1 U10086 ( .A(n8545), .B(n8546), .ZN(n8696) );
  NAND2_X1 U10087 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U10088 ( .A1(n8548), .A2(n10207), .ZN(n8549) );
  OR2_X1 U10089 ( .A1(n8550), .A2(n8549), .ZN(n8553) );
  AOI22_X1 U10090 ( .A1(n8551), .A2(n10202), .B1(n10204), .B2(n8578), .ZN(
        n8552) );
  NAND2_X1 U10091 ( .A1(n8553), .A2(n8552), .ZN(n8694) );
  MUX2_X1 U10092 ( .A(n8694), .B(P2_REG2_REG_19__SCAN_IN), .S(n10235), .Z(
        n8554) );
  INV_X1 U10093 ( .A(n8554), .ZN(n8558) );
  AOI22_X1 U10094 ( .A1(n8556), .A2(n10210), .B1(n10211), .B2(n8555), .ZN(
        n8557) );
  OAI211_X1 U10095 ( .C1(n8696), .C2(n8605), .A(n8558), .B(n8557), .ZN(
        P2_U3214) );
  NAND2_X1 U10096 ( .A1(n8559), .A2(n8563), .ZN(n8560) );
  INV_X1 U10097 ( .A(n8638), .ZN(n8574) );
  XNOR2_X1 U10098 ( .A(n8562), .B(n8563), .ZN(n8564) );
  OAI222_X1 U10099 ( .A1(n10221), .A2(n8566), .B1(n10220), .B2(n8565), .C1(
        n8564), .C2(n10225), .ZN(n8637) );
  NAND2_X1 U10100 ( .A1(n8637), .A2(n8601), .ZN(n8573) );
  INV_X1 U10101 ( .A(n8567), .ZN(n8568) );
  OAI22_X1 U10102 ( .A1(n8601), .A2(n8569), .B1(n8568), .B2(n10217), .ZN(n8570) );
  AOI21_X1 U10103 ( .B1(n8571), .B2(n10210), .A(n8570), .ZN(n8572) );
  OAI211_X1 U10104 ( .C1(n8574), .C2(n8605), .A(n8573), .B(n8572), .ZN(
        P2_U3215) );
  XNOR2_X1 U10105 ( .A(n8575), .B(n8576), .ZN(n8709) );
  INV_X1 U10106 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8580) );
  XNOR2_X1 U10107 ( .A(n8577), .B(n8576), .ZN(n8579) );
  AOI222_X1 U10108 ( .A1(n10207), .A2(n8579), .B1(n8578), .B2(n10202), .C1(
        n8599), .C2(n10204), .ZN(n8704) );
  MUX2_X1 U10109 ( .A(n8580), .B(n8704), .S(n8601), .Z(n8583) );
  AOI22_X1 U10110 ( .A1(n8706), .A2(n10210), .B1(n10211), .B2(n8581), .ZN(
        n8582) );
  OAI211_X1 U10111 ( .C1(n8709), .C2(n8605), .A(n8583), .B(n8582), .ZN(
        P2_U3216) );
  XNOR2_X1 U10112 ( .A(n8584), .B(n8585), .ZN(n8715) );
  INV_X1 U10113 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8590) );
  XOR2_X1 U10114 ( .A(n8586), .B(n8585), .Z(n8589) );
  AOI222_X1 U10115 ( .A1(n10207), .A2(n8589), .B1(n8588), .B2(n10202), .C1(
        n8587), .C2(n10204), .ZN(n8710) );
  MUX2_X1 U10116 ( .A(n8590), .B(n8710), .S(n8601), .Z(n8593) );
  AOI22_X1 U10117 ( .A1(n8712), .A2(n10210), .B1(n10211), .B2(n8591), .ZN(
        n8592) );
  OAI211_X1 U10118 ( .C1(n8715), .C2(n8605), .A(n8593), .B(n8592), .ZN(
        P2_U3217) );
  XNOR2_X1 U10119 ( .A(n8595), .B(n8596), .ZN(n8722) );
  XNOR2_X1 U10120 ( .A(n8597), .B(n8596), .ZN(n8600) );
  AOI222_X1 U10121 ( .A1(n10207), .A2(n8600), .B1(n8599), .B2(n10202), .C1(
        n8598), .C2(n10204), .ZN(n8716) );
  MUX2_X1 U10122 ( .A(n8341), .B(n8716), .S(n8601), .Z(n8604) );
  AOI22_X1 U10123 ( .A1(n8718), .A2(n10210), .B1(n10211), .B2(n8602), .ZN(
        n8603) );
  OAI211_X1 U10124 ( .C1(n8722), .C2(n8605), .A(n8604), .B(n8603), .ZN(
        P2_U3218) );
  INV_X1 U10125 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8608) );
  NAND2_X1 U10126 ( .A1(n8606), .A2(n8646), .ZN(n8607) );
  NAND2_X1 U10127 ( .A1(n8650), .A2(n10325), .ZN(n8609) );
  OAI211_X1 U10128 ( .C1(n10325), .C2(n8608), .A(n8607), .B(n8609), .ZN(
        P2_U3490) );
  NAND2_X1 U10129 ( .A1(n10323), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8610) );
  OAI211_X1 U10130 ( .C1(n8655), .C2(n8640), .A(n8610), .B(n8609), .ZN(
        P2_U3489) );
  INV_X1 U10131 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8611) );
  MUX2_X1 U10132 ( .A(n8611), .B(n8656), .S(n10325), .Z(n8613) );
  NAND2_X1 U10133 ( .A1(n8658), .A2(n8646), .ZN(n8612) );
  OAI211_X1 U10134 ( .C1(n8661), .C2(n8649), .A(n8613), .B(n8612), .ZN(
        P2_U3486) );
  INV_X1 U10135 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8616) );
  AOI21_X1 U10136 ( .B1(n8615), .B2(n10275), .A(n8614), .ZN(n8662) );
  OAI21_X1 U10137 ( .B1(n8665), .B2(n8640), .A(n8617), .ZN(P2_U3485) );
  INV_X1 U10138 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8618) );
  MUX2_X1 U10139 ( .A(n8618), .B(n8666), .S(n10325), .Z(n8620) );
  NAND2_X1 U10140 ( .A1(n8667), .A2(n8646), .ZN(n8619) );
  OAI211_X1 U10141 ( .C1(n8670), .C2(n8649), .A(n8620), .B(n8619), .ZN(
        P2_U3484) );
  MUX2_X1 U10142 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8671), .S(n10325), .Z(
        n8622) );
  OAI22_X1 U10143 ( .A1(n8673), .A2(n8649), .B1(n8672), .B2(n8640), .ZN(n8621)
         );
  OR2_X1 U10144 ( .A1(n8622), .A2(n8621), .ZN(P2_U3483) );
  MUX2_X1 U10145 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8676), .S(n10325), .Z(
        n8624) );
  OAI22_X1 U10146 ( .A1(n8678), .A2(n8649), .B1(n8677), .B2(n8640), .ZN(n8623)
         );
  OR2_X1 U10147 ( .A1(n8624), .A2(n8623), .ZN(P2_U3482) );
  INV_X1 U10148 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8627) );
  AOI21_X1 U10149 ( .B1(n10275), .B2(n8626), .A(n8625), .ZN(n8681) );
  MUX2_X1 U10150 ( .A(n8627), .B(n8681), .S(n10325), .Z(n8628) );
  OAI21_X1 U10151 ( .B1(n8684), .B2(n8640), .A(n8628), .ZN(P2_U3481) );
  INV_X1 U10152 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8966) );
  MUX2_X1 U10153 ( .A(n8966), .B(n8685), .S(n10325), .Z(n8630) );
  NAND2_X1 U10154 ( .A1(n8687), .A2(n8646), .ZN(n8629) );
  OAI211_X1 U10155 ( .C1(n8649), .C2(n8690), .A(n8630), .B(n8629), .ZN(
        P2_U3480) );
  INV_X1 U10156 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8633) );
  AOI21_X1 U10157 ( .B1(n10299), .B2(n8632), .A(n8631), .ZN(n8691) );
  MUX2_X1 U10158 ( .A(n8633), .B(n8691), .S(n10325), .Z(n8634) );
  OAI21_X1 U10159 ( .B1(n8649), .B2(n8693), .A(n8634), .ZN(P2_U3479) );
  MUX2_X1 U10160 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8694), .S(n10325), .Z(
        n8636) );
  OAI22_X1 U10161 ( .A1(n8696), .A2(n8649), .B1(n8695), .B2(n8640), .ZN(n8635)
         );
  OR2_X1 U10162 ( .A1(n8636), .A2(n8635), .ZN(P2_U3478) );
  AOI21_X1 U10163 ( .B1(n8638), .B2(n10275), .A(n8637), .ZN(n8699) );
  MUX2_X1 U10164 ( .A(n8918), .B(n8699), .S(n10325), .Z(n8639) );
  OAI21_X1 U10165 ( .B1(n8703), .B2(n8640), .A(n8639), .ZN(P2_U3477) );
  MUX2_X1 U10166 ( .A(n8857), .B(n8704), .S(n10325), .Z(n8642) );
  NAND2_X1 U10167 ( .A1(n8706), .A2(n8646), .ZN(n8641) );
  OAI211_X1 U10168 ( .C1(n8709), .C2(n8649), .A(n8642), .B(n8641), .ZN(
        P2_U3476) );
  MUX2_X1 U10169 ( .A(n8643), .B(n8710), .S(n10325), .Z(n8645) );
  NAND2_X1 U10170 ( .A1(n8712), .A2(n8646), .ZN(n8644) );
  OAI211_X1 U10171 ( .C1(n8715), .C2(n8649), .A(n8645), .B(n8644), .ZN(
        P2_U3475) );
  MUX2_X1 U10172 ( .A(n8892), .B(n8716), .S(n10325), .Z(n8648) );
  NAND2_X1 U10173 ( .A1(n8718), .A2(n8646), .ZN(n8647) );
  OAI211_X1 U10174 ( .C1(n8649), .C2(n8722), .A(n8648), .B(n8647), .ZN(
        P2_U3474) );
  NAND2_X1 U10175 ( .A1(n8650), .A2(n10300), .ZN(n8653) );
  NAND2_X1 U10176 ( .A1(n10302), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8651) );
  OAI211_X1 U10177 ( .C1(n8652), .C2(n8702), .A(n8653), .B(n8651), .ZN(
        P2_U3458) );
  NAND2_X1 U10178 ( .A1(n10302), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8654) );
  OAI211_X1 U10179 ( .C1(n8655), .C2(n8702), .A(n8654), .B(n8653), .ZN(
        P2_U3457) );
  MUX2_X1 U10180 ( .A(n8657), .B(n8656), .S(n10300), .Z(n8660) );
  NAND2_X1 U10181 ( .A1(n8658), .A2(n5662), .ZN(n8659) );
  OAI211_X1 U10182 ( .C1(n8661), .C2(n8721), .A(n8660), .B(n8659), .ZN(
        P2_U3454) );
  OAI21_X1 U10183 ( .B1(n8665), .B2(n8702), .A(n8664), .ZN(P2_U3453) );
  MUX2_X1 U10184 ( .A(n8803), .B(n8666), .S(n10300), .Z(n8669) );
  NAND2_X1 U10185 ( .A1(n8667), .A2(n5662), .ZN(n8668) );
  OAI211_X1 U10186 ( .C1(n8670), .C2(n8721), .A(n8669), .B(n8668), .ZN(
        P2_U3452) );
  MUX2_X1 U10187 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8671), .S(n10300), .Z(
        n8675) );
  OAI22_X1 U10188 ( .A1(n8673), .A2(n8721), .B1(n8672), .B2(n8702), .ZN(n8674)
         );
  OR2_X1 U10189 ( .A1(n8675), .A2(n8674), .ZN(P2_U3451) );
  MUX2_X1 U10190 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8676), .S(n10300), .Z(
        n8680) );
  OAI22_X1 U10191 ( .A1(n8678), .A2(n8721), .B1(n8677), .B2(n8702), .ZN(n8679)
         );
  OR2_X1 U10192 ( .A1(n8680), .A2(n8679), .ZN(P2_U3450) );
  MUX2_X1 U10193 ( .A(n8682), .B(n8681), .S(n10300), .Z(n8683) );
  OAI21_X1 U10194 ( .B1(n8684), .B2(n8702), .A(n8683), .ZN(P2_U3449) );
  INV_X1 U10195 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8686) );
  MUX2_X1 U10196 ( .A(n8686), .B(n8685), .S(n10300), .Z(n8689) );
  NAND2_X1 U10197 ( .A1(n8687), .A2(n5662), .ZN(n8688) );
  OAI211_X1 U10198 ( .C1(n8690), .C2(n8721), .A(n8689), .B(n8688), .ZN(
        P2_U3448) );
  INV_X1 U10199 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8815) );
  MUX2_X1 U10200 ( .A(n8815), .B(n8691), .S(n10300), .Z(n8692) );
  OAI21_X1 U10201 ( .B1(n8693), .B2(n8721), .A(n8692), .ZN(P2_U3447) );
  MUX2_X1 U10202 ( .A(n8694), .B(P2_REG0_REG_19__SCAN_IN), .S(n10302), .Z(
        n8698) );
  OAI22_X1 U10203 ( .A1(n8696), .A2(n8721), .B1(n8695), .B2(n8702), .ZN(n8697)
         );
  OR2_X1 U10204 ( .A1(n8698), .A2(n8697), .ZN(P2_U3446) );
  INV_X1 U10205 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8700) );
  MUX2_X1 U10206 ( .A(n8700), .B(n8699), .S(n10300), .Z(n8701) );
  OAI21_X1 U10207 ( .B1(n8703), .B2(n8702), .A(n8701), .ZN(P2_U3444) );
  INV_X1 U10208 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8705) );
  MUX2_X1 U10209 ( .A(n8705), .B(n8704), .S(n10300), .Z(n8708) );
  NAND2_X1 U10210 ( .A1(n8706), .A2(n5662), .ZN(n8707) );
  OAI211_X1 U10211 ( .C1(n8709), .C2(n8721), .A(n8708), .B(n8707), .ZN(
        P2_U3441) );
  INV_X1 U10212 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8711) );
  MUX2_X1 U10213 ( .A(n8711), .B(n8710), .S(n10300), .Z(n8714) );
  NAND2_X1 U10214 ( .A1(n8712), .A2(n5662), .ZN(n8713) );
  OAI211_X1 U10215 ( .C1(n8715), .C2(n8721), .A(n8714), .B(n8713), .ZN(
        P2_U3438) );
  INV_X1 U10216 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8717) );
  MUX2_X1 U10217 ( .A(n8717), .B(n8716), .S(n10300), .Z(n8720) );
  NAND2_X1 U10218 ( .A1(n8718), .A2(n5662), .ZN(n8719) );
  OAI211_X1 U10219 ( .C1(n8722), .C2(n8721), .A(n8720), .B(n8719), .ZN(
        P2_U3435) );
  INV_X1 U10220 ( .A(n8723), .ZN(n9864) );
  NOR4_X1 U10221 ( .A1(n8724), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8725), .A4(
        P2_U3151), .ZN(n8726) );
  AOI21_X1 U10222 ( .B1(n9020), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8726), .ZN(
        n8727) );
  OAI21_X1 U10223 ( .B1(n9864), .B2(n8733), .A(n8727), .ZN(P2_U3264) );
  INV_X1 U10224 ( .A(n8728), .ZN(n9866) );
  AOI22_X1 U10225 ( .A1(n8729), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9020), .ZN(n8730) );
  OAI21_X1 U10226 ( .B1(n9866), .B2(n8733), .A(n8730), .ZN(P2_U3265) );
  AOI22_X1 U10227 ( .A1(n8731), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9020), .ZN(n8732) );
  OAI21_X1 U10228 ( .B1(n9871), .B2(n8733), .A(n8732), .ZN(P2_U3266) );
  NAND4_X1 U10229 ( .A1(keyinput78), .A2(keyinput10), .A3(keyinput12), .A4(
        keyinput21), .ZN(n8734) );
  NOR3_X1 U10230 ( .A1(keyinput86), .A2(keyinput29), .A3(n8734), .ZN(n8735) );
  NAND3_X1 U10231 ( .A1(keyinput34), .A2(keyinput6), .A3(n8735), .ZN(n8748) );
  INV_X1 U10232 ( .A(keyinput11), .ZN(n8736) );
  NAND4_X1 U10233 ( .A1(keyinput96), .A2(keyinput112), .A3(keyinput22), .A4(
        n8736), .ZN(n8747) );
  NOR2_X1 U10234 ( .A1(keyinput115), .A2(keyinput108), .ZN(n8737) );
  NAND3_X1 U10235 ( .A1(keyinput100), .A2(keyinput126), .A3(n8737), .ZN(n8746)
         );
  INV_X1 U10236 ( .A(keyinput51), .ZN(n8738) );
  NOR4_X1 U10237 ( .A1(keyinput79), .A2(keyinput75), .A3(keyinput106), .A4(
        n8738), .ZN(n8744) );
  NOR4_X1 U10238 ( .A1(keyinput56), .A2(keyinput25), .A3(keyinput90), .A4(
        keyinput89), .ZN(n8743) );
  INV_X1 U10239 ( .A(keyinput76), .ZN(n8739) );
  NOR4_X1 U10240 ( .A1(keyinput70), .A2(keyinput16), .A3(keyinput60), .A4(
        n8739), .ZN(n8742) );
  NAND2_X1 U10241 ( .A1(keyinput45), .A2(keyinput105), .ZN(n8740) );
  NOR3_X1 U10242 ( .A1(keyinput42), .A2(keyinput27), .A3(n8740), .ZN(n8741) );
  NAND4_X1 U10243 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n8745)
         );
  NOR4_X1 U10244 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n8796)
         );
  NOR2_X1 U10245 ( .A1(keyinput57), .A2(keyinput24), .ZN(n8749) );
  NAND3_X1 U10246 ( .A1(keyinput124), .A2(keyinput54), .A3(n8749), .ZN(n8794)
         );
  NAND4_X1 U10247 ( .A1(keyinput123), .A2(keyinput47), .A3(keyinput73), .A4(
        keyinput37), .ZN(n8793) );
  INV_X1 U10248 ( .A(keyinput97), .ZN(n8751) );
  NAND4_X1 U10249 ( .A1(keyinput41), .A2(keyinput119), .A3(keyinput36), .A4(
        keyinput63), .ZN(n8750) );
  NOR4_X1 U10250 ( .A1(keyinput93), .A2(keyinput32), .A3(n8751), .A4(n8750), 
        .ZN(n8760) );
  NAND2_X1 U10251 ( .A1(keyinput26), .A2(keyinput8), .ZN(n8752) );
  NOR3_X1 U10252 ( .A1(keyinput67), .A2(keyinput48), .A3(n8752), .ZN(n8759) );
  NAND2_X1 U10253 ( .A1(keyinput33), .A2(keyinput71), .ZN(n8753) );
  NOR3_X1 U10254 ( .A1(keyinput87), .A2(keyinput53), .A3(n8753), .ZN(n8758) );
  NAND2_X1 U10255 ( .A1(keyinput66), .A2(keyinput84), .ZN(n8754) );
  NOR3_X1 U10256 ( .A1(keyinput2), .A2(keyinput82), .A3(n8754), .ZN(n8755) );
  NAND3_X1 U10257 ( .A1(keyinput80), .A2(keyinput31), .A3(n8755), .ZN(n8756)
         );
  NOR3_X1 U10258 ( .A1(keyinput88), .A2(keyinput17), .A3(n8756), .ZN(n8757) );
  NAND4_X1 U10259 ( .A1(n8760), .A2(n8759), .A3(n8758), .A4(n8757), .ZN(n8792)
         );
  NAND2_X1 U10260 ( .A1(keyinput117), .A2(keyinput114), .ZN(n8761) );
  NOR3_X1 U10261 ( .A1(keyinput81), .A2(keyinput72), .A3(n8761), .ZN(n8762) );
  NAND3_X1 U10262 ( .A1(keyinput116), .A2(keyinput18), .A3(n8762), .ZN(n8774)
         );
  NOR2_X1 U10263 ( .A1(keyinput111), .A2(keyinput30), .ZN(n8763) );
  NAND3_X1 U10264 ( .A1(keyinput38), .A2(keyinput58), .A3(n8763), .ZN(n8764)
         );
  NOR3_X1 U10265 ( .A1(keyinput59), .A2(keyinput118), .A3(n8764), .ZN(n8772)
         );
  NAND4_X1 U10266 ( .A1(keyinput46), .A2(keyinput110), .A3(keyinput40), .A4(
        keyinput15), .ZN(n8770) );
  NAND4_X1 U10267 ( .A1(keyinput39), .A2(keyinput44), .A3(keyinput4), .A4(
        keyinput50), .ZN(n8769) );
  INV_X1 U10268 ( .A(keyinput74), .ZN(n8765) );
  NAND4_X1 U10269 ( .A1(keyinput49), .A2(keyinput120), .A3(keyinput113), .A4(
        n8765), .ZN(n8768) );
  NOR3_X1 U10270 ( .A1(keyinput43), .A2(keyinput7), .A3(keyinput85), .ZN(n8766) );
  NAND2_X1 U10271 ( .A1(keyinput35), .A2(n8766), .ZN(n8767) );
  NOR4_X1 U10272 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8771)
         );
  NAND4_X1 U10273 ( .A1(keyinput14), .A2(keyinput62), .A3(n8772), .A4(n8771), 
        .ZN(n8773) );
  NOR4_X1 U10274 ( .A1(keyinput9), .A2(keyinput94), .A3(n8774), .A4(n8773), 
        .ZN(n8790) );
  AND4_X1 U10275 ( .A1(keyinput122), .A2(keyinput55), .A3(keyinput64), .A4(
        keyinput0), .ZN(n8789) );
  INV_X1 U10276 ( .A(keyinput83), .ZN(n8775) );
  NOR4_X1 U10277 ( .A1(keyinput13), .A2(keyinput3), .A3(keyinput52), .A4(n8775), .ZN(n8788) );
  NAND2_X1 U10278 ( .A1(keyinput95), .A2(keyinput19), .ZN(n8776) );
  NOR3_X1 U10279 ( .A1(keyinput99), .A2(keyinput127), .A3(n8776), .ZN(n8777)
         );
  NAND3_X1 U10280 ( .A1(keyinput103), .A2(keyinput92), .A3(n8777), .ZN(n8786)
         );
  NAND3_X1 U10281 ( .A1(keyinput104), .A2(keyinput20), .A3(keyinput69), .ZN(
        n8778) );
  NOR2_X1 U10282 ( .A1(keyinput91), .A2(n8778), .ZN(n8784) );
  INV_X1 U10283 ( .A(keyinput102), .ZN(n8779) );
  NOR4_X1 U10284 ( .A1(keyinput125), .A2(keyinput5), .A3(keyinput23), .A4(
        n8779), .ZN(n8783) );
  NOR4_X1 U10285 ( .A1(keyinput107), .A2(keyinput77), .A3(keyinput98), .A4(
        keyinput61), .ZN(n8782) );
  NAND3_X1 U10286 ( .A1(keyinput1), .A2(keyinput121), .A3(keyinput101), .ZN(
        n8780) );
  NOR2_X1 U10287 ( .A1(keyinput28), .A2(n8780), .ZN(n8781) );
  NAND4_X1 U10288 ( .A1(n8784), .A2(n8783), .A3(n8782), .A4(n8781), .ZN(n8785)
         );
  NOR4_X1 U10289 ( .A1(keyinput109), .A2(keyinput65), .A3(n8786), .A4(n8785), 
        .ZN(n8787) );
  NAND4_X1 U10290 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n8791)
         );
  NOR4_X1 U10291 ( .A1(n8794), .A2(n8793), .A3(n8792), .A4(n8791), .ZN(n8795)
         );
  AOI21_X1 U10292 ( .B1(n8796), .B2(n8795), .A(keyinput68), .ZN(n9019) );
  AOI22_X1 U10293 ( .A1(n10328), .A2(keyinput44), .B1(n8798), .B2(keyinput4), 
        .ZN(n8797) );
  OAI221_X1 U10294 ( .B1(n10328), .B2(keyinput44), .C1(n8798), .C2(keyinput4), 
        .A(n8797), .ZN(n8808) );
  AOI22_X1 U10295 ( .A1(n9835), .A2(keyinput50), .B1(n8800), .B2(keyinput46), 
        .ZN(n8799) );
  OAI221_X1 U10296 ( .B1(n9835), .B2(keyinput50), .C1(n8800), .C2(keyinput46), 
        .A(n8799), .ZN(n8807) );
  INV_X1 U10297 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8802) );
  AOI22_X1 U10298 ( .A1(n8803), .A2(keyinput110), .B1(keyinput40), .B2(n8802), 
        .ZN(n8801) );
  OAI221_X1 U10299 ( .B1(n8803), .B2(keyinput110), .C1(n8802), .C2(keyinput40), 
        .A(n8801), .ZN(n8806) );
  AOI22_X1 U10300 ( .A1(n9791), .A2(keyinput15), .B1(n10215), .B2(keyinput116), 
        .ZN(n8804) );
  OAI221_X1 U10301 ( .B1(n9791), .B2(keyinput15), .C1(n10215), .C2(keyinput116), .A(n8804), .ZN(n8805) );
  NOR4_X1 U10302 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n8850)
         );
  INV_X1 U10303 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10075) );
  AOI22_X1 U10304 ( .A1(n10075), .A2(keyinput72), .B1(keyinput59), .B2(n8810), 
        .ZN(n8809) );
  OAI221_X1 U10305 ( .B1(n10075), .B2(keyinput72), .C1(n8810), .C2(keyinput59), 
        .A(n8809), .ZN(n8821) );
  INV_X1 U10306 ( .A(P2_B_REG_SCAN_IN), .ZN(n8812) );
  AOI22_X1 U10307 ( .A1(n5208), .A2(keyinput81), .B1(keyinput117), .B2(n8812), 
        .ZN(n8811) );
  OAI221_X1 U10308 ( .B1(n5208), .B2(keyinput81), .C1(n8812), .C2(keyinput117), 
        .A(n8811), .ZN(n8820) );
  AOI22_X1 U10309 ( .A1(n8815), .A2(keyinput18), .B1(n8814), .B2(keyinput9), 
        .ZN(n8813) );
  OAI221_X1 U10310 ( .B1(n8815), .B2(keyinput18), .C1(n8814), .C2(keyinput9), 
        .A(n8813), .ZN(n8819) );
  XOR2_X1 U10311 ( .A(n6447), .B(keyinput94), .Z(n8817) );
  XNOR2_X1 U10312 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput114), .ZN(n8816) );
  NAND2_X1 U10313 ( .A1(n8817), .A2(n8816), .ZN(n8818) );
  NOR4_X1 U10314 ( .A1(n8821), .A2(n8820), .A3(n8819), .A4(n8818), .ZN(n8849)
         );
  INV_X1 U10315 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8823) );
  INV_X1 U10316 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U10317 ( .A1(n8823), .A2(keyinput118), .B1(keyinput111), .B2(n10247), .ZN(n8822) );
  OAI221_X1 U10318 ( .B1(n8823), .B2(keyinput118), .C1(n10247), .C2(
        keyinput111), .A(n8822), .ZN(n8835) );
  AOI22_X1 U10319 ( .A1(n8826), .A2(keyinput38), .B1(keyinput58), .B2(n8825), 
        .ZN(n8824) );
  OAI221_X1 U10320 ( .B1(n8826), .B2(keyinput38), .C1(n8825), .C2(keyinput58), 
        .A(n8824), .ZN(n8834) );
  AOI22_X1 U10321 ( .A1(n8829), .A2(keyinput30), .B1(keyinput14), .B2(n8828), 
        .ZN(n8827) );
  OAI221_X1 U10322 ( .B1(n8829), .B2(keyinput30), .C1(n8828), .C2(keyinput14), 
        .A(n8827), .ZN(n8833) );
  INV_X1 U10323 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U10324 ( .A1(n10099), .A2(keyinput62), .B1(keyinput43), .B2(n8831), 
        .ZN(n8830) );
  OAI221_X1 U10325 ( .B1(n10099), .B2(keyinput62), .C1(n8831), .C2(keyinput43), 
        .A(n8830), .ZN(n8832) );
  NOR4_X1 U10326 ( .A1(n8835), .A2(n8834), .A3(n8833), .A4(n8832), .ZN(n8848)
         );
  INV_X1 U10327 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n8837) );
  AOI22_X1 U10328 ( .A1(n8837), .A2(keyinput113), .B1(n7550), .B2(keyinput99), 
        .ZN(n8836) );
  OAI221_X1 U10329 ( .B1(n8837), .B2(keyinput113), .C1(n7550), .C2(keyinput99), 
        .A(n8836), .ZN(n8846) );
  AOI22_X1 U10330 ( .A1(n5588), .A2(keyinput7), .B1(n6000), .B2(keyinput49), 
        .ZN(n8838) );
  OAI221_X1 U10331 ( .B1(n5588), .B2(keyinput7), .C1(n6000), .C2(keyinput49), 
        .A(n8838), .ZN(n8845) );
  AOI22_X1 U10332 ( .A1(n8840), .A2(keyinput85), .B1(keyinput35), .B2(n9356), 
        .ZN(n8839) );
  OAI221_X1 U10333 ( .B1(n8840), .B2(keyinput85), .C1(n9356), .C2(keyinput35), 
        .A(n8839), .ZN(n8844) );
  XOR2_X1 U10334 ( .A(n5627), .B(keyinput120), .Z(n8842) );
  XNOR2_X1 U10335 ( .A(P2_IR_REG_18__SCAN_IN), .B(keyinput74), .ZN(n8841) );
  NAND2_X1 U10336 ( .A1(n8842), .A2(n8841), .ZN(n8843) );
  NOR4_X1 U10337 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n8847)
         );
  NAND4_X1 U10338 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n9017)
         );
  AOI22_X1 U10339 ( .A1(n6333), .A2(keyinput65), .B1(keyinput125), .B2(n10212), 
        .ZN(n8851) );
  OAI221_X1 U10340 ( .B1(n6333), .B2(keyinput65), .C1(n10212), .C2(keyinput125), .A(n8851), .ZN(n8863) );
  AOI22_X1 U10341 ( .A1(n8854), .A2(keyinput19), .B1(keyinput103), .B2(n8853), 
        .ZN(n8852) );
  OAI221_X1 U10342 ( .B1(n8854), .B2(keyinput19), .C1(n8853), .C2(keyinput103), 
        .A(n8852), .ZN(n8862) );
  INV_X1 U10343 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8856) );
  AOI22_X1 U10344 ( .A1(n8857), .A2(keyinput92), .B1(n8856), .B2(keyinput95), 
        .ZN(n8855) );
  OAI221_X1 U10345 ( .B1(n8857), .B2(keyinput92), .C1(n8856), .C2(keyinput95), 
        .A(n8855), .ZN(n8861) );
  XOR2_X1 U10346 ( .A(n7094), .B(keyinput109), .Z(n8859) );
  XNOR2_X1 U10347 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput127), .ZN(n8858)
         );
  NAND2_X1 U10348 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  NOR4_X1 U10349 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n8905)
         );
  AOI22_X1 U10350 ( .A1(n8866), .A2(keyinput91), .B1(n8865), .B2(keyinput13), 
        .ZN(n8864) );
  OAI221_X1 U10351 ( .B1(n8866), .B2(keyinput91), .C1(n8865), .C2(keyinput13), 
        .A(n8864), .ZN(n8877) );
  INV_X1 U10352 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9942) );
  INV_X1 U10353 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8868) );
  AOI22_X1 U10354 ( .A1(n9942), .A2(keyinput69), .B1(n8868), .B2(keyinput104), 
        .ZN(n8867) );
  OAI221_X1 U10355 ( .B1(n9942), .B2(keyinput69), .C1(n8868), .C2(keyinput104), 
        .A(n8867), .ZN(n8876) );
  AOI22_X1 U10356 ( .A1(n8871), .A2(keyinput5), .B1(keyinput23), .B2(n8870), 
        .ZN(n8869) );
  OAI221_X1 U10357 ( .B1(n8871), .B2(keyinput5), .C1(n8870), .C2(keyinput23), 
        .A(n8869), .ZN(n8875) );
  XNOR2_X1 U10358 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput102), .ZN(n8873) );
  XNOR2_X1 U10359 ( .A(SI_30_), .B(keyinput20), .ZN(n8872) );
  NAND2_X1 U10360 ( .A1(n8873), .A2(n8872), .ZN(n8874) );
  NOR4_X1 U10361 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8904)
         );
  AOI22_X1 U10362 ( .A1(n5155), .A2(keyinput0), .B1(keyinput121), .B2(n10311), 
        .ZN(n8878) );
  OAI221_X1 U10363 ( .B1(n5155), .B2(keyinput0), .C1(n10311), .C2(keyinput121), 
        .A(n8878), .ZN(n8889) );
  AOI22_X1 U10364 ( .A1(n8880), .A2(keyinput55), .B1(keyinput64), .B2(n8580), 
        .ZN(n8879) );
  OAI221_X1 U10365 ( .B1(n8880), .B2(keyinput55), .C1(n8580), .C2(keyinput64), 
        .A(n8879), .ZN(n8888) );
  AOI22_X1 U10366 ( .A1(n8883), .A2(keyinput83), .B1(keyinput3), .B2(n8882), 
        .ZN(n8881) );
  OAI221_X1 U10367 ( .B1(n8883), .B2(keyinput83), .C1(n8882), .C2(keyinput3), 
        .A(n8881), .ZN(n8887) );
  XNOR2_X1 U10368 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput52), .ZN(n8885) );
  XNOR2_X1 U10369 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput122), .ZN(n8884)
         );
  NAND2_X1 U10370 ( .A1(n8885), .A2(n8884), .ZN(n8886) );
  NOR4_X1 U10371 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n8903)
         );
  AOI22_X1 U10372 ( .A1(n8892), .A2(keyinput101), .B1(n8891), .B2(keyinput107), 
        .ZN(n8890) );
  OAI221_X1 U10373 ( .B1(n8892), .B2(keyinput101), .C1(n8891), .C2(keyinput107), .A(n8890), .ZN(n8901) );
  INV_X1 U10374 ( .A(SI_7_), .ZN(n8895) );
  INV_X1 U10375 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8894) );
  AOI22_X1 U10376 ( .A1(n8895), .A2(keyinput77), .B1(keyinput1), .B2(n8894), 
        .ZN(n8893) );
  OAI221_X1 U10377 ( .B1(n8895), .B2(keyinput77), .C1(n8894), .C2(keyinput1), 
        .A(n8893), .ZN(n8900) );
  INV_X1 U10378 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10071) );
  AOI22_X1 U10379 ( .A1(n10071), .A2(keyinput28), .B1(keyinput98), .B2(n6712), 
        .ZN(n8896) );
  OAI221_X1 U10380 ( .B1(n10071), .B2(keyinput28), .C1(n6712), .C2(keyinput98), 
        .A(n8896), .ZN(n8899) );
  INV_X1 U10381 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10281) );
  AOI22_X1 U10382 ( .A1(n6563), .A2(keyinput93), .B1(keyinput61), .B2(n10281), 
        .ZN(n8897) );
  OAI221_X1 U10383 ( .B1(n6563), .B2(keyinput93), .C1(n10281), .C2(keyinput61), 
        .A(n8897), .ZN(n8898) );
  NOR4_X1 U10384 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n8902)
         );
  NAND4_X1 U10385 ( .A1(n8905), .A2(n8904), .A3(n8903), .A4(n8902), .ZN(n9016)
         );
  INV_X1 U10386 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10072) );
  AOI22_X1 U10387 ( .A1(n10072), .A2(keyinput60), .B1(keyinput34), .B2(n6613), 
        .ZN(n8906) );
  OAI221_X1 U10388 ( .B1(n10072), .B2(keyinput60), .C1(n6613), .C2(keyinput34), 
        .A(n8906), .ZN(n8916) );
  INV_X1 U10389 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10069) );
  AOI22_X1 U10390 ( .A1(n10069), .A2(keyinput27), .B1(keyinput76), .B2(n6713), 
        .ZN(n8907) );
  OAI221_X1 U10391 ( .B1(n10069), .B2(keyinput27), .C1(n6713), .C2(keyinput76), 
        .A(n8907), .ZN(n8915) );
  INV_X1 U10392 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8909) );
  AOI22_X1 U10393 ( .A1(n8910), .A2(keyinput42), .B1(keyinput45), .B2(n8909), 
        .ZN(n8908) );
  OAI221_X1 U10394 ( .B1(n8910), .B2(keyinput42), .C1(n8909), .C2(keyinput45), 
        .A(n8908), .ZN(n8914) );
  XNOR2_X1 U10395 ( .A(P2_REG2_REG_25__SCAN_IN), .B(keyinput16), .ZN(n8912) );
  XNOR2_X1 U10396 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput70), .ZN(n8911) );
  NAND2_X1 U10397 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  NOR4_X1 U10398 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n8960)
         );
  AOI22_X1 U10399 ( .A1(n8918), .A2(keyinput51), .B1(n6399), .B2(keyinput75), 
        .ZN(n8917) );
  OAI221_X1 U10400 ( .B1(n8918), .B2(keyinput51), .C1(n6399), .C2(keyinput75), 
        .A(n8917), .ZN(n8928) );
  AOI22_X1 U10401 ( .A1(n10070), .A2(keyinput106), .B1(keyinput105), .B2(n8920), .ZN(n8919) );
  OAI221_X1 U10402 ( .B1(n10070), .B2(keyinput106), .C1(n8920), .C2(
        keyinput105), .A(n8919), .ZN(n8927) );
  AOI22_X1 U10403 ( .A1(n10076), .A2(keyinput89), .B1(keyinput79), .B2(n8922), 
        .ZN(n8921) );
  OAI221_X1 U10404 ( .B1(n10076), .B2(keyinput89), .C1(n8922), .C2(keyinput79), 
        .A(n8921), .ZN(n8926) );
  XNOR2_X1 U10405 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput90), .ZN(n8924) );
  XNOR2_X1 U10406 ( .A(SI_28_), .B(keyinput25), .ZN(n8923) );
  NAND2_X1 U10407 ( .A1(n8924), .A2(n8923), .ZN(n8925) );
  NOR4_X1 U10408 ( .A1(n8928), .A2(n8927), .A3(n8926), .A4(n8925), .ZN(n8959)
         );
  INV_X1 U10409 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8930) );
  AOI22_X1 U10410 ( .A1(n9299), .A2(keyinput108), .B1(keyinput11), .B2(n8930), 
        .ZN(n8929) );
  OAI221_X1 U10411 ( .B1(n9299), .B2(keyinput108), .C1(n8930), .C2(keyinput11), 
        .A(n8929), .ZN(n8941) );
  AOI22_X1 U10412 ( .A1(n8932), .A2(keyinput115), .B1(keyinput126), .B2(n9799), 
        .ZN(n8931) );
  OAI221_X1 U10413 ( .B1(n8932), .B2(keyinput115), .C1(n9799), .C2(keyinput126), .A(n8931), .ZN(n8940) );
  AOI22_X1 U10414 ( .A1(n8935), .A2(keyinput22), .B1(keyinput39), .B2(n8934), 
        .ZN(n8933) );
  OAI221_X1 U10415 ( .B1(n8935), .B2(keyinput22), .C1(n8934), .C2(keyinput39), 
        .A(n8933), .ZN(n8939) );
  AOI22_X1 U10416 ( .A1(n8937), .A2(keyinput96), .B1(keyinput112), .B2(n10023), 
        .ZN(n8936) );
  OAI221_X1 U10417 ( .B1(n8937), .B2(keyinput96), .C1(n10023), .C2(keyinput112), .A(n8936), .ZN(n8938) );
  NOR4_X1 U10418 ( .A1(n8941), .A2(n8940), .A3(n8939), .A4(n8938), .ZN(n8958)
         );
  AOI22_X1 U10419 ( .A1(n8944), .A2(keyinput21), .B1(keyinput86), .B2(n8943), 
        .ZN(n8942) );
  OAI221_X1 U10420 ( .B1(n8944), .B2(keyinput21), .C1(n8943), .C2(keyinput86), 
        .A(n8942), .ZN(n8950) );
  AOI22_X1 U10421 ( .A1(n8947), .A2(keyinput6), .B1(n8946), .B2(keyinput78), 
        .ZN(n8945) );
  OAI221_X1 U10422 ( .B1(n8947), .B2(keyinput6), .C1(n8946), .C2(keyinput78), 
        .A(n8945), .ZN(n8949) );
  XOR2_X1 U10423 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput29), .Z(n8948) );
  OR3_X1 U10424 ( .A1(n8950), .A2(n8949), .A3(n8948), .ZN(n8956) );
  AOI22_X1 U10425 ( .A1(n8953), .A2(keyinput10), .B1(keyinput12), .B2(n8952), 
        .ZN(n8951) );
  OAI221_X1 U10426 ( .B1(n8953), .B2(keyinput10), .C1(n8952), .C2(keyinput12), 
        .A(n8951), .ZN(n8955) );
  INV_X1 U10427 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10040) );
  XNOR2_X1 U10428 ( .A(n10040), .B(keyinput100), .ZN(n8954) );
  NOR3_X1 U10429 ( .A1(n8956), .A2(n8955), .A3(n8954), .ZN(n8957) );
  NAND4_X1 U10430 ( .A1(n8960), .A2(n8959), .A3(n8958), .A4(n8957), .ZN(n9015)
         );
  INV_X1 U10431 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8962) );
  AOI22_X1 U10432 ( .A1(n5750), .A2(keyinput57), .B1(keyinput73), .B2(n8962), 
        .ZN(n8961) );
  OAI221_X1 U10433 ( .B1(n5750), .B2(keyinput57), .C1(n8962), .C2(keyinput73), 
        .A(n8961), .ZN(n8973) );
  AOI22_X1 U10434 ( .A1(n8964), .A2(keyinput24), .B1(n6204), .B2(keyinput87), 
        .ZN(n8963) );
  OAI221_X1 U10435 ( .B1(n8964), .B2(keyinput24), .C1(n6204), .C2(keyinput87), 
        .A(n8963), .ZN(n8972) );
  AOI22_X1 U10436 ( .A1(n8967), .A2(keyinput47), .B1(keyinput124), .B2(n8966), 
        .ZN(n8965) );
  OAI221_X1 U10437 ( .B1(n8967), .B2(keyinput47), .C1(n8966), .C2(keyinput124), 
        .A(n8965), .ZN(n8971) );
  XOR2_X1 U10438 ( .A(n9546), .B(keyinput54), .Z(n8969) );
  XNOR2_X1 U10439 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput37), .ZN(n8968) );
  NAND2_X1 U10440 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  NOR4_X1 U10441 ( .A1(n8973), .A2(n8972), .A3(n8971), .A4(n8970), .ZN(n9013)
         );
  NAND2_X1 U10442 ( .A1(n9850), .A2(keyinput97), .ZN(n8974) );
  OAI221_X1 U10443 ( .B1(n9595), .B2(keyinput68), .C1(n9850), .C2(keyinput97), 
        .A(n8974), .ZN(n8985) );
  INV_X1 U10444 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8976) );
  AOI22_X1 U10445 ( .A1(n8977), .A2(keyinput41), .B1(n8976), .B2(keyinput119), 
        .ZN(n8975) );
  OAI221_X1 U10446 ( .B1(n8977), .B2(keyinput41), .C1(n8976), .C2(keyinput119), 
        .A(n8975), .ZN(n8984) );
  AOI22_X1 U10447 ( .A1(n7619), .A2(keyinput63), .B1(n5685), .B2(keyinput123), 
        .ZN(n8978) );
  OAI221_X1 U10448 ( .B1(n7619), .B2(keyinput63), .C1(n5685), .C2(keyinput123), 
        .A(n8978), .ZN(n8983) );
  AOI22_X1 U10449 ( .A1(n8981), .A2(keyinput32), .B1(keyinput36), .B2(n8980), 
        .ZN(n8979) );
  OAI221_X1 U10450 ( .B1(n8981), .B2(keyinput32), .C1(n8980), .C2(keyinput36), 
        .A(n8979), .ZN(n8982) );
  NOR4_X1 U10451 ( .A1(n8985), .A2(n8984), .A3(n8983), .A4(n8982), .ZN(n9012)
         );
  AOI22_X1 U10452 ( .A1(n7266), .A2(keyinput82), .B1(keyinput88), .B2(n5785), 
        .ZN(n8986) );
  OAI221_X1 U10453 ( .B1(n7266), .B2(keyinput82), .C1(n5785), .C2(keyinput88), 
        .A(n8986), .ZN(n8997) );
  INV_X1 U10454 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U10455 ( .A1(n9467), .A2(keyinput84), .B1(n8988), .B2(keyinput66), 
        .ZN(n8987) );
  OAI221_X1 U10456 ( .B1(n9467), .B2(keyinput84), .C1(n8988), .C2(keyinput66), 
        .A(n8987), .ZN(n8996) );
  AOI22_X1 U10457 ( .A1(n6065), .A2(keyinput31), .B1(n8990), .B2(keyinput56), 
        .ZN(n8989) );
  OAI221_X1 U10458 ( .B1(n6065), .B2(keyinput31), .C1(n8990), .C2(keyinput56), 
        .A(n8989), .ZN(n8995) );
  AOI22_X1 U10459 ( .A1(n8993), .A2(keyinput17), .B1(n8992), .B2(keyinput80), 
        .ZN(n8991) );
  OAI221_X1 U10460 ( .B1(n8993), .B2(keyinput17), .C1(n8992), .C2(keyinput80), 
        .A(n8991), .ZN(n8994) );
  NOR4_X1 U10461 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n8994), .ZN(n9011)
         );
  AOI22_X1 U10462 ( .A1(n6266), .A2(keyinput53), .B1(keyinput67), .B2(n8999), 
        .ZN(n8998) );
  OAI221_X1 U10463 ( .B1(n6266), .B2(keyinput53), .C1(n8999), .C2(keyinput67), 
        .A(n8998), .ZN(n9009) );
  AOI22_X1 U10464 ( .A1(n10074), .A2(keyinput71), .B1(keyinput33), .B2(n10073), 
        .ZN(n9000) );
  OAI221_X1 U10465 ( .B1(n10074), .B2(keyinput71), .C1(n10073), .C2(keyinput33), .A(n9000), .ZN(n9008) );
  INV_X1 U10466 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U10467 ( .A1(n9941), .A2(keyinput48), .B1(keyinput2), .B2(n9002), 
        .ZN(n9001) );
  OAI221_X1 U10468 ( .B1(n9941), .B2(keyinput48), .C1(n9002), .C2(keyinput2), 
        .A(n9001), .ZN(n9007) );
  INV_X1 U10469 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9005) );
  INV_X1 U10470 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9004) );
  AOI22_X1 U10471 ( .A1(n9005), .A2(keyinput8), .B1(n9004), .B2(keyinput26), 
        .ZN(n9003) );
  OAI221_X1 U10472 ( .B1(n9005), .B2(keyinput8), .C1(n9004), .C2(keyinput26), 
        .A(n9003), .ZN(n9006) );
  NOR4_X1 U10473 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n9010)
         );
  NAND4_X1 U10474 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n9014)
         );
  NOR4_X1 U10475 ( .A1(n9017), .A2(n9016), .A3(n9015), .A4(n9014), .ZN(n9018)
         );
  OAI21_X1 U10476 ( .B1(P1_REG2_REG_22__SCAN_IN), .B2(n9019), .A(n9018), .ZN(
        n9025) );
  AOI222_X1 U10477 ( .A1(n9023), .A2(n9022), .B1(n9021), .B2(
        P2_STATE_REG_SCAN_IN), .C1(P1_DATAO_REG_9__SCAN_IN), .C2(n9020), .ZN(
        n9024) );
  XOR2_X1 U10478 ( .A(n9025), .B(n9024), .Z(P2_U3286) );
  MUX2_X1 U10479 ( .A(n9026), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI22_X1 U10480 ( .A1(n9034), .A2(n4514), .B1(n9137), .B2(n9389), .ZN(n9032)
         );
  XOR2_X1 U10481 ( .A(n9140), .B(n9032), .Z(n9033) );
  AOI22_X1 U10482 ( .A1(n9034), .A2(n9082), .B1(n9081), .B2(n9389), .ZN(n9922)
         );
  NAND2_X1 U10483 ( .A1(n9920), .A2(n4915), .ZN(n9324) );
  NAND2_X1 U10484 ( .A1(n9333), .A2(n4514), .ZN(n9036) );
  OR2_X1 U10485 ( .A1(n9038), .A2(n9207), .ZN(n9035) );
  NAND2_X1 U10486 ( .A1(n9036), .A2(n9035), .ZN(n9037) );
  XNOR2_X1 U10487 ( .A(n9037), .B(n9204), .ZN(n9041) );
  NOR2_X1 U10488 ( .A1(n9038), .A2(n9201), .ZN(n9039) );
  AOI21_X1 U10489 ( .B1(n9333), .B2(n9137), .A(n9039), .ZN(n9040) );
  OR2_X1 U10490 ( .A1(n9041), .A2(n9040), .ZN(n9325) );
  NAND2_X1 U10491 ( .A1(n9324), .A2(n9325), .ZN(n9323) );
  NAND2_X1 U10492 ( .A1(n9041), .A2(n9040), .ZN(n9327) );
  NAND2_X1 U10493 ( .A1(n9241), .A2(n4514), .ZN(n9044) );
  OR2_X1 U10494 ( .A1(n9042), .A2(n9207), .ZN(n9043) );
  NAND2_X1 U10495 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  XNOR2_X1 U10496 ( .A(n9045), .B(n9140), .ZN(n9048) );
  AOI22_X1 U10497 ( .A1(n9241), .A2(n9082), .B1(n9081), .B2(n9387), .ZN(n9046)
         );
  XNOR2_X1 U10498 ( .A(n9048), .B(n9046), .ZN(n9235) );
  INV_X1 U10499 ( .A(n9046), .ZN(n9047) );
  NAND2_X1 U10500 ( .A1(n9309), .A2(n4514), .ZN(n9052) );
  OR2_X1 U10501 ( .A1(n9050), .A2(n9207), .ZN(n9051) );
  NAND2_X1 U10502 ( .A1(n9052), .A2(n9051), .ZN(n9053) );
  XNOR2_X1 U10503 ( .A(n9053), .B(n9140), .ZN(n9054) );
  AOI22_X1 U10504 ( .A1(n9309), .A2(n9082), .B1(n9081), .B2(n9386), .ZN(n9055)
         );
  XNOR2_X1 U10505 ( .A(n9054), .B(n9055), .ZN(n9303) );
  INV_X1 U10506 ( .A(n9054), .ZN(n9056) );
  NAND2_X1 U10507 ( .A1(n9172), .A2(n4514), .ZN(n9059) );
  OR2_X1 U10508 ( .A1(n9057), .A2(n9207), .ZN(n9058) );
  NAND2_X1 U10509 ( .A1(n9059), .A2(n9058), .ZN(n9060) );
  XNOR2_X1 U10510 ( .A(n9060), .B(n9140), .ZN(n9062) );
  AOI22_X1 U10511 ( .A1(n9172), .A2(n9082), .B1(n9081), .B2(n9385), .ZN(n9171)
         );
  INV_X1 U10512 ( .A(n9062), .ZN(n9063) );
  NAND2_X1 U10513 ( .A1(n9061), .A2(n9063), .ZN(n9064) );
  NAND2_X1 U10514 ( .A1(n9169), .A2(n9064), .ZN(n9256) );
  NAND2_X1 U10515 ( .A1(n9846), .A2(n4514), .ZN(n9066) );
  NAND2_X1 U10516 ( .A1(n9383), .A2(n6752), .ZN(n9065) );
  NAND2_X1 U10517 ( .A1(n9066), .A2(n9065), .ZN(n9067) );
  XNOR2_X1 U10518 ( .A(n9067), .B(n9140), .ZN(n9260) );
  AOI22_X1 U10519 ( .A1(n9846), .A2(n9082), .B1(n9081), .B2(n9383), .ZN(n9259)
         );
  INV_X1 U10520 ( .A(n9259), .ZN(n9073) );
  NOR2_X1 U10521 ( .A1(n9068), .A2(n9201), .ZN(n9069) );
  AOI21_X1 U10522 ( .B1(n9708), .B2(n9137), .A(n9069), .ZN(n9074) );
  INV_X1 U10523 ( .A(n9074), .ZN(n9363) );
  NAND2_X1 U10524 ( .A1(n9708), .A2(n4514), .ZN(n9071) );
  NAND2_X1 U10525 ( .A1(n9384), .A2(n6752), .ZN(n9070) );
  NAND2_X1 U10526 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  XNOR2_X1 U10527 ( .A(n9072), .B(n9204), .ZN(n9258) );
  INV_X1 U10528 ( .A(n9258), .ZN(n9076) );
  AOI22_X1 U10529 ( .A1(n9260), .A2(n9073), .B1(n9363), .B2(n9076), .ZN(n9079)
         );
  AOI21_X1 U10530 ( .B1(n9258), .B2(n9074), .A(n9259), .ZN(n9077) );
  NAND2_X1 U10531 ( .A1(n9259), .A2(n9074), .ZN(n9075) );
  OAI22_X1 U10532 ( .A1(n9077), .A2(n9260), .B1(n9076), .B2(n9075), .ZN(n9078)
         );
  OAI22_X1 U10533 ( .A1(n9681), .A2(n9112), .B1(n9340), .B2(n9207), .ZN(n9080)
         );
  XOR2_X1 U10534 ( .A(n9140), .B(n9080), .Z(n9084) );
  AOI22_X1 U10535 ( .A1(n9840), .A2(n9082), .B1(n9081), .B2(n9382), .ZN(n9083)
         );
  NOR2_X1 U10536 ( .A1(n9084), .A2(n9083), .ZN(n9270) );
  NAND2_X1 U10537 ( .A1(n9766), .A2(n4514), .ZN(n9086) );
  OR2_X1 U10538 ( .A1(n9272), .A2(n9207), .ZN(n9085) );
  NAND2_X1 U10539 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  XNOR2_X1 U10540 ( .A(n9087), .B(n9204), .ZN(n9089) );
  NOR2_X1 U10541 ( .A1(n9272), .A2(n9201), .ZN(n9088) );
  AOI21_X1 U10542 ( .B1(n9766), .B2(n9137), .A(n9088), .ZN(n9090) );
  AND2_X1 U10543 ( .A1(n9089), .A2(n9090), .ZN(n9336) );
  INV_X1 U10544 ( .A(n9089), .ZN(n9092) );
  INV_X1 U10545 ( .A(n9090), .ZN(n9091) );
  NAND2_X1 U10546 ( .A1(n9092), .A2(n9091), .ZN(n9337) );
  NAND2_X1 U10547 ( .A1(n9648), .A2(n4514), .ZN(n9094) );
  NAND2_X1 U10548 ( .A1(n9381), .A2(n6752), .ZN(n9093) );
  NAND2_X1 U10549 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  XNOR2_X1 U10550 ( .A(n9095), .B(n9204), .ZN(n9098) );
  NOR2_X1 U10551 ( .A1(n9341), .A2(n9201), .ZN(n9096) );
  AOI21_X1 U10552 ( .B1(n9648), .B2(n9137), .A(n9096), .ZN(n9097) );
  NOR2_X1 U10553 ( .A1(n9098), .A2(n9097), .ZN(n9194) );
  AOI22_X1 U10554 ( .A1(n9627), .A2(n4514), .B1(n9137), .B2(n9380), .ZN(n9099)
         );
  XOR2_X1 U10555 ( .A(n9140), .B(n9099), .Z(n9101) );
  OAI22_X1 U10556 ( .A1(n9828), .A2(n9207), .B1(n9227), .B2(n9201), .ZN(n9100)
         );
  NOR2_X1 U10557 ( .A1(n9101), .A2(n9100), .ZN(n9102) );
  AOI21_X1 U10558 ( .B1(n9101), .B2(n9100), .A(n9102), .ZN(n9294) );
  NAND2_X1 U10559 ( .A1(n9293), .A2(n9294), .ZN(n9292) );
  INV_X1 U10560 ( .A(n9102), .ZN(n9103) );
  OAI22_X1 U10561 ( .A1(n9614), .A2(n9207), .B1(n9316), .B2(n9201), .ZN(n9108)
         );
  NAND2_X1 U10562 ( .A1(n9752), .A2(n4514), .ZN(n9105) );
  OR2_X1 U10563 ( .A1(n9316), .A2(n9207), .ZN(n9104) );
  NAND2_X1 U10564 ( .A1(n9105), .A2(n9104), .ZN(n9106) );
  XNOR2_X1 U10565 ( .A(n9106), .B(n9140), .ZN(n9107) );
  XOR2_X1 U10566 ( .A(n9108), .B(n9107), .Z(n9225) );
  INV_X1 U10567 ( .A(n9107), .ZN(n9110) );
  INV_X1 U10568 ( .A(n9108), .ZN(n9109) );
  NAND2_X1 U10569 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  OAI22_X1 U10570 ( .A1(n9747), .A2(n9112), .B1(n9180), .B2(n9207), .ZN(n9113)
         );
  XOR2_X1 U10571 ( .A(n9140), .B(n9113), .Z(n9115) );
  INV_X1 U10572 ( .A(n9115), .ZN(n9114) );
  OAI22_X1 U10573 ( .A1(n9747), .A2(n9207), .B1(n9180), .B2(n9201), .ZN(n9314)
         );
  NAND2_X1 U10574 ( .A1(n9742), .A2(n4514), .ZN(n9119) );
  OR2_X1 U10575 ( .A1(n9315), .A2(n9207), .ZN(n9118) );
  NAND2_X1 U10576 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  XNOR2_X1 U10577 ( .A(n9120), .B(n9204), .ZN(n9123) );
  NOR2_X1 U10578 ( .A1(n9315), .A2(n9201), .ZN(n9121) );
  AOI21_X1 U10579 ( .B1(n9742), .B2(n9137), .A(n9121), .ZN(n9122) );
  NAND2_X1 U10580 ( .A1(n9123), .A2(n9122), .ZN(n9286) );
  OR2_X1 U10581 ( .A1(n9123), .A2(n9122), .ZN(n9124) );
  NAND2_X1 U10582 ( .A1(n9813), .A2(n4514), .ZN(n9126) );
  OR2_X1 U10583 ( .A1(n9247), .A2(n9207), .ZN(n9125) );
  NAND2_X1 U10584 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  XNOR2_X1 U10585 ( .A(n9127), .B(n9204), .ZN(n9130) );
  NOR2_X1 U10586 ( .A1(n9247), .A2(n9201), .ZN(n9128) );
  AOI21_X1 U10587 ( .B1(n9813), .B2(n9137), .A(n9128), .ZN(n9129) );
  NAND2_X1 U10588 ( .A1(n9130), .A2(n9129), .ZN(n9132) );
  OR2_X1 U10589 ( .A1(n9130), .A2(n9129), .ZN(n9131) );
  INV_X1 U10590 ( .A(n9808), .ZN(n9549) );
  OAI22_X1 U10591 ( .A1(n9549), .A2(n9207), .B1(n9351), .B2(n9201), .ZN(n9142)
         );
  NAND2_X1 U10592 ( .A1(n9808), .A2(n4514), .ZN(n9134) );
  OR2_X1 U10593 ( .A1(n9351), .A2(n9207), .ZN(n9133) );
  NAND2_X1 U10594 ( .A1(n9134), .A2(n9133), .ZN(n9135) );
  XNOR2_X1 U10595 ( .A(n9135), .B(n9140), .ZN(n9143) );
  XOR2_X1 U10596 ( .A(n9142), .B(n9143), .Z(n9246) );
  NOR2_X1 U10597 ( .A1(n9248), .A2(n9201), .ZN(n9136) );
  AOI21_X1 U10598 ( .B1(n9729), .B2(n9137), .A(n9136), .ZN(n9145) );
  NAND2_X1 U10599 ( .A1(n9729), .A2(n4514), .ZN(n9139) );
  OR2_X1 U10600 ( .A1(n9248), .A2(n9207), .ZN(n9138) );
  NAND2_X1 U10601 ( .A1(n9139), .A2(n9138), .ZN(n9141) );
  XNOR2_X1 U10602 ( .A(n9141), .B(n9140), .ZN(n9147) );
  XOR2_X1 U10603 ( .A(n9145), .B(n9147), .Z(n9347) );
  NOR2_X1 U10604 ( .A1(n9143), .A2(n9142), .ZN(n9348) );
  NOR2_X1 U10605 ( .A1(n9347), .A2(n9348), .ZN(n9144) );
  INV_X1 U10606 ( .A(n9145), .ZN(n9146) );
  NAND2_X1 U10607 ( .A1(n9147), .A2(n9146), .ZN(n9157) );
  NAND2_X1 U10608 ( .A1(n9724), .A2(n4514), .ZN(n9149) );
  OR2_X1 U10609 ( .A1(n9353), .A2(n9207), .ZN(n9148) );
  NAND2_X1 U10610 ( .A1(n9149), .A2(n9148), .ZN(n9150) );
  XNOR2_X1 U10611 ( .A(n9150), .B(n9204), .ZN(n9153) );
  INV_X1 U10612 ( .A(n9153), .ZN(n9155) );
  NOR2_X1 U10613 ( .A1(n9353), .A2(n9201), .ZN(n9151) );
  AOI21_X1 U10614 ( .B1(n9724), .B2(n9137), .A(n9151), .ZN(n9152) );
  INV_X1 U10615 ( .A(n9152), .ZN(n9154) );
  AOI21_X1 U10616 ( .B1(n9155), .B2(n9154), .A(n9217), .ZN(n9156) );
  AOI21_X1 U10617 ( .B1(n9160), .B2(n9157), .A(n9156), .ZN(n9161) );
  INV_X1 U10618 ( .A(n9156), .ZN(n9159) );
  INV_X1 U10619 ( .A(n9157), .ZN(n9158) );
  INV_X1 U10620 ( .A(n9162), .ZN(n9515) );
  OR2_X1 U10621 ( .A1(n9208), .A2(n9352), .ZN(n9164) );
  OR2_X1 U10622 ( .A1(n9248), .A2(n9350), .ZN(n9163) );
  AND2_X1 U10623 ( .A1(n9164), .A2(n9163), .ZN(n9512) );
  OAI22_X1 U10624 ( .A1(n9357), .A2(n9512), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9165), .ZN(n9166) );
  AOI21_X1 U10625 ( .B1(n9359), .B2(n9515), .A(n9166), .ZN(n9167) );
  OAI211_X1 U10626 ( .C1(n9518), .C2(n9928), .A(n9168), .B(n9167), .ZN(
        P1_U3214) );
  OAI21_X1 U10627 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9178) );
  NAND2_X1 U10628 ( .A1(n9172), .A2(n9368), .ZN(n9175) );
  AOI22_X1 U10629 ( .A1(n9926), .A2(n9173), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n9174) );
  OAI211_X1 U10630 ( .C1(n9935), .C2(n9176), .A(n9175), .B(n9174), .ZN(n9177)
         );
  AOI21_X1 U10631 ( .B1(n9178), .B2(n9931), .A(n9177), .ZN(n9179) );
  INV_X1 U10632 ( .A(n9179), .ZN(P1_U3215) );
  OR2_X1 U10633 ( .A1(n9247), .A2(n9352), .ZN(n9182) );
  INV_X1 U10634 ( .A(n9180), .ZN(n9378) );
  NAND2_X1 U10635 ( .A1(n9378), .A2(n9296), .ZN(n9181) );
  NAND2_X1 U10636 ( .A1(n9182), .A2(n9181), .ZN(n9576) );
  AOI22_X1 U10637 ( .A1(n9576), .A2(n9926), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9183) );
  OAI21_X1 U10638 ( .B1(n9935), .B2(n9184), .A(n9183), .ZN(n9192) );
  INV_X1 U10639 ( .A(n9187), .ZN(n9188) );
  NAND3_X1 U10640 ( .A1(n9186), .A2(n9189), .A3(n9188), .ZN(n9190) );
  AOI21_X1 U10641 ( .B1(n9185), .B2(n9190), .A(n9370), .ZN(n9191) );
  AOI211_X1 U10642 ( .C1(n9742), .C2(n9368), .A(n9192), .B(n9191), .ZN(n9193)
         );
  INV_X1 U10643 ( .A(n9193), .ZN(P1_U3216) );
  NOR2_X1 U10644 ( .A1(n9194), .A2(n4500), .ZN(n9195) );
  XNOR2_X1 U10645 ( .A(n9196), .B(n9195), .ZN(n9200) );
  OAI22_X1 U10646 ( .A1(n9227), .A2(n9352), .B1(n9272), .B2(n9350), .ZN(n9637)
         );
  AOI22_X1 U10647 ( .A1(n9637), .A2(n9926), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9197) );
  OAI21_X1 U10648 ( .B1(n9935), .B2(n9642), .A(n9197), .ZN(n9198) );
  AOI21_X1 U10649 ( .B1(n9648), .B2(n9368), .A(n9198), .ZN(n9199) );
  OAI21_X1 U10650 ( .B1(n9200), .B2(n9370), .A(n9199), .ZN(P1_U3219) );
  NAND2_X1 U10651 ( .A1(n9719), .A2(n6752), .ZN(n9203) );
  OR2_X1 U10652 ( .A1(n9208), .A2(n9201), .ZN(n9202) );
  NAND2_X1 U10653 ( .A1(n9203), .A2(n9202), .ZN(n9205) );
  XNOR2_X1 U10654 ( .A(n9205), .B(n9204), .ZN(n9210) );
  NAND2_X1 U10655 ( .A1(n9719), .A2(n4514), .ZN(n9206) );
  OAI21_X1 U10656 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9209) );
  XNOR2_X1 U10657 ( .A(n9210), .B(n9209), .ZN(n9218) );
  NAND3_X1 U10658 ( .A1(n9211), .A2(n9931), .A3(n9218), .ZN(n9221) );
  OR2_X1 U10659 ( .A1(n9212), .A2(n9352), .ZN(n9214) );
  OR2_X1 U10660 ( .A1(n9353), .A2(n9350), .ZN(n9213) );
  NAND2_X1 U10661 ( .A1(n9214), .A2(n9213), .ZN(n9495) );
  AOI22_X1 U10662 ( .A1(n9926), .A2(n9495), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9215) );
  OAI21_X1 U10663 ( .B1(n9935), .B2(n9501), .A(n9215), .ZN(n9216) );
  AOI21_X1 U10664 ( .B1(n9719), .B2(n9368), .A(n9216), .ZN(n9220) );
  NAND3_X1 U10665 ( .A1(n9218), .A2(n9931), .A3(n9217), .ZN(n9219) );
  NAND4_X1 U10666 ( .A1(n9222), .A2(n9221), .A3(n9220), .A4(n9219), .ZN(
        P1_U3220) );
  OAI21_X1 U10667 ( .B1(n9225), .B2(n9224), .A(n9223), .ZN(n9226) );
  NAND2_X1 U10668 ( .A1(n9226), .A2(n9931), .ZN(n9233) );
  NOR2_X1 U10669 ( .A1(n9227), .A2(n9350), .ZN(n9228) );
  AOI21_X1 U10670 ( .B1(n9378), .B2(n9229), .A(n9228), .ZN(n9608) );
  OAI22_X1 U10671 ( .A1(n9608), .A2(n9357), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9230), .ZN(n9231) );
  AOI21_X1 U10672 ( .B1(n9611), .B2(n9359), .A(n9231), .ZN(n9232) );
  OAI211_X1 U10673 ( .C1(n9614), .C2(n9928), .A(n9233), .B(n9232), .ZN(
        P1_U3223) );
  XOR2_X1 U10674 ( .A(n9234), .B(n9235), .Z(n9243) );
  NAND2_X1 U10675 ( .A1(n9926), .A2(n9236), .ZN(n9237) );
  OAI211_X1 U10676 ( .C1(n9935), .C2(n9239), .A(n9238), .B(n9237), .ZN(n9240)
         );
  AOI21_X1 U10677 ( .B1(n9241), .B2(n9368), .A(n9240), .ZN(n9242) );
  OAI21_X1 U10678 ( .B1(n9243), .B2(n9370), .A(n9242), .ZN(P1_U3224) );
  OAI21_X1 U10679 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9254) );
  NAND2_X1 U10680 ( .A1(n9808), .A2(n9368), .ZN(n9252) );
  OR2_X1 U10681 ( .A1(n9247), .A2(n9350), .ZN(n9250) );
  OR2_X1 U10682 ( .A1(n9248), .A2(n9352), .ZN(n9249) );
  NAND2_X1 U10683 ( .A1(n9250), .A2(n9249), .ZN(n9539) );
  AOI22_X1 U10684 ( .A1(n9539), .A2(n9926), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9251) );
  OAI211_X1 U10685 ( .C1(n9935), .C2(n9545), .A(n9252), .B(n9251), .ZN(n9253)
         );
  AOI21_X1 U10686 ( .B1(n9254), .B2(n9931), .A(n9253), .ZN(n9255) );
  INV_X1 U10687 ( .A(n9255), .ZN(P1_U3225) );
  XNOR2_X1 U10688 ( .A(n9257), .B(n9258), .ZN(n9364) );
  NOR2_X1 U10689 ( .A1(n9364), .A2(n9363), .ZN(n9362) );
  AOI21_X1 U10690 ( .B1(n9258), .B2(n9257), .A(n9362), .ZN(n9262) );
  XNOR2_X1 U10691 ( .A(n9260), .B(n9259), .ZN(n9261) );
  XNOR2_X1 U10692 ( .A(n9262), .B(n9261), .ZN(n9268) );
  OR2_X1 U10693 ( .A1(n9340), .A2(n9352), .ZN(n9264) );
  NAND2_X1 U10694 ( .A1(n9384), .A2(n9296), .ZN(n9263) );
  NAND2_X1 U10695 ( .A1(n9264), .A2(n9263), .ZN(n9696) );
  AOI22_X1 U10696 ( .A1(n9926), .A2(n9696), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3086), .ZN(n9265) );
  OAI21_X1 U10697 ( .B1(n9935), .B2(n9689), .A(n9265), .ZN(n9266) );
  AOI21_X1 U10698 ( .B1(n9846), .B2(n9368), .A(n9266), .ZN(n9267) );
  OAI21_X1 U10699 ( .B1(n9268), .B2(n9370), .A(n9267), .ZN(P1_U3226) );
  NOR2_X1 U10700 ( .A1(n9270), .A2(n4499), .ZN(n9271) );
  XNOR2_X1 U10701 ( .A(n9269), .B(n9271), .ZN(n9279) );
  OR2_X1 U10702 ( .A1(n9272), .A2(n9352), .ZN(n9274) );
  NAND2_X1 U10703 ( .A1(n9383), .A2(n9296), .ZN(n9273) );
  AND2_X1 U10704 ( .A1(n9274), .A2(n9273), .ZN(n9677) );
  NAND2_X1 U10705 ( .A1(n9359), .A2(n9682), .ZN(n9276) );
  OAI211_X1 U10706 ( .C1(n9677), .C2(n9357), .A(n9276), .B(n9275), .ZN(n9277)
         );
  AOI21_X1 U10707 ( .B1(n9840), .B2(n9368), .A(n9277), .ZN(n9278) );
  OAI21_X1 U10708 ( .B1(n9279), .B2(n9370), .A(n9278), .ZN(P1_U3228) );
  OR2_X1 U10709 ( .A1(n9315), .A2(n9350), .ZN(n9281) );
  OR2_X1 U10710 ( .A1(n9351), .A2(n9352), .ZN(n9280) );
  NAND2_X1 U10711 ( .A1(n9281), .A2(n9280), .ZN(n9563) );
  AOI22_X1 U10712 ( .A1(n9563), .A2(n9926), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9282) );
  OAI21_X1 U10713 ( .B1(n9935), .B2(n9283), .A(n9282), .ZN(n9290) );
  INV_X1 U10714 ( .A(n9284), .ZN(n9285) );
  NAND3_X1 U10715 ( .A1(n9185), .A2(n9286), .A3(n9285), .ZN(n9287) );
  AOI21_X1 U10716 ( .B1(n9288), .B2(n9287), .A(n9370), .ZN(n9289) );
  AOI211_X1 U10717 ( .C1(n9813), .C2(n9368), .A(n9290), .B(n9289), .ZN(n9291)
         );
  INV_X1 U10718 ( .A(n9291), .ZN(P1_U3229) );
  OAI21_X1 U10719 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9295) );
  NAND2_X1 U10720 ( .A1(n9295), .A2(n9931), .ZN(n9302) );
  OR2_X1 U10721 ( .A1(n9316), .A2(n9352), .ZN(n9298) );
  NAND2_X1 U10722 ( .A1(n9381), .A2(n9296), .ZN(n9297) );
  AND2_X1 U10723 ( .A1(n9298), .A2(n9297), .ZN(n9622) );
  OAI22_X1 U10724 ( .A1(n9622), .A2(n9357), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9299), .ZN(n9300) );
  AOI21_X1 U10725 ( .B1(n9629), .B2(n9359), .A(n9300), .ZN(n9301) );
  OAI211_X1 U10726 ( .C1(n9828), .C2(n9928), .A(n9302), .B(n9301), .ZN(
        P1_U3233) );
  XOR2_X1 U10727 ( .A(n9304), .B(n9303), .Z(n9311) );
  AOI22_X1 U10728 ( .A1(n9926), .A2(n9305), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n9306) );
  OAI21_X1 U10729 ( .B1(n9935), .B2(n9307), .A(n9306), .ZN(n9308) );
  AOI21_X1 U10730 ( .B1(n9309), .B2(n9368), .A(n9308), .ZN(n9310) );
  OAI21_X1 U10731 ( .B1(n9311), .B2(n9370), .A(n9310), .ZN(P1_U3234) );
  INV_X1 U10732 ( .A(n9186), .ZN(n9312) );
  AOI21_X1 U10733 ( .B1(n9314), .B2(n9313), .A(n9312), .ZN(n9322) );
  OR2_X1 U10734 ( .A1(n9315), .A2(n9352), .ZN(n9318) );
  OR2_X1 U10735 ( .A1(n9316), .A2(n9350), .ZN(n9317) );
  NAND2_X1 U10736 ( .A1(n9318), .A2(n9317), .ZN(n9590) );
  AOI22_X1 U10737 ( .A1(n9590), .A2(n9926), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9319) );
  OAI21_X1 U10738 ( .B1(n9935), .B2(n9596), .A(n9319), .ZN(n9320) );
  AOI21_X1 U10739 ( .B1(n9600), .B2(n9368), .A(n9320), .ZN(n9321) );
  OAI21_X1 U10740 ( .B1(n9322), .B2(n9370), .A(n9321), .ZN(P1_U3235) );
  INV_X1 U10741 ( .A(n9323), .ZN(n9328) );
  AOI21_X1 U10742 ( .B1(n9325), .B2(n9327), .A(n9324), .ZN(n9326) );
  AOI21_X1 U10743 ( .B1(n9328), .B2(n9327), .A(n9326), .ZN(n9335) );
  AOI22_X1 U10744 ( .A1(n9926), .A2(n9329), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9330) );
  OAI21_X1 U10745 ( .B1(n9935), .B2(n9331), .A(n9330), .ZN(n9332) );
  AOI21_X1 U10746 ( .B1(n9333), .B2(n9368), .A(n9332), .ZN(n9334) );
  OAI21_X1 U10747 ( .B1(n9335), .B2(n9370), .A(n9334), .ZN(P1_U3236) );
  NAND2_X1 U10748 ( .A1(n4660), .A2(n9337), .ZN(n9338) );
  XNOR2_X1 U10749 ( .A(n9339), .B(n9338), .ZN(n9346) );
  INV_X1 U10750 ( .A(n9666), .ZN(n9343) );
  OAI22_X1 U10751 ( .A1(n9341), .A2(n9352), .B1(n9340), .B2(n9350), .ZN(n9659)
         );
  AOI22_X1 U10752 ( .A1(n9926), .A2(n9659), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9342) );
  OAI21_X1 U10753 ( .B1(n9935), .B2(n9343), .A(n9342), .ZN(n9344) );
  AOI21_X1 U10754 ( .B1(n9766), .B2(n9368), .A(n9344), .ZN(n9345) );
  OAI21_X1 U10755 ( .B1(n9346), .B2(n9370), .A(n9345), .ZN(P1_U3238) );
  INV_X1 U10756 ( .A(n9349), .ZN(n9531) );
  OR2_X1 U10757 ( .A1(n9351), .A2(n9350), .ZN(n9355) );
  OR2_X1 U10758 ( .A1(n9353), .A2(n9352), .ZN(n9354) );
  AND2_X1 U10759 ( .A1(n9355), .A2(n9354), .ZN(n9526) );
  OAI22_X1 U10760 ( .A1(n9357), .A2(n9526), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9356), .ZN(n9358) );
  AOI21_X1 U10761 ( .B1(n9359), .B2(n9531), .A(n9358), .ZN(n9360) );
  OAI211_X1 U10762 ( .C1(n9534), .C2(n9928), .A(n9361), .B(n9360), .ZN(
        P1_U3240) );
  AOI21_X1 U10763 ( .B1(n9364), .B2(n9363), .A(n9362), .ZN(n9371) );
  AOI22_X1 U10764 ( .A1(n9926), .A2(n9365), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9366) );
  OAI21_X1 U10765 ( .B1(n9935), .B2(n9704), .A(n9366), .ZN(n9367) );
  AOI21_X1 U10766 ( .B1(n9708), .B2(n9368), .A(n9367), .ZN(n9369) );
  OAI21_X1 U10767 ( .B1(n9371), .B2(n9370), .A(n9369), .ZN(P1_U3241) );
  MUX2_X1 U10768 ( .A(n9372), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9398), .Z(
        P1_U3584) );
  MUX2_X1 U10769 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9373), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10770 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9374), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10771 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9375), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10772 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9376), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10773 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9377), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10774 ( .A(n9378), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9398), .Z(
        P1_U3576) );
  MUX2_X1 U10775 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9379), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10776 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9380), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10777 ( .A(n9381), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9398), .Z(
        P1_U3573) );
  MUX2_X1 U10778 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9382), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10779 ( .A(n9383), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9398), .Z(
        P1_U3570) );
  MUX2_X1 U10780 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9384), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10781 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9385), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10782 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9386), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10783 ( .A(n9387), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9398), .Z(
        P1_U3566) );
  MUX2_X1 U10784 ( .A(n9388), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9398), .Z(
        P1_U3565) );
  MUX2_X1 U10785 ( .A(n9389), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9398), .Z(
        P1_U3564) );
  MUX2_X1 U10786 ( .A(n9390), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9398), .Z(
        P1_U3563) );
  MUX2_X1 U10787 ( .A(n9391), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9398), .Z(
        P1_U3562) );
  MUX2_X1 U10788 ( .A(n9392), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9398), .Z(
        P1_U3561) );
  MUX2_X1 U10789 ( .A(n9393), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9398), .Z(
        P1_U3560) );
  MUX2_X1 U10790 ( .A(n9394), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9398), .Z(
        P1_U3559) );
  MUX2_X1 U10791 ( .A(n9395), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9398), .Z(
        P1_U3558) );
  MUX2_X1 U10792 ( .A(n9396), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9398), .Z(
        P1_U3557) );
  MUX2_X1 U10793 ( .A(n9397), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9398), .Z(
        P1_U3556) );
  MUX2_X1 U10794 ( .A(n9399), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9398), .Z(
        P1_U3555) );
  OAI211_X1 U10795 ( .C1(n9402), .C2(n9401), .A(n9474), .B(n9400), .ZN(n9410)
         );
  AOI22_X1 U10796 ( .A1(n9948), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9409) );
  NAND2_X1 U10797 ( .A1(n10031), .A2(n9403), .ZN(n9408) );
  OAI211_X1 U10798 ( .C1(n9406), .C2(n9405), .A(n10024), .B(n9404), .ZN(n9407)
         );
  NAND4_X1 U10799 ( .A1(n9410), .A2(n9409), .A3(n9408), .A4(n9407), .ZN(
        P1_U3244) );
  INV_X1 U10800 ( .A(n9411), .ZN(n9415) );
  NAND2_X1 U10801 ( .A1(n9948), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n9412) );
  OAI21_X1 U10802 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9413), .A(n9412), .ZN(
        n9414) );
  AOI21_X1 U10803 ( .B1(n9415), .B2(n10031), .A(n9414), .ZN(n9424) );
  OAI211_X1 U10804 ( .C1(n9418), .C2(n9417), .A(n9474), .B(n9416), .ZN(n9423)
         );
  OAI211_X1 U10805 ( .C1(n9421), .C2(n9420), .A(n10024), .B(n9419), .ZN(n9422)
         );
  NAND4_X1 U10806 ( .A1(n9425), .A2(n9424), .A3(n9423), .A4(n9422), .ZN(
        P1_U3245) );
  INV_X1 U10807 ( .A(n9426), .ZN(n9430) );
  INV_X1 U10808 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U10809 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9427) );
  OAI21_X1 U10810 ( .B1(n10039), .B2(n9428), .A(n9427), .ZN(n9429) );
  AOI21_X1 U10811 ( .B1(n9430), .B2(n10031), .A(n9429), .ZN(n9439) );
  OAI211_X1 U10812 ( .C1(n9433), .C2(n9432), .A(n9474), .B(n9431), .ZN(n9438)
         );
  OAI211_X1 U10813 ( .C1(n9436), .C2(n9435), .A(n10024), .B(n9434), .ZN(n9437)
         );
  NAND3_X1 U10814 ( .A1(n9439), .A2(n9438), .A3(n9437), .ZN(P1_U3246) );
  INV_X1 U10815 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9441) );
  NAND2_X1 U10816 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9440) );
  OAI21_X1 U10817 ( .B1(n10039), .B2(n9441), .A(n9440), .ZN(n9442) );
  AOI21_X1 U10818 ( .B1(n9443), .B2(n10031), .A(n9442), .ZN(n9452) );
  OAI211_X1 U10819 ( .C1(n9446), .C2(n9445), .A(n9474), .B(n9444), .ZN(n9451)
         );
  OAI211_X1 U10820 ( .C1(n9449), .C2(n9448), .A(n10024), .B(n9447), .ZN(n9450)
         );
  NAND3_X1 U10821 ( .A1(n9452), .A2(n9451), .A3(n9450), .ZN(P1_U3248) );
  INV_X1 U10822 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9454) );
  NAND2_X1 U10823 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9453) );
  OAI21_X1 U10824 ( .B1(n10039), .B2(n9454), .A(n9453), .ZN(n9455) );
  AOI21_X1 U10825 ( .B1(n9456), .B2(n10031), .A(n9455), .ZN(n9465) );
  OAI211_X1 U10826 ( .C1(n9459), .C2(n9458), .A(n9474), .B(n9457), .ZN(n9464)
         );
  OAI211_X1 U10827 ( .C1(n9462), .C2(n9461), .A(n10024), .B(n9460), .ZN(n9463)
         );
  NAND3_X1 U10828 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(P1_U3249) );
  OAI21_X1 U10829 ( .B1(n10039), .B2(n9467), .A(n9466), .ZN(n9468) );
  AOI21_X1 U10830 ( .B1(n9469), .B2(n10031), .A(n9468), .ZN(n9479) );
  OAI211_X1 U10831 ( .C1(n9472), .C2(n9471), .A(n10024), .B(n9470), .ZN(n9478)
         );
  OAI211_X1 U10832 ( .C1(n9476), .C2(n9475), .A(n9474), .B(n9473), .ZN(n9477)
         );
  NAND3_X1 U10833 ( .A1(n9479), .A2(n9478), .A3(n9477), .ZN(P1_U3250) );
  NAND2_X1 U10834 ( .A1(n9714), .A2(n9665), .ZN(n9486) );
  INV_X1 U10835 ( .A(n9482), .ZN(n9483) );
  AND2_X1 U10836 ( .A1(n9484), .A2(n9483), .ZN(n9713) );
  INV_X1 U10837 ( .A(n9713), .ZN(n9936) );
  NOR2_X1 U10838 ( .A1(n9581), .A2(n9936), .ZN(n9489) );
  AOI21_X1 U10839 ( .B1(n9712), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9489), .ZN(
        n9485) );
  OAI211_X1 U10840 ( .C1(n9793), .C2(n10062), .A(n9486), .B(n9485), .ZN(
        P1_U3263) );
  XNOR2_X1 U10841 ( .A(n9488), .B(n9487), .ZN(n9940) );
  NAND2_X1 U10842 ( .A1(n9940), .A2(n10060), .ZN(n9491) );
  AOI21_X1 U10843 ( .B1(n9712), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9489), .ZN(
        n9490) );
  OAI211_X1 U10844 ( .C1(n9937), .C2(n10062), .A(n9491), .B(n9490), .ZN(
        P1_U3264) );
  XNOR2_X1 U10845 ( .A(n9494), .B(n9493), .ZN(n9497) );
  INV_X1 U10846 ( .A(n9495), .ZN(n9496) );
  OAI21_X1 U10847 ( .B1(n9497), .B2(n9578), .A(n9496), .ZN(n9717) );
  INV_X1 U10848 ( .A(n9514), .ZN(n9500) );
  INV_X1 U10849 ( .A(n9498), .ZN(n9499) );
  AOI211_X1 U10850 ( .C1(n9719), .C2(n9500), .A(n9664), .B(n9499), .ZN(n9718)
         );
  NAND2_X1 U10851 ( .A1(n9718), .A2(n9665), .ZN(n9504) );
  INV_X1 U10852 ( .A(n9501), .ZN(n9502) );
  AOI22_X1 U10853 ( .A1(n9581), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9502), .B2(
        n10065), .ZN(n9503) );
  OAI211_X1 U10854 ( .C1(n9505), .C2(n10062), .A(n9504), .B(n9503), .ZN(n9506)
         );
  AOI21_X1 U10855 ( .B1(n10067), .B2(n9717), .A(n9506), .ZN(n9507) );
  OAI21_X1 U10856 ( .B1(n9797), .B2(n9701), .A(n9507), .ZN(P1_U3265) );
  XNOR2_X1 U10857 ( .A(n9509), .B(n9508), .ZN(n9801) );
  XNOR2_X1 U10858 ( .A(n9511), .B(n9510), .ZN(n9513) );
  OAI21_X1 U10859 ( .B1(n9513), .B2(n9578), .A(n9512), .ZN(n9723) );
  AOI211_X1 U10860 ( .C1(n9724), .C2(n9529), .A(n9664), .B(n9514), .ZN(n9722)
         );
  NAND2_X1 U10861 ( .A1(n9722), .A2(n9665), .ZN(n9517) );
  AOI22_X1 U10862 ( .A1(n9581), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9515), .B2(
        n10065), .ZN(n9516) );
  OAI211_X1 U10863 ( .C1(n9518), .C2(n10062), .A(n9517), .B(n9516), .ZN(n9519)
         );
  AOI21_X1 U10864 ( .B1(n10067), .B2(n9723), .A(n9519), .ZN(n9520) );
  OAI21_X1 U10865 ( .B1(n9801), .B2(n9701), .A(n9520), .ZN(P1_U3266) );
  NAND2_X1 U10866 ( .A1(n9537), .A2(n9522), .ZN(n9524) );
  XNOR2_X1 U10867 ( .A(n9524), .B(n9523), .ZN(n9525) );
  NAND2_X1 U10868 ( .A1(n9527), .A2(n9526), .ZN(n9728) );
  INV_X1 U10869 ( .A(n9528), .ZN(n9547) );
  INV_X1 U10870 ( .A(n9529), .ZN(n9530) );
  AOI211_X1 U10871 ( .C1(n9729), .C2(n9547), .A(n9664), .B(n9530), .ZN(n9727)
         );
  NAND2_X1 U10872 ( .A1(n9727), .A2(n9665), .ZN(n9533) );
  AOI22_X1 U10873 ( .A1(n9581), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9531), .B2(
        n10065), .ZN(n9532) );
  OAI211_X1 U10874 ( .C1(n9534), .C2(n10062), .A(n9533), .B(n9532), .ZN(n9535)
         );
  AOI21_X1 U10875 ( .B1(n10067), .B2(n9728), .A(n9535), .ZN(n9536) );
  OAI21_X1 U10876 ( .B1(n9805), .B2(n9701), .A(n9536), .ZN(P1_U3267) );
  OAI211_X1 U10877 ( .C1(n9542), .C2(n9538), .A(n9537), .B(n9697), .ZN(n9541)
         );
  INV_X1 U10878 ( .A(n9539), .ZN(n9540) );
  XNOR2_X1 U10879 ( .A(n9543), .B(n9542), .ZN(n9810) );
  INV_X1 U10880 ( .A(n9810), .ZN(n9544) );
  NAND2_X1 U10881 ( .A1(n9544), .A2(n10053), .ZN(n9553) );
  OAI22_X1 U10882 ( .A1(n10067), .A2(n9546), .B1(n9545), .B2(n10042), .ZN(
        n9551) );
  INV_X1 U10883 ( .A(n9555), .ZN(n9548) );
  OAI211_X1 U10884 ( .C1(n9549), .C2(n9548), .A(n9547), .B(n9939), .ZN(n9732)
         );
  NOR2_X1 U10885 ( .A1(n9732), .A2(n10049), .ZN(n9550) );
  AOI211_X1 U10886 ( .C1(n10047), .C2(n9808), .A(n9551), .B(n9550), .ZN(n9552)
         );
  OAI211_X1 U10887 ( .C1(n9712), .C2(n9733), .A(n9553), .B(n9552), .ZN(
        P1_U3268) );
  XNOR2_X1 U10888 ( .A(n9554), .B(n9559), .ZN(n9815) );
  OAI211_X1 U10889 ( .C1(n9558), .C2(n9580), .A(n9939), .B(n9555), .ZN(n9736)
         );
  INV_X1 U10890 ( .A(n9736), .ZN(n9568) );
  AOI22_X1 U10891 ( .A1(n9556), .A2(n10065), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n9581), .ZN(n9557) );
  OAI21_X1 U10892 ( .B1(n9558), .B2(n10062), .A(n9557), .ZN(n9567) );
  OAI21_X1 U10893 ( .B1(n9573), .B2(n9560), .A(n9559), .ZN(n9562) );
  NAND3_X1 U10894 ( .A1(n9562), .A2(n9697), .A3(n9561), .ZN(n9565) );
  INV_X1 U10895 ( .A(n9563), .ZN(n9564) );
  AND2_X1 U10896 ( .A1(n9565), .A2(n9564), .ZN(n9737) );
  NOR2_X1 U10897 ( .A1(n9737), .A2(n9581), .ZN(n9566) );
  AOI211_X1 U10898 ( .C1(n9568), .C2(n9628), .A(n9567), .B(n9566), .ZN(n9569)
         );
  OAI21_X1 U10899 ( .B1(n9815), .B2(n9701), .A(n9569), .ZN(P1_U3269) );
  XNOR2_X1 U10900 ( .A(n9571), .B(n9570), .ZN(n9819) );
  INV_X1 U10901 ( .A(n9572), .ZN(n9575) );
  AOI21_X1 U10902 ( .B1(n9575), .B2(n9574), .A(n9573), .ZN(n9579) );
  INV_X1 U10903 ( .A(n9576), .ZN(n9577) );
  OAI21_X1 U10904 ( .B1(n9579), .B2(n9578), .A(n9577), .ZN(n9740) );
  INV_X1 U10905 ( .A(n9742), .ZN(n9585) );
  AOI211_X1 U10906 ( .C1(n9742), .C2(n9597), .A(n9664), .B(n9580), .ZN(n9741)
         );
  NAND2_X1 U10907 ( .A1(n9741), .A2(n9665), .ZN(n9584) );
  AOI22_X1 U10908 ( .A1(n9582), .A2(n10065), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n9581), .ZN(n9583) );
  OAI211_X1 U10909 ( .C1(n9585), .C2(n10062), .A(n9584), .B(n9583), .ZN(n9586)
         );
  AOI21_X1 U10910 ( .B1(n10067), .B2(n9740), .A(n9586), .ZN(n9587) );
  OAI21_X1 U10911 ( .B1(n9819), .B2(n9701), .A(n9587), .ZN(P1_U3270) );
  XNOR2_X1 U10912 ( .A(n9589), .B(n9588), .ZN(n9591) );
  AOI21_X1 U10913 ( .B1(n9591), .B2(n9697), .A(n9590), .ZN(n9746) );
  XNOR2_X1 U10914 ( .A(n9593), .B(n9592), .ZN(n9823) );
  INV_X1 U10915 ( .A(n9823), .ZN(n9594) );
  NAND2_X1 U10916 ( .A1(n9594), .A2(n10053), .ZN(n9602) );
  OAI22_X1 U10917 ( .A1(n9596), .A2(n10042), .B1(n9595), .B2(n10067), .ZN(
        n9599) );
  OAI211_X1 U10918 ( .C1(n9747), .C2(n9610), .A(n9939), .B(n9597), .ZN(n9745)
         );
  NOR2_X1 U10919 ( .A1(n9745), .A2(n10049), .ZN(n9598) );
  AOI211_X1 U10920 ( .C1(n10047), .C2(n9600), .A(n9599), .B(n9598), .ZN(n9601)
         );
  OAI211_X1 U10921 ( .C1(n9712), .C2(n9746), .A(n9602), .B(n9601), .ZN(
        P1_U3271) );
  XNOR2_X1 U10922 ( .A(n4509), .B(n9604), .ZN(n9754) );
  AOI21_X1 U10923 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  OAI21_X1 U10924 ( .B1(n9607), .B2(n4471), .A(n9697), .ZN(n9609) );
  NAND2_X1 U10925 ( .A1(n9609), .A2(n9608), .ZN(n9750) );
  AOI211_X1 U10926 ( .C1(n9752), .C2(n9625), .A(n9664), .B(n9610), .ZN(n9751)
         );
  NAND2_X1 U10927 ( .A1(n9751), .A2(n9665), .ZN(n9613) );
  AOI22_X1 U10928 ( .A1(n9712), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9611), .B2(
        n10065), .ZN(n9612) );
  OAI211_X1 U10929 ( .C1(n9614), .C2(n10062), .A(n9613), .B(n9612), .ZN(n9615)
         );
  AOI21_X1 U10930 ( .B1(n10067), .B2(n9750), .A(n9615), .ZN(n9616) );
  OAI21_X1 U10931 ( .B1(n9754), .B2(n9701), .A(n9616), .ZN(P1_U3272) );
  XOR2_X1 U10932 ( .A(n9618), .B(n9617), .Z(n9757) );
  INV_X1 U10933 ( .A(n9757), .ZN(n9634) );
  INV_X1 U10934 ( .A(n9618), .ZN(n9619) );
  XNOR2_X1 U10935 ( .A(n9620), .B(n9619), .ZN(n9621) );
  NAND2_X1 U10936 ( .A1(n9621), .A2(n9697), .ZN(n9623) );
  NAND2_X1 U10937 ( .A1(n9623), .A2(n9622), .ZN(n9755) );
  INV_X1 U10938 ( .A(n9624), .ZN(n9645) );
  INV_X1 U10939 ( .A(n9625), .ZN(n9626) );
  AOI211_X1 U10940 ( .C1(n9627), .C2(n9645), .A(n9664), .B(n9626), .ZN(n9756)
         );
  NAND2_X1 U10941 ( .A1(n9756), .A2(n9628), .ZN(n9631) );
  AOI22_X1 U10942 ( .A1(n9712), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9629), .B2(
        n10065), .ZN(n9630) );
  OAI211_X1 U10943 ( .C1(n9828), .C2(n10062), .A(n9631), .B(n9630), .ZN(n9632)
         );
  AOI21_X1 U10944 ( .B1(n10067), .B2(n9755), .A(n9632), .ZN(n9633) );
  OAI21_X1 U10945 ( .B1(n9634), .B2(n9701), .A(n9633), .ZN(P1_U3273) );
  XNOR2_X1 U10946 ( .A(n9636), .B(n9635), .ZN(n9638) );
  AOI21_X1 U10947 ( .B1(n9638), .B2(n9697), .A(n9637), .ZN(n9761) );
  XNOR2_X1 U10948 ( .A(n9640), .B(n9639), .ZN(n9830) );
  INV_X1 U10949 ( .A(n9830), .ZN(n9641) );
  NAND2_X1 U10950 ( .A1(n9641), .A2(n10053), .ZN(n9650) );
  INV_X1 U10951 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9643) );
  OAI22_X1 U10952 ( .A1(n10067), .A2(n9643), .B1(n9642), .B2(n10042), .ZN(
        n9647) );
  INV_X1 U10953 ( .A(n9644), .ZN(n9663) );
  OAI211_X1 U10954 ( .C1(n9829), .C2(n9663), .A(n9645), .B(n9939), .ZN(n9760)
         );
  NOR2_X1 U10955 ( .A1(n9760), .A2(n10049), .ZN(n9646) );
  AOI211_X1 U10956 ( .C1(n10047), .C2(n9648), .A(n9647), .B(n9646), .ZN(n9649)
         );
  OAI211_X1 U10957 ( .C1(n9712), .C2(n9761), .A(n9650), .B(n9649), .ZN(
        P1_U3274) );
  OAI21_X1 U10958 ( .B1(n9652), .B2(n9654), .A(n9651), .ZN(n9837) );
  NAND2_X1 U10959 ( .A1(n9676), .A2(n9653), .ZN(n9655) );
  NAND2_X1 U10960 ( .A1(n9655), .A2(n9654), .ZN(n9656) );
  NAND2_X1 U10961 ( .A1(n9657), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U10962 ( .A1(n9658), .A2(n9697), .ZN(n9661) );
  INV_X1 U10963 ( .A(n9659), .ZN(n9660) );
  NAND2_X1 U10964 ( .A1(n9661), .A2(n9660), .ZN(n9765) );
  INV_X1 U10965 ( .A(n9662), .ZN(n9679) );
  AOI211_X1 U10966 ( .C1(n9766), .C2(n9679), .A(n9664), .B(n9663), .ZN(n9764)
         );
  NAND2_X1 U10967 ( .A1(n9764), .A2(n9665), .ZN(n9668) );
  AOI22_X1 U10968 ( .A1(n9712), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9666), .B2(
        n10065), .ZN(n9667) );
  OAI211_X1 U10969 ( .C1(n9669), .C2(n10062), .A(n9668), .B(n9667), .ZN(n9670)
         );
  AOI21_X1 U10970 ( .B1(n10067), .B2(n9765), .A(n9670), .ZN(n9671) );
  OAI21_X1 U10971 ( .B1(n9837), .B2(n9701), .A(n9671), .ZN(P1_U3275) );
  XNOR2_X1 U10972 ( .A(n9672), .B(n9673), .ZN(n9843) );
  NAND2_X1 U10973 ( .A1(n9674), .A2(n9673), .ZN(n9675) );
  NAND3_X1 U10974 ( .A1(n9676), .A2(n9697), .A3(n9675), .ZN(n9678) );
  AND2_X1 U10975 ( .A1(n9678), .A2(n9677), .ZN(n9771) );
  INV_X1 U10976 ( .A(n9771), .ZN(n9686) );
  INV_X1 U10977 ( .A(n9690), .ZN(n9680) );
  OAI211_X1 U10978 ( .C1(n9681), .C2(n9680), .A(n9679), .B(n9939), .ZN(n9770)
         );
  AOI22_X1 U10979 ( .A1(n9712), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9682), .B2(
        n10065), .ZN(n9684) );
  NAND2_X1 U10980 ( .A1(n9840), .A2(n10047), .ZN(n9683) );
  OAI211_X1 U10981 ( .C1(n9770), .C2(n10049), .A(n9684), .B(n9683), .ZN(n9685)
         );
  AOI21_X1 U10982 ( .B1(n9686), .B2(n10067), .A(n9685), .ZN(n9687) );
  OAI21_X1 U10983 ( .B1(n9843), .B2(n9701), .A(n9687), .ZN(P1_U3276) );
  XNOR2_X1 U10984 ( .A(n9688), .B(n9694), .ZN(n9779) );
  OAI22_X1 U10985 ( .A1(n10067), .A2(n8962), .B1(n9689), .B2(n10042), .ZN(
        n9693) );
  OAI211_X1 U10986 ( .C1(n9783), .C2(n9691), .A(n9690), .B(n9939), .ZN(n9776)
         );
  NOR2_X1 U10987 ( .A1(n9776), .A2(n10049), .ZN(n9692) );
  AOI211_X1 U10988 ( .C1(n10047), .C2(n9846), .A(n9693), .B(n9692), .ZN(n9700)
         );
  XNOR2_X1 U10989 ( .A(n9695), .B(n9694), .ZN(n9698) );
  AOI21_X1 U10990 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9777) );
  OR2_X1 U10991 ( .A1(n9777), .A2(n9581), .ZN(n9699) );
  OAI211_X1 U10992 ( .C1(n9779), .C2(n9701), .A(n9700), .B(n9699), .ZN(
        P1_U3277) );
  INV_X1 U10993 ( .A(n9702), .ZN(n9703) );
  NAND2_X1 U10994 ( .A1(n9703), .A2(n10053), .ZN(n9710) );
  OAI22_X1 U10995 ( .A1(n10067), .A2(n10002), .B1(n9704), .B2(n10042), .ZN(
        n9707) );
  NOR2_X1 U10996 ( .A1(n9705), .A2(n10049), .ZN(n9706) );
  AOI211_X1 U10997 ( .C1(n10047), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9709)
         );
  OAI211_X1 U10998 ( .C1(n9712), .C2(n9711), .A(n9710), .B(n9709), .ZN(
        P1_U3278) );
  INV_X1 U10999 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9715) );
  NOR2_X1 U11000 ( .A1(n9714), .A2(n9713), .ZN(n9790) );
  MUX2_X1 U11001 ( .A(n9715), .B(n9790), .S(n10106), .Z(n9716) );
  OAI21_X1 U11002 ( .B1(n9793), .B2(n9789), .A(n9716), .ZN(P1_U3553) );
  AOI211_X1 U11003 ( .C1(n9767), .C2(n9719), .A(n9718), .B(n9717), .ZN(n9794)
         );
  MUX2_X1 U11004 ( .A(n9720), .B(n9794), .S(n10106), .Z(n9721) );
  OAI21_X1 U11005 ( .B1(n9797), .B2(n9775), .A(n9721), .ZN(P1_U3550) );
  INV_X1 U11006 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9725) );
  AOI211_X1 U11007 ( .C1(n9767), .C2(n9724), .A(n9723), .B(n9722), .ZN(n9798)
         );
  MUX2_X1 U11008 ( .A(n9725), .B(n9798), .S(n10106), .Z(n9726) );
  OAI21_X1 U11009 ( .B1(n9801), .B2(n9775), .A(n9726), .ZN(P1_U3549) );
  AOI211_X1 U11010 ( .C1(n9767), .C2(n9729), .A(n9728), .B(n9727), .ZN(n9802)
         );
  MUX2_X1 U11011 ( .A(n9730), .B(n9802), .S(n10106), .Z(n9731) );
  OAI21_X1 U11012 ( .B1(n9805), .B2(n9775), .A(n9731), .ZN(P1_U3548) );
  NAND2_X1 U11013 ( .A1(n9733), .A2(n9732), .ZN(n9806) );
  MUX2_X1 U11014 ( .A(n9806), .B(P1_REG1_REG_25__SCAN_IN), .S(n4826), .Z(n9734) );
  AOI21_X1 U11015 ( .B1(n9773), .B2(n9808), .A(n9734), .ZN(n9735) );
  OAI21_X1 U11016 ( .B1(n9810), .B2(n9775), .A(n9735), .ZN(P1_U3547) );
  NAND2_X1 U11017 ( .A1(n9737), .A2(n9736), .ZN(n9811) );
  MUX2_X1 U11018 ( .A(n9811), .B(P1_REG1_REG_24__SCAN_IN), .S(n4826), .Z(n9738) );
  AOI21_X1 U11019 ( .B1(n9773), .B2(n9813), .A(n9738), .ZN(n9739) );
  OAI21_X1 U11020 ( .B1(n9815), .B2(n9775), .A(n9739), .ZN(P1_U3546) );
  INV_X1 U11021 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9743) );
  AOI211_X1 U11022 ( .C1(n9767), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9816)
         );
  MUX2_X1 U11023 ( .A(n9743), .B(n9816), .S(n10106), .Z(n9744) );
  OAI21_X1 U11024 ( .B1(n9819), .B2(n9775), .A(n9744), .ZN(P1_U3545) );
  OAI211_X1 U11025 ( .C1(n9747), .C2(n10094), .A(n9746), .B(n9745), .ZN(n9820)
         );
  MUX2_X1 U11026 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9820), .S(n10106), .Z(
        n9748) );
  INV_X1 U11027 ( .A(n9748), .ZN(n9749) );
  OAI21_X1 U11028 ( .B1(n9823), .B2(n9775), .A(n9749), .ZN(P1_U3544) );
  AOI211_X1 U11029 ( .C1(n9767), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9753)
         );
  OAI21_X1 U11030 ( .B1(n9754), .B2(n9778), .A(n9753), .ZN(n9824) );
  MUX2_X1 U11031 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9824), .S(n10106), .Z(
        P1_U3543) );
  INV_X1 U11032 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9758) );
  AOI211_X1 U11033 ( .C1(n9757), .C2(n10096), .A(n9756), .B(n9755), .ZN(n9825)
         );
  MUX2_X1 U11034 ( .A(n9758), .B(n9825), .S(n10106), .Z(n9759) );
  OAI21_X1 U11035 ( .B1(n9828), .B2(n9789), .A(n9759), .ZN(P1_U3542) );
  OAI22_X1 U11036 ( .A1(n9830), .A2(n9775), .B1(n9829), .B2(n9789), .ZN(n9763)
         );
  NAND2_X1 U11037 ( .A1(n9761), .A2(n9760), .ZN(n9831) );
  MUX2_X1 U11038 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9831), .S(n10106), .Z(
        n9762) );
  OR2_X1 U11039 ( .A1(n9763), .A2(n9762), .ZN(P1_U3541) );
  INV_X1 U11040 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9768) );
  AOI211_X1 U11041 ( .C1(n9767), .C2(n9766), .A(n9765), .B(n9764), .ZN(n9834)
         );
  MUX2_X1 U11042 ( .A(n9768), .B(n9834), .S(n10106), .Z(n9769) );
  OAI21_X1 U11043 ( .B1(n9837), .B2(n9775), .A(n9769), .ZN(P1_U3540) );
  NAND2_X1 U11044 ( .A1(n9771), .A2(n9770), .ZN(n9838) );
  MUX2_X1 U11045 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9838), .S(n10106), .Z(
        n9772) );
  AOI21_X1 U11046 ( .B1(n9773), .B2(n9840), .A(n9772), .ZN(n9774) );
  OAI21_X1 U11047 ( .B1(n9843), .B2(n9775), .A(n9774), .ZN(P1_U3539) );
  OAI211_X1 U11048 ( .C1(n9779), .C2(n9778), .A(n9777), .B(n9776), .ZN(n9844)
         );
  INV_X1 U11049 ( .A(n9844), .ZN(n9780) );
  MUX2_X1 U11050 ( .A(n9781), .B(n9780), .S(n10106), .Z(n9782) );
  OAI21_X1 U11051 ( .B1(n9783), .B2(n9789), .A(n9782), .ZN(P1_U3538) );
  AOI211_X1 U11052 ( .C1(n9786), .C2(n10096), .A(n9785), .B(n9784), .ZN(n9849)
         );
  MUX2_X1 U11053 ( .A(n9787), .B(n9849), .S(n10106), .Z(n9788) );
  OAI21_X1 U11054 ( .B1(n4588), .B2(n9789), .A(n9788), .ZN(P1_U3536) );
  MUX2_X1 U11055 ( .A(n9791), .B(n9790), .S(n10100), .Z(n9792) );
  OAI21_X1 U11056 ( .B1(n9793), .B2(n9852), .A(n9792), .ZN(P1_U3521) );
  MUX2_X1 U11057 ( .A(n9795), .B(n9794), .S(n10100), .Z(n9796) );
  OAI21_X1 U11058 ( .B1(n9797), .B2(n9842), .A(n9796), .ZN(P1_U3518) );
  MUX2_X1 U11059 ( .A(n9799), .B(n9798), .S(n10100), .Z(n9800) );
  OAI21_X1 U11060 ( .B1(n9801), .B2(n9842), .A(n9800), .ZN(P1_U3517) );
  MUX2_X1 U11061 ( .A(n9803), .B(n9802), .S(n10100), .Z(n9804) );
  OAI21_X1 U11062 ( .B1(n9805), .B2(n9842), .A(n9804), .ZN(P1_U3516) );
  MUX2_X1 U11063 ( .A(n9806), .B(P1_REG0_REG_25__SCAN_IN), .S(n10098), .Z(
        n9807) );
  AOI21_X1 U11064 ( .B1(n9847), .B2(n9808), .A(n9807), .ZN(n9809) );
  OAI21_X1 U11065 ( .B1(n9810), .B2(n9842), .A(n9809), .ZN(P1_U3515) );
  MUX2_X1 U11066 ( .A(n9811), .B(P1_REG0_REG_24__SCAN_IN), .S(n10098), .Z(
        n9812) );
  AOI21_X1 U11067 ( .B1(n9847), .B2(n9813), .A(n9812), .ZN(n9814) );
  OAI21_X1 U11068 ( .B1(n9815), .B2(n9842), .A(n9814), .ZN(P1_U3514) );
  MUX2_X1 U11069 ( .A(n9817), .B(n9816), .S(n10100), .Z(n9818) );
  OAI21_X1 U11070 ( .B1(n9819), .B2(n9842), .A(n9818), .ZN(P1_U3513) );
  MUX2_X1 U11071 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9820), .S(n10100), .Z(
        n9821) );
  INV_X1 U11072 ( .A(n9821), .ZN(n9822) );
  OAI21_X1 U11073 ( .B1(n9823), .B2(n9842), .A(n9822), .ZN(P1_U3512) );
  MUX2_X1 U11074 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9824), .S(n10100), .Z(
        P1_U3511) );
  INV_X1 U11075 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9826) );
  MUX2_X1 U11076 ( .A(n9826), .B(n9825), .S(n10100), .Z(n9827) );
  OAI21_X1 U11077 ( .B1(n9828), .B2(n9852), .A(n9827), .ZN(P1_U3510) );
  OAI22_X1 U11078 ( .A1(n9830), .A2(n9842), .B1(n9829), .B2(n9852), .ZN(n9833)
         );
  MUX2_X1 U11079 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9831), .S(n10100), .Z(
        n9832) );
  OR2_X1 U11080 ( .A1(n9833), .A2(n9832), .ZN(P1_U3509) );
  MUX2_X1 U11081 ( .A(n9835), .B(n9834), .S(n10100), .Z(n9836) );
  OAI21_X1 U11082 ( .B1(n9837), .B2(n9842), .A(n9836), .ZN(P1_U3507) );
  MUX2_X1 U11083 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9838), .S(n10100), .Z(
        n9839) );
  AOI21_X1 U11084 ( .B1(n9847), .B2(n9840), .A(n9839), .ZN(n9841) );
  OAI21_X1 U11085 ( .B1(n9843), .B2(n9842), .A(n9841), .ZN(P1_U3504) );
  MUX2_X1 U11086 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9844), .S(n10100), .Z(
        n9845) );
  AOI21_X1 U11087 ( .B1(n9847), .B2(n9846), .A(n9845), .ZN(n9848) );
  INV_X1 U11088 ( .A(n9848), .ZN(P1_U3501) );
  MUX2_X1 U11089 ( .A(n9850), .B(n9849), .S(n10100), .Z(n9851) );
  OAI21_X1 U11090 ( .B1(n4588), .B2(n9852), .A(n9851), .ZN(P1_U3495) );
  AND2_X1 U11091 ( .A1(n9854), .A2(n9853), .ZN(n10077) );
  MUX2_X1 U11092 ( .A(P1_D_REG_1__SCAN_IN), .B(n9855), .S(n10077), .Z(P1_U3440) );
  MUX2_X1 U11093 ( .A(P1_D_REG_0__SCAN_IN), .B(n9856), .S(n10077), .Z(P1_U3439) );
  OR2_X1 U11094 ( .A1(n9857), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9861) );
  INV_X1 U11095 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9858) );
  NAND3_X1 U11096 ( .A1(n9858), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9860) );
  OAI22_X1 U11097 ( .A1(n9861), .A2(n9860), .B1(n9859), .B2(n9868), .ZN(n9862)
         );
  INV_X1 U11098 ( .A(n9862), .ZN(n9863) );
  OAI21_X1 U11099 ( .B1(n9864), .B2(n9872), .A(n9863), .ZN(P1_U3324) );
  OAI222_X1 U11100 ( .A1(n9868), .A2(n9867), .B1(n9872), .B2(n9866), .C1(
        P1_U3086), .C2(n9865), .ZN(P1_U3325) );
  OAI222_X1 U11101 ( .A1(n9872), .A2(n9871), .B1(n9870), .B2(P1_U3086), .C1(
        n9869), .C2(n9868), .ZN(P1_U3326) );
  INV_X1 U11102 ( .A(n9873), .ZN(n9874) );
  MUX2_X1 U11103 ( .A(n9874), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11104 ( .A(n9875), .ZN(n9876) );
  AOI21_X1 U11105 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(n9893) );
  INV_X1 U11106 ( .A(n9890), .ZN(n9880) );
  NAND3_X1 U11107 ( .A1(n9880), .A2(P2_U3893), .A3(n9887), .ZN(n9881) );
  AOI21_X1 U11108 ( .B1(n9881), .B2(n10185), .A(n9888), .ZN(n9884) );
  OAI21_X1 U11109 ( .B1(n10183), .B2(n10332), .A(n9882), .ZN(n9883) );
  AOI211_X1 U11110 ( .C1(n9886), .C2(n9885), .A(n9884), .B(n9883), .ZN(n9892)
         );
  INV_X1 U11111 ( .A(n9887), .ZN(n9889) );
  OAI211_X1 U11112 ( .C1(n9890), .C2(n9889), .A(n10167), .B(n9888), .ZN(n9891)
         );
  OAI211_X1 U11113 ( .C1(n9893), .C2(n10199), .A(n9892), .B(n9891), .ZN(
        P2_U3200) );
  INV_X1 U11114 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9905) );
  AOI211_X1 U11115 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n10028), .ZN(n9901)
         );
  INV_X1 U11116 ( .A(n10024), .ZN(n10010) );
  AOI211_X1 U11117 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n10010), .ZN(n9900)
         );
  AOI211_X1 U11118 ( .C1(n10031), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9904)
         );
  NAND2_X1 U11119 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9923) );
  OAI211_X1 U11120 ( .C1(n9905), .C2(n10039), .A(n9904), .B(n9923), .ZN(
        P1_U3253) );
  INV_X1 U11121 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9919) );
  INV_X1 U11122 ( .A(n9906), .ZN(n9909) );
  AOI211_X1 U11123 ( .C1(n9909), .C2(n9908), .A(n9907), .B(n10028), .ZN(n9915)
         );
  INV_X1 U11124 ( .A(n9910), .ZN(n9913) );
  AOI211_X1 U11125 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n10010), .ZN(n9914)
         );
  AOI211_X1 U11126 ( .C1(n10031), .C2(n9916), .A(n9915), .B(n9914), .ZN(n9918)
         );
  OAI211_X1 U11127 ( .C1(n9919), .C2(n10039), .A(n9918), .B(n9917), .ZN(
        P1_U3251) );
  OAI21_X1 U11128 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9932) );
  INV_X1 U11129 ( .A(n9923), .ZN(n9924) );
  AOI21_X1 U11130 ( .B1(n9926), .B2(n9925), .A(n9924), .ZN(n9927) );
  OAI21_X1 U11131 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  AOI21_X1 U11132 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9933) );
  OAI21_X1 U11133 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(P1_U3217) );
  OAI21_X1 U11134 ( .B1(n9937), .B2(n10094), .A(n9936), .ZN(n9938) );
  AOI21_X1 U11135 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n9943) );
  AOI22_X1 U11136 ( .A1(n10106), .A2(n9943), .B1(n9941), .B2(n4826), .ZN(
        P1_U3552) );
  AOI22_X1 U11137 ( .A1(n10100), .A2(n9943), .B1(n9942), .B2(n10098), .ZN(
        P1_U3520) );
  XNOR2_X1 U11138 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11139 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11140 ( .B1(n4416), .B2(n9945), .A(n9944), .ZN(n9947) );
  XNOR2_X1 U11141 ( .A(n9947), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U11142 ( .A1(n9948), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9949) );
  OAI21_X1 U11143 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(P1_U3243) );
  AOI211_X1 U11144 ( .C1(n9954), .C2(n9953), .A(n9952), .B(n10028), .ZN(n9959)
         );
  AOI211_X1 U11145 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n10010), .ZN(n9958)
         );
  AOI211_X1 U11146 ( .C1(n10031), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9962)
         );
  NAND2_X1 U11147 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9961) );
  OAI211_X1 U11148 ( .C1(n9963), .C2(n10039), .A(n9962), .B(n9961), .ZN(
        P1_U3254) );
  NAND2_X1 U11149 ( .A1(n9965), .A2(n9964), .ZN(n9968) );
  INV_X1 U11150 ( .A(n9966), .ZN(n9967) );
  NAND2_X1 U11151 ( .A1(n9968), .A2(n9967), .ZN(n9976) );
  NAND2_X1 U11152 ( .A1(n10031), .A2(n9969), .ZN(n9975) );
  AOI21_X1 U11153 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(n9973) );
  NAND2_X1 U11154 ( .A1(n10024), .A2(n9973), .ZN(n9974) );
  OAI211_X1 U11155 ( .C1(n10028), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9977)
         );
  INV_X1 U11156 ( .A(n9977), .ZN(n9979) );
  NAND2_X1 U11157 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9978) );
  OAI211_X1 U11158 ( .C1(n9980), .C2(n10039), .A(n9979), .B(n9978), .ZN(
        P1_U3256) );
  NAND2_X1 U11159 ( .A1(n9982), .A2(n9981), .ZN(n9985) );
  INV_X1 U11160 ( .A(n9983), .ZN(n9984) );
  NAND2_X1 U11161 ( .A1(n9985), .A2(n9984), .ZN(n9993) );
  NAND2_X1 U11162 ( .A1(n10031), .A2(n9986), .ZN(n9992) );
  AOI21_X1 U11163 ( .B1(n9989), .B2(n9988), .A(n9987), .ZN(n9990) );
  NAND2_X1 U11164 ( .A1(n10024), .A2(n9990), .ZN(n9991) );
  OAI211_X1 U11165 ( .C1(n10028), .C2(n9993), .A(n9992), .B(n9991), .ZN(n9994)
         );
  INV_X1 U11166 ( .A(n9994), .ZN(n9996) );
  NAND2_X1 U11167 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9995) );
  OAI211_X1 U11168 ( .C1(n9997), .C2(n10039), .A(n9996), .B(n9995), .ZN(
        P1_U3257) );
  AOI211_X1 U11169 ( .C1(n10000), .C2(n9999), .A(n9998), .B(n10028), .ZN(
        n10005) );
  AOI211_X1 U11170 ( .C1(n10003), .C2(n10002), .A(n10001), .B(n10010), .ZN(
        n10004) );
  AOI211_X1 U11171 ( .C1(n10031), .C2(n10006), .A(n10005), .B(n10004), .ZN(
        n10008) );
  NAND2_X1 U11172 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n10007)
         );
  OAI211_X1 U11173 ( .C1(n10009), .C2(n10039), .A(n10008), .B(n10007), .ZN(
        P1_U3258) );
  AOI21_X1 U11174 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(n10020) );
  XOR2_X1 U11175 ( .A(n10014), .B(n10013), .Z(n10017) );
  OAI22_X1 U11176 ( .A1(n10017), .A2(n10028), .B1(n10016), .B2(n10015), .ZN(
        n10018) );
  AOI21_X1 U11177 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10022) );
  NAND2_X1 U11178 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n10021)
         );
  OAI211_X1 U11179 ( .C1(n10023), .C2(n10039), .A(n10022), .B(n10021), .ZN(
        P1_U3259) );
  OAI211_X1 U11180 ( .C1(n10027), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        n10036) );
  AOI21_X1 U11181 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10034) );
  AOI22_X1 U11182 ( .A1(n10034), .A2(n10033), .B1(n10032), .B2(n10031), .ZN(
        n10035) );
  AND2_X1 U11183 ( .A1(n10036), .A2(n10035), .ZN(n10038) );
  NAND2_X1 U11184 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n10037)
         );
  OAI211_X1 U11185 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        P1_U3261) );
  INV_X1 U11186 ( .A(n10041), .ZN(n10050) );
  OAI22_X1 U11187 ( .A1(n10067), .A2(n10044), .B1(n10043), .B2(n10042), .ZN(
        n10045) );
  AOI21_X1 U11188 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(n10048) );
  OAI21_X1 U11189 ( .B1(n10050), .B2(n10049), .A(n10048), .ZN(n10051) );
  AOI21_X1 U11190 ( .B1(n10053), .B2(n10052), .A(n10051), .ZN(n10054) );
  OAI21_X1 U11191 ( .B1(n9581), .B2(n10055), .A(n10054), .ZN(P1_U3289) );
  INV_X1 U11192 ( .A(n10056), .ZN(n10059) );
  AOI21_X1 U11193 ( .B1(n10059), .B2(n10058), .A(n10057), .ZN(n10068) );
  INV_X1 U11194 ( .A(n10060), .ZN(n10063) );
  AOI21_X1 U11195 ( .B1(n10063), .B2(n10062), .A(n10061), .ZN(n10064) );
  AOI21_X1 U11196 ( .B1(n10065), .B2(P1_REG3_REG_0__SCAN_IN), .A(n10064), .ZN(
        n10066) );
  OAI221_X1 U11197 ( .B1(n9581), .B2(n10068), .C1(n10067), .C2(n5726), .A(
        n10066), .ZN(P1_U3293) );
  AND2_X1 U11198 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10078), .ZN(P1_U3294) );
  AND2_X1 U11199 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10078), .ZN(P1_U3295) );
  AND2_X1 U11200 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10078), .ZN(P1_U3296) );
  AND2_X1 U11201 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10078), .ZN(P1_U3297) );
  AND2_X1 U11202 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10078), .ZN(P1_U3298) );
  NOR2_X1 U11203 ( .A1(n10077), .A2(n10069), .ZN(P1_U3299) );
  AND2_X1 U11204 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10078), .ZN(P1_U3300) );
  AND2_X1 U11205 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10078), .ZN(P1_U3301) );
  AND2_X1 U11206 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10078), .ZN(P1_U3302) );
  NOR2_X1 U11207 ( .A1(n10077), .A2(n10070), .ZN(P1_U3303) );
  AND2_X1 U11208 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10078), .ZN(P1_U3304) );
  AND2_X1 U11209 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10078), .ZN(P1_U3305) );
  AND2_X1 U11210 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10078), .ZN(P1_U3306) );
  AND2_X1 U11211 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10078), .ZN(P1_U3307) );
  NOR2_X1 U11212 ( .A1(n10077), .A2(n10071), .ZN(P1_U3308) );
  AND2_X1 U11213 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10078), .ZN(P1_U3309) );
  AND2_X1 U11214 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10078), .ZN(P1_U3310) );
  NOR2_X1 U11215 ( .A1(n10077), .A2(n10072), .ZN(P1_U3311) );
  AND2_X1 U11216 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10078), .ZN(P1_U3312) );
  NOR2_X1 U11217 ( .A1(n10077), .A2(n10073), .ZN(P1_U3313) );
  AND2_X1 U11218 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10078), .ZN(P1_U3314) );
  AND2_X1 U11219 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10078), .ZN(P1_U3315) );
  AND2_X1 U11220 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10078), .ZN(P1_U3316) );
  AND2_X1 U11221 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10078), .ZN(P1_U3317) );
  NOR2_X1 U11222 ( .A1(n10077), .A2(n10074), .ZN(P1_U3318) );
  AND2_X1 U11223 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10078), .ZN(P1_U3319) );
  NOR2_X1 U11224 ( .A1(n10077), .A2(n10075), .ZN(P1_U3320) );
  AND2_X1 U11225 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10078), .ZN(P1_U3321) );
  NOR2_X1 U11226 ( .A1(n10077), .A2(n10076), .ZN(P1_U3322) );
  AND2_X1 U11227 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10078), .ZN(P1_U3323) );
  OAI21_X1 U11228 ( .B1(n10080), .B2(n10094), .A(n10079), .ZN(n10081) );
  AOI21_X1 U11229 ( .B1(n10083), .B2(n10082), .A(n10081), .ZN(n10084) );
  AND2_X1 U11230 ( .A1(n10085), .A2(n10084), .ZN(n10102) );
  AOI22_X1 U11231 ( .A1(n10100), .A2(n10102), .B1(n5927), .B2(n10098), .ZN(
        P1_U3456) );
  OAI21_X1 U11232 ( .B1(n10087), .B2(n10094), .A(n10086), .ZN(n10088) );
  AOI211_X1 U11233 ( .C1(n10090), .C2(n10096), .A(n10089), .B(n10088), .ZN(
        n10103) );
  AOI22_X1 U11234 ( .A1(n10100), .A2(n10103), .B1(n6304), .B2(n10098), .ZN(
        P1_U3474) );
  OAI211_X1 U11235 ( .C1(n4591), .C2(n10094), .A(n10093), .B(n10092), .ZN(
        n10095) );
  AOI21_X1 U11236 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10105) );
  AOI22_X1 U11237 ( .A1(n10100), .A2(n10105), .B1(n10099), .B2(n10098), .ZN(
        P1_U3480) );
  AOI22_X1 U11238 ( .A1(n10106), .A2(n10102), .B1(n10101), .B2(n4826), .ZN(
        P1_U3523) );
  AOI22_X1 U11239 ( .A1(n10106), .A2(n10103), .B1(n6308), .B2(n4826), .ZN(
        P1_U3529) );
  AOI22_X1 U11240 ( .A1(n10106), .A2(n10105), .B1(n10104), .B2(n4826), .ZN(
        P1_U3531) );
  AOI22_X1 U11241 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10175), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10111) );
  XNOR2_X1 U11242 ( .A(n10107), .B(P2_IR_REG_0__SCAN_IN), .ZN(n10108) );
  OAI21_X1 U11243 ( .B1(n10167), .B2(n10109), .A(n10108), .ZN(n10110) );
  OAI211_X1 U11244 ( .C1(n10185), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        P2_U3182) );
  AOI21_X1 U11245 ( .B1(n10115), .B2(n10114), .A(n10113), .ZN(n10117) );
  OAI22_X1 U11246 ( .A1(n10191), .A2(n10117), .B1(n10185), .B2(n10116), .ZN(
        n10122) );
  AOI211_X1 U11247 ( .C1(n10120), .C2(n10119), .A(n10193), .B(n10118), .ZN(
        n10121) );
  AOI211_X1 U11248 ( .C1(n10175), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10122), .B(
        n10121), .ZN(n10131) );
  INV_X1 U11249 ( .A(n10123), .ZN(n10126) );
  INV_X1 U11250 ( .A(n10124), .ZN(n10125) );
  AND2_X1 U11251 ( .A1(n10126), .A2(n10125), .ZN(n10128) );
  OAI21_X1 U11252 ( .B1(n10129), .B2(n10128), .A(n10127), .ZN(n10130) );
  OAI211_X1 U11253 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6190), .A(n10131), .B(
        n10130), .ZN(P2_U3184) );
  AOI21_X1 U11254 ( .B1(n10305), .B2(n10133), .A(n10132), .ZN(n10146) );
  OAI21_X1 U11255 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(n10137) );
  AND2_X1 U11256 ( .A1(n10137), .A2(n10167), .ZN(n10143) );
  AOI21_X1 U11257 ( .B1(n10139), .B2(n10215), .A(n10138), .ZN(n10141) );
  OAI22_X1 U11258 ( .A1(n10191), .A2(n10141), .B1(n10185), .B2(n10140), .ZN(
        n10142) );
  AOI211_X1 U11259 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10175), .A(n10143), .B(
        n10142), .ZN(n10145) );
  OAI211_X1 U11260 ( .C1(n10146), .C2(n10199), .A(n10145), .B(n10144), .ZN(
        P2_U3185) );
  AOI21_X1 U11261 ( .B1(n4507), .B2(n10148), .A(n10147), .ZN(n10161) );
  OAI21_X1 U11262 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10152) );
  AND2_X1 U11263 ( .A1(n10152), .A2(n10167), .ZN(n10158) );
  AOI21_X1 U11264 ( .B1(n4508), .B2(n10154), .A(n10153), .ZN(n10156) );
  OAI22_X1 U11265 ( .A1(n10156), .A2(n10191), .B1(n10185), .B2(n10155), .ZN(
        n10157) );
  AOI211_X1 U11266 ( .C1(P2_ADDR_REG_6__SCAN_IN), .C2(n10175), .A(n10158), .B(
        n10157), .ZN(n10160) );
  OAI211_X1 U11267 ( .C1(n10161), .C2(n10199), .A(n10160), .B(n10159), .ZN(
        P2_U3188) );
  AOI21_X1 U11268 ( .B1(n4506), .B2(n10163), .A(n10162), .ZN(n10179) );
  OAI21_X1 U11269 ( .B1(n10166), .B2(n10165), .A(n10164), .ZN(n10168) );
  AND2_X1 U11270 ( .A1(n10168), .A2(n10167), .ZN(n10174) );
  AOI21_X1 U11271 ( .B1(n4501), .B2(n10170), .A(n10169), .ZN(n10172) );
  OAI22_X1 U11272 ( .A1(n10172), .A2(n10191), .B1(n10185), .B2(n10171), .ZN(
        n10173) );
  AOI211_X1 U11273 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10175), .A(n10174), .B(
        n10173), .ZN(n10178) );
  INV_X1 U11274 ( .A(n10176), .ZN(n10177) );
  OAI211_X1 U11275 ( .C1(n10179), .C2(n10199), .A(n10178), .B(n10177), .ZN(
        P2_U3190) );
  AOI21_X1 U11276 ( .B1(n4505), .B2(n10181), .A(n10180), .ZN(n10200) );
  INV_X1 U11277 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10182) );
  OAI22_X1 U11278 ( .A1(n10185), .A2(n10184), .B1(n10183), .B2(n10182), .ZN(
        n10196) );
  AOI21_X1 U11279 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(n10194) );
  AOI21_X1 U11280 ( .B1(n4502), .B2(n10190), .A(n10189), .ZN(n10192) );
  OAI22_X1 U11281 ( .A1(n10194), .A2(n10193), .B1(n10192), .B2(n10191), .ZN(
        n10195) );
  NOR3_X1 U11282 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n10198) );
  OAI21_X1 U11283 ( .B1(n10200), .B2(n10199), .A(n10198), .ZN(P2_U3192) );
  XOR2_X1 U11284 ( .A(n10201), .B(n10208), .Z(n10206) );
  AOI222_X1 U11285 ( .A1(n10207), .A2(n10206), .B1(n10205), .B2(n10204), .C1(
        n10203), .C2(n10202), .ZN(n10246) );
  XNOR2_X1 U11286 ( .A(n10209), .B(n10208), .ZN(n10244) );
  AOI222_X1 U11287 ( .A1(n10244), .A2(n10213), .B1(n10212), .B2(n10211), .C1(
        n10243), .C2(n10210), .ZN(n10214) );
  OAI221_X1 U11288 ( .B1(n10235), .B2(n10246), .C1(n8601), .C2(n10215), .A(
        n10214), .ZN(P2_U3230) );
  XNOR2_X1 U11289 ( .A(n10216), .B(n10224), .ZN(n10239) );
  OAI22_X1 U11290 ( .A1(n10219), .A2(n10218), .B1(n6190), .B2(n10217), .ZN(
        n10232) );
  OAI22_X1 U11291 ( .A1(n10222), .A2(n10221), .B1(n6061), .B2(n10220), .ZN(
        n10229) );
  NAND3_X1 U11292 ( .A1(n6195), .A2(n10224), .A3(n10223), .ZN(n10226) );
  AOI21_X1 U11293 ( .B1(n10227), .B2(n10226), .A(n10225), .ZN(n10228) );
  AOI211_X1 U11294 ( .C1(n10239), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10241) );
  INV_X1 U11295 ( .A(n10241), .ZN(n10231) );
  AOI211_X1 U11296 ( .C1(n10233), .C2(n10239), .A(n10232), .B(n10231), .ZN(
        n10234) );
  AOI22_X1 U11297 ( .A1(n10235), .A2(n6374), .B1(n10234), .B2(n8601), .ZN(
        P2_U3231) );
  INV_X1 U11298 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U11299 ( .A1(n10302), .A2(n10237), .B1(n10236), .B2(n10300), .ZN(
        P2_U3393) );
  INV_X1 U11300 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11301 ( .A1(n10239), .A2(n10255), .B1(n10299), .B2(n10238), .ZN(
        n10240) );
  AND2_X1 U11302 ( .A1(n10241), .A2(n10240), .ZN(n10304) );
  AOI22_X1 U11303 ( .A1(n10302), .A2(n10242), .B1(n10304), .B2(n10300), .ZN(
        P2_U3396) );
  AOI22_X1 U11304 ( .A1(n10244), .A2(n10275), .B1(n10299), .B2(n10243), .ZN(
        n10245) );
  AND2_X1 U11305 ( .A1(n10246), .A2(n10245), .ZN(n10306) );
  AOI22_X1 U11306 ( .A1(n10302), .A2(n10247), .B1(n10306), .B2(n10300), .ZN(
        P2_U3399) );
  INV_X1 U11307 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10253) );
  OR2_X1 U11308 ( .A1(n10248), .A2(n10294), .ZN(n10251) );
  NAND2_X1 U11309 ( .A1(n10249), .A2(n10299), .ZN(n10250) );
  AND3_X1 U11310 ( .A1(n10252), .A2(n10251), .A3(n10250), .ZN(n10308) );
  AOI22_X1 U11311 ( .A1(n10302), .A2(n10253), .B1(n10308), .B2(n10300), .ZN(
        P2_U3402) );
  INV_X1 U11312 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U11313 ( .A1(n10256), .A2(n10255), .B1(n10299), .B2(n10254), .ZN(
        n10257) );
  AND2_X1 U11314 ( .A1(n10258), .A2(n10257), .ZN(n10310) );
  AOI22_X1 U11315 ( .A1(n10302), .A2(n10259), .B1(n10310), .B2(n10300), .ZN(
        P2_U3405) );
  INV_X1 U11316 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11317 ( .A1(n10261), .A2(n10275), .B1(n10299), .B2(n10260), .ZN(
        n10262) );
  AND2_X1 U11318 ( .A1(n10263), .A2(n10262), .ZN(n10312) );
  AOI22_X1 U11319 ( .A1(n10302), .A2(n10264), .B1(n10312), .B2(n10300), .ZN(
        P2_U3408) );
  INV_X1 U11320 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10269) );
  OAI22_X1 U11321 ( .A1(n10266), .A2(n10284), .B1(n10265), .B2(n10282), .ZN(
        n10267) );
  NOR2_X1 U11322 ( .A1(n10268), .A2(n10267), .ZN(n10314) );
  AOI22_X1 U11323 ( .A1(n10302), .A2(n10269), .B1(n10314), .B2(n10300), .ZN(
        P2_U3411) );
  INV_X1 U11324 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10276) );
  INV_X1 U11325 ( .A(n10270), .ZN(n10274) );
  OAI21_X1 U11326 ( .B1(n10272), .B2(n10282), .A(n10271), .ZN(n10273) );
  AOI21_X1 U11327 ( .B1(n10275), .B2(n10274), .A(n10273), .ZN(n10316) );
  AOI22_X1 U11328 ( .A1(n10302), .A2(n10276), .B1(n10316), .B2(n10300), .ZN(
        P2_U3414) );
  OAI22_X1 U11329 ( .A1(n10278), .A2(n10284), .B1(n10277), .B2(n10282), .ZN(
        n10279) );
  NOR2_X1 U11330 ( .A1(n10280), .A2(n10279), .ZN(n10318) );
  AOI22_X1 U11331 ( .A1(n10302), .A2(n10281), .B1(n10318), .B2(n10300), .ZN(
        P2_U3417) );
  INV_X1 U11332 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10288) );
  OAI22_X1 U11333 ( .A1(n10285), .A2(n10284), .B1(n10283), .B2(n10282), .ZN(
        n10286) );
  NOR2_X1 U11334 ( .A1(n10287), .A2(n10286), .ZN(n10320) );
  AOI22_X1 U11335 ( .A1(n10302), .A2(n10288), .B1(n10320), .B2(n10300), .ZN(
        P2_U3420) );
  INV_X1 U11336 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10293) );
  NOR2_X1 U11337 ( .A1(n10289), .A2(n10294), .ZN(n10291) );
  AOI211_X1 U11338 ( .C1(n10299), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10322) );
  AOI22_X1 U11339 ( .A1(n10302), .A2(n10293), .B1(n10322), .B2(n10300), .ZN(
        P2_U3423) );
  INV_X1 U11340 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10301) );
  NOR2_X1 U11341 ( .A1(n10295), .A2(n10294), .ZN(n10297) );
  AOI211_X1 U11342 ( .C1(n10299), .C2(n10298), .A(n10297), .B(n10296), .ZN(
        n10324) );
  AOI22_X1 U11343 ( .A1(n10302), .A2(n10301), .B1(n10324), .B2(n10300), .ZN(
        P2_U3426) );
  INV_X1 U11344 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U11345 ( .A1(n10325), .A2(n10304), .B1(n10303), .B2(n10323), .ZN(
        P2_U3461) );
  AOI22_X1 U11346 ( .A1(n10325), .A2(n10306), .B1(n10305), .B2(n10323), .ZN(
        P2_U3462) );
  INV_X1 U11347 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U11348 ( .A1(n10325), .A2(n10308), .B1(n10307), .B2(n10323), .ZN(
        P2_U3463) );
  AOI22_X1 U11349 ( .A1(n10325), .A2(n10310), .B1(n10309), .B2(n10323), .ZN(
        P2_U3464) );
  AOI22_X1 U11350 ( .A1(n10325), .A2(n10312), .B1(n10311), .B2(n10323), .ZN(
        P2_U3465) );
  AOI22_X1 U11351 ( .A1(n10325), .A2(n10314), .B1(n10313), .B2(n10323), .ZN(
        P2_U3466) );
  AOI22_X1 U11352 ( .A1(n10325), .A2(n10316), .B1(n10315), .B2(n10323), .ZN(
        P2_U3467) );
  AOI22_X1 U11353 ( .A1(n10325), .A2(n10318), .B1(n10317), .B2(n10323), .ZN(
        P2_U3468) );
  AOI22_X1 U11354 ( .A1(n10325), .A2(n10320), .B1(n10319), .B2(n10323), .ZN(
        P2_U3469) );
  AOI22_X1 U11355 ( .A1(n10325), .A2(n10322), .B1(n10321), .B2(n10323), .ZN(
        P2_U3470) );
  AOI22_X1 U11356 ( .A1(n10325), .A2(n10324), .B1(n7337), .B2(n10323), .ZN(
        P2_U3471) );
  NOR2_X1 U11357 ( .A1(n10327), .A2(n10326), .ZN(n10329) );
  XNOR2_X1 U11358 ( .A(n10329), .B(n10328), .ZN(ADD_1068_U5) );
  XOR2_X1 U11359 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  AOI21_X1 U11360 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10331), .A(n10330), 
        .ZN(n10333) );
  XNOR2_X1 U11361 ( .A(n10333), .B(n10332), .ZN(ADD_1068_U55) );
  XNOR2_X1 U11362 ( .A(n10335), .B(n10334), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11363 ( .A(n10337), .B(n10336), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11364 ( .A(n10339), .B(n10338), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11365 ( .A(n10341), .B(n10340), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11366 ( .A(n10343), .B(n10342), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11367 ( .A(n10345), .B(n10344), .ZN(ADD_1068_U61) );
  XOR2_X1 U11368 ( .A(n10347), .B(n10346), .Z(ADD_1068_U62) );
  XOR2_X1 U11369 ( .A(n10349), .B(n10348), .Z(ADD_1068_U63) );
  NOR2_X1 U11370 ( .A1(n10351), .A2(n10350), .ZN(n10352) );
  XOR2_X1 U11371 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10352), .Z(ADD_1068_U51) );
  XOR2_X1 U11372 ( .A(n10353), .B(P2_ADDR_REG_9__SCAN_IN), .Z(ADD_1068_U47) );
  XOR2_X1 U11373 ( .A(n10354), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11374 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10355), .Z(ADD_1068_U48) );
  XOR2_X1 U11375 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10356), .Z(ADD_1068_U50) );
  XOR2_X1 U11376 ( .A(n10358), .B(n10357), .Z(ADD_1068_U54) );
  XOR2_X1 U11377 ( .A(n10360), .B(n10359), .Z(ADD_1068_U53) );
  XNOR2_X1 U11378 ( .A(n10362), .B(n10361), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4928 ( .A(n5187), .Z(n5200) );
  CLKBUF_X1 U4932 ( .A(n5256), .Z(n5447) );
  CLKBUF_X1 U4935 ( .A(n7932), .Z(n4415) );
  CLKBUF_X1 U5143 ( .A(n5189), .Z(n5209) );
endmodule

