

module b14_C_SARLock_k_64_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713;

  CLKBUF_X2 U2275 ( .A(n2359), .Z(n3851) );
  INV_X1 U2277 ( .A(n2700), .ZN(n2761) );
  CLKBUF_X2 U2278 ( .A(n2295), .Z(n2577) );
  INV_X1 U2279 ( .A(n2761), .ZN(n2861) );
  INV_X2 U2280 ( .A(n3856), .ZN(n3857) );
  BUF_X1 U2281 ( .A(n2294), .Z(n3852) );
  AND2_X1 U2282 ( .A1(n2677), .A2(n2963), .ZN(n4693) );
  NOR2_X2 U2283 ( .A1(n2496), .A2(IR_REG_17__SCAN_IN), .ZN(n2508) );
  AND2_X4 U2284 ( .A1(n2682), .A2(n2683), .ZN(n2762) );
  INV_X2 U2285 ( .A(n2763), .ZN(n2856) );
  OAI22_X2 U2286 ( .A1(n3211), .A2(n2397), .B1(n3343), .B2(n3962), .ZN(n3350)
         );
  OAI21_X2 U2287 ( .B1(n3242), .B2(n2169), .A(n2167), .ZN(n3211) );
  NOR2_X1 U2288 ( .A1(n3007), .A2(n3009), .ZN(n3008) );
  OAI21_X2 U2289 ( .B1(n3408), .B2(n3409), .A(n3410), .ZN(n2765) );
  MUX2_X1 U2290 ( .A(REG1_REG_29__SCAN_IN), .B(n2680), .S(n4713), .Z(n2675) );
  NAND2_X1 U2291 ( .A1(n3200), .A2(n2072), .ZN(n2186) );
  AOI21_X1 U2292 ( .B1(n2696), .B2(n2700), .A(n2699), .ZN(n2702) );
  AND2_X1 U2293 ( .A1(n3180), .A2(n2303), .ZN(n3077) );
  INV_X1 U2294 ( .A(n2865), .ZN(n2697) );
  INV_X1 U2295 ( .A(n4102), .ZN(n3256) );
  NOR2_X1 U2296 ( .A1(n2651), .A2(n2650), .ZN(n2924) );
  XNOR2_X1 U2297 ( .A(n2269), .B(IR_REG_29__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U2298 ( .A1(n2291), .A2(n2309), .ZN(n2317) );
  INV_X2 U2299 ( .A(IR_REG_31__SCAN_IN), .ZN(n2649) );
  OR2_X1 U2300 ( .A1(n2905), .A2(n2876), .ZN(n2907) );
  NAND2_X1 U2301 ( .A1(n2799), .A2(n2798), .ZN(n3704) );
  OAI21_X1 U2302 ( .B1(n4207), .B2(n4214), .A(n2244), .ZN(n2584) );
  NAND2_X1 U2303 ( .A1(n2075), .A2(n2199), .ZN(n2785) );
  NAND2_X1 U2304 ( .A1(n2161), .A2(n2159), .ZN(n2247) );
  NAND2_X1 U2305 ( .A1(n4576), .A2(n3314), .ZN(n4581) );
  AOI22_X1 U2306 ( .A1(n2184), .A2(n2192), .B1(n2189), .B2(n2037), .ZN(n2183)
         );
  OR2_X1 U2307 ( .A1(n2064), .A2(n2185), .ZN(n2037) );
  OR2_X1 U2308 ( .A1(n3063), .A2(n3062), .ZN(n3312) );
  NOR2_X1 U2309 ( .A1(n3262), .A2(n2188), .ZN(n2184) );
  AND2_X2 U2310 ( .A1(n3166), .A2(n4634), .ZN(n4664) );
  NOR2_X1 U2311 ( .A1(n2690), .A2(n2689), .ZN(n3007) );
  NAND4_X1 U2312 ( .A1(n2339), .A2(n2338), .A3(n2337), .A4(n2336), .ZN(n4102)
         );
  NAND4_X2 U2313 ( .A1(n2325), .A2(n2324), .A3(n2323), .A4(n2322), .ZN(n4103)
         );
  INV_X1 U2314 ( .A(n2725), .ZN(n3694) );
  INV_X1 U2315 ( .A(n4190), .ZN(n4196) );
  NAND4_X2 U2316 ( .A1(n2308), .A2(n2307), .A3(n2306), .A4(n2305), .ZN(n3182)
         );
  OR2_X1 U2317 ( .A1(n2641), .A2(n2640), .ZN(n2919) );
  INV_X1 U2318 ( .A(n2927), .ZN(n2032) );
  NAND2_X1 U2319 ( .A1(n3620), .A2(IR_REG_31__SCAN_IN), .ZN(n2268) );
  NAND4_X1 U2320 ( .A1(n2391), .A2(n2257), .A3(n2256), .A4(n2255), .ZN(n2258)
         );
  NOR2_X1 U2321 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2257)
         );
  NOR2_X1 U2322 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2256)
         );
  NOR2_X1 U2323 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2255)
         );
  INV_X1 U2324 ( .A(IR_REG_3__SCAN_IN), .ZN(n2326) );
  INV_X1 U2325 ( .A(IR_REG_4__SCAN_IN), .ZN(n2329) );
  INV_X4 U2326 ( .A(n2762), .ZN(n2763) );
  INV_X1 U2327 ( .A(n2297), .ZN(n2350) );
  CLKBUF_X1 U2328 ( .A(n2296), .Z(n2359) );
  NAND2_X1 U2329 ( .A1(n2036), .A2(n3724), .ZN(n2180) );
  AND3_X1 U2330 ( .A1(n2081), .A2(n2083), .A3(n2062), .ZN(n3054) );
  AND2_X1 U2331 ( .A1(n3879), .A2(n2407), .ZN(n2156) );
  OR2_X1 U2332 ( .A1(n2696), .A2(n3185), .ZN(n3794) );
  AND2_X1 U2333 ( .A1(n2236), .A2(n2266), .ZN(n2235) );
  NOR2_X1 U2334 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2259)
         );
  NAND2_X1 U2335 ( .A1(n2625), .A2(IR_REG_28__SCAN_IN), .ZN(n2277) );
  OR2_X1 U2336 ( .A1(n2930), .A2(n2927), .ZN(n2294) );
  OR2_X1 U2337 ( .A1(n2294), .A2(n2286), .ZN(n2287) );
  NAND2_X1 U2338 ( .A1(n2930), .A2(n2927), .ZN(n2295) );
  NOR2_X1 U2339 ( .A1(n2930), .A2(n2032), .ZN(n2296) );
  AND2_X1 U2340 ( .A1(n2930), .A2(n2032), .ZN(n2297) );
  NAND2_X1 U2341 ( .A1(n4581), .A2(n4582), .ZN(n4580) );
  XNOR2_X1 U2342 ( .A(n3333), .B(n2176), .ZN(n4594) );
  AOI21_X1 U2343 ( .B1(n2565), .B2(n2173), .A(n2566), .ZN(n4207) );
  AND2_X1 U2344 ( .A1(n4412), .A2(n4418), .ZN(n2566) );
  NAND2_X1 U2345 ( .A1(n4430), .A2(n4231), .ZN(n2173) );
  AND2_X1 U2346 ( .A1(n2559), .A2(REG3_REG_27__SCAN_IN), .ZN(n2567) );
  NOR2_X1 U2347 ( .A1(n2548), .A2(n2280), .ZN(n2557) );
  OR2_X1 U2348 ( .A1(n2540), .A2(n3642), .ZN(n2546) );
  OR2_X1 U2349 ( .A1(n3380), .A2(n2439), .ZN(n2441) );
  NAND2_X1 U2350 ( .A1(n2157), .A2(n2156), .ZN(n3417) );
  AND2_X1 U2351 ( .A1(n2684), .A2(n2897), .ZN(n2963) );
  AOI22_X1 U2352 ( .A1(n2634), .A2(n4329), .B1(n4202), .B2(n3954), .ZN(n3623)
         );
  AOI21_X1 U2353 ( .B1(n4215), .B2(n2621), .A(n3850), .ZN(n2622) );
  AND2_X1 U2354 ( .A1(n2263), .A2(n2264), .ZN(n2234) );
  INV_X1 U2355 ( .A(IR_REG_21__SCAN_IN), .ZN(n2264) );
  AND2_X1 U2356 ( .A1(n3015), .A2(n3014), .ZN(n3047) );
  NAND2_X1 U2357 ( .A1(n2233), .A2(n2232), .ZN(n2231) );
  INV_X1 U2358 ( .A(n3752), .ZN(n2232) );
  INV_X1 U2359 ( .A(n3753), .ZN(n2233) );
  AOI21_X1 U2360 ( .B1(n2034), .B2(n2202), .A(n2200), .ZN(n2199) );
  NAND2_X1 U2361 ( .A1(n2774), .A2(n2034), .ZN(n2075) );
  INV_X1 U2362 ( .A(n3596), .ZN(n2200) );
  INV_X1 U2363 ( .A(IR_REG_19__SCAN_IN), .ZN(n2585) );
  OAI21_X1 U2364 ( .B1(n2983), .B2(n2051), .A(n2104), .ZN(n2985) );
  AND2_X1 U2365 ( .A1(n2107), .A2(n2977), .ZN(n2105) );
  NAND2_X1 U2366 ( .A1(n3055), .A2(n4559), .ZN(n2099) );
  NOR2_X1 U2367 ( .A1(n3866), .A2(n3886), .ZN(n2127) );
  AND2_X1 U2368 ( .A1(n4353), .A2(n2607), .ZN(n2608) );
  INV_X1 U2369 ( .A(n2462), .ZN(n2166) );
  AOI21_X1 U2370 ( .B1(n3210), .B2(n3816), .A(n2125), .ZN(n2124) );
  INV_X1 U2371 ( .A(n3821), .ZN(n2125) );
  NAND2_X1 U2372 ( .A1(n2382), .A2(n2170), .ZN(n2169) );
  INV_X1 U2373 ( .A(n3807), .ZN(n2135) );
  INV_X1 U2374 ( .A(n3803), .ZN(n2131) );
  NOR2_X1 U2375 ( .A1(n2145), .A2(n2146), .ZN(n2144) );
  NAND2_X1 U2376 ( .A1(n3367), .A2(n2597), .ZN(n2146) );
  AND2_X1 U2377 ( .A1(n3950), .A2(n3941), .ZN(n2942) );
  AND2_X1 U2378 ( .A1(n2240), .A2(n2265), .ZN(n2236) );
  INV_X1 U2379 ( .A(IR_REG_14__SCAN_IN), .ZN(n2448) );
  NOR2_X1 U2380 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2102)
         );
  NAND2_X1 U2381 ( .A1(n3202), .A2(n3201), .ZN(n2193) );
  NAND2_X1 U2382 ( .A1(n3753), .A2(n3752), .ZN(n2230) );
  NAND2_X1 U2383 ( .A1(n3755), .A2(n2231), .ZN(n2229) );
  NAND2_X1 U2384 ( .A1(n2737), .A2(n2738), .ZN(n2197) );
  AND2_X1 U2385 ( .A1(n2464), .A2(REG3_REG_16__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U2386 ( .A1(n2207), .A2(n2208), .ZN(n3711) );
  AOI21_X1 U2387 ( .B1(n2211), .B2(n2842), .A(n2038), .ZN(n2208) );
  OR2_X1 U2388 ( .A1(n3662), .A2(n2060), .ZN(n2207) );
  NAND2_X1 U2389 ( .A1(n2071), .A2(n2846), .ZN(n3712) );
  INV_X1 U2390 ( .A(n2180), .ZN(n2181) );
  AND2_X1 U2391 ( .A1(n2194), .A2(n3224), .ZN(n2072) );
  INV_X1 U2392 ( .A(n2193), .ZN(n2192) );
  AOI22_X1 U2393 ( .A1(n2762), .A2(n3197), .B1(IR_REG_0__SCAN_IN), .B2(n2692), 
        .ZN(n2693) );
  INV_X1 U2394 ( .A(n2231), .ZN(n2225) );
  NOR2_X1 U2395 ( .A1(n3648), .A2(n2228), .ZN(n2227) );
  INV_X1 U2396 ( .A(n2230), .ZN(n2228) );
  AND3_X1 U2397 ( .A1(n3164), .A2(n2872), .A3(n2871), .ZN(n2896) );
  OR2_X1 U2398 ( .A1(n2294), .A2(n2293), .ZN(n2301) );
  NAND2_X1 U2399 ( .A1(n4140), .A2(n2976), .ZN(n2990) );
  XNOR2_X1 U2400 ( .A(n2985), .B(n4561), .ZN(n4149) );
  NAND2_X1 U2401 ( .A1(n3034), .A2(n2997), .ZN(n3013) );
  AOI21_X1 U2402 ( .B1(n2099), .B2(n2096), .A(n3057), .ZN(n2095) );
  INV_X1 U2403 ( .A(n2099), .ZN(n2097) );
  OR2_X1 U2404 ( .A1(n2395), .A2(IR_REG_9__SCAN_IN), .ZN(n2415) );
  XNOR2_X1 U2405 ( .A(n3330), .B(n2177), .ZN(n4572) );
  NAND2_X1 U2406 ( .A1(n4598), .A2(n3317), .ZN(n3320) );
  NAND2_X1 U2407 ( .A1(n3320), .A2(n3319), .ZN(n3519) );
  NAND2_X1 U2408 ( .A1(n4583), .A2(n3332), .ZN(n3333) );
  NAND2_X1 U2409 ( .A1(n4594), .A2(REG2_REG_12__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U2410 ( .A1(n2091), .A2(n2090), .ZN(n4172) );
  INV_X1 U2411 ( .A(n2088), .ZN(n2090) );
  OAI21_X1 U2412 ( .B1(n3533), .B2(REG2_REG_14__SCAN_IN), .A(n2089), .ZN(n2088) );
  AND2_X1 U2413 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  NOR2_X1 U2414 ( .A1(n4419), .A2(n4426), .ZN(n2564) );
  INV_X1 U2415 ( .A(n3931), .ZN(n4222) );
  OR2_X1 U2416 ( .A1(n4263), .A2(n4280), .ZN(n2554) );
  NOR2_X1 U2417 ( .A1(n2164), .A2(n2047), .ZN(n2163) );
  NOR2_X1 U2418 ( .A1(n2039), .A2(n2530), .ZN(n2164) );
  OR2_X1 U2419 ( .A1(n3606), .A2(n2055), .ZN(n2161) );
  NOR2_X1 U2420 ( .A1(n2502), .A2(n2501), .ZN(n2510) );
  NOR2_X1 U2421 ( .A1(n3875), .A2(n2118), .ZN(n2117) );
  INV_X1 U2422 ( .A(n3824), .ZN(n2118) );
  NAND2_X1 U2423 ( .A1(n3913), .A2(n3872), .ZN(n2119) );
  NAND2_X1 U2424 ( .A1(n2441), .A2(n2041), .ZN(n3436) );
  OAI21_X1 U2425 ( .B1(n3350), .B2(n2050), .A(n2153), .ZN(n2152) );
  INV_X1 U2426 ( .A(n2154), .ZN(n2153) );
  NAND2_X1 U2427 ( .A1(n2158), .A2(n2035), .ZN(n2157) );
  AND2_X1 U2428 ( .A1(n3810), .A2(n3812), .ZN(n2243) );
  NAND2_X1 U2429 ( .A1(n2593), .A2(n3809), .ZN(n3234) );
  OR2_X1 U2430 ( .A1(n3148), .A2(n3806), .ZN(n2593) );
  NAND2_X1 U2431 ( .A1(n3181), .A2(n3868), .ZN(n3180) );
  AOI21_X1 U2432 ( .B1(n2674), .B2(n2939), .A(n2938), .ZN(n2872) );
  NAND2_X1 U2433 ( .A1(n4208), .A2(n3859), .ZN(n4399) );
  NOR2_X1 U2434 ( .A1(n4279), .A2(n2139), .ZN(n4208) );
  OR3_X1 U2435 ( .A1(n4210), .A2(n4418), .A3(n2140), .ZN(n2139) );
  NOR2_X1 U2436 ( .A1(n2141), .A2(n4418), .ZN(n4227) );
  INV_X1 U2437 ( .A(n4252), .ZN(n2141) );
  NOR2_X1 U2438 ( .A1(n4279), .A2(n2140), .ZN(n4252) );
  INV_X1 U2439 ( .A(n4412), .ZN(n4430) );
  OR2_X1 U2440 ( .A1(n4303), .A2(n4439), .ZN(n4279) );
  OR2_X1 U2441 ( .A1(n2042), .A2(n3575), .ZN(n3438) );
  NAND2_X1 U2442 ( .A1(n4702), .A2(n2370), .ZN(n3272) );
  AND3_X1 U2443 ( .A1(n2671), .A2(n2870), .A3(n2670), .ZN(n2679) );
  AND2_X1 U2444 ( .A1(n2683), .A2(n4675), .ZN(n3160) );
  NAND2_X1 U2445 ( .A1(n2234), .A2(n2235), .ZN(n2111) );
  OR2_X1 U2446 ( .A1(n2647), .A2(IR_REG_27__SCAN_IN), .ZN(n2627) );
  NOR2_X1 U2447 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2262)
         );
  NOR2_X1 U2448 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2261)
         );
  NOR2_X1 U2449 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2260)
         );
  CLKBUF_X1 U2450 ( .A(n2340), .Z(n2341) );
  NAND2_X1 U2451 ( .A1(n2652), .A2(n2924), .ZN(n2683) );
  NOR2_X1 U2452 ( .A1(n2919), .A2(n2672), .ZN(n2652) );
  OR2_X1 U2453 ( .A1(n2567), .A2(n2253), .ZN(n4228) );
  NAND2_X1 U2454 ( .A1(n2705), .A2(n2686), .ZN(n2707) );
  OAI211_X1 U2455 ( .C1(n2350), .C2(n4306), .A(n2543), .B(n2542), .ZN(n4441)
         );
  OR2_X1 U2456 ( .A1(n2295), .A2(n3094), .ZN(n2289) );
  XNOR2_X1 U2457 ( .A(n3059), .B(n2070), .ZN(n3060) );
  NAND2_X1 U2458 ( .A1(n4584), .A2(n4585), .ZN(n4583) );
  XNOR2_X1 U2459 ( .A(n4173), .B(n4159), .ZN(n4613) );
  NAND2_X1 U2460 ( .A1(n4613), .A2(n4611), .ZN(n4612) );
  NAND2_X1 U2461 ( .A1(n4621), .A2(n4623), .ZN(n4622) );
  NOR2_X1 U2462 ( .A1(n4629), .A2(n4628), .ZN(n4630) );
  NAND2_X1 U2463 ( .A1(n3623), .A2(n2137), .ZN(n2680) );
  INV_X1 U2464 ( .A(n2138), .ZN(n2137) );
  OAI21_X1 U2465 ( .B1(n3630), .B2(n4498), .A(n2637), .ZN(n2138) );
  AOI21_X1 U2466 ( .B1(n2773), .B2(n2206), .A(n2205), .ZN(n2204) );
  INV_X1 U2467 ( .A(n3570), .ZN(n2205) );
  INV_X1 U2468 ( .A(n2842), .ZN(n2209) );
  INV_X1 U2469 ( .A(n3537), .ZN(n2089) );
  OAI21_X1 U2470 ( .B1(n2156), .B2(n2155), .A(n2048), .ZN(n2154) );
  INV_X1 U2471 ( .A(n2428), .ZN(n2155) );
  OR2_X1 U2472 ( .A1(n4103), .A2(n3176), .ZN(n3801) );
  OR2_X1 U2473 ( .A1(n3182), .A2(n3072), .ZN(n3795) );
  AND2_X1 U2474 ( .A1(n4233), .A2(n4408), .ZN(n3844) );
  NAND2_X1 U2475 ( .A1(n4267), .A2(n4250), .ZN(n2140) );
  NAND2_X1 U2476 ( .A1(n2150), .A2(n4387), .ZN(n2149) );
  NOR2_X1 U2477 ( .A1(n3757), .A2(n4478), .ZN(n2150) );
  OR2_X1 U2478 ( .A1(n3544), .A2(n4487), .ZN(n3543) );
  INV_X1 U2479 ( .A(n3251), .ZN(n2730) );
  INV_X1 U2480 ( .A(n3125), .ZN(n2708) );
  INV_X1 U2481 ( .A(IR_REG_24__SCAN_IN), .ZN(n2645) );
  INV_X1 U2482 ( .A(IR_REG_23__SCAN_IN), .ZN(n2653) );
  AOI21_X1 U2483 ( .B1(n2586), .B2(n2585), .A(n2649), .ZN(n2076) );
  INV_X1 U2484 ( .A(IR_REG_18__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U2485 ( .A1(n2482), .A2(n2481), .ZN(n2496) );
  NOR2_X1 U2486 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2481)
         );
  INV_X1 U2487 ( .A(IR_REG_6__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U2488 ( .A1(n2196), .A2(n2195), .ZN(n2194) );
  INV_X1 U2489 ( .A(n3201), .ZN(n2196) );
  INV_X1 U2490 ( .A(n3202), .ZN(n2195) );
  NAND2_X1 U2491 ( .A1(n2204), .A2(n3571), .ZN(n2201) );
  NOR2_X1 U2492 ( .A1(n2204), .A2(n2203), .ZN(n2202) );
  NOR2_X1 U2493 ( .A1(n2773), .A2(n2206), .ZN(n2203) );
  NOR2_X1 U2494 ( .A1(n2222), .A2(n2221), .ZN(n2220) );
  INV_X1 U2495 ( .A(n2059), .ZN(n2222) );
  NAND2_X1 U2496 ( .A1(n3764), .A2(n2219), .ZN(n2218) );
  INV_X1 U2497 ( .A(n3669), .ZN(n2219) );
  INV_X1 U2498 ( .A(n2815), .ZN(n2867) );
  INV_X1 U2499 ( .A(n2197), .ZN(n2185) );
  INV_X1 U2500 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2384) );
  AND2_X1 U2501 ( .A1(n2692), .A2(REG1_REG_0__SCAN_IN), .ZN(n2689) );
  NOR2_X1 U2502 ( .A1(n3857), .A2(n2516), .ZN(n3890) );
  AOI22_X1 U2503 ( .A1(n2696), .A2(n2762), .B1(n3196), .B2(n2815), .ZN(n2698)
         );
  AOI22_X1 U2504 ( .A1(n3182), .A2(n2762), .B1(n3102), .B2(n2815), .ZN(n2685)
         );
  NAND2_X1 U2505 ( .A1(n2074), .A2(n2073), .ZN(n3690) );
  NAND2_X1 U2506 ( .A1(n2723), .A2(n2180), .ZN(n2179) );
  AND3_X1 U2507 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2352) );
  INV_X1 U2508 ( .A(n2786), .ZN(n2787) );
  INV_X1 U2509 ( .A(n2785), .ZN(n2788) );
  NOR2_X1 U2510 ( .A1(n2452), .A2(n2251), .ZN(n2464) );
  OR2_X1 U2511 ( .A1(n2763), .A2(n2884), .ZN(n2893) );
  NAND2_X1 U2512 ( .A1(n2992), .A2(n2991), .ZN(n2994) );
  AND2_X1 U2513 ( .A1(n2108), .A2(n2109), .ZN(n3029) );
  NAND2_X1 U2514 ( .A1(n3018), .A2(n2084), .ZN(n2081) );
  NOR2_X1 U2515 ( .A1(n3040), .A2(n2085), .ZN(n2084) );
  INV_X1 U2516 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2085) );
  OR2_X1 U2517 ( .A1(n2086), .A2(n3040), .ZN(n2083) );
  NAND2_X1 U2518 ( .A1(n2094), .A2(n2058), .ZN(n3330) );
  NAND2_X1 U2519 ( .A1(n4580), .A2(n3315), .ZN(n3316) );
  NAND2_X1 U2520 ( .A1(n3519), .A2(n3520), .ZN(n3522) );
  NAND2_X1 U2521 ( .A1(n4157), .A2(n4158), .ZN(n4160) );
  NAND2_X1 U2522 ( .A1(n4622), .A2(n2100), .ZN(n4176) );
  OR2_X1 U2523 ( .A1(n4175), .A2(REG2_REG_17__SCAN_IN), .ZN(n2100) );
  NOR2_X1 U2524 ( .A1(n4176), .A2(n4177), .ZN(n4188) );
  NAND2_X1 U2525 ( .A1(n2128), .A2(n2126), .ZN(n2619) );
  AND2_X1 U2526 ( .A1(n2129), .A2(n2127), .ZN(n2126) );
  OR2_X1 U2527 ( .A1(n4223), .A2(n4222), .ZN(n4225) );
  NAND2_X1 U2528 ( .A1(n2128), .A2(n2127), .ZN(n4260) );
  NAND2_X1 U2529 ( .A1(n2531), .A2(n2252), .ZN(n2540) );
  NAND2_X1 U2530 ( .A1(n2611), .A2(n3918), .ZN(n4328) );
  NAND2_X1 U2531 ( .A1(n2474), .A2(REG3_REG_17__SCAN_IN), .ZN(n2490) );
  OR2_X1 U2532 ( .A1(n2490), .A2(n2489), .ZN(n2502) );
  AND2_X1 U2533 ( .A1(n4376), .A2(n4377), .ZN(n3873) );
  AOI21_X1 U2534 ( .B1(n2117), .B2(n3437), .A(n2115), .ZN(n2114) );
  OR2_X1 U2535 ( .A1(n3913), .A2(n2116), .ZN(n2113) );
  INV_X1 U2536 ( .A(n2117), .ZN(n2116) );
  NAND2_X1 U2537 ( .A1(n3548), .A2(n3878), .ZN(n3582) );
  OAI21_X1 U2538 ( .B1(n2451), .B2(n2166), .A(n2043), .ZN(n2165) );
  NAND2_X1 U2539 ( .A1(n2417), .A2(REG3_REG_12__SCAN_IN), .ZN(n2429) );
  AOI21_X1 U2540 ( .B1(n2124), .B2(n2122), .A(n2121), .ZN(n2120) );
  INV_X1 U2541 ( .A(n2124), .ZN(n2123) );
  INV_X1 U2542 ( .A(n3816), .ZN(n2122) );
  INV_X1 U2543 ( .A(n2168), .ZN(n2167) );
  OAI21_X1 U2544 ( .B1(n2169), .B2(n2370), .A(n2383), .ZN(n2168) );
  OAI21_X1 U2545 ( .B1(n3234), .B2(n2594), .A(n3812), .ZN(n3273) );
  NOR2_X1 U2546 ( .A1(n2361), .A2(n3048), .ZN(n2372) );
  AOI21_X1 U2547 ( .B1(n2134), .B2(n2132), .A(n2131), .ZN(n2130) );
  INV_X1 U2548 ( .A(n2134), .ZN(n2133) );
  INV_X1 U2549 ( .A(n3804), .ZN(n2132) );
  INV_X1 U2550 ( .A(n4251), .ZN(n4338) );
  NAND2_X1 U2551 ( .A1(n3795), .A2(n3798), .ZN(n3076) );
  NOR2_X1 U2552 ( .A1(n4399), .A2(n4400), .ZN(n4398) );
  AND2_X1 U2553 ( .A1(n2575), .A2(n2574), .ZN(n4421) );
  OR2_X1 U2554 ( .A1(n4213), .A2(n2577), .ZN(n2575) );
  INV_X1 U2555 ( .A(n4280), .ZN(n4439) );
  NAND2_X1 U2556 ( .A1(n4320), .A2(n4304), .ZN(n4303) );
  AND2_X1 U2557 ( .A1(n4334), .A2(n4318), .ZN(n4320) );
  NOR2_X1 U2558 ( .A1(n4365), .A2(n4459), .ZN(n4334) );
  INV_X1 U2559 ( .A(n3891), .ZN(n4387) );
  NOR2_X1 U2560 ( .A1(n3543), .A2(n2148), .ZN(n4388) );
  INV_X1 U2561 ( .A(n2150), .ZN(n2148) );
  NOR2_X1 U2562 ( .A1(n3543), .A2(n4478), .ZN(n3610) );
  INV_X1 U2563 ( .A(n3781), .ZN(n3498) );
  NAND2_X1 U2564 ( .A1(n3499), .A2(n3498), .ZN(n3544) );
  NOR2_X1 U2565 ( .A1(n3438), .A2(n3599), .ZN(n3499) );
  NAND2_X1 U2566 ( .A1(n2144), .A2(n2601), .ZN(n2143) );
  INV_X1 U2567 ( .A(n2144), .ZN(n2142) );
  NOR2_X1 U2568 ( .A1(n3282), .A2(n2146), .ZN(n3430) );
  INV_X1 U2569 ( .A(n3455), .ZN(n3367) );
  NOR2_X1 U2570 ( .A1(n3282), .A2(n3343), .ZN(n3354) );
  OR2_X1 U2571 ( .A1(n3280), .A2(n3279), .ZN(n3282) );
  NAND2_X1 U2572 ( .A1(n2172), .A2(n2171), .ZN(n4702) );
  INV_X1 U2573 ( .A(n2243), .ZN(n2171) );
  AND2_X1 U2574 ( .A1(n3152), .A2(n2730), .ZN(n3233) );
  NAND2_X1 U2575 ( .A1(n2066), .A2(n3176), .ZN(n3175) );
  NOR2_X1 U2576 ( .A1(n3175), .A2(n3694), .ZN(n3152) );
  OR2_X1 U2577 ( .A1(n4564), .A2(n2635), .ZN(n4492) );
  NOR2_X1 U2578 ( .A1(n3102), .A2(n3194), .ZN(n3117) );
  INV_X1 U2579 ( .A(n4688), .ZN(n4698) );
  NAND2_X1 U2580 ( .A1(n2627), .A2(n2275), .ZN(n2626) );
  INV_X1 U2581 ( .A(IR_REG_27__SCAN_IN), .ZN(n2274) );
  AND2_X1 U2582 ( .A1(n2647), .A2(n2276), .ZN(n2625) );
  AND2_X1 U2583 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2276)
         );
  CLKBUF_X1 U2584 ( .A(n2677), .Z(n2655) );
  INV_X1 U2585 ( .A(IR_REG_13__SCAN_IN), .ZN(n2437) );
  INV_X1 U2586 ( .A(IR_REG_7__SCAN_IN), .ZN(n2378) );
  NOR2_X1 U2587 ( .A1(n2291), .A2(n2649), .ZN(n2178) );
  NAND2_X1 U2588 ( .A1(n2103), .A2(n2101), .ZN(n2974) );
  NAND2_X1 U2589 ( .A1(n2052), .A2(IR_REG_1__SCAN_IN), .ZN(n2103) );
  NOR2_X1 U2590 ( .A1(n2291), .A2(n2102), .ZN(n2101) );
  NAND2_X1 U2591 ( .A1(n2191), .A2(n2193), .ZN(n3225) );
  NAND2_X1 U2592 ( .A1(n3200), .A2(n2194), .ZN(n2191) );
  AOI21_X1 U2593 ( .B1(n3671), .B2(n2220), .A(n2080), .ZN(n2079) );
  NAND2_X1 U2594 ( .A1(n2198), .A2(n2201), .ZN(n3598) );
  OR2_X1 U2595 ( .A1(n2774), .A2(n2202), .ZN(n2198) );
  NAND2_X1 U2596 ( .A1(n3637), .A2(n2842), .ZN(n3640) );
  NAND2_X1 U2597 ( .A1(n2229), .A2(n2230), .ZN(n3649) );
  OAI21_X1 U2598 ( .B1(n3671), .B2(n2080), .A(n2214), .ZN(n2905) );
  AND2_X1 U2599 ( .A1(n2215), .A2(n3631), .ZN(n2214) );
  NAND2_X1 U2600 ( .A1(n2216), .A2(n2217), .ZN(n2215) );
  INV_X1 U2601 ( .A(n2220), .ZN(n2216) );
  NAND2_X1 U2602 ( .A1(n2903), .A2(n2902), .ZN(n2904) );
  NOR2_X1 U2603 ( .A1(n2190), .A2(n2187), .ZN(n3264) );
  AND2_X1 U2604 ( .A1(n2192), .A2(n3224), .ZN(n2187) );
  INV_X1 U2605 ( .A(n3185), .ZN(n3196) );
  INV_X1 U2606 ( .A(n4336), .ZN(n4459) );
  AND2_X1 U2607 ( .A1(n2182), .A2(n2036), .ZN(n3725) );
  INV_X1 U2608 ( .A(n2227), .ZN(n2226) );
  AOI21_X1 U2609 ( .B1(n2225), .B2(n2227), .A(n2224), .ZN(n2223) );
  INV_X1 U2610 ( .A(n2814), .ZN(n2224) );
  NAND2_X1 U2611 ( .A1(n3658), .A2(n3733), .ZN(n3737) );
  NAND2_X1 U2612 ( .A1(n2213), .A2(n3656), .ZN(n3744) );
  INV_X1 U2613 ( .A(n3072), .ZN(n3102) );
  AND2_X1 U2614 ( .A1(n2896), .A2(n2874), .ZN(n3787) );
  OAI21_X1 U2615 ( .B1(n4270), .B2(n2577), .A(n2285), .ZN(n4427) );
  NAND2_X1 U2616 ( .A1(n2553), .A2(n2552), .ZN(n4300) );
  OR2_X1 U2617 ( .A1(n2515), .A2(n2514), .ZN(n3955) );
  OR2_X1 U2618 ( .A1(n2506), .A2(n2505), .ZN(n3956) );
  NAND4_X1 U2619 ( .A1(n2469), .A2(n2468), .A3(n2467), .A4(n2466), .ZN(n3957)
         );
  NAND4_X1 U2620 ( .A1(n2316), .A2(n2315), .A3(n2314), .A4(n2313), .ZN(n4104)
         );
  OR2_X1 U2621 ( .A1(n2295), .A2(n3012), .ZN(n2300) );
  NAND2_X1 U2622 ( .A1(n4118), .A2(n4124), .ZN(n4137) );
  XNOR2_X1 U2623 ( .A(n2994), .B(n2993), .ZN(n4152) );
  NAND2_X1 U2624 ( .A1(n4152), .A2(REG1_REG_4__SCAN_IN), .ZN(n4151) );
  XNOR2_X1 U2625 ( .A(n3013), .B(n2998), .ZN(n2999) );
  NAND2_X1 U2626 ( .A1(n2999), .A2(REG1_REG_6__SCAN_IN), .ZN(n3015) );
  XNOR2_X1 U2627 ( .A(n3017), .B(n4560), .ZN(n3018) );
  NAND2_X1 U2628 ( .A1(n2081), .A2(n2083), .ZN(n3039) );
  AND2_X1 U2629 ( .A1(n2082), .A2(n2086), .ZN(n3041) );
  NAND2_X1 U2630 ( .A1(n3018), .A2(REG2_REG_6__SCAN_IN), .ZN(n2082) );
  AND2_X1 U2631 ( .A1(n2069), .A2(n2068), .ZN(n3063) );
  INV_X1 U2632 ( .A(n3312), .ZN(n3311) );
  AOI21_X1 U2633 ( .B1(n3056), .B2(REG2_REG_8__SCAN_IN), .A(n2097), .ZN(n3058)
         );
  XOR2_X1 U2634 ( .A(n3316), .B(n4591), .Z(n4599) );
  NAND2_X1 U2635 ( .A1(n4599), .A2(REG1_REG_12__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U2636 ( .A1(n4592), .A2(n3334), .ZN(n3531) );
  XOR2_X1 U2637 ( .A(n3522), .B(n3521), .Z(n4608) );
  OR2_X1 U2638 ( .A1(n4603), .A2(n4604), .ZN(n2093) );
  XNOR2_X1 U2639 ( .A(n4160), .B(n4159), .ZN(n4616) );
  NOR2_X1 U2640 ( .A1(n4616), .A2(REG1_REG_16__SCAN_IN), .ZN(n4617) );
  NAND2_X1 U2641 ( .A1(n4612), .A2(n4174), .ZN(n4621) );
  NOR2_X1 U2642 ( .A1(n4163), .A2(n4630), .ZN(n4184) );
  INV_X1 U2643 ( .A(n2565), .ZN(n4221) );
  OAI21_X1 U2644 ( .B1(n4228), .B2(n2577), .A(n2273), .ZN(n4412) );
  AND2_X1 U2645 ( .A1(n4566), .A2(n4489), .ZN(n4337) );
  NAND2_X1 U2646 ( .A1(n2128), .A2(n2616), .ZN(n4275) );
  NOR2_X1 U2647 ( .A1(n2160), .A2(n4316), .ZN(n2159) );
  INV_X1 U2648 ( .A(n2163), .ZN(n2160) );
  NAND2_X1 U2649 ( .A1(n2161), .A2(n2163), .ZN(n4317) );
  AND2_X1 U2650 ( .A1(n2162), .A2(n2039), .ZN(n4332) );
  OR2_X1 U2651 ( .A1(n3606), .A2(n2517), .ZN(n2162) );
  NAND2_X1 U2652 ( .A1(n2119), .A2(n2117), .ZN(n3495) );
  NAND2_X1 U2653 ( .A1(n2119), .A2(n3824), .ZN(n3494) );
  NAND2_X1 U2654 ( .A1(n3436), .A2(n2451), .ZN(n3497) );
  NAND2_X1 U2655 ( .A1(n4566), .A2(n3193), .ZN(n4389) );
  NAND2_X1 U2656 ( .A1(n2157), .A2(n2407), .ZN(n3419) );
  NAND4_X1 U2657 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n3961)
         );
  INV_X1 U2658 ( .A(n4394), .ZN(n4333) );
  NAND3_X1 U2659 ( .A1(n3160), .A2(n4698), .A3(n2897), .ZN(n4634) );
  INV_X1 U2660 ( .A(n4389), .ZN(n4651) );
  INV_X1 U2661 ( .A(n4713), .ZN(n4711) );
  OR2_X1 U2662 ( .A1(n4227), .A2(n4226), .ZN(n4515) );
  NAND2_X1 U2663 ( .A1(n3160), .A2(n2935), .ZN(n4674) );
  INV_X1 U2664 ( .A(IR_REG_29__SCAN_IN), .ZN(n2267) );
  OR2_X1 U2665 ( .A1(n2054), .A2(n2649), .ZN(n2269) );
  MUX2_X1 U2666 ( .A(n2649), .B(n2648), .S(IR_REG_26__SCAN_IN), .Z(n2650) );
  XNOR2_X1 U2667 ( .A(n2589), .B(IR_REG_22__SCAN_IN), .ZN(n3950) );
  XNOR2_X1 U2668 ( .A(n2587), .B(IR_REG_21__SCAN_IN), .ZN(n3941) );
  INV_X1 U2669 ( .A(n4175), .ZN(n4677) );
  INV_X1 U2670 ( .A(n3327), .ZN(n4683) );
  INV_X1 U2671 ( .A(IR_REG_5__SCAN_IN), .ZN(n2342) );
  OAI21_X1 U2672 ( .B1(n2680), .B2(n2136), .A(n2067), .ZN(n2681) );
  INV_X1 U2673 ( .A(n2302), .ZN(n3856) );
  NAND2_X1 U2674 ( .A1(n2278), .A2(n2277), .ZN(n2302) );
  AND2_X1 U2675 ( .A1(n2201), .A2(n2063), .ZN(n2034) );
  OR2_X1 U2676 ( .A1(n3961), .A2(n3455), .ZN(n2035) );
  NAND2_X1 U2677 ( .A1(n2715), .A2(n2714), .ZN(n2036) );
  NAND2_X1 U2678 ( .A1(n2720), .A2(n2722), .ZN(n2723) );
  INV_X1 U2679 ( .A(n3830), .ZN(n2115) );
  NAND2_X1 U2680 ( .A1(n2449), .A2(n2448), .ZN(n2480) );
  NAND2_X1 U2681 ( .A1(n2848), .A2(n2847), .ZN(n2038) );
  INV_X1 U2682 ( .A(n4418), .ZN(n4231) );
  NOR2_X1 U2683 ( .A1(n3857), .A2(n2279), .ZN(n4418) );
  NAND4_X1 U2684 ( .A1(n2301), .A2(n2300), .A3(n2299), .A4(n2298), .ZN(n2691)
         );
  NAND2_X1 U2685 ( .A1(n2615), .A2(n2614), .ZN(n2128) );
  OR2_X1 U2686 ( .A1(n2522), .A2(n2521), .ZN(n2039) );
  OR2_X1 U2687 ( .A1(n2729), .A2(n2728), .ZN(n2040) );
  AND2_X1 U2688 ( .A1(n3437), .A2(n2440), .ZN(n2041) );
  OR2_X1 U2689 ( .A1(n3282), .A2(n2143), .ZN(n2042) );
  INV_X1 U2690 ( .A(IR_REG_2__SCAN_IN), .ZN(n2309) );
  OR2_X1 U2691 ( .A1(n3681), .A2(n3781), .ZN(n2043) );
  NAND2_X1 U2692 ( .A1(n2229), .A2(n2227), .ZN(n3647) );
  AND2_X1 U2693 ( .A1(n2723), .A2(n3123), .ZN(n2044) );
  NOR2_X1 U2694 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2045)
         );
  NAND2_X1 U2695 ( .A1(n2435), .A2(n2234), .ZN(n2588) );
  AND2_X1 U2696 ( .A1(n2041), .A2(n2462), .ZN(n2046) );
  NOR2_X1 U2697 ( .A1(n4361), .A2(n4459), .ZN(n2047) );
  INV_X1 U2698 ( .A(n3262), .ZN(n2189) );
  OAI21_X1 U2699 ( .B1(n3755), .B2(n2226), .A(n2223), .ZN(n3658) );
  NAND2_X1 U2700 ( .A1(n3574), .A2(n3487), .ZN(n2048) );
  AND3_X1 U2701 ( .A1(n2174), .A2(n2234), .A3(n2175), .ZN(n2642) );
  NAND2_X1 U2702 ( .A1(n2435), .A2(n2263), .ZN(n2049) );
  NAND2_X1 U2703 ( .A1(n2428), .A2(n2035), .ZN(n2050) );
  NOR2_X1 U2704 ( .A1(n2977), .A2(n2106), .ZN(n2051) );
  XNOR2_X1 U2705 ( .A(n2685), .B(n2033), .ZN(n2705) );
  AND2_X1 U2706 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2052)
         );
  OR2_X1 U2707 ( .A1(n4279), .A2(n2676), .ZN(n2053) );
  NOR2_X1 U2708 ( .A1(n2110), .A2(n2111), .ZN(n2054) );
  INV_X1 U2709 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3190) );
  OR2_X1 U2710 ( .A1(n2517), .A2(n2530), .ZN(n2055) );
  INV_X1 U2711 ( .A(IR_REG_28__SCAN_IN), .ZN(n2628) );
  NOR2_X1 U2712 ( .A1(n2774), .A2(n2773), .ZN(n2056) );
  INV_X1 U2713 ( .A(n3668), .ZN(n2221) );
  INV_X1 U2714 ( .A(n3928), .ZN(n2129) );
  AND2_X1 U2715 ( .A1(n2441), .A2(n2440), .ZN(n2057) );
  NOR3_X1 U2716 ( .A1(n3543), .A2(n2149), .A3(n3890), .ZN(n2151) );
  OR2_X1 U2717 ( .A1(n3329), .A2(n3300), .ZN(n2058) );
  INV_X1 U2718 ( .A(n2147), .ZN(n4386) );
  NOR2_X1 U2719 ( .A1(n3543), .A2(n2149), .ZN(n2147) );
  NAND2_X1 U2720 ( .A1(n2863), .A2(n2862), .ZN(n2059) );
  NAND2_X1 U2721 ( .A1(n2059), .A2(n2218), .ZN(n2217) );
  INV_X1 U2722 ( .A(n2211), .ZN(n2210) );
  NAND2_X1 U2723 ( .A1(n2212), .A2(n3656), .ZN(n2211) );
  INV_X1 U2724 ( .A(n2480), .ZN(n2482) );
  OR2_X1 U2725 ( .A1(n2209), .A2(n3655), .ZN(n2060) );
  AND2_X1 U2726 ( .A1(n2093), .A2(n2092), .ZN(n2061) );
  OR2_X1 U2727 ( .A1(n3050), .A2(n3241), .ZN(n2062) );
  AND2_X2 U2728 ( .A1(n2679), .A2(n3165), .ZN(n4706) );
  INV_X1 U2729 ( .A(n4706), .ZN(n2136) );
  NAND2_X1 U2730 ( .A1(n3690), .A2(n2040), .ZN(n3200) );
  OR2_X1 U2731 ( .A1(n2781), .A2(n2780), .ZN(n2063) );
  NOR2_X1 U2732 ( .A1(n2743), .A2(n2742), .ZN(n2064) );
  OR2_X1 U2733 ( .A1(n4190), .A2(n2684), .ZN(n2882) );
  NAND2_X1 U2734 ( .A1(n3723), .A2(n2723), .ZN(n3689) );
  INV_X1 U2735 ( .A(n3818), .ZN(n2121) );
  NAND2_X1 U2736 ( .A1(n2182), .A2(n2181), .ZN(n3723) );
  OR2_X1 U2737 ( .A1(n3282), .A2(n2142), .ZN(n2065) );
  AND2_X1 U2738 ( .A1(n2708), .A2(n3117), .ZN(n2066) );
  INV_X1 U2739 ( .A(n3429), .ZN(n2145) );
  INV_X1 U2740 ( .A(n4159), .ZN(n4679) );
  INV_X1 U2741 ( .A(n4210), .ZN(n4408) );
  OR2_X1 U2742 ( .A1(REG0_REG_29__SCAN_IN), .A2(n4706), .ZN(n2067) );
  INV_X1 U2743 ( .A(n4591), .ZN(n2176) );
  INV_X1 U2744 ( .A(n4570), .ZN(n2177) );
  INV_X1 U2745 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2106) );
  INV_X1 U2746 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2096) );
  NAND2_X1 U2747 ( .A1(n3059), .A2(n4559), .ZN(n2068) );
  NAND2_X1 U2748 ( .A1(n3060), .A2(REG1_REG_8__SCAN_IN), .ZN(n2069) );
  INV_X1 U2749 ( .A(n4559), .ZN(n2070) );
  NAND2_X1 U2750 ( .A1(n2979), .A2(REG1_REG_3__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U2751 ( .A1(n3526), .A2(n3525), .ZN(n4157) );
  NAND2_X1 U2752 ( .A1(n4577), .A2(REG1_REG_10__SCAN_IN), .ZN(n4576) );
  NOR2_X2 U2753 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2291)
         );
  NAND2_X1 U2754 ( .A1(n3640), .A2(n2848), .ZN(n2071) );
  NAND2_X1 U2755 ( .A1(n2213), .A2(n2210), .ZN(n3637) );
  NAND2_X1 U2756 ( .A1(n3122), .A2(n2044), .ZN(n2073) );
  AND2_X1 U2757 ( .A1(n2179), .A2(n3691), .ZN(n2074) );
  AOI21_X2 U2758 ( .B1(n3704), .B2(n3700), .A(n3702), .ZN(n3755) );
  NOR2_X2 U2759 ( .A1(n3485), .A2(n3481), .ZN(n2774) );
  XNOR2_X2 U2760 ( .A(n2076), .B(IR_REG_20__SCAN_IN), .ZN(n2677) );
  NAND2_X2 U2761 ( .A1(n2509), .A2(IR_REG_31__SCAN_IN), .ZN(n2586) );
  OAI21_X1 U2762 ( .B1(n2077), .B2(n3771), .A(n3636), .ZN(U3211) );
  XNOR2_X1 U2763 ( .A(n2079), .B(n2078), .ZN(n2077) );
  INV_X1 U2764 ( .A(n3631), .ZN(n2078) );
  INV_X1 U2765 ( .A(n2217), .ZN(n2080) );
  AND2_X2 U2766 ( .A1(n2435), .A2(n2437), .ZN(n2449) );
  NAND2_X1 U2767 ( .A1(n2087), .A2(n4560), .ZN(n2086) );
  INV_X1 U2768 ( .A(n3017), .ZN(n2087) );
  INV_X1 U2769 ( .A(n3533), .ZN(n2092) );
  NAND2_X1 U2770 ( .A1(n2092), .A2(n4603), .ZN(n2091) );
  INV_X1 U2771 ( .A(n2093), .ZN(n4602) );
  OAI21_X1 U2772 ( .B1(n2097), .B2(n3056), .A(n2095), .ZN(n2094) );
  OAI21_X1 U2773 ( .B1(n2097), .B2(n3056), .A(n2095), .ZN(n2098) );
  INV_X1 U2774 ( .A(n2098), .ZN(n3328) );
  MUX2_X1 U2775 ( .A(n3190), .B(REG2_REG_1__SCAN_IN), .S(n2974), .Z(n4118) );
  NAND2_X1 U2776 ( .A1(n2983), .A2(n2105), .ZN(n2104) );
  NAND2_X1 U2777 ( .A1(n4149), .A2(REG2_REG_4__SCAN_IN), .ZN(n2108) );
  NAND2_X1 U2778 ( .A1(n2977), .A2(REG2_REG_3__SCAN_IN), .ZN(n2107) );
  XNOR2_X1 U2779 ( .A(n2983), .B(n2977), .ZN(n2984) );
  NAND2_X1 U2780 ( .A1(n2986), .A2(n4561), .ZN(n2109) );
  NAND3_X1 U2781 ( .A1(n2174), .A2(n2175), .A3(n2045), .ZN(n2110) );
  OR2_X1 U2782 ( .A1(n2112), .A2(n2111), .ZN(n3620) );
  NAND4_X1 U2783 ( .A1(n2174), .A2(n2175), .A3(n2045), .A4(n2267), .ZN(n2112)
         );
  NAND4_X1 U2784 ( .A1(n2174), .A2(n2234), .A3(n2235), .A4(n2175), .ZN(n2647)
         );
  NAND2_X1 U2785 ( .A1(n2113), .A2(n2114), .ZN(n3548) );
  NAND2_X2 U2786 ( .A1(n3794), .A2(n3791), .ZN(n3868) );
  OAI21_X1 U2787 ( .B1(n3212), .B2(n2123), .A(n2120), .ZN(n3421) );
  OAI21_X1 U2788 ( .B1(n3212), .B2(n3210), .A(n3816), .ZN(n3352) );
  OAI21_X1 U2789 ( .B1(n3168), .B2(n2133), .A(n2130), .ZN(n3148) );
  OAI21_X1 U2790 ( .B1(n3168), .B2(n2592), .A(n3804), .ZN(n3134) );
  AOI21_X1 U2791 ( .B1(n2592), .B2(n3804), .A(n2135), .ZN(n2134) );
  NAND2_X1 U2792 ( .A1(n3068), .A2(n3795), .ZN(n3111) );
  AOI21_X2 U2793 ( .B1(n3047), .B2(n3043), .A(n3042), .ZN(n3059) );
  NAND2_X1 U2794 ( .A1(n2619), .A2(n2618), .ZN(n4223) );
  XNOR2_X1 U2795 ( .A(n3532), .B(n4681), .ZN(n4603) );
  INV_X1 U2796 ( .A(n2151), .ZN(n4365) );
  INV_X1 U2797 ( .A(n3350), .ZN(n2158) );
  INV_X1 U2798 ( .A(n2152), .ZN(n3380) );
  AOI21_X2 U2799 ( .B1(n2441), .B2(n2046), .A(n2165), .ZN(n3542) );
  NAND2_X1 U2800 ( .A1(n2243), .A2(n2370), .ZN(n2170) );
  INV_X1 U2801 ( .A(n3242), .ZN(n2172) );
  INV_X1 U2802 ( .A(n2340), .ZN(n2174) );
  NOR2_X2 U2803 ( .A1(n2258), .A2(IR_REG_22__SCAN_IN), .ZN(n2175) );
  NOR2_X2 U2804 ( .A1(n2340), .A2(n2258), .ZN(n2435) );
  XNOR2_X2 U2805 ( .A(n2178), .B(IR_REG_2__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U2806 ( .A1(n3122), .A2(n3123), .ZN(n2182) );
  INV_X1 U2807 ( .A(n3224), .ZN(n2188) );
  OAI21_X2 U2808 ( .B1(n2186), .B2(n3262), .A(n2183), .ZN(n3340) );
  NAND2_X1 U2809 ( .A1(n2186), .A2(n2197), .ZN(n2190) );
  INV_X1 U2810 ( .A(n3571), .ZN(n2206) );
  OR2_X1 U2811 ( .A1(n3662), .A2(n3655), .ZN(n2213) );
  INV_X1 U2812 ( .A(n3745), .ZN(n2212) );
  AOI21_X1 U2813 ( .B1(n3671), .B2(n3668), .A(n3669), .ZN(n3766) );
  AND2_X1 U2814 ( .A1(n2642), .A2(n2236), .ZN(n2640) );
  AND2_X1 U2815 ( .A1(n2642), .A2(n2240), .ZN(n2638) );
  OAI21_X2 U2816 ( .B1(n3340), .B2(n3339), .A(n2750), .ZN(n3450) );
  INV_X2 U2817 ( .A(n4664), .ZN(n4566) );
  AND3_X1 U2818 ( .A1(n2879), .A2(n2880), .A3(n3787), .ZN(n2237) );
  INV_X1 U2819 ( .A(n4552), .ZN(n4505) );
  AND2_X1 U2820 ( .A1(n2704), .A2(n2703), .ZN(n2238) );
  AND2_X1 U2821 ( .A1(n2326), .A2(n2329), .ZN(n2239) );
  AND2_X1 U2822 ( .A1(n2653), .A2(n2645), .ZN(n2240) );
  OR2_X1 U2823 ( .A1(n4300), .A2(n4439), .ZN(n2241) );
  AND2_X1 U2824 ( .A1(n4441), .A2(n2544), .ZN(n2242) );
  OR2_X1 U2825 ( .A1(n4421), .A2(n4408), .ZN(n2244) );
  OAI21_X1 U2826 ( .B1(n3131), .B2(n2349), .A(n2348), .ZN(n3147) );
  OR2_X1 U2827 ( .A1(n3625), .A2(n4552), .ZN(n2245) );
  OR2_X1 U2828 ( .A1(n3625), .A2(n4486), .ZN(n2246) );
  OR2_X1 U2829 ( .A1(n4298), .A2(n4318), .ZN(n2248) );
  AND2_X1 U2830 ( .A1(n3956), .A2(n3891), .ZN(n2249) );
  OR2_X1 U2831 ( .A1(n3633), .A2(n4250), .ZN(n2250) );
  AND4_X1 U2832 ( .A1(n2262), .A2(n2261), .A3(n2260), .A4(n2259), .ZN(n2263)
         );
  AND2_X1 U2833 ( .A1(n3256), .A2(n2725), .ZN(n2347) );
  INV_X1 U2834 ( .A(n3453), .ZN(n2754) );
  INV_X1 U2835 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2408) );
  OR2_X1 U2836 ( .A1(n3871), .A2(n2347), .ZN(n2349) );
  INV_X1 U2837 ( .A(IR_REG_25__SCAN_IN), .ZN(n2265) );
  INV_X1 U2838 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2399) );
  OR2_X1 U2839 ( .A1(n2385), .A2(n2384), .ZN(n2400) );
  INV_X1 U2840 ( .A(n3482), .ZN(n2773) );
  NAND2_X1 U2841 ( .A1(n2352), .A2(REG3_REG_6__SCAN_IN), .ZN(n2361) );
  AND2_X1 U2842 ( .A1(n2557), .A2(REG3_REG_26__SCAN_IN), .ZN(n2559) );
  AND2_X1 U2843 ( .A1(n2510), .A2(REG3_REG_20__SCAN_IN), .ZN(n2531) );
  INV_X1 U2844 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3048) );
  INV_X1 U2845 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3321) );
  AND2_X1 U2846 ( .A1(n2610), .A2(n2609), .ZN(n3918) );
  OR2_X1 U2847 ( .A1(n2429), .A2(n3321), .ZN(n2452) );
  NOR2_X1 U2848 ( .A1(n2409), .A2(n2408), .ZN(n2417) );
  NAND2_X1 U2849 ( .A1(n2372), .A2(REG3_REG_8__SCAN_IN), .ZN(n2385) );
  INV_X1 U2850 ( .A(n3587), .ZN(n4478) );
  AND2_X1 U2851 ( .A1(n3944), .A2(n2963), .ZN(n4488) );
  INV_X1 U2852 ( .A(IR_REG_26__SCAN_IN), .ZN(n2266) );
  INV_X1 U2853 ( .A(n2642), .ZN(n2643) );
  OR2_X1 U2854 ( .A1(n2393), .A2(n2392), .ZN(n2395) );
  INV_X1 U2855 ( .A(n4300), .ZN(n4263) );
  OR2_X1 U2856 ( .A1(n2400), .A2(n2399), .ZN(n2409) );
  OR2_X1 U2857 ( .A1(n2546), .A2(n3716), .ZN(n2548) );
  XNOR2_X1 U2858 ( .A(n2705), .B(n2706), .ZN(n3097) );
  OR2_X1 U2859 ( .A1(n2559), .A2(n2558), .ZN(n4245) );
  INV_X1 U2860 ( .A(n4444), .ZN(n4489) );
  AND2_X1 U2861 ( .A1(n4294), .A2(n2612), .ZN(n4316) );
  OR2_X1 U2862 ( .A1(n3606), .A2(n3873), .ZN(n4374) );
  INV_X1 U2863 ( .A(n2472), .ZN(n4487) );
  INV_X1 U2864 ( .A(n4247), .ZN(n4342) );
  INV_X1 U2865 ( .A(n2935), .ZN(n2674) );
  INV_X1 U2866 ( .A(n4488), .ZN(n4409) );
  INV_X1 U2867 ( .A(n4250), .ZN(n4426) );
  INV_X1 U2868 ( .A(n3507), .ZN(n3599) );
  INV_X1 U2869 ( .A(n4492), .ZN(n4440) );
  INV_X1 U2870 ( .A(n4329), .ZN(n4384) );
  INV_X1 U2871 ( .A(n3715), .ZN(n3778) );
  NAND2_X1 U2872 ( .A1(n2898), .A2(n4634), .ZN(n3780) );
  NAND4_X1 U2873 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n3681)
         );
  NOR2_X1 U2874 ( .A1(n2978), .A2(n2971), .ZN(n4593) );
  NOR2_X1 U2875 ( .A1(n3850), .A2(n3844), .ZN(n4214) );
  AND2_X1 U2876 ( .A1(n4566), .A2(n4440), .ZN(n4247) );
  NAND2_X1 U2877 ( .A1(n2624), .A2(n2623), .ZN(n4329) );
  INV_X1 U2878 ( .A(n4486), .ZN(n4401) );
  AND2_X1 U2879 ( .A1(n4363), .A2(n4688), .ZN(n4498) );
  INV_X1 U2880 ( .A(n4498), .ZN(n4700) );
  NAND2_X1 U2881 ( .A1(n2666), .A2(n2924), .ZN(n2935) );
  XNOR2_X1 U2882 ( .A(n2646), .B(n2645), .ZN(n2672) );
  AND2_X1 U2883 ( .A1(n2470), .A2(n2461), .ZN(n3534) );
  INV_X1 U2884 ( .A(n4167), .ZN(n4626) );
  INV_X1 U2885 ( .A(n3787), .ZN(n3771) );
  INV_X1 U2886 ( .A(n4421), .ZN(n4233) );
  NAND2_X1 U2887 ( .A1(n2529), .A2(n2528), .ZN(n4361) );
  INV_X1 U2888 ( .A(n4593), .ZN(n4620) );
  NAND2_X1 U2889 ( .A1(n4109), .A2(n4564), .ZN(n4633) );
  NAND2_X1 U2890 ( .A1(n4566), .A2(n3244), .ZN(n4394) );
  NAND2_X1 U2891 ( .A1(n4713), .A2(n4693), .ZN(n4486) );
  AND2_X2 U2892 ( .A1(n2679), .A2(n2872), .ZN(n4713) );
  NAND2_X1 U2893 ( .A1(n4706), .A2(n4693), .ZN(n4552) );
  AND3_X1 U2894 ( .A1(n4705), .A2(n4704), .A3(n4703), .ZN(n4712) );
  INV_X1 U2895 ( .A(n4674), .ZN(n4673) );
  XNOR2_X1 U2896 ( .A(n2629), .B(n2628), .ZN(n4564) );
  AND2_X1 U2897 ( .A1(n2941), .A2(STATE_REG_SCAN_IN), .ZN(n4675) );
  OR2_X1 U2898 ( .A1(n2450), .A2(n2482), .ZN(n4681) );
  NAND2_X1 U2899 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n2251) );
  INV_X1 U2900 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2489) );
  INV_X1 U2901 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2501) );
  AND2_X1 U2902 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2252) );
  INV_X1 U2903 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3642) );
  INV_X1 U2904 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3716) );
  INV_X1 U2905 ( .A(REG3_REG_25__SCAN_IN), .ZN(n2280) );
  NOR2_X1 U2906 ( .A1(n2559), .A2(REG3_REG_27__SCAN_IN), .ZN(n2253) );
  INV_X1 U2907 ( .A(n2317), .ZN(n2254) );
  NAND2_X1 U2908 ( .A1(n2254), .A2(n2239), .ZN(n2340) );
  NOR2_X2 U2909 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2391)
         );
  XNOR2_X2 U2910 ( .A(n2268), .B(IR_REG_30__SCAN_IN), .ZN(n2930) );
  INV_X1 U2911 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4513) );
  NAND2_X1 U2912 ( .A1(n2630), .A2(REG2_REG_27__SCAN_IN), .ZN(n2271) );
  NAND2_X1 U2913 ( .A1(n3851), .A2(REG1_REG_27__SCAN_IN), .ZN(n2270) );
  OAI211_X1 U2914 ( .C1(n3852), .C2(n4513), .A(n2271), .B(n2270), .ZN(n2272)
         );
  INV_X1 U2915 ( .A(n2272), .ZN(n2273) );
  NAND2_X1 U2916 ( .A1(n2274), .A2(n2649), .ZN(n2275) );
  NAND2_X1 U2917 ( .A1(n2626), .A2(n2628), .ZN(n2278) );
  INV_X1 U2918 ( .A(DATAI_27_), .ZN(n2279) );
  NAND2_X1 U2919 ( .A1(n3856), .A2(DATAI_25_), .ZN(n4267) );
  INV_X1 U2920 ( .A(n4267), .ZN(n2676) );
  AND2_X1 U2921 ( .A1(n2548), .A2(n2280), .ZN(n2281) );
  OR2_X1 U2922 ( .A1(n2281), .A2(n2557), .ZN(n4270) );
  INV_X1 U2923 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U2924 ( .A1(n3851), .A2(REG1_REG_25__SCAN_IN), .ZN(n2283) );
  NAND2_X1 U2925 ( .A1(n2630), .A2(REG2_REG_25__SCAN_IN), .ZN(n2282) );
  OAI211_X1 U2926 ( .C1(n3852), .C2(n4521), .A(n2283), .B(n2282), .ZN(n2284)
         );
  INV_X1 U2927 ( .A(n2284), .ZN(n2285) );
  INV_X1 U2928 ( .A(n4427), .ZN(n4445) );
  NAND2_X1 U2929 ( .A1(n2296), .A2(REG1_REG_1__SCAN_IN), .ZN(n2290) );
  INV_X1 U2930 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3094) );
  NAND2_X1 U2931 ( .A1(n2297), .A2(REG2_REG_1__SCAN_IN), .ZN(n2288) );
  INV_X1 U2932 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2286) );
  NAND4_X2 U2933 ( .A1(n2290), .A2(n2289), .A3(n2288), .A4(n2287), .ZN(n2696)
         );
  INV_X1 U2934 ( .A(DATAI_1_), .ZN(n2292) );
  MUX2_X1 U2935 ( .A(n2292), .B(n2974), .S(n2302), .Z(n3185) );
  NAND2_X1 U2936 ( .A1(n2696), .A2(n3185), .ZN(n3791) );
  INV_X1 U2937 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2293) );
  INV_X1 U2938 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3012) );
  NAND2_X1 U2939 ( .A1(n2296), .A2(REG1_REG_0__SCAN_IN), .ZN(n2299) );
  NAND2_X1 U2940 ( .A1(n2297), .A2(REG2_REG_0__SCAN_IN), .ZN(n2298) );
  MUX2_X1 U2941 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2302), .Z(n3197) );
  AND2_X1 U2942 ( .A1(n2691), .A2(n3197), .ZN(n3181) );
  NAND2_X1 U2943 ( .A1(n2696), .A2(n3196), .ZN(n2303) );
  NAND2_X1 U2944 ( .A1(n2297), .A2(REG2_REG_2__SCAN_IN), .ZN(n2308) );
  NAND2_X1 U2945 ( .A1(n2359), .A2(REG1_REG_2__SCAN_IN), .ZN(n2307) );
  INV_X1 U2946 ( .A(REG3_REG_2__SCAN_IN), .ZN(n4129) );
  OR2_X1 U2947 ( .A1(n2577), .A2(n4129), .ZN(n2306) );
  INV_X1 U2948 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2304) );
  OR2_X1 U2949 ( .A1(n2294), .A2(n2304), .ZN(n2305) );
  INV_X1 U2950 ( .A(DATAI_2_), .ZN(n2310) );
  MUX2_X1 U2951 ( .A(n2310), .B(n4133), .S(n2302), .Z(n3072) );
  NAND2_X1 U2952 ( .A1(n3182), .A2(n3072), .ZN(n3798) );
  NAND2_X1 U2953 ( .A1(n3077), .A2(n3076), .ZN(n3075) );
  OR2_X1 U2954 ( .A1(n3182), .A2(n3102), .ZN(n2311) );
  NAND2_X1 U2955 ( .A1(n3075), .A2(n2311), .ZN(n3110) );
  NAND2_X1 U2956 ( .A1(n2630), .A2(REG2_REG_3__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2957 ( .A1(n2359), .A2(REG1_REG_3__SCAN_IN), .ZN(n2315) );
  OR2_X1 U2958 ( .A1(n2577), .A2(REG3_REG_3__SCAN_IN), .ZN(n2314) );
  INV_X1 U2959 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2312) );
  OR2_X1 U2960 ( .A1(n2294), .A2(n2312), .ZN(n2313) );
  NAND2_X1 U2961 ( .A1(n2317), .A2(IR_REG_31__SCAN_IN), .ZN(n2327) );
  XNOR2_X1 U2962 ( .A(n2327), .B(IR_REG_3__SCAN_IN), .ZN(n2989) );
  MUX2_X1 U2963 ( .A(DATAI_3_), .B(n2989), .S(n3857), .Z(n3125) );
  NAND2_X1 U2964 ( .A1(n4104), .A2(n3125), .ZN(n2318) );
  NAND2_X1 U2965 ( .A1(n3110), .A2(n2318), .ZN(n2320) );
  INV_X1 U2966 ( .A(n4104), .ZN(n3100) );
  NAND2_X1 U2967 ( .A1(n3100), .A2(n2708), .ZN(n2319) );
  NAND2_X1 U2968 ( .A1(n2320), .A2(n2319), .ZN(n3131) );
  NAND2_X1 U2969 ( .A1(n2359), .A2(REG1_REG_4__SCAN_IN), .ZN(n2325) );
  NAND2_X1 U2970 ( .A1(n2630), .A2(REG2_REG_4__SCAN_IN), .ZN(n2324) );
  INV_X1 U2971 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2321) );
  OR2_X1 U2972 ( .A1(n2294), .A2(n2321), .ZN(n2323) );
  XNOR2_X1 U2973 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3728) );
  OR2_X1 U2974 ( .A1(n2577), .A2(n3728), .ZN(n2322) );
  INV_X1 U2975 ( .A(DATAI_4_), .ZN(n2331) );
  NAND2_X1 U2976 ( .A1(n2327), .A2(n2326), .ZN(n2328) );
  NAND2_X1 U2977 ( .A1(n2328), .A2(IR_REG_31__SCAN_IN), .ZN(n2330) );
  XNOR2_X1 U2978 ( .A(n2330), .B(n2329), .ZN(n2993) );
  MUX2_X1 U2979 ( .A(n2331), .B(n2993), .S(n2302), .Z(n3176) );
  NAND2_X1 U2980 ( .A1(n4103), .A2(n3176), .ZN(n3804) );
  NAND2_X1 U2981 ( .A1(n3801), .A2(n3804), .ZN(n3169) );
  INV_X1 U2982 ( .A(n3169), .ZN(n3871) );
  NAND2_X1 U2983 ( .A1(n2359), .A2(REG1_REG_5__SCAN_IN), .ZN(n2339) );
  NAND2_X1 U2984 ( .A1(n2630), .A2(REG2_REG_5__SCAN_IN), .ZN(n2338) );
  INV_X1 U2985 ( .A(REG0_REG_5__SCAN_IN), .ZN(n3140) );
  OR2_X1 U2986 ( .A1(n2294), .A2(n3140), .ZN(n2337) );
  INV_X1 U2987 ( .A(n2352), .ZN(n2335) );
  INV_X1 U2988 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U2989 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2332) );
  NAND2_X1 U2990 ( .A1(n2333), .A2(n2332), .ZN(n2334) );
  NAND2_X1 U2991 ( .A1(n2335), .A2(n2334), .ZN(n3695) );
  OR2_X1 U2992 ( .A1(n2577), .A2(n3695), .ZN(n2336) );
  INV_X1 U2993 ( .A(DATAI_5_), .ZN(n2344) );
  NAND2_X1 U2994 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2343) );
  XNOR2_X1 U2995 ( .A(n2343), .B(n2342), .ZN(n3031) );
  MUX2_X1 U2996 ( .A(n2344), .B(n3031), .S(n3857), .Z(n2725) );
  INV_X1 U2997 ( .A(n3176), .ZN(n3727) );
  NAND2_X1 U2998 ( .A1(n4103), .A2(n3727), .ZN(n3132) );
  NAND2_X1 U2999 ( .A1(n4102), .A2(n3694), .ZN(n2345) );
  AND2_X1 U3000 ( .A1(n3132), .A2(n2345), .ZN(n2346) );
  OR2_X1 U3001 ( .A1(n2347), .A2(n2346), .ZN(n2348) );
  NAND2_X1 U3002 ( .A1(n3851), .A2(REG1_REG_6__SCAN_IN), .ZN(n2356) );
  INV_X4 U3003 ( .A(n2350), .ZN(n2630) );
  NAND2_X1 U3004 ( .A1(n2630), .A2(REG2_REG_6__SCAN_IN), .ZN(n2355) );
  INV_X1 U3005 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2351) );
  OR2_X1 U3006 ( .A1(n3852), .A2(n2351), .ZN(n2354) );
  OAI21_X1 U3007 ( .B1(n2352), .B2(REG3_REG_6__SCAN_IN), .A(n2361), .ZN(n3252)
         );
  OR2_X1 U3008 ( .A1(n2577), .A2(n3252), .ZN(n2353) );
  NAND4_X1 U3009 ( .A1(n2356), .A2(n2355), .A3(n2354), .A4(n2353), .ZN(n3693)
         );
  NOR2_X1 U3010 ( .A1(n2341), .A2(IR_REG_5__SCAN_IN), .ZN(n2368) );
  OR2_X1 U3011 ( .A1(n2368), .A2(n2649), .ZN(n2357) );
  XNOR2_X1 U3012 ( .A(n2357), .B(IR_REG_6__SCAN_IN), .ZN(n4560) );
  MUX2_X1 U3013 ( .A(DATAI_6_), .B(n4560), .S(n3857), .Z(n3251) );
  AND2_X1 U3014 ( .A1(n3693), .A2(n3251), .ZN(n2358) );
  OAI22_X1 U3015 ( .A1(n3147), .A2(n2358), .B1(n3251), .B2(n3693), .ZN(n3242)
         );
  NAND2_X1 U3016 ( .A1(n2359), .A2(REG1_REG_7__SCAN_IN), .ZN(n2366) );
  NAND2_X1 U3017 ( .A1(n2630), .A2(REG2_REG_7__SCAN_IN), .ZN(n2365) );
  INV_X1 U3018 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2360) );
  OR2_X1 U3019 ( .A1(n2294), .A2(n2360), .ZN(n2364) );
  AND2_X1 U3020 ( .A1(n2361), .A2(n3048), .ZN(n2362) );
  OR2_X1 U3021 ( .A1(n2362), .A2(n2372), .ZN(n3240) );
  OR2_X1 U3022 ( .A1(n2577), .A2(n3240), .ZN(n2363) );
  NAND4_X1 U3023 ( .A1(n2366), .A2(n2365), .A3(n2364), .A4(n2363), .ZN(n3274)
         );
  INV_X1 U3024 ( .A(DATAI_7_), .ZN(n2369) );
  NAND2_X1 U3025 ( .A1(n2368), .A2(n2367), .ZN(n2393) );
  NAND2_X1 U3026 ( .A1(n2393), .A2(IR_REG_31__SCAN_IN), .ZN(n2379) );
  XNOR2_X1 U3027 ( .A(n2379), .B(n2378), .ZN(n3050) );
  MUX2_X1 U3028 ( .A(n2369), .B(n3050), .S(n3857), .Z(n3237) );
  OR2_X1 U3029 ( .A1(n3274), .A2(n3237), .ZN(n3810) );
  NAND2_X1 U3030 ( .A1(n3274), .A2(n3237), .ZN(n3812) );
  INV_X1 U3031 ( .A(n3237), .ZN(n3227) );
  NAND2_X1 U3032 ( .A1(n3274), .A2(n3227), .ZN(n2370) );
  NAND2_X1 U3033 ( .A1(n3851), .A2(REG1_REG_8__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U3034 ( .A1(n2630), .A2(REG2_REG_8__SCAN_IN), .ZN(n2376) );
  INV_X1 U3035 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3036 ( .A1(n3852), .A2(n2371), .ZN(n2375) );
  OR2_X1 U3037 ( .A1(n2372), .A2(REG3_REG_8__SCAN_IN), .ZN(n2373) );
  NAND2_X1 U3038 ( .A1(n2385), .A2(n2373), .ZN(n4635) );
  OR2_X1 U3039 ( .A1(n2577), .A2(n4635), .ZN(n2374) );
  NAND4_X1 U3040 ( .A1(n2377), .A2(n2376), .A3(n2375), .A4(n2374), .ZN(n3342)
         );
  NAND2_X1 U3041 ( .A1(n2379), .A2(n2378), .ZN(n2380) );
  NAND2_X1 U3042 ( .A1(n2380), .A2(IR_REG_31__SCAN_IN), .ZN(n2381) );
  XNOR2_X1 U3043 ( .A(n2381), .B(IR_REG_8__SCAN_IN), .ZN(n4559) );
  MUX2_X1 U3044 ( .A(DATAI_8_), .B(n4559), .S(n3857), .Z(n3279) );
  OR2_X1 U3045 ( .A1(n3342), .A2(n3279), .ZN(n2382) );
  NAND2_X1 U3046 ( .A1(n3342), .A2(n3279), .ZN(n2383) );
  NAND2_X1 U3047 ( .A1(n2630), .A2(REG2_REG_9__SCAN_IN), .ZN(n2390) );
  NAND2_X1 U3048 ( .A1(n3851), .A2(REG1_REG_9__SCAN_IN), .ZN(n2389) );
  NAND2_X1 U3049 ( .A1(n2385), .A2(n2384), .ZN(n2386) );
  NAND2_X1 U3050 ( .A1(n2400), .A2(n2386), .ZN(n3346) );
  OR2_X1 U3051 ( .A1(n2577), .A2(n3346), .ZN(n2388) );
  INV_X1 U3052 ( .A(REG0_REG_9__SCAN_IN), .ZN(n3218) );
  OR2_X1 U3053 ( .A1(n3852), .A2(n3218), .ZN(n2387) );
  NAND4_X1 U3054 ( .A1(n2390), .A2(n2389), .A3(n2388), .A4(n2387), .ZN(n3962)
         );
  INV_X1 U3055 ( .A(n2391), .ZN(n2392) );
  NAND2_X1 U3056 ( .A1(n2395), .A2(IR_REG_31__SCAN_IN), .ZN(n2394) );
  MUX2_X1 U3057 ( .A(IR_REG_31__SCAN_IN), .B(n2394), .S(IR_REG_9__SCAN_IN), 
        .Z(n2396) );
  NAND2_X1 U3058 ( .A1(n2396), .A2(n2415), .ZN(n3329) );
  INV_X1 U3059 ( .A(n3329), .ZN(n4558) );
  MUX2_X1 U3060 ( .A(DATAI_9_), .B(n4558), .S(n3857), .Z(n3343) );
  AND2_X1 U3061 ( .A1(n3962), .A2(n3343), .ZN(n2397) );
  NAND2_X1 U3062 ( .A1(n3851), .A2(REG1_REG_10__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3063 ( .A1(n2630), .A2(REG2_REG_10__SCAN_IN), .ZN(n2404) );
  INV_X1 U3064 ( .A(REG0_REG_10__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3065 ( .A1(n3852), .A2(n2398), .ZN(n2403) );
  NAND2_X1 U3066 ( .A1(n2400), .A2(n2399), .ZN(n2401) );
  NAND2_X1 U3067 ( .A1(n2409), .A2(n2401), .ZN(n3458) );
  OR2_X1 U3068 ( .A1(n2577), .A2(n3458), .ZN(n2402) );
  NAND2_X1 U3069 ( .A1(n2415), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  XNOR2_X1 U3070 ( .A(n2406), .B(IR_REG_10__SCAN_IN), .ZN(n4570) );
  MUX2_X1 U3071 ( .A(DATAI_10_), .B(n4570), .S(n3857), .Z(n3455) );
  NAND2_X1 U3072 ( .A1(n3961), .A2(n3455), .ZN(n2407) );
  NAND2_X1 U3073 ( .A1(n3851), .A2(REG1_REG_11__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3074 ( .A1(n2630), .A2(REG2_REG_11__SCAN_IN), .ZN(n2413) );
  INV_X1 U3075 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3557) );
  OR2_X1 U3076 ( .A1(n3852), .A2(n3557), .ZN(n2412) );
  AND2_X1 U3077 ( .A1(n2409), .A2(n2408), .ZN(n2410) );
  OR2_X1 U3078 ( .A1(n2410), .A2(n2417), .ZN(n3428) );
  OR2_X1 U3079 ( .A1(n2577), .A2(n3428), .ZN(n2411) );
  NAND4_X1 U3080 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n3959)
         );
  INV_X1 U3081 ( .A(DATAI_11_), .ZN(n2416) );
  OAI21_X1 U3082 ( .B1(n2415), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2424) );
  XNOR2_X1 U3083 ( .A(n2424), .B(IR_REG_11__SCAN_IN), .ZN(n3327) );
  MUX2_X1 U3084 ( .A(n2416), .B(n4683), .S(n3857), .Z(n3429) );
  OR2_X1 U3085 ( .A1(n3959), .A2(n3429), .ZN(n3381) );
  NAND2_X1 U3086 ( .A1(n3959), .A2(n3429), .ZN(n3822) );
  NAND2_X1 U3087 ( .A1(n3381), .A2(n3822), .ZN(n3879) );
  INV_X1 U3088 ( .A(n3879), .ZN(n3420) );
  INV_X1 U3089 ( .A(n3959), .ZN(n3470) );
  NAND2_X1 U3090 ( .A1(n3470), .A2(n3429), .ZN(n3394) );
  NAND2_X1 U3091 ( .A1(n3851), .A2(REG1_REG_12__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U3092 ( .A1(n2630), .A2(REG2_REG_12__SCAN_IN), .ZN(n2421) );
  INV_X1 U3093 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3478) );
  OR2_X1 U3094 ( .A1(n3852), .A2(n3478), .ZN(n2420) );
  OR2_X1 U3095 ( .A1(n2417), .A2(REG3_REG_12__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3096 ( .A1(n2429), .A2(n2418), .ZN(n3490) );
  OR2_X1 U3097 ( .A1(n2577), .A2(n3490), .ZN(n2419) );
  NAND4_X1 U3098 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(n3574)
         );
  INV_X1 U3099 ( .A(n3574), .ZN(n3422) );
  INV_X1 U3100 ( .A(IR_REG_11__SCAN_IN), .ZN(n2423) );
  NAND2_X1 U3101 ( .A1(n2424), .A2(n2423), .ZN(n2425) );
  NAND2_X1 U3102 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3103 ( .A(n2426), .B(IR_REG_12__SCAN_IN), .ZN(n4591) );
  MUX2_X1 U3104 ( .A(DATAI_12_), .B(n4591), .S(n3857), .Z(n3487) );
  INV_X1 U3105 ( .A(n3487), .ZN(n2601) );
  NAND2_X1 U3106 ( .A1(n3422), .A2(n2601), .ZN(n2427) );
  AND2_X1 U3107 ( .A1(n3394), .A2(n2427), .ZN(n2428) );
  NAND2_X1 U3108 ( .A1(n3851), .A2(REG1_REG_13__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3109 ( .A1(n2630), .A2(REG2_REG_13__SCAN_IN), .ZN(n2433) );
  INV_X1 U3110 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3465) );
  OR2_X1 U3111 ( .A1(n3852), .A2(n3465), .ZN(n2432) );
  NAND2_X1 U3112 ( .A1(n2429), .A2(n3321), .ZN(n2430) );
  NAND2_X1 U3113 ( .A1(n2452), .A2(n2430), .ZN(n3578) );
  OR2_X1 U3114 ( .A1(n2577), .A2(n3578), .ZN(n2431) );
  NAND4_X1 U3115 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(n3958)
         );
  NOR2_X1 U3116 ( .A1(n2435), .A2(n2649), .ZN(n2436) );
  MUX2_X1 U3117 ( .A(n2649), .B(n2436), .S(IR_REG_13__SCAN_IN), .Z(n2438) );
  OR2_X1 U3118 ( .A1(n2438), .A2(n2449), .ZN(n3324) );
  INV_X1 U3119 ( .A(n3324), .ZN(n4557) );
  MUX2_X1 U3120 ( .A(DATAI_13_), .B(n4557), .S(n3857), .Z(n3575) );
  NOR2_X1 U3121 ( .A1(n3958), .A2(n3575), .ZN(n2439) );
  NAND2_X1 U3122 ( .A1(n3958), .A2(n3575), .ZN(n2440) );
  NAND2_X1 U3123 ( .A1(n3851), .A2(REG1_REG_14__SCAN_IN), .ZN(n2446) );
  NAND2_X1 U3124 ( .A1(n2630), .A2(REG2_REG_14__SCAN_IN), .ZN(n2445) );
  INV_X1 U3125 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3514) );
  OR2_X1 U3126 ( .A1(n3852), .A2(n3514), .ZN(n2444) );
  INV_X1 U3127 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2442) );
  XNOR2_X1 U3128 ( .A(n2452), .B(n2442), .ZN(n3602) );
  OR2_X1 U3129 ( .A1(n2577), .A2(n3602), .ZN(n2443) );
  NAND4_X1 U3130 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n3777)
         );
  INV_X1 U3131 ( .A(DATAI_14_), .ZN(n4680) );
  NOR2_X1 U3132 ( .A1(n2449), .A2(n2649), .ZN(n2447) );
  MUX2_X1 U3133 ( .A(n2649), .B(n2447), .S(IR_REG_14__SCAN_IN), .Z(n2450) );
  MUX2_X1 U3134 ( .A(n4680), .B(n4681), .S(n3857), .Z(n3507) );
  OR2_X1 U3135 ( .A1(n3777), .A2(n3507), .ZN(n3824) );
  NAND2_X1 U3136 ( .A1(n3777), .A2(n3507), .ZN(n3829) );
  NAND2_X1 U3137 ( .A1(n3824), .A2(n3829), .ZN(n3437) );
  INV_X1 U3138 ( .A(n3777), .ZN(n3562) );
  NAND2_X1 U3139 ( .A1(n3562), .A2(n3507), .ZN(n2451) );
  NAND2_X1 U3140 ( .A1(n3851), .A2(REG1_REG_15__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3141 ( .A1(n2630), .A2(REG2_REG_15__SCAN_IN), .ZN(n2457) );
  INV_X1 U3142 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3565) );
  OR2_X1 U3143 ( .A1(n3852), .A2(n3565), .ZN(n2456) );
  INV_X1 U3144 ( .A(n2452), .ZN(n2453) );
  AOI21_X1 U3145 ( .B1(n2453), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n2454) );
  OR2_X1 U3146 ( .A1(n2454), .A2(n2464), .ZN(n3784) );
  OR2_X1 U3147 ( .A1(n2577), .A2(n3784), .ZN(n2455) );
  NAND2_X1 U31480 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2460) );
  INV_X1 U31490 ( .A(IR_REG_15__SCAN_IN), .ZN(n2459) );
  NAND2_X1 U3150 ( .A1(n2460), .A2(n2459), .ZN(n2470) );
  OR2_X1 U3151 ( .A1(n2460), .A2(n2459), .ZN(n2461) );
  MUX2_X1 U3152 ( .A(DATAI_15_), .B(n3534), .S(n3857), .Z(n3781) );
  NAND2_X1 U3153 ( .A1(n3681), .A2(n3781), .ZN(n2462) );
  NAND2_X1 U3154 ( .A1(n3851), .A2(REG1_REG_16__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3155 ( .A1(n2630), .A2(REG2_REG_16__SCAN_IN), .ZN(n2468) );
  INV_X1 U3156 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2463) );
  OR2_X1 U3157 ( .A1(n3852), .A2(n2463), .ZN(n2467) );
  NOR2_X1 U3158 ( .A1(n2464), .A2(REG3_REG_16__SCAN_IN), .ZN(n2465) );
  OR2_X1 U3159 ( .A1(n2474), .A2(n2465), .ZN(n3685) );
  OR2_X1 U3160 ( .A1(n2577), .A2(n3685), .ZN(n2466) );
  INV_X1 U3161 ( .A(DATAI_16_), .ZN(n4678) );
  NAND2_X1 U3162 ( .A1(n2470), .A2(IR_REG_31__SCAN_IN), .ZN(n2471) );
  XNOR2_X1 U3163 ( .A(n2471), .B(IR_REG_16__SCAN_IN), .ZN(n4159) );
  MUX2_X1 U3164 ( .A(n4678), .B(n4679), .S(n3857), .Z(n2472) );
  OR2_X1 U3165 ( .A1(n3957), .A2(n2472), .ZN(n3916) );
  NAND2_X1 U3166 ( .A1(n3957), .A2(n2472), .ZN(n3833) );
  NAND2_X1 U3167 ( .A1(n3916), .A2(n3833), .ZN(n3541) );
  NAND2_X1 U3168 ( .A1(n3542), .A2(n3541), .ZN(n3540) );
  NAND2_X1 U3169 ( .A1(n3957), .A2(n4487), .ZN(n2473) );
  NAND2_X1 U3170 ( .A1(n3540), .A2(n2473), .ZN(n3585) );
  NAND2_X1 U3171 ( .A1(n3851), .A2(REG1_REG_17__SCAN_IN), .ZN(n2479) );
  NAND2_X1 U3172 ( .A1(n2630), .A2(REG2_REG_17__SCAN_IN), .ZN(n2478) );
  INV_X1 U3173 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4550) );
  OR2_X1 U3174 ( .A1(n3852), .A2(n4550), .ZN(n2477) );
  OR2_X1 U3175 ( .A1(n2474), .A2(REG3_REG_17__SCAN_IN), .ZN(n2475) );
  NAND2_X1 U3176 ( .A1(n2490), .A2(n2475), .ZN(n3707) );
  OR2_X1 U3177 ( .A1(n2577), .A2(n3707), .ZN(n2476) );
  NAND4_X1 U3178 ( .A1(n2479), .A2(n2478), .A3(n2477), .A4(n2476), .ZN(n4490)
         );
  INV_X1 U3179 ( .A(n4490), .ZN(n3613) );
  INV_X1 U3180 ( .A(DATAI_17_), .ZN(n2484) );
  NAND2_X1 U3181 ( .A1(n2496), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  XNOR2_X1 U3182 ( .A(n2483), .B(IR_REG_17__SCAN_IN), .ZN(n4175) );
  MUX2_X1 U3183 ( .A(n2484), .B(n4677), .S(n3857), .Z(n3587) );
  NAND2_X1 U3184 ( .A1(n3613), .A2(n3587), .ZN(n2485) );
  NAND2_X1 U3185 ( .A1(n3585), .A2(n2485), .ZN(n2487) );
  NAND2_X1 U3186 ( .A1(n4490), .A2(n4478), .ZN(n2486) );
  NAND2_X1 U3187 ( .A1(n2487), .A2(n2486), .ZN(n3606) );
  NAND2_X1 U3188 ( .A1(n3851), .A2(REG1_REG_18__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U3189 ( .A1(n2630), .A2(REG2_REG_18__SCAN_IN), .ZN(n2494) );
  INV_X1 U3190 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2488) );
  OR2_X1 U3191 ( .A1(n3852), .A2(n2488), .ZN(n2493) );
  NAND2_X1 U3192 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U3193 ( .A1(n2502), .A2(n2491), .ZN(n3760) );
  OR2_X1 U3194 ( .A1(n2577), .A2(n3760), .ZN(n2492) );
  NAND4_X1 U3195 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n4479)
         );
  INV_X1 U3196 ( .A(DATAI_18_), .ZN(n2499) );
  INV_X1 U3197 ( .A(n2508), .ZN(n2497) );
  NAND2_X1 U3198 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U3199 ( .A(n2498), .B(n2507), .ZN(n4164) );
  MUX2_X1 U3200 ( .A(n2499), .B(n4164), .S(n3857), .Z(n3609) );
  OR2_X1 U3201 ( .A1(n4479), .A2(n3609), .ZN(n4376) );
  NAND2_X1 U3202 ( .A1(n4479), .A2(n3609), .ZN(n4377) );
  INV_X1 U3203 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4545) );
  NAND2_X1 U3204 ( .A1(n3851), .A2(REG1_REG_19__SCAN_IN), .ZN(n2500) );
  OAI21_X1 U3205 ( .B1(n3852), .B2(n4545), .A(n2500), .ZN(n2506) );
  AND2_X1 U3206 ( .A1(n2502), .A2(n2501), .ZN(n2503) );
  OR2_X1 U3207 ( .A1(n2503), .A2(n2510), .ZN(n4390) );
  NAND2_X1 U3208 ( .A1(n2630), .A2(REG2_REG_19__SCAN_IN), .ZN(n2504) );
  OAI21_X1 U3209 ( .B1(n4390), .B2(n2577), .A(n2504), .ZN(n2505) );
  NAND2_X1 U32100 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  XNOR2_X2 U32110 ( .A(n2586), .B(IR_REG_19__SCAN_IN), .ZN(n4190) );
  MUX2_X1 U32120 ( .A(DATAI_19_), .B(n4190), .S(n3857), .Z(n3891) );
  OR2_X1 U32130 ( .A1(n3873), .A2(n2249), .ZN(n4347) );
  NOR2_X1 U32140 ( .A1(n2510), .A2(REG3_REG_20__SCAN_IN), .ZN(n2511) );
  OR2_X1 U32150 ( .A1(n2531), .A2(n2511), .ZN(n4367) );
  NAND2_X1 U32160 ( .A1(n2630), .A2(REG2_REG_20__SCAN_IN), .ZN(n2512) );
  OAI21_X1 U32170 ( .B1(n4367), .B2(n2577), .A(n2512), .ZN(n2515) );
  INV_X1 U32180 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U32190 ( .A1(n3851), .A2(REG1_REG_20__SCAN_IN), .ZN(n2513) );
  OAI21_X1 U32200 ( .B1(n3852), .B2(n4541), .A(n2513), .ZN(n2514) );
  INV_X1 U32210 ( .A(DATAI_20_), .ZN(n2516) );
  AND2_X1 U32220 ( .A1(n3955), .A2(n3890), .ZN(n2522) );
  OR2_X1 U32230 ( .A1(n4347), .A2(n2522), .ZN(n2517) );
  OR2_X1 U32240 ( .A1(n3955), .A2(n3890), .ZN(n2520) );
  INV_X1 U32250 ( .A(n3609), .ZN(n3757) );
  OR2_X1 U32260 ( .A1(n4479), .A2(n3757), .ZN(n4373) );
  INV_X1 U32270 ( .A(n3956), .ZN(n4351) );
  NAND2_X1 U32280 ( .A1(n4351), .A2(n4387), .ZN(n2518) );
  AND2_X1 U32290 ( .A1(n4373), .A2(n2518), .ZN(n2519) );
  OR2_X1 U32300 ( .A1(n2249), .A2(n2519), .ZN(n4348) );
  AND2_X1 U32310 ( .A1(n2520), .A2(n4348), .ZN(n2521) );
  INV_X1 U32320 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U32330 ( .A1(n3851), .A2(REG1_REG_21__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32340 ( .A1(n2630), .A2(REG2_REG_21__SCAN_IN), .ZN(n2523) );
  OAI211_X1 U32350 ( .C1(n3852), .C2(n4537), .A(n2524), .B(n2523), .ZN(n2525)
         );
  INV_X1 U32360 ( .A(n2525), .ZN(n2529) );
  INV_X1 U32370 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2526) );
  XNOR2_X1 U32380 ( .A(n2531), .B(n2526), .ZN(n4339) );
  INV_X1 U32390 ( .A(n2577), .ZN(n2527) );
  NAND2_X1 U32400 ( .A1(n4339), .A2(n2527), .ZN(n2528) );
  NAND2_X1 U32410 ( .A1(n3856), .A2(DATAI_21_), .ZN(n4336) );
  AND2_X1 U32420 ( .A1(n4361), .A2(n4459), .ZN(n2530) );
  INV_X1 U32430 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U32440 ( .A1(n2531), .A2(REG3_REG_21__SCAN_IN), .ZN(n2533) );
  INV_X1 U32450 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32460 ( .A1(n2533), .A2(n2532), .ZN(n2534) );
  NAND2_X1 U32470 ( .A1(n2534), .A2(n2540), .ZN(n4321) );
  OR2_X1 U32480 ( .A1(n4321), .A2(n2577), .ZN(n2538) );
  NAND2_X1 U32490 ( .A1(n2630), .A2(REG2_REG_22__SCAN_IN), .ZN(n2536) );
  NAND2_X1 U32500 ( .A1(n3851), .A2(REG1_REG_22__SCAN_IN), .ZN(n2535) );
  AND2_X1 U32510 ( .A1(n2536), .A2(n2535), .ZN(n2537) );
  OAI211_X1 U32520 ( .C1(n3852), .C2(n2539), .A(n2538), .B(n2537), .ZN(n4460)
         );
  NAND2_X1 U32530 ( .A1(n3856), .A2(DATAI_22_), .ZN(n4318) );
  OR2_X1 U32540 ( .A1(n4460), .A2(n4318), .ZN(n4294) );
  NAND2_X1 U32550 ( .A1(n4460), .A2(n4318), .ZN(n2612) );
  INV_X1 U32560 ( .A(n4460), .ZN(n4298) );
  NAND2_X1 U32570 ( .A1(n2247), .A2(n2248), .ZN(n4290) );
  INV_X1 U32580 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U32590 ( .A1(n2540), .A2(n3642), .ZN(n2541) );
  NAND2_X1 U32600 ( .A1(n2546), .A2(n2541), .ZN(n4305) );
  OR2_X1 U32610 ( .A1(n4305), .A2(n2577), .ZN(n2543) );
  INV_X1 U32620 ( .A(n3852), .ZN(n2578) );
  AOI22_X1 U32630 ( .A1(n2578), .A2(REG0_REG_23__SCAN_IN), .B1(n3851), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n2542) );
  INV_X1 U32640 ( .A(n4441), .ZN(n4285) );
  NAND2_X1 U32650 ( .A1(n3856), .A2(DATAI_23_), .ZN(n4304) );
  NAND2_X1 U32660 ( .A1(n4285), .A2(n4304), .ZN(n2545) );
  INV_X1 U32670 ( .A(n4304), .ZN(n2544) );
  AOI21_X1 U32680 ( .B1(n4290), .B2(n2545), .A(n2242), .ZN(n4277) );
  NAND2_X1 U32690 ( .A1(n2546), .A2(n3716), .ZN(n2547) );
  AND2_X1 U32700 ( .A1(n2548), .A2(n2547), .ZN(n4282) );
  NAND2_X1 U32710 ( .A1(n4282), .A2(n2527), .ZN(n2553) );
  INV_X1 U32720 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4525) );
  NAND2_X1 U32730 ( .A1(n3851), .A2(REG1_REG_24__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32740 ( .A1(n2630), .A2(REG2_REG_24__SCAN_IN), .ZN(n2549) );
  OAI211_X1 U32750 ( .C1(n3852), .C2(n4525), .A(n2550), .B(n2549), .ZN(n2551)
         );
  INV_X1 U32760 ( .A(n2551), .ZN(n2552) );
  NAND2_X1 U32770 ( .A1(n3856), .A2(DATAI_24_), .ZN(n4280) );
  NAND2_X1 U32780 ( .A1(n4277), .A2(n2554), .ZN(n2555) );
  NAND2_X1 U32790 ( .A1(n2555), .A2(n2241), .ZN(n4258) );
  AOI21_X1 U32800 ( .B1(n4445), .B2(n4267), .A(n4258), .ZN(n2556) );
  AOI21_X1 U32810 ( .B1(n2676), .B2(n4427), .A(n2556), .ZN(n4244) );
  NOR2_X1 U32820 ( .A1(n2557), .A2(REG3_REG_26__SCAN_IN), .ZN(n2558) );
  INV_X1 U32830 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U32840 ( .A1(n3851), .A2(REG1_REG_26__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32850 ( .A1(n2630), .A2(REG2_REG_26__SCAN_IN), .ZN(n2560) );
  OAI211_X1 U32860 ( .C1(n3852), .C2(n4517), .A(n2561), .B(n2560), .ZN(n2562)
         );
  INV_X1 U32870 ( .A(n2562), .ZN(n2563) );
  OAI21_X2 U32880 ( .B1(n4245), .B2(n2577), .A(n2563), .ZN(n4419) );
  INV_X1 U32890 ( .A(n4419), .ZN(n3633) );
  NAND2_X1 U32900 ( .A1(n3856), .A2(DATAI_26_), .ZN(n4250) );
  AOI21_X1 U32910 ( .B1(n4244), .B2(n2250), .A(n2564), .ZN(n2565) );
  NAND2_X1 U32920 ( .A1(n2567), .A2(REG3_REG_28__SCAN_IN), .ZN(n3624) );
  INV_X1 U32930 ( .A(n2567), .ZN(n2569) );
  INV_X1 U32940 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2568) );
  NAND2_X1 U32950 ( .A1(n2569), .A2(n2568), .ZN(n2570) );
  NAND2_X1 U32960 ( .A1(n3624), .A2(n2570), .ZN(n4213) );
  INV_X1 U32970 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3969) );
  NAND2_X1 U32980 ( .A1(n3851), .A2(REG1_REG_28__SCAN_IN), .ZN(n2572) );
  NAND2_X1 U32990 ( .A1(n2297), .A2(REG2_REG_28__SCAN_IN), .ZN(n2571) );
  OAI211_X1 U33000 ( .C1(n3852), .C2(n3969), .A(n2572), .B(n2571), .ZN(n2573)
         );
  INV_X1 U33010 ( .A(n2573), .ZN(n2574) );
  INV_X1 U33020 ( .A(DATAI_28_), .ZN(n2576) );
  NOR2_X1 U33030 ( .A1(n3857), .A2(n2576), .ZN(n4210) );
  AND2_X1 U33040 ( .A1(n4421), .A2(n4210), .ZN(n3850) );
  OR2_X1 U33050 ( .A1(n3624), .A2(n2577), .ZN(n2583) );
  INV_X1 U33060 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U33070 ( .A1(n3851), .A2(REG1_REG_29__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U33080 ( .A1(n2578), .A2(REG0_REG_29__SCAN_IN), .ZN(n2579) );
  OAI211_X1 U33090 ( .C1(n3621), .C2(n2350), .A(n2580), .B(n2579), .ZN(n2581)
         );
  INV_X1 U33100 ( .A(n2581), .ZN(n2582) );
  NAND2_X1 U33110 ( .A1(n2583), .A2(n2582), .ZN(n4407) );
  NAND2_X1 U33120 ( .A1(n3856), .A2(DATAI_29_), .ZN(n3859) );
  XNOR2_X1 U33130 ( .A(n4407), .B(n3859), .ZN(n3909) );
  XNOR2_X1 U33140 ( .A(n2584), .B(n3909), .ZN(n3630) );
  NAND2_X1 U33150 ( .A1(n2049), .A2(IR_REG_31__SCAN_IN), .ZN(n2587) );
  NAND2_X2 U33160 ( .A1(n2677), .A2(n3941), .ZN(n3167) );
  NAND2_X1 U33170 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2589) );
  XNOR2_X1 U33180 ( .A(n3167), .B(n3950), .ZN(n2590) );
  NAND2_X1 U33190 ( .A1(n2590), .A2(n4196), .ZN(n4363) );
  NAND2_X1 U33200 ( .A1(n2655), .A2(n4190), .ZN(n4657) );
  OR2_X1 U33210 ( .A1(n4657), .A2(n3950), .ZN(n4688) );
  INV_X1 U33220 ( .A(n3197), .ZN(n2962) );
  OR2_X1 U33230 ( .A1(n2691), .A2(n2962), .ZN(n3790) );
  OAI21_X1 U33240 ( .B1(n3868), .B2(n3790), .A(n3794), .ZN(n3069) );
  INV_X1 U33250 ( .A(n3076), .ZN(n3870) );
  NAND2_X1 U33260 ( .A1(n3069), .A2(n3870), .ZN(n3068) );
  OR2_X1 U33270 ( .A1(n4104), .A2(n2708), .ZN(n3800) );
  NAND2_X1 U33280 ( .A1(n4104), .A2(n2708), .ZN(n3797) );
  NAND2_X1 U33290 ( .A1(n3800), .A2(n3797), .ZN(n3109) );
  INV_X1 U33300 ( .A(n3109), .ZN(n3877) );
  NAND2_X1 U33310 ( .A1(n3111), .A2(n3877), .ZN(n2591) );
  NAND2_X1 U33320 ( .A1(n2591), .A2(n3800), .ZN(n3168) );
  INV_X1 U33330 ( .A(n3801), .ZN(n2592) );
  OR2_X1 U33340 ( .A1(n4102), .A2(n2725), .ZN(n3807) );
  NAND2_X1 U33350 ( .A1(n4102), .A2(n2725), .ZN(n3803) );
  AND2_X1 U33360 ( .A1(n3693), .A2(n2730), .ZN(n3806) );
  OR2_X1 U33370 ( .A1(n3693), .A2(n2730), .ZN(n3809) );
  INV_X1 U33380 ( .A(n3810), .ZN(n2594) );
  INV_X1 U33390 ( .A(n3279), .ZN(n2595) );
  OR2_X1 U33400 ( .A1(n3342), .A2(n2595), .ZN(n3815) );
  NAND2_X1 U33410 ( .A1(n3273), .A2(n3815), .ZN(n2596) );
  NAND2_X1 U33420 ( .A1(n3342), .A2(n2595), .ZN(n3811) );
  NAND2_X1 U33430 ( .A1(n2596), .A2(n3811), .ZN(n3212) );
  INV_X1 U33440 ( .A(n3343), .ZN(n2597) );
  AND2_X1 U33450 ( .A1(n3962), .A2(n2597), .ZN(n3210) );
  OR2_X1 U33460 ( .A1(n3962), .A2(n2597), .ZN(n3816) );
  NAND2_X1 U33470 ( .A1(n3961), .A2(n3367), .ZN(n3821) );
  OR2_X1 U33480 ( .A1(n3961), .A2(n3367), .ZN(n3818) );
  NAND2_X1 U33490 ( .A1(n3574), .A2(n2601), .ZN(n3395) );
  INV_X1 U33500 ( .A(n3575), .ZN(n3385) );
  NAND2_X1 U33510 ( .A1(n3958), .A2(n3385), .ZN(n3377) );
  NAND2_X1 U33520 ( .A1(n3395), .A2(n3377), .ZN(n2600) );
  INV_X1 U3353 ( .A(n3822), .ZN(n2598) );
  NOR2_X1 U33540 ( .A1(n2600), .A2(n2598), .ZN(n2599) );
  NAND2_X1 U3355 ( .A1(n3421), .A2(n2599), .ZN(n2603) );
  INV_X1 U3356 ( .A(n2600), .ZN(n3823) );
  OR2_X1 U3357 ( .A1(n3574), .A2(n2601), .ZN(n3396) );
  NAND2_X1 U3358 ( .A1(n3381), .A2(n3396), .ZN(n2602) );
  NOR2_X1 U3359 ( .A1(n3958), .A2(n3385), .ZN(n3378) );
  AOI21_X1 U3360 ( .B1(n3823), .B2(n2602), .A(n3378), .ZN(n3825) );
  NAND2_X1 U3361 ( .A1(n2603), .A2(n3825), .ZN(n3913) );
  INV_X1 U3362 ( .A(n3437), .ZN(n3872) );
  OR2_X1 U3363 ( .A1(n3681), .A2(n3498), .ZN(n3831) );
  NAND2_X1 U3364 ( .A1(n3681), .A2(n3498), .ZN(n3830) );
  NAND2_X1 U3365 ( .A1(n3831), .A2(n3830), .ZN(n3875) );
  INV_X1 U3366 ( .A(n3541), .ZN(n3878) );
  NAND2_X1 U3367 ( .A1(n4490), .A2(n3587), .ZN(n3835) );
  AND2_X1 U3368 ( .A1(n3833), .A2(n3835), .ZN(n3914) );
  NAND2_X1 U3369 ( .A1(n3582), .A2(n3914), .ZN(n4355) );
  NAND2_X1 U3370 ( .A1(n3956), .A2(n4387), .ZN(n2604) );
  AND2_X1 U3371 ( .A1(n2604), .A2(n4377), .ZN(n4352) );
  OR2_X1 U3372 ( .A1(n4490), .A2(n3587), .ZN(n3611) );
  NAND2_X1 U3373 ( .A1(n4376), .A2(n3611), .ZN(n2606) );
  NOR2_X1 U3374 ( .A1(n3956), .A2(n4387), .ZN(n2605) );
  AOI21_X1 U3375 ( .B1(n4352), .B2(n2606), .A(n2605), .ZN(n4353) );
  INV_X1 U3376 ( .A(n3955), .ZN(n4463) );
  NAND2_X1 U3377 ( .A1(n4463), .A2(n3890), .ZN(n2607) );
  NAND2_X1 U3378 ( .A1(n4355), .A2(n2608), .ZN(n2611) );
  INV_X1 U3379 ( .A(n2608), .ZN(n3919) );
  OR2_X1 U3380 ( .A1(n3919), .A2(n4352), .ZN(n2610) );
  INV_X1 U3381 ( .A(n3890), .ZN(n4366) );
  NAND2_X1 U3382 ( .A1(n3955), .A2(n4366), .ZN(n2609) );
  OR2_X1 U3383 ( .A1(n4361), .A2(n4336), .ZN(n4292) );
  AND2_X1 U3384 ( .A1(n4294), .A2(n4292), .ZN(n3923) );
  NAND2_X1 U3385 ( .A1(n4328), .A2(n3923), .ZN(n2615) );
  NAND2_X1 U3386 ( .A1(n4441), .A2(n4304), .ZN(n3884) );
  AND2_X1 U3387 ( .A1(n3884), .A2(n2612), .ZN(n3842) );
  AND2_X1 U3388 ( .A1(n4361), .A2(n4336), .ZN(n4291) );
  NAND2_X1 U3389 ( .A1(n4291), .A2(n4294), .ZN(n2613) );
  NAND2_X1 U3390 ( .A1(n3842), .A2(n2613), .ZN(n3924) );
  INV_X1 U3391 ( .A(n3924), .ZN(n2614) );
  NOR2_X1 U3392 ( .A1(n4441), .A2(n4304), .ZN(n3886) );
  INV_X1 U3393 ( .A(n3886), .ZN(n2616) );
  NOR2_X1 U3394 ( .A1(n4300), .A2(n4280), .ZN(n3866) );
  OR2_X1 U3395 ( .A1(n4419), .A2(n4250), .ZN(n2617) );
  OR2_X1 U3396 ( .A1(n4427), .A2(n4267), .ZN(n4238) );
  NAND2_X1 U3397 ( .A1(n2617), .A2(n4238), .ZN(n3928) );
  NAND2_X1 U3398 ( .A1(n4427), .A2(n4267), .ZN(n3883) );
  NAND2_X1 U3399 ( .A1(n4300), .A2(n4280), .ZN(n4259) );
  AND2_X1 U3400 ( .A1(n3883), .A2(n4259), .ZN(n4240) );
  NAND2_X1 U3401 ( .A1(n4419), .A2(n4250), .ZN(n3929) );
  OAI21_X1 U3402 ( .B1(n3928), .B2(n4240), .A(n3929), .ZN(n3846) );
  INV_X1 U3403 ( .A(n3846), .ZN(n2618) );
  XNOR2_X1 U3404 ( .A(n4412), .B(n4418), .ZN(n3931) );
  NOR2_X1 U3405 ( .A1(n4412), .A2(n4231), .ZN(n3849) );
  INV_X1 U3406 ( .A(n3849), .ZN(n2620) );
  NAND2_X1 U3407 ( .A1(n4225), .A2(n2620), .ZN(n4215) );
  INV_X1 U3408 ( .A(n3844), .ZN(n2621) );
  XNOR2_X1 U3409 ( .A(n2622), .B(n3909), .ZN(n2634) );
  INV_X1 U3410 ( .A(n2655), .ZN(n3944) );
  NAND2_X1 U3411 ( .A1(n3944), .A2(n3941), .ZN(n2624) );
  NAND2_X1 U3412 ( .A1(n4190), .A2(n3950), .ZN(n2623) );
  NOR2_X1 U3413 ( .A1(n2626), .A2(n2625), .ZN(n4555) );
  NAND2_X1 U3414 ( .A1(n2627), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  NAND2_X1 U3415 ( .A1(n4564), .A2(n2942), .ZN(n4444) );
  AOI21_X1 U3416 ( .B1(B_REG_SCAN_IN), .B2(n4555), .A(n4444), .ZN(n4202) );
  INV_X1 U3417 ( .A(REG0_REG_30__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U3418 ( .A1(n2630), .A2(REG2_REG_30__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U3419 ( .A1(n3851), .A2(REG1_REG_30__SCAN_IN), .ZN(n2631) );
  OAI211_X1 U3420 ( .C1(n3852), .C2(n2633), .A(n2632), .B(n2631), .ZN(n3954)
         );
  INV_X1 U3421 ( .A(n2942), .ZN(n2635) );
  INV_X1 U3422 ( .A(n3950), .ZN(n2684) );
  INV_X1 U3423 ( .A(n3941), .ZN(n2897) );
  INV_X1 U3424 ( .A(n3859), .ZN(n2636) );
  AOI22_X1 U3425 ( .A1(n4233), .A2(n4440), .B1(n4488), .B2(n2636), .ZN(n2637)
         );
  NOR2_X1 U3426 ( .A1(n2638), .A2(n2649), .ZN(n2639) );
  MUX2_X1 U3427 ( .A(n2649), .B(n2639), .S(IR_REG_25__SCAN_IN), .Z(n2641) );
  NAND2_X1 U3428 ( .A1(n2643), .A2(IR_REG_31__SCAN_IN), .ZN(n2654) );
  NAND2_X1 U3429 ( .A1(n2654), .A2(n2653), .ZN(n2644) );
  NAND2_X1 U3430 ( .A1(n2644), .A2(IR_REG_31__SCAN_IN), .ZN(n2646) );
  INV_X1 U3431 ( .A(n2647), .ZN(n2651) );
  NOR2_X1 U3432 ( .A1(n2640), .A2(n2649), .ZN(n2648) );
  XNOR2_X1 U3433 ( .A(n2654), .B(n2653), .ZN(n2941) );
  NAND2_X1 U3434 ( .A1(n2655), .A2(n4196), .ZN(n2873) );
  NAND2_X1 U3435 ( .A1(n2873), .A2(n2942), .ZN(n3163) );
  OAI211_X1 U3436 ( .C1(n3941), .C2(n4688), .A(n3160), .B(n3163), .ZN(n2656)
         );
  INV_X1 U3437 ( .A(n2656), .ZN(n2671) );
  NOR4_X1 U3438 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_14__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2660) );
  NOR4_X1 U3439 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_10__SCAN_IN), .ZN(n2659) );
  NOR4_X1 U3440 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_24__SCAN_IN), .A3(
        D_REG_26__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2658) );
  NOR4_X1 U3441 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2657) );
  NAND4_X1 U3442 ( .A1(n2660), .A2(n2659), .A3(n2658), .A4(n2657), .ZN(n2668)
         );
  NOR2_X1 U3443 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_23__SCAN_IN), .ZN(n2664)
         );
  NOR4_X1 U3444 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2663) );
  NOR4_X1 U3445 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2662) );
  NOR4_X1 U3446 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2661) );
  NAND4_X1 U3447 ( .A1(n2664), .A2(n2663), .A3(n2662), .A4(n2661), .ZN(n2667)
         );
  NAND2_X1 U3448 ( .A1(n2919), .A2(B_REG_SCAN_IN), .ZN(n2665) );
  INV_X1 U3449 ( .A(n2672), .ZN(n4556) );
  MUX2_X1 U3450 ( .A(n2665), .B(B_REG_SCAN_IN), .S(n4556), .Z(n2666) );
  OAI21_X1 U3451 ( .B1(n2668), .B2(n2667), .A(n2674), .ZN(n2870) );
  INV_X1 U3452 ( .A(D_REG_1__SCAN_IN), .ZN(n2669) );
  NAND2_X1 U3453 ( .A1(n2674), .A2(n2669), .ZN(n2871) );
  INV_X1 U3454 ( .A(n2924), .ZN(n2673) );
  NAND2_X1 U3455 ( .A1(n2673), .A2(n2919), .ZN(n2936) );
  NAND2_X1 U3456 ( .A1(n2871), .A2(n2936), .ZN(n2670) );
  INV_X1 U3457 ( .A(D_REG_0__SCAN_IN), .ZN(n2939) );
  AND2_X1 U34580 ( .A1(n2673), .A2(n2672), .ZN(n2938) );
  INV_X1 U34590 ( .A(n2675), .ZN(n2678) );
  NAND2_X1 U3460 ( .A1(n3185), .A2(n2962), .ZN(n3194) );
  NAND2_X1 U3461 ( .A1(n3233), .A2(n3237), .ZN(n3280) );
  OAI21_X1 U3462 ( .B1(n4208), .B2(n3859), .A(n4399), .ZN(n3625) );
  NAND2_X1 U3463 ( .A1(n2678), .A2(n2246), .ZN(U3547) );
  INV_X1 U3464 ( .A(n2872), .ZN(n3165) );
  NAND2_X1 U3465 ( .A1(n2681), .A2(n2245), .ZN(U3515) );
  INV_X2 U3466 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U34670 ( .A(n3167), .ZN(n2682) );
  AND2_X4 U3468 ( .A1(n2683), .A2(n3167), .ZN(n2815) );
  AND2_X2 U34690 ( .A1(n3167), .A2(n2882), .ZN(n2865) );
  NAND2_X1 U3470 ( .A1(n4693), .A2(n4196), .ZN(n3192) );
  AND2_X2 U34710 ( .A1(n2815), .A2(n3192), .ZN(n2700) );
  AOI22_X1 U3472 ( .A1(n3182), .A2(n2700), .B1(n2856), .B2(n3102), .ZN(n2686)
         );
  INV_X1 U34730 ( .A(n2686), .ZN(n2706) );
  NAND2_X1 U3474 ( .A1(n2691), .A2(n2762), .ZN(n2688) );
  NAND2_X1 U34750 ( .A1(n3197), .A2(n2815), .ZN(n2687) );
  NAND2_X1 U3476 ( .A1(n2688), .A2(n2687), .ZN(n2690) );
  INV_X1 U34770 ( .A(n2690), .ZN(n2695) );
  INV_X1 U3478 ( .A(n2683), .ZN(n2692) );
  NAND2_X1 U34790 ( .A1(n2691), .A2(n2700), .ZN(n2694) );
  AND2_X1 U3480 ( .A1(n2694), .A2(n2693), .ZN(n3009) );
  AOI21_X1 U34810 ( .B1(n2695), .B2(n2865), .A(n3008), .ZN(n3086) );
  XNOR2_X1 U3482 ( .A(n2698), .B(n2697), .ZN(n2701) );
  NOR2_X1 U34830 ( .A1(n3185), .A2(n2760), .ZN(n2699) );
  XNOR2_X1 U3484 ( .A(n2701), .B(n2702), .ZN(n3084) );
  NOR2_X1 U34850 ( .A1(n3086), .A2(n3084), .ZN(n3085) );
  INV_X1 U3486 ( .A(n2701), .ZN(n2704) );
  INV_X1 U34870 ( .A(n2702), .ZN(n2703) );
  NOR2_X1 U3488 ( .A1(n3085), .A2(n2238), .ZN(n3096) );
  NAND2_X1 U34890 ( .A1(n3097), .A2(n3096), .ZN(n3095) );
  NAND2_X1 U3490 ( .A1(n3095), .A2(n2707), .ZN(n3122) );
  OAI22_X1 U34910 ( .A1(n3100), .A2(n2761), .B1(n2763), .B2(n2708), .ZN(n2713)
         );
  NAND2_X1 U3492 ( .A1(n4104), .A2(n2762), .ZN(n2710) );
  NAND2_X1 U34930 ( .A1(n3125), .A2(n2815), .ZN(n2709) );
  NAND2_X1 U3494 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  XNOR2_X1 U34950 ( .A(n2711), .B(n2033), .ZN(n2712) );
  XOR2_X1 U3496 ( .A(n2713), .B(n2712), .Z(n3123) );
  INV_X1 U34970 ( .A(n2712), .ZN(n2715) );
  INV_X1 U3498 ( .A(n2713), .ZN(n2714) );
  NAND2_X1 U34990 ( .A1(n4103), .A2(n2762), .ZN(n2717) );
  NAND2_X1 U3500 ( .A1(n3727), .A2(n2815), .ZN(n2716) );
  NAND2_X1 U35010 ( .A1(n2717), .A2(n2716), .ZN(n2718) );
  XNOR2_X1 U3502 ( .A(n2718), .B(n2033), .ZN(n2720) );
  NOR2_X1 U35030 ( .A1(n3176), .A2(n2763), .ZN(n2719) );
  AOI21_X1 U3504 ( .B1(n4103), .B2(n2700), .A(n2719), .ZN(n2721) );
  XNOR2_X1 U35050 ( .A(n2720), .B(n2721), .ZN(n3724) );
  INV_X1 U35060 ( .A(n2721), .ZN(n2722) );
  OAI22_X1 U35070 ( .A1(n3256), .A2(n2763), .B1(n2867), .B2(n2725), .ZN(n2724)
         );
  XNOR2_X1 U35080 ( .A(n2724), .B(n2033), .ZN(n2727) );
  NOR2_X1 U35090 ( .A1(n2725), .A2(n2763), .ZN(n2726) );
  AOI21_X1 U35100 ( .B1(n4102), .B2(n2861), .A(n2726), .ZN(n2728) );
  XNOR2_X1 U35110 ( .A(n2727), .B(n2728), .ZN(n3691) );
  INV_X1 U35120 ( .A(n2727), .ZN(n2729) );
  INV_X1 U35130 ( .A(n3693), .ZN(n2731) );
  OAI22_X1 U35140 ( .A1(n2731), .A2(n2761), .B1(n2763), .B2(n2730), .ZN(n3201)
         );
  AOI22_X1 U35150 ( .A1(n3693), .A2(n2856), .B1(n2815), .B2(n3251), .ZN(n2732)
         );
  XOR2_X1 U35160 ( .A(n2033), .B(n2732), .Z(n3202) );
  NOR2_X1 U35170 ( .A1(n3237), .A2(n2763), .ZN(n2733) );
  AOI21_X1 U35180 ( .B1(n3274), .B2(n2700), .A(n2733), .ZN(n2735) );
  AOI22_X1 U35190 ( .A1(n3274), .A2(n2856), .B1(n2815), .B2(n3227), .ZN(n2734)
         );
  XNOR2_X1 U35200 ( .A(n2734), .B(n2033), .ZN(n2736) );
  XOR2_X1 U35210 ( .A(n2735), .B(n2736), .Z(n3224) );
  INV_X1 U35220 ( .A(n2735), .ZN(n2738) );
  INV_X1 U35230 ( .A(n2736), .ZN(n2737) );
  NAND2_X1 U35240 ( .A1(n3342), .A2(n2856), .ZN(n2740) );
  NAND2_X1 U35250 ( .A1(n3279), .A2(n2815), .ZN(n2739) );
  NAND2_X1 U35260 ( .A1(n2740), .A2(n2739), .ZN(n2741) );
  XNOR2_X1 U35270 ( .A(n2741), .B(n2865), .ZN(n2743) );
  AOI22_X1 U35280 ( .A1(n3342), .A2(n2861), .B1(n2856), .B2(n3279), .ZN(n2742)
         );
  AND2_X1 U35290 ( .A1(n2743), .A2(n2742), .ZN(n3262) );
  AOI22_X1 U35300 ( .A1(n3962), .A2(n2861), .B1(n2856), .B2(n3343), .ZN(n2747)
         );
  NAND2_X1 U35310 ( .A1(n3962), .A2(n2856), .ZN(n2745) );
  NAND2_X1 U35320 ( .A1(n3343), .A2(n2815), .ZN(n2744) );
  NAND2_X1 U35330 ( .A1(n2745), .A2(n2744), .ZN(n2746) );
  XNOR2_X1 U35340 ( .A(n2746), .B(n2033), .ZN(n2749) );
  XOR2_X1 U35350 ( .A(n2747), .B(n2749), .Z(n3339) );
  INV_X1 U35360 ( .A(n2747), .ZN(n2748) );
  OR2_X1 U35370 ( .A1(n2749), .A2(n2748), .ZN(n2750) );
  INV_X1 U35380 ( .A(n3450), .ZN(n2755) );
  AOI22_X1 U35390 ( .A1(n3961), .A2(n2861), .B1(n2762), .B2(n3455), .ZN(n2757)
         );
  NAND2_X1 U35400 ( .A1(n3961), .A2(n2762), .ZN(n2752) );
  NAND2_X1 U35410 ( .A1(n3455), .A2(n2815), .ZN(n2751) );
  NAND2_X1 U35420 ( .A1(n2752), .A2(n2751), .ZN(n2753) );
  XNOR2_X1 U35430 ( .A(n2753), .B(n2033), .ZN(n2756) );
  XOR2_X1 U35440 ( .A(n2757), .B(n2756), .Z(n3453) );
  NAND2_X1 U35450 ( .A1(n2755), .A2(n2754), .ZN(n3451) );
  INV_X1 U35460 ( .A(n2756), .ZN(n2758) );
  OR2_X1 U35470 ( .A1(n2758), .A2(n2757), .ZN(n2759) );
  NAND2_X1 U35480 ( .A1(n3451), .A2(n2759), .ZN(n3408) );
  INV_X1 U35490 ( .A(n3408), .ZN(n2767) );
  INV_X1 U35500 ( .A(n2762), .ZN(n2760) );
  OAI22_X1 U35510 ( .A1(n3470), .A2(n2761), .B1(n2763), .B2(n3429), .ZN(n3409)
         );
  INV_X1 U35520 ( .A(n3409), .ZN(n2766) );
  OAI22_X1 U35530 ( .A1(n3470), .A2(n2763), .B1(n2867), .B2(n3429), .ZN(n2764)
         );
  XNOR2_X1 U35540 ( .A(n2764), .B(n2033), .ZN(n3410) );
  OAI21_X1 U35550 ( .B1(n2767), .B2(n2766), .A(n2765), .ZN(n3485) );
  NAND2_X1 U35560 ( .A1(n3574), .A2(n2762), .ZN(n2769) );
  NAND2_X1 U35570 ( .A1(n3487), .A2(n2815), .ZN(n2768) );
  NAND2_X1 U35580 ( .A1(n2769), .A2(n2768), .ZN(n2770) );
  XNOR2_X1 U35590 ( .A(n2770), .B(n2865), .ZN(n2772) );
  AOI22_X1 U35600 ( .A1(n3574), .A2(n2700), .B1(n2762), .B2(n3487), .ZN(n2771)
         );
  NOR2_X1 U35610 ( .A1(n2772), .A2(n2771), .ZN(n3481) );
  NAND2_X1 U35620 ( .A1(n2772), .A2(n2771), .ZN(n3482) );
  AOI22_X1 U35630 ( .A1(n3958), .A2(n2762), .B1(n2815), .B2(n3575), .ZN(n2775)
         );
  XOR2_X1 U35640 ( .A(n2033), .B(n2775), .Z(n3571) );
  INV_X1 U35650 ( .A(n3958), .ZN(n3444) );
  OAI22_X1 U35660 ( .A1(n3444), .A2(n2761), .B1(n2763), .B2(n3385), .ZN(n3570)
         );
  NAND2_X1 U35670 ( .A1(n3777), .A2(n2762), .ZN(n2777) );
  NAND2_X1 U35680 ( .A1(n3599), .A2(n2815), .ZN(n2776) );
  NAND2_X1 U35690 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  XNOR2_X1 U35700 ( .A(n2778), .B(n2865), .ZN(n2781) );
  NOR2_X1 U35710 ( .A1(n3507), .A2(n2763), .ZN(n2779) );
  AOI21_X1 U35720 ( .B1(n3777), .B2(n2700), .A(n2779), .ZN(n2780) );
  NAND2_X1 U35730 ( .A1(n2781), .A2(n2780), .ZN(n3596) );
  AOI22_X1 U35740 ( .A1(n3681), .A2(n2762), .B1(n2815), .B2(n3781), .ZN(n2782)
         );
  XNOR2_X1 U35750 ( .A(n2782), .B(n2033), .ZN(n2786) );
  NAND2_X1 U35760 ( .A1(n2785), .A2(n2786), .ZN(n3677) );
  NAND2_X1 U35770 ( .A1(n3681), .A2(n2861), .ZN(n2784) );
  NAND2_X1 U35780 ( .A1(n3781), .A2(n2762), .ZN(n2783) );
  NAND2_X1 U35790 ( .A1(n2784), .A2(n2783), .ZN(n3774) );
  NAND2_X1 U35800 ( .A1(n3677), .A2(n3774), .ZN(n2796) );
  NAND2_X1 U35810 ( .A1(n2788), .A2(n2787), .ZN(n3773) );
  NAND2_X1 U3582 ( .A1(n3957), .A2(n2762), .ZN(n2790) );
  NAND2_X1 U3583 ( .A1(n4487), .A2(n2815), .ZN(n2789) );
  NAND2_X1 U3584 ( .A1(n2790), .A2(n2789), .ZN(n2791) );
  XNOR2_X1 U3585 ( .A(n2791), .B(n2033), .ZN(n2795) );
  NAND2_X1 U3586 ( .A1(n3957), .A2(n2861), .ZN(n2793) );
  NAND2_X1 U3587 ( .A1(n4487), .A2(n2762), .ZN(n2792) );
  NAND2_X1 U3588 ( .A1(n2793), .A2(n2792), .ZN(n2794) );
  NOR2_X1 U3589 ( .A1(n2795), .A2(n2794), .ZN(n2797) );
  AOI21_X1 U3590 ( .B1(n2795), .B2(n2794), .A(n2797), .ZN(n3679) );
  NAND3_X1 U3591 ( .A1(n2796), .A2(n3773), .A3(n3679), .ZN(n2799) );
  INV_X1 U3592 ( .A(n2797), .ZN(n2798) );
  NAND2_X1 U3593 ( .A1(n4490), .A2(n2762), .ZN(n2801) );
  NAND2_X1 U3594 ( .A1(n4478), .A2(n2815), .ZN(n2800) );
  NAND2_X1 U3595 ( .A1(n2801), .A2(n2800), .ZN(n2802) );
  XNOR2_X1 U3596 ( .A(n2802), .B(n2033), .ZN(n2806) );
  NAND2_X1 U3597 ( .A1(n4490), .A2(n2861), .ZN(n2804) );
  NAND2_X1 U3598 ( .A1(n4478), .A2(n2762), .ZN(n2803) );
  NAND2_X1 U3599 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  NAND2_X1 U3600 ( .A1(n2806), .A2(n2805), .ZN(n3700) );
  NOR2_X1 U3601 ( .A1(n2806), .A2(n2805), .ZN(n3702) );
  INV_X1 U3602 ( .A(n4479), .ZN(n2807) );
  OAI22_X1 U3603 ( .A1(n2807), .A2(n2761), .B1(n2763), .B2(n3609), .ZN(n3752)
         );
  AOI22_X1 U3604 ( .A1(n4479), .A2(n2762), .B1(n2815), .B2(n3757), .ZN(n2808)
         );
  XOR2_X1 U3605 ( .A(n2033), .B(n2808), .Z(n3753) );
  NAND2_X1 U3606 ( .A1(n3956), .A2(n2762), .ZN(n2810) );
  NAND2_X1 U3607 ( .A1(n3891), .A2(n2815), .ZN(n2809) );
  NAND2_X1 U3608 ( .A1(n2810), .A2(n2809), .ZN(n2811) );
  XNOR2_X1 U3609 ( .A(n2811), .B(n2865), .ZN(n2813) );
  AOI22_X1 U3610 ( .A1(n3956), .A2(n2861), .B1(n2762), .B2(n3891), .ZN(n2812)
         );
  NAND2_X1 U3611 ( .A1(n2813), .A2(n2812), .ZN(n2814) );
  OAI21_X1 U3612 ( .B1(n2813), .B2(n2812), .A(n2814), .ZN(n3648) );
  NAND2_X1 U3613 ( .A1(n3955), .A2(n2762), .ZN(n2817) );
  NAND2_X1 U3614 ( .A1(n3890), .A2(n2815), .ZN(n2816) );
  NAND2_X1 U3615 ( .A1(n2817), .A2(n2816), .ZN(n2818) );
  XNOR2_X1 U3616 ( .A(n2818), .B(n2033), .ZN(n2821) );
  NAND2_X1 U3617 ( .A1(n3955), .A2(n2861), .ZN(n2820) );
  NAND2_X1 U3618 ( .A1(n3890), .A2(n2762), .ZN(n2819) );
  NAND2_X1 U3619 ( .A1(n2820), .A2(n2819), .ZN(n2822) );
  NAND2_X1 U3620 ( .A1(n2821), .A2(n2822), .ZN(n3733) );
  INV_X1 U3621 ( .A(n2821), .ZN(n2824) );
  INV_X1 U3622 ( .A(n2822), .ZN(n2823) );
  NAND2_X1 U3623 ( .A1(n2824), .A2(n2823), .ZN(n3659) );
  NAND2_X1 U3624 ( .A1(n3737), .A2(n3659), .ZN(n3662) );
  NAND2_X1 U3625 ( .A1(n4361), .A2(n2762), .ZN(n2826) );
  OR2_X1 U3626 ( .A1(n4336), .A2(n2867), .ZN(n2825) );
  NAND2_X1 U3627 ( .A1(n2826), .A2(n2825), .ZN(n2827) );
  XNOR2_X1 U3628 ( .A(n2827), .B(n2865), .ZN(n2829) );
  NOR2_X1 U3629 ( .A1(n4336), .A2(n2763), .ZN(n2828) );
  AOI21_X1 U3630 ( .B1(n4361), .B2(n2861), .A(n2828), .ZN(n2830) );
  AND2_X1 U3631 ( .A1(n2829), .A2(n2830), .ZN(n3655) );
  INV_X1 U3632 ( .A(n2829), .ZN(n2832) );
  INV_X1 U3633 ( .A(n2830), .ZN(n2831) );
  NAND2_X1 U3634 ( .A1(n2832), .A2(n2831), .ZN(n3656) );
  NAND2_X1 U3635 ( .A1(n4460), .A2(n2762), .ZN(n2834) );
  OR2_X1 U3636 ( .A1(n4318), .A2(n2867), .ZN(n2833) );
  NAND2_X1 U3637 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  XNOR2_X1 U3638 ( .A(n2835), .B(n2033), .ZN(n2841) );
  OAI22_X1 U3639 ( .A1(n4298), .A2(n2761), .B1(n2763), .B2(n4318), .ZN(n2840)
         );
  XNOR2_X1 U3640 ( .A(n2841), .B(n2840), .ZN(n3745) );
  NAND2_X1 U3641 ( .A1(n4441), .A2(n2762), .ZN(n2837) );
  OR2_X1 U3642 ( .A1(n4304), .A2(n2867), .ZN(n2836) );
  NAND2_X1 U3643 ( .A1(n2837), .A2(n2836), .ZN(n2838) );
  XNOR2_X1 U3644 ( .A(n2838), .B(n2865), .ZN(n2844) );
  NOR2_X1 U3645 ( .A1(n4304), .A2(n2763), .ZN(n2839) );
  AOI21_X1 U3646 ( .B1(n4441), .B2(n2861), .A(n2839), .ZN(n2843) );
  XNOR2_X1 U3647 ( .A(n2844), .B(n2843), .ZN(n3638) );
  NOR2_X1 U3648 ( .A1(n2841), .A2(n2840), .ZN(n3639) );
  NOR2_X1 U3649 ( .A1(n3638), .A2(n3639), .ZN(n2842) );
  OR2_X1 U3650 ( .A1(n2844), .A2(n2843), .ZN(n2848) );
  NOR2_X1 U3651 ( .A1(n4280), .A2(n2763), .ZN(n2845) );
  AOI21_X1 U3652 ( .B1(n4300), .B2(n2861), .A(n2845), .ZN(n2847) );
  INV_X1 U3653 ( .A(n2847), .ZN(n2846) );
  OAI22_X1 U3654 ( .A1(n4263), .A2(n2763), .B1(n2867), .B2(n4280), .ZN(n2849)
         );
  XNOR2_X1 U3655 ( .A(n2849), .B(n2033), .ZN(n3714) );
  NAND2_X1 U3656 ( .A1(n3711), .A2(n3714), .ZN(n2850) );
  NAND2_X1 U3657 ( .A1(n3712), .A2(n2850), .ZN(n3671) );
  NOR2_X1 U3658 ( .A1(n4267), .A2(n2867), .ZN(n2851) );
  AOI21_X1 U3659 ( .B1(n4427), .B2(n2762), .A(n2851), .ZN(n2852) );
  XNOR2_X1 U3660 ( .A(n2852), .B(n2033), .ZN(n2855) );
  NOR2_X1 U3661 ( .A1(n4267), .A2(n2763), .ZN(n2853) );
  AOI21_X1 U3662 ( .B1(n4427), .B2(n2861), .A(n2853), .ZN(n2854) );
  NAND2_X1 U3663 ( .A1(n2855), .A2(n2854), .ZN(n3668) );
  NOR2_X1 U3664 ( .A1(n2855), .A2(n2854), .ZN(n3669) );
  NAND2_X1 U3665 ( .A1(n4419), .A2(n2762), .ZN(n2858) );
  OR2_X1 U3666 ( .A1(n4250), .A2(n2867), .ZN(n2857) );
  NAND2_X1 U3667 ( .A1(n2858), .A2(n2857), .ZN(n2859) );
  XNOR2_X1 U3668 ( .A(n2859), .B(n2865), .ZN(n2863) );
  NOR2_X1 U3669 ( .A1(n4250), .A2(n2763), .ZN(n2860) );
  AOI21_X1 U3670 ( .B1(n4419), .B2(n2861), .A(n2860), .ZN(n2862) );
  OR2_X1 U3671 ( .A1(n2863), .A2(n2862), .ZN(n3764) );
  OAI22_X1 U3672 ( .A1(n4430), .A2(n2761), .B1(n4231), .B2(n2763), .ZN(n2877)
         );
  OAI22_X1 U3673 ( .A1(n4430), .A2(n2763), .B1(n4231), .B2(n2867), .ZN(n2864)
         );
  XNOR2_X1 U3674 ( .A(n2864), .B(n2033), .ZN(n2878) );
  XOR2_X1 U3675 ( .A(n2877), .B(n2878), .Z(n3631) );
  OAI22_X1 U3676 ( .A1(n4421), .A2(n2761), .B1(n2763), .B2(n4408), .ZN(n2866)
         );
  XNOR2_X1 U3677 ( .A(n2866), .B(n2865), .ZN(n2869) );
  OAI22_X1 U3678 ( .A1(n4421), .A2(n2763), .B1(n2867), .B2(n4408), .ZN(n2868)
         );
  XNOR2_X1 U3679 ( .A(n2869), .B(n2868), .ZN(n2880) );
  INV_X1 U3680 ( .A(n2880), .ZN(n2875) );
  AND2_X1 U3681 ( .A1(n2870), .A2(n2936), .ZN(n3164) );
  AOI21_X1 U3682 ( .B1(n2873), .B2(n2963), .A(n2942), .ZN(n2886) );
  AND2_X1 U3683 ( .A1(n3160), .A2(n2886), .ZN(n2874) );
  NAND2_X1 U3684 ( .A1(n2875), .A2(n3787), .ZN(n2876) );
  NAND2_X1 U3685 ( .A1(n2878), .A2(n2877), .ZN(n2879) );
  INV_X1 U3686 ( .A(n2879), .ZN(n2881) );
  NAND3_X1 U3687 ( .A1(n2881), .A2(n3787), .A3(n2875), .ZN(n2903) );
  INV_X1 U3688 ( .A(n2882), .ZN(n2883) );
  NAND2_X1 U3689 ( .A1(n2883), .A2(n4675), .ZN(n2884) );
  INV_X1 U3690 ( .A(n4564), .ZN(n2970) );
  NOR2_X1 U3691 ( .A1(n2893), .A2(n2970), .ZN(n2885) );
  AND2_X2 U3692 ( .A1(n2896), .A2(n2885), .ZN(n3779) );
  INV_X1 U3693 ( .A(n2896), .ZN(n2891) );
  INV_X1 U3694 ( .A(n2886), .ZN(n2887) );
  NAND2_X1 U3695 ( .A1(n2887), .A2(n4409), .ZN(n2888) );
  NAND2_X1 U3696 ( .A1(n2891), .A2(n2888), .ZN(n2889) );
  NAND2_X1 U3697 ( .A1(n2889), .A2(n3163), .ZN(n3005) );
  NAND2_X1 U3698 ( .A1(n2683), .A2(n2941), .ZN(n2890) );
  OAI21_X1 U3699 ( .B1(n3005), .B2(n2890), .A(STATE_REG_SCAN_IN), .ZN(n2892)
         );
  INV_X1 U3700 ( .A(n2893), .ZN(n3948) );
  NAND2_X1 U3701 ( .A1(n2891), .A2(n3948), .ZN(n3003) );
  AND2_X2 U3702 ( .A1(n2892), .A2(n3003), .ZN(n3785) );
  NOR2_X1 U3703 ( .A1(n4213), .A2(n3785), .ZN(n2901) );
  NOR2_X1 U3704 ( .A1(n2893), .A2(n4564), .ZN(n2894) );
  NAND2_X1 U3705 ( .A1(n2896), .A2(n2894), .ZN(n3715) );
  AND2_X1 U3706 ( .A1(n3160), .A2(n4488), .ZN(n2895) );
  NAND2_X1 U3707 ( .A1(n2896), .A2(n2895), .ZN(n2898) );
  AOI22_X1 U3708 ( .A1(n3780), .A2(n4210), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2899) );
  OAI21_X1 U3709 ( .B1(n4430), .B2(n3715), .A(n2899), .ZN(n2900) );
  AOI211_X1 U3710 ( .C1(n3779), .C2(n4407), .A(n2901), .B(n2900), .ZN(n2902)
         );
  AOI21_X1 U3711 ( .B1(n2905), .B2(n2237), .A(n2904), .ZN(n2906) );
  NAND2_X1 U3712 ( .A1(n2907), .A2(n2906), .ZN(U3217) );
  INV_X1 U3713 ( .A(n4675), .ZN(n2908) );
  NOR2_X1 U3714 ( .A1(n2683), .A2(n2908), .ZN(U4043) );
  MUX2_X1 U3715 ( .A(n3031), .B(n2344), .S(U3149), .Z(n2909) );
  INV_X1 U3716 ( .A(n2909), .ZN(U3347) );
  INV_X1 U3717 ( .A(DATAI_3_), .ZN(n2910) );
  INV_X1 U3718 ( .A(n2989), .ZN(n2977) );
  MUX2_X1 U3719 ( .A(n2910), .B(n2977), .S(STATE_REG_SCAN_IN), .Z(n2911) );
  INV_X1 U3720 ( .A(n2911), .ZN(U3349) );
  MUX2_X1 U3721 ( .A(n2369), .B(n3050), .S(STATE_REG_SCAN_IN), .Z(n2912) );
  INV_X1 U3722 ( .A(n2912), .ZN(U3345) );
  INV_X1 U3723 ( .A(DATAI_21_), .ZN(n2914) );
  NAND2_X1 U3724 ( .A1(n3941), .A2(STATE_REG_SCAN_IN), .ZN(n2913) );
  OAI21_X1 U3725 ( .B1(STATE_REG_SCAN_IN), .B2(n2914), .A(n2913), .ZN(U3331)
         );
  INV_X1 U3726 ( .A(DATAI_22_), .ZN(n2916) );
  NAND2_X1 U3727 ( .A1(n3950), .A2(STATE_REG_SCAN_IN), .ZN(n2915) );
  OAI21_X1 U3728 ( .B1(STATE_REG_SCAN_IN), .B2(n2916), .A(n2915), .ZN(U3330)
         );
  INV_X1 U3729 ( .A(DATAI_15_), .ZN(n2918) );
  NAND2_X1 U3730 ( .A1(n3534), .A2(STATE_REG_SCAN_IN), .ZN(n2917) );
  OAI21_X1 U3731 ( .B1(STATE_REG_SCAN_IN), .B2(n2918), .A(n2917), .ZN(U3337)
         );
  INV_X1 U3732 ( .A(DATAI_25_), .ZN(n2922) );
  INV_X1 U3733 ( .A(n2919), .ZN(n2920) );
  NAND2_X1 U3734 ( .A1(n2920), .A2(STATE_REG_SCAN_IN), .ZN(n2921) );
  OAI21_X1 U3735 ( .B1(STATE_REG_SCAN_IN), .B2(n2922), .A(n2921), .ZN(U3327)
         );
  INV_X1 U3736 ( .A(n4164), .ZN(n4189) );
  NAND2_X1 U3737 ( .A1(n4189), .A2(STATE_REG_SCAN_IN), .ZN(n2923) );
  OAI21_X1 U3738 ( .B1(STATE_REG_SCAN_IN), .B2(n2499), .A(n2923), .ZN(U3334)
         );
  INV_X1 U3739 ( .A(DATAI_26_), .ZN(n2926) );
  NAND2_X1 U3740 ( .A1(n2924), .A2(STATE_REG_SCAN_IN), .ZN(n2925) );
  OAI21_X1 U3741 ( .B1(STATE_REG_SCAN_IN), .B2(n2926), .A(n2925), .ZN(U3326)
         );
  INV_X1 U3742 ( .A(DATAI_29_), .ZN(n4008) );
  NAND2_X1 U3743 ( .A1(n2927), .A2(STATE_REG_SCAN_IN), .ZN(n2928) );
  OAI21_X1 U3744 ( .B1(STATE_REG_SCAN_IN), .B2(n4008), .A(n2928), .ZN(U3323)
         );
  NAND2_X1 U3745 ( .A1(n3944), .A2(STATE_REG_SCAN_IN), .ZN(n2929) );
  OAI21_X1 U3746 ( .B1(STATE_REG_SCAN_IN), .B2(n2516), .A(n2929), .ZN(U3332)
         );
  INV_X1 U3747 ( .A(DATAI_30_), .ZN(n2932) );
  NAND2_X1 U3748 ( .A1(n2930), .A2(STATE_REG_SCAN_IN), .ZN(n2931) );
  OAI21_X1 U3749 ( .B1(STATE_REG_SCAN_IN), .B2(n2932), .A(n2931), .ZN(U3322)
         );
  INV_X1 U3750 ( .A(DATAI_19_), .ZN(n2933) );
  MUX2_X1 U3751 ( .A(n2933), .B(n4196), .S(STATE_REG_SCAN_IN), .Z(n2934) );
  INV_X1 U3752 ( .A(n2934), .ZN(U3333) );
  INV_X1 U3753 ( .A(n2936), .ZN(n2937) );
  AOI22_X1 U3754 ( .A1(n4674), .A2(n2669), .B1(n2937), .B2(n4675), .ZN(U3459)
         );
  AOI22_X1 U3755 ( .A1(n4674), .A2(n2939), .B1(n2938), .B2(n4675), .ZN(U3458)
         );
  OR2_X1 U3756 ( .A1(n2941), .A2(U3149), .ZN(n3952) );
  INV_X1 U3757 ( .A(n3952), .ZN(n2940) );
  OR2_X1 U3758 ( .A1(n3160), .A2(n2940), .ZN(n2969) );
  AND2_X1 U3759 ( .A1(n2942), .A2(n2941), .ZN(n2943) );
  NOR2_X1 U3760 ( .A1(n3857), .A2(n2943), .ZN(n2968) );
  INV_X1 U3761 ( .A(n2968), .ZN(n2944) );
  NAND2_X1 U3762 ( .A1(n2969), .A2(n2944), .ZN(n4167) );
  NOR2_X1 U3763 ( .A1(n4626), .A2(n3960), .ZN(U3148) );
  CLKBUF_X2 U3764 ( .A(U4043), .Z(n3960) );
  INV_X1 U3765 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n2947) );
  NAND2_X1 U3766 ( .A1(n3182), .A2(n3960), .ZN(n2946) );
  OAI21_X1 U3767 ( .B1(n3960), .B2(n2947), .A(n2946), .ZN(U3552) );
  INV_X1 U3768 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n2949) );
  NAND2_X1 U3769 ( .A1(n3777), .A2(n3960), .ZN(n2948) );
  OAI21_X1 U3770 ( .B1(n3960), .B2(n2949), .A(n2948), .ZN(U3564) );
  INV_X1 U3771 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n2951) );
  NAND2_X1 U3772 ( .A1(n4479), .A2(n3960), .ZN(n2950) );
  OAI21_X1 U3773 ( .B1(n3960), .B2(n2951), .A(n2950), .ZN(U3568) );
  INV_X1 U3774 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n2953) );
  NAND2_X1 U3775 ( .A1(n3574), .A2(n3960), .ZN(n2952) );
  OAI21_X1 U3776 ( .B1(n3960), .B2(n2953), .A(n2952), .ZN(U3562) );
  INV_X1 U3777 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n2955) );
  NAND2_X1 U3778 ( .A1(n3681), .A2(n3960), .ZN(n2954) );
  OAI21_X1 U3779 ( .B1(n3960), .B2(n2955), .A(n2954), .ZN(U3565) );
  INV_X1 U3780 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n2957) );
  NAND2_X1 U3781 ( .A1(n3342), .A2(n3960), .ZN(n2956) );
  OAI21_X1 U3782 ( .B1(n3960), .B2(n2957), .A(n2956), .ZN(U3558) );
  INV_X1 U3783 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n2959) );
  NAND2_X1 U3784 ( .A1(n3274), .A2(n3960), .ZN(n2958) );
  OAI21_X1 U3785 ( .B1(n3960), .B2(n2959), .A(n2958), .ZN(U3557) );
  INV_X1 U3786 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n2961) );
  NAND2_X1 U3787 ( .A1(n3693), .A2(n3960), .ZN(n2960) );
  OAI21_X1 U3788 ( .B1(n3960), .B2(n2961), .A(n2960), .ZN(U3556) );
  NAND2_X1 U3789 ( .A1(n2691), .A2(n2962), .ZN(n3792) );
  NAND2_X1 U3790 ( .A1(n3790), .A2(n3792), .ZN(n4660) );
  AND2_X1 U3791 ( .A1(n3197), .A2(n2963), .ZN(n4658) );
  INV_X1 U3792 ( .A(n2696), .ZN(n3099) );
  INV_X1 U3793 ( .A(n4363), .ZN(n3424) );
  OAI21_X1 U3794 ( .B1(n3424), .B2(n4329), .A(n4660), .ZN(n2964) );
  OAI21_X1 U3795 ( .B1(n3099), .B2(n4444), .A(n2964), .ZN(n4656) );
  AOI211_X1 U3796 ( .C1(n4698), .C2(n4660), .A(n4658), .B(n4656), .ZN(n4687)
         );
  NAND2_X1 U3797 ( .A1(n4711), .A2(REG1_REG_0__SCAN_IN), .ZN(n2965) );
  OAI21_X1 U3798 ( .B1(n4687), .B2(n4711), .A(n2965), .ZN(U3518) );
  INV_X1 U3799 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4134) );
  AND2_X1 U3800 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4124)
         );
  INV_X1 U3801 ( .A(n2974), .ZN(n4563) );
  NAND2_X1 U3802 ( .A1(n4563), .A2(REG2_REG_1__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U3803 ( .A1(n4137), .A2(n4136), .ZN(n2967) );
  MUX2_X1 U3804 ( .A(n4134), .B(REG2_REG_2__SCAN_IN), .S(n4133), .Z(n2966) );
  NAND2_X1 U3805 ( .A1(n2967), .A2(n2966), .ZN(n4139) );
  OAI21_X1 U3806 ( .B1(n4134), .B2(n4133), .A(n4139), .ZN(n2983) );
  XNOR2_X1 U3807 ( .A(n2984), .B(REG2_REG_3__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U3808 ( .A1(n2969), .A2(n2968), .ZN(n2978) );
  AND2_X1 U3809 ( .A1(n2970), .A2(n4555), .ZN(n4125) );
  INV_X1 U3810 ( .A(n4125), .ZN(n2971) );
  INV_X1 U3811 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4644) );
  NOR2_X1 U3812 ( .A1(STATE_REG_SCAN_IN), .A2(n4644), .ZN(n3124) );
  INV_X1 U3813 ( .A(n2978), .ZN(n4109) );
  NOR2_X1 U3814 ( .A1(n4633), .A2(n2977), .ZN(n2972) );
  AOI211_X1 U3815 ( .C1(n4626), .C2(ADDR_REG_3__SCAN_IN), .A(n3124), .B(n2972), 
        .ZN(n2981) );
  INV_X1 U3816 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2973) );
  MUX2_X1 U3817 ( .A(n2973), .B(REG1_REG_2__SCAN_IN), .S(n4133), .Z(n4142) );
  XNOR2_X1 U3818 ( .A(n2974), .B(REG1_REG_1__SCAN_IN), .ZN(n4117) );
  AND2_X1 U3819 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4116)
         );
  NAND2_X1 U3820 ( .A1(n4117), .A2(n4116), .ZN(n4115) );
  NAND2_X1 U3821 ( .A1(n4563), .A2(REG1_REG_1__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3822 ( .A1(n4115), .A2(n2975), .ZN(n4141) );
  NAND2_X1 U3823 ( .A1(n4142), .A2(n4141), .ZN(n4140) );
  INV_X1 U3824 ( .A(n4133), .ZN(n4562) );
  NAND2_X1 U3825 ( .A1(n4562), .A2(REG1_REG_2__SCAN_IN), .ZN(n2976) );
  XNOR2_X1 U3826 ( .A(n2990), .B(n2977), .ZN(n2979) );
  NOR2_X2 U3827 ( .A1(n2978), .A2(n4555), .ZN(n4627) );
  OAI211_X1 U3828 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2979), .A(n4627), .B(n2992), 
        .ZN(n2980) );
  OAI211_X1 U3829 ( .C1(n2982), .C2(n4620), .A(n2981), .B(n2980), .ZN(U3243)
         );
  INV_X1 U3830 ( .A(n3031), .ZN(n2987) );
  INV_X1 U3831 ( .A(n2993), .ZN(n4561) );
  INV_X1 U3832 ( .A(n2985), .ZN(n2986) );
  INV_X1 U3833 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4019) );
  MUX2_X1 U3834 ( .A(REG2_REG_5__SCAN_IN), .B(n4019), .S(n3031), .Z(n3028) );
  NOR2_X1 U3835 ( .A1(n3029), .A2(n3028), .ZN(n3027) );
  AOI21_X1 U3836 ( .B1(n2987), .B2(REG2_REG_5__SCAN_IN), .A(n3027), .ZN(n3017)
         );
  XNOR2_X1 U3837 ( .A(n3018), .B(REG2_REG_6__SCAN_IN), .ZN(n3002) );
  AND2_X1 U3838 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3204) );
  INV_X1 U3839 ( .A(n4560), .ZN(n2998) );
  NOR2_X1 U3840 ( .A1(n4633), .A2(n2998), .ZN(n2988) );
  AOI211_X1 U3841 ( .C1(n4626), .C2(ADDR_REG_6__SCAN_IN), .A(n3204), .B(n2988), 
        .ZN(n3001) );
  NAND2_X1 U3842 ( .A1(n2990), .A2(n2989), .ZN(n2991) );
  NAND2_X1 U3843 ( .A1(n2994), .A2(n4561), .ZN(n2995) );
  NAND2_X1 U3844 ( .A1(n4151), .A2(n2995), .ZN(n3035) );
  XNOR2_X1 U3845 ( .A(n3031), .B(REG1_REG_5__SCAN_IN), .ZN(n3036) );
  NAND2_X1 U3846 ( .A1(n3035), .A2(n3036), .ZN(n3034) );
  INV_X1 U3847 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2996) );
  OR2_X1 U3848 ( .A1(n3031), .A2(n2996), .ZN(n2997) );
  OAI211_X1 U3849 ( .C1(n2999), .C2(REG1_REG_6__SCAN_IN), .A(n4627), .B(n3015), 
        .ZN(n3000) );
  OAI211_X1 U3850 ( .C1(n3002), .C2(n4620), .A(n3001), .B(n3000), .ZN(U3246)
         );
  INV_X1 U3851 ( .A(n3003), .ZN(n3006) );
  INV_X1 U3852 ( .A(n3160), .ZN(n3004) );
  NOR3_X1 U3853 ( .A1(n3006), .A2(n3005), .A3(n3004), .ZN(n3105) );
  AOI21_X1 U3854 ( .B1(n3009), .B2(n3007), .A(n3008), .ZN(n4123) );
  NAND2_X1 U3855 ( .A1(n4123), .A2(n3787), .ZN(n3011) );
  AOI22_X1 U3856 ( .A1(n3197), .A2(n3780), .B1(n3779), .B2(n2696), .ZN(n3010)
         );
  OAI211_X1 U3857 ( .C1(n3105), .C2(n3012), .A(n3011), .B(n3010), .ZN(U3229)
         );
  NAND2_X1 U3858 ( .A1(n3013), .A2(n4560), .ZN(n3014) );
  INV_X1 U3859 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3016) );
  OR2_X1 U3860 ( .A1(n3050), .A2(n3016), .ZN(n3043) );
  AND2_X1 U3861 ( .A1(n3050), .A2(n3016), .ZN(n3042) );
  XNOR2_X1 U3862 ( .A(n3060), .B(REG1_REG_8__SCAN_IN), .ZN(n3024) );
  INV_X1 U3863 ( .A(n4627), .ZN(n4200) );
  INV_X1 U3864 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3241) );
  MUX2_X1 U3865 ( .A(REG2_REG_7__SCAN_IN), .B(n3241), .S(n3050), .Z(n3040) );
  XNOR2_X1 U3866 ( .A(n3054), .B(n4559), .ZN(n3056) );
  XOR2_X1 U3867 ( .A(REG2_REG_8__SCAN_IN), .B(n3056), .Z(n3019) );
  NAND2_X1 U3868 ( .A1(n4593), .A2(n3019), .ZN(n3020) );
  NAND2_X1 U3869 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3265) );
  NAND2_X1 U3870 ( .A1(n3020), .A2(n3265), .ZN(n3021) );
  AOI21_X1 U3871 ( .B1(n4626), .B2(ADDR_REG_8__SCAN_IN), .A(n3021), .ZN(n3023)
         );
  INV_X1 U3872 ( .A(n4633), .ZN(n4180) );
  NAND2_X1 U3873 ( .A1(n4180), .A2(n4559), .ZN(n3022) );
  OAI211_X1 U3874 ( .C1(n3024), .C2(n4200), .A(n3023), .B(n3022), .ZN(U3248)
         );
  INV_X1 U3875 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n3026) );
  NAND2_X1 U3876 ( .A1(n4419), .A2(n3960), .ZN(n3025) );
  OAI21_X1 U3877 ( .B1(n3960), .B2(n3026), .A(n3025), .ZN(U3576) );
  AOI211_X1 U3878 ( .C1(n3029), .C2(n3028), .A(n3027), .B(n4620), .ZN(n3033)
         );
  AND2_X1 U3879 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3692) );
  AOI21_X1 U3880 ( .B1(n4626), .B2(ADDR_REG_5__SCAN_IN), .A(n3692), .ZN(n3030)
         );
  OAI21_X1 U3881 ( .B1(n4633), .B2(n3031), .A(n3030), .ZN(n3032) );
  NOR2_X1 U3882 ( .A1(n3033), .A2(n3032), .ZN(n3038) );
  OAI211_X1 U3883 ( .C1(n3036), .C2(n3035), .A(n4627), .B(n3034), .ZN(n3037)
         );
  NAND2_X1 U3884 ( .A1(n3038), .A2(n3037), .ZN(U3245) );
  AOI211_X1 U3885 ( .C1(n3041), .C2(n3040), .A(n4620), .B(n3039), .ZN(n3053)
         );
  INV_X1 U3886 ( .A(n3042), .ZN(n3044) );
  NAND2_X1 U3887 ( .A1(n3044), .A2(n3043), .ZN(n3046) );
  OAI21_X1 U3888 ( .B1(n3047), .B2(n3046), .A(n4627), .ZN(n3045) );
  AOI21_X1 U3889 ( .B1(n3047), .B2(n3046), .A(n3045), .ZN(n3052) );
  NOR2_X1 U3890 ( .A1(STATE_REG_SCAN_IN), .A2(n3048), .ZN(n3226) );
  AOI21_X1 U3891 ( .B1(n4626), .B2(ADDR_REG_7__SCAN_IN), .A(n3226), .ZN(n3049)
         );
  OAI21_X1 U3892 ( .B1(n4633), .B2(n3050), .A(n3049), .ZN(n3051) );
  OR3_X1 U3893 ( .A1(n3053), .A2(n3052), .A3(n3051), .ZN(U3247) );
  INV_X1 U3894 ( .A(n3054), .ZN(n3055) );
  INV_X1 U3895 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3300) );
  MUX2_X1 U3896 ( .A(REG2_REG_9__SCAN_IN), .B(n3300), .S(n3329), .Z(n3057) );
  AOI211_X1 U3897 ( .C1(n3058), .C2(n3057), .A(n4620), .B(n3328), .ZN(n3067)
         );
  INV_X1 U3898 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3061) );
  MUX2_X1 U3899 ( .A(REG1_REG_9__SCAN_IN), .B(n3061), .S(n3329), .Z(n3062) );
  AOI211_X1 U3900 ( .C1(n3063), .C2(n3062), .A(n4200), .B(n3311), .ZN(n3066)
         );
  AND2_X1 U3901 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3341) );
  AOI21_X1 U3902 ( .B1(n4626), .B2(ADDR_REG_9__SCAN_IN), .A(n3341), .ZN(n3064)
         );
  OAI21_X1 U3903 ( .B1(n4633), .B2(n3329), .A(n3064), .ZN(n3065) );
  OR3_X1 U3904 ( .A1(n3067), .A2(n3066), .A3(n3065), .ZN(U3249) );
  OAI21_X1 U3905 ( .B1(n3870), .B2(n3069), .A(n3068), .ZN(n3074) );
  NAND2_X1 U3906 ( .A1(n4104), .A2(n4489), .ZN(n3071) );
  NAND2_X1 U3907 ( .A1(n2696), .A2(n4440), .ZN(n3070) );
  OAI211_X1 U3908 ( .C1(n4409), .C2(n3072), .A(n3071), .B(n3070), .ZN(n3073)
         );
  AOI21_X1 U3909 ( .B1(n3074), .B2(n4329), .A(n3073), .ZN(n3079) );
  OAI21_X1 U3910 ( .B1(n3077), .B2(n3076), .A(n3075), .ZN(n4652) );
  NAND2_X1 U3911 ( .A1(n4652), .A2(n3424), .ZN(n3078) );
  AND2_X1 U3912 ( .A1(n3079), .A2(n3078), .ZN(n4655) );
  NAND2_X1 U3913 ( .A1(n4652), .A2(n4698), .ZN(n3080) );
  NAND2_X1 U3914 ( .A1(n4655), .A2(n3080), .ZN(n3106) );
  INV_X1 U3915 ( .A(n3106), .ZN(n3083) );
  AND2_X1 U3916 ( .A1(n3194), .A2(n3102), .ZN(n3081) );
  NOR2_X1 U3917 ( .A1(n3117), .A2(n3081), .ZN(n4650) );
  AOI22_X1 U3918 ( .A1(n4505), .A2(n4650), .B1(REG0_REG_2__SCAN_IN), .B2(n2136), .ZN(n3082) );
  OAI21_X1 U3919 ( .B1(n3083), .B2(n2136), .A(n3082), .ZN(U3471) );
  AOI211_X1 U3920 ( .C1(n3086), .C2(n3084), .A(n3771), .B(n3085), .ZN(n3087)
         );
  INV_X1 U3921 ( .A(n3087), .ZN(n3093) );
  INV_X1 U3922 ( .A(n3780), .ZN(n3088) );
  INV_X1 U3923 ( .A(n3088), .ZN(n3682) );
  INV_X1 U3924 ( .A(n3779), .ZN(n3717) );
  INV_X1 U3925 ( .A(n3182), .ZN(n3090) );
  INV_X1 U3926 ( .A(n2691), .ZN(n3089) );
  OAI22_X1 U3927 ( .A1(n3717), .A2(n3090), .B1(n3089), .B2(n3715), .ZN(n3091)
         );
  AOI21_X1 U3928 ( .B1(n3196), .B2(n3682), .A(n3091), .ZN(n3092) );
  OAI211_X1 U3929 ( .C1(n3105), .C2(n3094), .A(n3093), .B(n3092), .ZN(U3219)
         );
  OAI21_X1 U3930 ( .B1(n3097), .B2(n3096), .A(n3095), .ZN(n3098) );
  NAND2_X1 U3931 ( .A1(n3098), .A2(n3787), .ZN(n3104) );
  OAI22_X1 U3932 ( .A1(n3717), .A2(n3100), .B1(n3099), .B2(n3715), .ZN(n3101)
         );
  AOI21_X1 U3933 ( .B1(n3102), .B2(n3780), .A(n3101), .ZN(n3103) );
  OAI211_X1 U3934 ( .C1(n3105), .C2(n4129), .A(n3104), .B(n3103), .ZN(U3234)
         );
  MUX2_X1 U3935 ( .A(n3106), .B(REG1_REG_2__SCAN_IN), .S(n4711), .Z(n3107) );
  AOI21_X1 U3936 ( .B1(n4401), .B2(n4650), .A(n3107), .ZN(n3108) );
  INV_X1 U3937 ( .A(n3108), .ZN(U3520) );
  XNOR2_X1 U3938 ( .A(n3110), .B(n3109), .ZN(n4646) );
  INV_X1 U3939 ( .A(n4103), .ZN(n3137) );
  XNOR2_X1 U3940 ( .A(n3111), .B(n3877), .ZN(n3112) );
  NAND2_X1 U3941 ( .A1(n3112), .A2(n4329), .ZN(n3114) );
  AOI22_X1 U3942 ( .A1(n3182), .A2(n4440), .B1(n4488), .B2(n3125), .ZN(n3113)
         );
  OAI211_X1 U3943 ( .C1(n3137), .C2(n4444), .A(n3114), .B(n3113), .ZN(n3115)
         );
  AOI21_X1 U3944 ( .B1(n3424), .B2(n4646), .A(n3115), .ZN(n4649) );
  INV_X1 U3945 ( .A(n4649), .ZN(n3116) );
  AOI21_X1 U3946 ( .B1(n4698), .B2(n4646), .A(n3116), .ZN(n3121) );
  INV_X1 U3947 ( .A(n3117), .ZN(n3118) );
  AOI21_X1 U3948 ( .B1(n3125), .B2(n3118), .A(n2066), .ZN(n4645) );
  AOI22_X1 U3949 ( .A1(n4645), .A2(n4505), .B1(REG0_REG_3__SCAN_IN), .B2(n2136), .ZN(n3119) );
  OAI21_X1 U3950 ( .B1(n3121), .B2(n2136), .A(n3119), .ZN(U3473) );
  AOI22_X1 U3951 ( .A1(n4645), .A2(n4401), .B1(REG1_REG_3__SCAN_IN), .B2(n4711), .ZN(n3120) );
  OAI21_X1 U3952 ( .B1(n3121), .B2(n4711), .A(n3120), .ZN(U3521) );
  XNOR2_X1 U3953 ( .A(n3122), .B(n3123), .ZN(n3129) );
  AOI21_X1 U3954 ( .B1(n3778), .B2(n3182), .A(n3124), .ZN(n3127) );
  AOI22_X1 U3955 ( .A1(n3125), .A2(n3780), .B1(n3779), .B2(n4103), .ZN(n3126)
         );
  OAI211_X1 U3956 ( .C1(n3785), .C2(REG3_REG_3__SCAN_IN), .A(n3127), .B(n3126), 
        .ZN(n3128) );
  AOI21_X1 U3957 ( .B1(n3129), .B2(n3787), .A(n3128), .ZN(n3130) );
  INV_X1 U3958 ( .A(n3130), .ZN(U3215) );
  NAND2_X1 U3959 ( .A1(n3807), .A2(n3803), .ZN(n3894) );
  OR2_X1 U3960 ( .A1(n3131), .A2(n3871), .ZN(n3159) );
  NAND2_X1 U3961 ( .A1(n3159), .A2(n3132), .ZN(n3133) );
  XOR2_X1 U3962 ( .A(n3894), .B(n3133), .Z(n3297) );
  XNOR2_X1 U3963 ( .A(n3134), .B(n3894), .ZN(n3135) );
  NAND2_X1 U3964 ( .A1(n3135), .A2(n4329), .ZN(n3294) );
  AOI22_X1 U3965 ( .A1(n3693), .A2(n4489), .B1(n4488), .B2(n3694), .ZN(n3136)
         );
  OAI211_X1 U3966 ( .C1(n3137), .C2(n4492), .A(n3294), .B(n3136), .ZN(n3138)
         );
  AOI21_X1 U3967 ( .B1(n3297), .B2(n4700), .A(n3138), .ZN(n3145) );
  AND2_X1 U3968 ( .A1(n3175), .A2(n3694), .ZN(n3139) );
  NOR2_X1 U3969 ( .A1(n3152), .A2(n3139), .ZN(n3289) );
  NOR2_X1 U3970 ( .A1(n4706), .A2(n3140), .ZN(n3141) );
  AOI21_X1 U3971 ( .B1(n3289), .B2(n4505), .A(n3141), .ZN(n3142) );
  OAI21_X1 U3972 ( .B1(n3145), .B2(n2136), .A(n3142), .ZN(U3477) );
  NAND2_X1 U3973 ( .A1(n4711), .A2(REG1_REG_5__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U3974 ( .A1(n3289), .A2(n4401), .ZN(n3143) );
  OAI211_X1 U3975 ( .C1(n3145), .C2(n4711), .A(n3144), .B(n3143), .ZN(U3523)
         );
  INV_X1 U3976 ( .A(n3806), .ZN(n3146) );
  NAND2_X1 U3977 ( .A1(n3146), .A2(n3809), .ZN(n3895) );
  XOR2_X1 U3978 ( .A(n3895), .B(n3147), .Z(n3250) );
  XNOR2_X1 U3979 ( .A(n3148), .B(n3895), .ZN(n3249) );
  NAND2_X1 U3980 ( .A1(n3249), .A2(n4329), .ZN(n3150) );
  AOI22_X1 U3981 ( .A1(n3274), .A2(n4489), .B1(n3251), .B2(n4488), .ZN(n3149)
         );
  OAI211_X1 U3982 ( .C1(n3256), .C2(n4492), .A(n3150), .B(n3149), .ZN(n3151)
         );
  AOI21_X1 U3983 ( .B1(n3250), .B2(n4700), .A(n3151), .ZN(n3157) );
  INV_X1 U3984 ( .A(n3152), .ZN(n3153) );
  AOI21_X1 U3985 ( .B1(n3251), .B2(n3153), .A(n3233), .ZN(n3258) );
  NOR2_X1 U3986 ( .A1(n4706), .A2(n2351), .ZN(n3154) );
  AOI21_X1 U3987 ( .B1(n3258), .B2(n4505), .A(n3154), .ZN(n3155) );
  OAI21_X1 U3988 ( .B1(n3157), .B2(n2136), .A(n3155), .ZN(U3479) );
  AOI22_X1 U3989 ( .A1(n3258), .A2(n4401), .B1(n4711), .B2(REG1_REG_6__SCAN_IN), .ZN(n3156) );
  OAI21_X1 U3990 ( .B1(n3157), .B2(n4711), .A(n3156), .ZN(U3524) );
  NAND2_X1 U3991 ( .A1(n3131), .A2(n3871), .ZN(n3158) );
  NAND2_X1 U3992 ( .A1(n3159), .A2(n3158), .ZN(n4694) );
  NAND2_X1 U3993 ( .A1(n3160), .A2(D_REG_1__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U3994 ( .A1(n4674), .A2(n3161), .ZN(n3162) );
  NAND4_X1 U3995 ( .A1(n3165), .A2(n3164), .A3(n3163), .A4(n3162), .ZN(n3166)
         );
  OR2_X1 U3996 ( .A1(n3167), .A2(n4196), .ZN(n3243) );
  NOR2_X1 U3997 ( .A1(n4664), .A2(n3243), .ZN(n4661) );
  INV_X1 U3998 ( .A(n4661), .ZN(n3435) );
  XNOR2_X1 U3999 ( .A(n3169), .B(n3168), .ZN(n3174) );
  NAND2_X1 U4000 ( .A1(n4104), .A2(n4440), .ZN(n3170) );
  OAI21_X1 U4001 ( .B1(n4409), .B2(n3176), .A(n3170), .ZN(n3172) );
  NOR2_X1 U4002 ( .A1(n4694), .A2(n4363), .ZN(n3171) );
  AOI211_X1 U4003 ( .C1(n4489), .C2(n4102), .A(n3172), .B(n3171), .ZN(n3173)
         );
  OAI21_X1 U4004 ( .B1(n4384), .B2(n3174), .A(n3173), .ZN(n4696) );
  OAI211_X1 U4005 ( .C1(n2066), .C2(n3176), .A(n4693), .B(n3175), .ZN(n4695)
         );
  OAI22_X1 U4006 ( .A1(n4695), .A2(n4190), .B1(n4634), .B2(n3728), .ZN(n3177)
         );
  OAI21_X1 U4007 ( .B1(n4696), .B2(n3177), .A(n4566), .ZN(n3179) );
  NAND2_X1 U4008 ( .A1(n4664), .A2(REG2_REG_4__SCAN_IN), .ZN(n3178) );
  OAI211_X1 U4009 ( .C1(n4694), .C2(n3435), .A(n3179), .B(n3178), .ZN(U3286)
         );
  OAI21_X1 U4010 ( .B1(n3868), .B2(n3181), .A(n3180), .ZN(n4689) );
  NAND2_X1 U4011 ( .A1(n2691), .A2(n4440), .ZN(n3184) );
  NAND2_X1 U4012 ( .A1(n3182), .A2(n4489), .ZN(n3183) );
  OAI211_X1 U4013 ( .C1(n4409), .C2(n3185), .A(n3184), .B(n3183), .ZN(n3186)
         );
  INV_X1 U4014 ( .A(n3186), .ZN(n3189) );
  XNOR2_X1 U4015 ( .A(n3868), .B(n3790), .ZN(n3187) );
  NAND2_X1 U4016 ( .A1(n3187), .A2(n4329), .ZN(n3188) );
  OAI211_X1 U4017 ( .C1(n4689), .C2(n4363), .A(n3189), .B(n3188), .ZN(n4690)
         );
  INV_X1 U4018 ( .A(n4690), .ZN(n3191) );
  MUX2_X1 U4019 ( .A(n3191), .B(n3190), .S(n4664), .Z(n3199) );
  INV_X1 U4020 ( .A(n3192), .ZN(n3193) );
  INV_X1 U4021 ( .A(n3194), .ZN(n3195) );
  AOI21_X1 U4022 ( .B1(n3197), .B2(n3196), .A(n3195), .ZN(n4692) );
  INV_X1 U4023 ( .A(n4634), .ZN(n4659) );
  AOI22_X1 U4024 ( .A1(n4651), .A2(n4692), .B1(REG3_REG_1__SCAN_IN), .B2(n4659), .ZN(n3198) );
  OAI211_X1 U4025 ( .C1(n4689), .C2(n3435), .A(n3199), .B(n3198), .ZN(U3289)
         );
  XNOR2_X1 U4026 ( .A(n3202), .B(n3201), .ZN(n3203) );
  XNOR2_X1 U4027 ( .A(n3200), .B(n3203), .ZN(n3208) );
  AOI21_X1 U4028 ( .B1(n3779), .B2(n3274), .A(n3204), .ZN(n3206) );
  AOI22_X1 U4029 ( .A1(n3778), .A2(n4102), .B1(n3780), .B2(n3251), .ZN(n3205)
         );
  OAI211_X1 U4030 ( .C1(n3785), .C2(n3252), .A(n3206), .B(n3205), .ZN(n3207)
         );
  AOI21_X1 U4031 ( .B1(n3208), .B2(n3787), .A(n3207), .ZN(n3209) );
  INV_X1 U4032 ( .A(n3209), .ZN(U3236) );
  INV_X1 U4033 ( .A(n3210), .ZN(n3819) );
  NAND2_X1 U4034 ( .A1(n3819), .A2(n3816), .ZN(n3893) );
  XOR2_X1 U4035 ( .A(n3893), .B(n3211), .Z(n3308) );
  INV_X1 U4036 ( .A(n3342), .ZN(n3215) );
  XNOR2_X1 U4037 ( .A(n3212), .B(n3893), .ZN(n3213) );
  NAND2_X1 U4038 ( .A1(n3213), .A2(n4329), .ZN(n3305) );
  AOI22_X1 U4039 ( .A1(n3961), .A2(n4489), .B1(n4488), .B2(n3343), .ZN(n3214)
         );
  OAI211_X1 U4040 ( .C1(n3215), .C2(n4492), .A(n3305), .B(n3214), .ZN(n3216)
         );
  AOI21_X1 U4041 ( .B1(n3308), .B2(n4700), .A(n3216), .ZN(n3223) );
  AND2_X1 U4042 ( .A1(n3282), .A2(n3343), .ZN(n3217) );
  NOR2_X1 U40430 ( .A1(n3354), .A2(n3217), .ZN(n3299) );
  NOR2_X1 U4044 ( .A1(n4706), .A2(n3218), .ZN(n3219) );
  AOI21_X1 U4045 ( .B1(n3299), .B2(n4505), .A(n3219), .ZN(n3220) );
  OAI21_X1 U4046 ( .B1(n3223), .B2(n2136), .A(n3220), .ZN(U3485) );
  NAND2_X1 U4047 ( .A1(n4711), .A2(REG1_REG_9__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4048 ( .A1(n3299), .A2(n4401), .ZN(n3221) );
  OAI211_X1 U4049 ( .C1(n3223), .C2(n4711), .A(n3222), .B(n3221), .ZN(U3527)
         );
  XOR2_X1 U4050 ( .A(n3225), .B(n3224), .Z(n3231) );
  AOI21_X1 U4051 ( .B1(n3778), .B2(n3693), .A(n3226), .ZN(n3229) );
  AOI22_X1 U4052 ( .A1(n3227), .A2(n3682), .B1(n3779), .B2(n3342), .ZN(n3228)
         );
  OAI211_X1 U4053 ( .C1(n3785), .C2(n3240), .A(n3229), .B(n3228), .ZN(n3230)
         );
  AOI21_X1 U4054 ( .B1(n3231), .B2(n3787), .A(n3230), .ZN(n3232) );
  INV_X1 U4055 ( .A(n3232), .ZN(U3210) );
  OAI211_X1 U4056 ( .C1(n3233), .C2(n3237), .A(n4693), .B(n3280), .ZN(n4704)
         );
  XNOR2_X1 U4057 ( .A(n3234), .B(n2243), .ZN(n3239) );
  NAND2_X1 U4058 ( .A1(n3693), .A2(n4440), .ZN(n3236) );
  NAND2_X1 U4059 ( .A1(n3342), .A2(n4489), .ZN(n3235) );
  OAI211_X1 U4060 ( .C1(n4409), .C2(n3237), .A(n3236), .B(n3235), .ZN(n3238)
         );
  AOI21_X1 U4061 ( .B1(n3239), .B2(n4329), .A(n3238), .ZN(n4705) );
  OAI21_X1 U4062 ( .B1(n4190), .B2(n4704), .A(n4705), .ZN(n3247) );
  OAI22_X1 U4063 ( .A1(n4566), .A2(n3241), .B1(n3240), .B2(n4634), .ZN(n3246)
         );
  NAND2_X1 U4064 ( .A1(n3242), .A2(n2243), .ZN(n4701) );
  NAND2_X1 U4065 ( .A1(n4363), .A2(n3243), .ZN(n3244) );
  AND3_X1 U4066 ( .A1(n4702), .A2(n4701), .A3(n4333), .ZN(n3245) );
  AOI211_X1 U4067 ( .C1(n3247), .C2(n4566), .A(n3246), .B(n3245), .ZN(n3248)
         );
  INV_X1 U4068 ( .A(n3248), .ZN(U3283) );
  INV_X1 U4069 ( .A(n3249), .ZN(n3261) );
  NAND2_X1 U4070 ( .A1(n4566), .A2(n4329), .ZN(n3449) );
  NAND2_X1 U4071 ( .A1(n3250), .A2(n4333), .ZN(n3260) );
  NAND2_X1 U4072 ( .A1(n4566), .A2(n4488), .ZN(n4251) );
  AOI22_X1 U4073 ( .A1(n4338), .A2(n3251), .B1(n4337), .B2(n3274), .ZN(n3255)
         );
  INV_X1 U4074 ( .A(n3252), .ZN(n3253) );
  AOI22_X1 U4075 ( .A1(n4664), .A2(REG2_REG_6__SCAN_IN), .B1(n3253), .B2(n4659), .ZN(n3254) );
  OAI211_X1 U4076 ( .C1(n3256), .C2(n4342), .A(n3255), .B(n3254), .ZN(n3257)
         );
  AOI21_X1 U4077 ( .B1(n3258), .B2(n4651), .A(n3257), .ZN(n3259) );
  OAI211_X1 U4078 ( .C1(n3261), .C2(n3449), .A(n3260), .B(n3259), .ZN(U3284)
         );
  NOR2_X1 U4079 ( .A1(n2064), .A2(n3262), .ZN(n3263) );
  XNOR2_X1 U4080 ( .A(n3264), .B(n3263), .ZN(n3270) );
  INV_X1 U4081 ( .A(n3265), .ZN(n3266) );
  AOI21_X1 U4082 ( .B1(n3778), .B2(n3274), .A(n3266), .ZN(n3268) );
  AOI22_X1 U4083 ( .A1(n3279), .A2(n3780), .B1(n3779), .B2(n3962), .ZN(n3267)
         );
  OAI211_X1 U4084 ( .C1(n3785), .C2(n4635), .A(n3268), .B(n3267), .ZN(n3269)
         );
  AOI21_X1 U4085 ( .B1(n3270), .B2(n3787), .A(n3269), .ZN(n3271) );
  INV_X1 U4086 ( .A(n3271), .ZN(U3218) );
  NAND2_X1 U4087 ( .A1(n3815), .A2(n3811), .ZN(n3892) );
  XNOR2_X1 U4088 ( .A(n3272), .B(n3892), .ZN(n4637) );
  XNOR2_X1 U4089 ( .A(n3273), .B(n3892), .ZN(n3278) );
  INV_X1 U4090 ( .A(n3962), .ZN(n3358) );
  AOI22_X1 U4091 ( .A1(n3274), .A2(n4440), .B1(n3279), .B2(n4488), .ZN(n3275)
         );
  OAI21_X1 U4092 ( .B1(n3358), .B2(n4444), .A(n3275), .ZN(n3277) );
  NOR2_X1 U4093 ( .A1(n4637), .A2(n4363), .ZN(n3276) );
  AOI211_X1 U4094 ( .C1(n4329), .C2(n3278), .A(n3277), .B(n3276), .ZN(n4643)
         );
  OAI21_X1 U4095 ( .B1(n4688), .B2(n4637), .A(n4643), .ZN(n3287) );
  NAND2_X1 U4096 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  NAND2_X1 U4097 ( .A1(n3282), .A2(n3281), .ZN(n4638) );
  INV_X1 U4098 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3283) );
  OAI22_X1 U4099 ( .A1(n4638), .A2(n4486), .B1(n4713), .B2(n3283), .ZN(n3284)
         );
  AOI21_X1 U4100 ( .B1(n3287), .B2(n4713), .A(n3284), .ZN(n3285) );
  INV_X1 U4101 ( .A(n3285), .ZN(U3526) );
  OAI22_X1 U4102 ( .A1(n4638), .A2(n4552), .B1(n4706), .B2(n2371), .ZN(n3286)
         );
  AOI21_X1 U4103 ( .B1(n3287), .B2(n4706), .A(n3286), .ZN(n3288) );
  INV_X1 U4104 ( .A(n3288), .ZN(U3483) );
  NAND2_X1 U4105 ( .A1(n3289), .A2(n4651), .ZN(n3293) );
  OAI22_X1 U4106 ( .A1(n4566), .A2(n4019), .B1(n3695), .B2(n4634), .ZN(n3290)
         );
  AOI21_X1 U4107 ( .B1(n4247), .B2(n4103), .A(n3290), .ZN(n3292) );
  AOI22_X1 U4108 ( .A1(n4338), .A2(n3694), .B1(n4337), .B2(n3693), .ZN(n3291)
         );
  NAND3_X1 U4109 ( .A1(n3293), .A2(n3292), .A3(n3291), .ZN(n3296) );
  NOR2_X1 U4110 ( .A1(n3294), .A2(n4664), .ZN(n3295) );
  AOI211_X1 U4111 ( .C1(n3297), .C2(n4333), .A(n3296), .B(n3295), .ZN(n3298)
         );
  INV_X1 U4112 ( .A(n3298), .ZN(U3285) );
  NAND2_X1 U4113 ( .A1(n3299), .A2(n4651), .ZN(n3304) );
  OAI22_X1 U4114 ( .A1(n3346), .A2(n4634), .B1(n3300), .B2(n4566), .ZN(n3301)
         );
  AOI21_X1 U4115 ( .B1(n4247), .B2(n3342), .A(n3301), .ZN(n3303) );
  AOI22_X1 U4116 ( .A1(n4338), .A2(n3343), .B1(n4337), .B2(n3961), .ZN(n3302)
         );
  NAND3_X1 U4117 ( .A1(n3304), .A2(n3303), .A3(n3302), .ZN(n3307) );
  NOR2_X1 U4118 ( .A1(n3305), .A2(n4664), .ZN(n3306) );
  AOI211_X1 U4119 ( .C1(n3308), .C2(n4333), .A(n3307), .B(n3306), .ZN(n3309)
         );
  INV_X1 U4120 ( .A(n3309), .ZN(U3281) );
  NAND2_X1 U4121 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3327), .ZN(n3315) );
  INV_X1 U4122 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4123 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3327), .B1(n4683), .B2(
        n3310), .ZN(n4582) );
  OAI21_X1 U4124 ( .B1(n3061), .B2(n3329), .A(n3312), .ZN(n3313) );
  NAND2_X1 U4125 ( .A1(n4570), .A2(n3313), .ZN(n3314) );
  XOR2_X1 U4126 ( .A(n3313), .B(n4570), .Z(n4577) );
  NAND2_X1 U4127 ( .A1(n4591), .A2(n3316), .ZN(n3317) );
  INV_X1 U4128 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3318) );
  NOR2_X1 U4129 ( .A1(n3324), .A2(n3318), .ZN(n3518) );
  AOI21_X1 U4130 ( .B1(n3318), .B2(n3324), .A(n3518), .ZN(n3319) );
  OAI211_X1 U4131 ( .C1(n3320), .C2(n3319), .A(n4627), .B(n3519), .ZN(n3323)
         );
  NOR2_X1 U4132 ( .A1(STATE_REG_SCAN_IN), .A2(n3321), .ZN(n3573) );
  AOI21_X1 U4133 ( .B1(n4626), .B2(ADDR_REG_13__SCAN_IN), .A(n3573), .ZN(n3322) );
  OAI211_X1 U4134 ( .C1(n4633), .C2(n3324), .A(n3323), .B(n3322), .ZN(n3338)
         );
  INV_X1 U4135 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3325) );
  NOR2_X1 U4136 ( .A1(n3324), .A2(n3325), .ZN(n3530) );
  AOI21_X1 U4137 ( .B1(n3325), .B2(n3324), .A(n3530), .ZN(n3336) );
  NAND2_X1 U4138 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3327), .ZN(n3332) );
  INV_X1 U4139 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4140 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3327), .B1(n4683), .B2(
        n3326), .ZN(n4585) );
  NAND2_X1 U4141 ( .A1(n4570), .A2(n3330), .ZN(n3331) );
  NAND2_X1 U4142 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4572), .ZN(n4571) );
  NAND2_X1 U4143 ( .A1(n3331), .A2(n4571), .ZN(n4584) );
  NAND2_X1 U4144 ( .A1(n4591), .A2(n3333), .ZN(n3334) );
  OAI21_X1 U4145 ( .B1(n3336), .B2(n3531), .A(n4593), .ZN(n3335) );
  AOI21_X1 U4146 ( .B1(n3336), .B2(n3531), .A(n3335), .ZN(n3337) );
  OR2_X1 U4147 ( .A1(n3338), .A2(n3337), .ZN(U3253) );
  XNOR2_X1 U4148 ( .A(n3340), .B(n3339), .ZN(n3348) );
  AOI21_X1 U4149 ( .B1(n3778), .B2(n3342), .A(n3341), .ZN(n3345) );
  AOI22_X1 U4150 ( .A1(n3343), .A2(n3682), .B1(n3779), .B2(n3961), .ZN(n3344)
         );
  OAI211_X1 U4151 ( .C1(n3785), .C2(n3346), .A(n3345), .B(n3344), .ZN(n3347)
         );
  AOI21_X1 U4152 ( .B1(n3348), .B2(n3787), .A(n3347), .ZN(n3349) );
  INV_X1 U4153 ( .A(n3349), .ZN(U3228) );
  NAND2_X1 U4154 ( .A1(n3818), .A2(n3821), .ZN(n3898) );
  XNOR2_X1 U4155 ( .A(n3350), .B(n3898), .ZN(n3364) );
  INV_X1 U4156 ( .A(n3364), .ZN(n3363) );
  INV_X1 U4157 ( .A(n3898), .ZN(n3351) );
  XNOR2_X1 U4158 ( .A(n3352), .B(n3351), .ZN(n3369) );
  INV_X1 U4159 ( .A(n3449), .ZN(n3361) );
  INV_X1 U4160 ( .A(n3430), .ZN(n3353) );
  OAI21_X1 U4161 ( .B1(n3354), .B2(n3367), .A(n3353), .ZN(n3376) );
  NOR2_X1 U4162 ( .A1(n3376), .A2(n4389), .ZN(n3360) );
  AOI22_X1 U4163 ( .A1(n4338), .A2(n3455), .B1(n4337), .B2(n3959), .ZN(n3357)
         );
  INV_X1 U4164 ( .A(n3458), .ZN(n3355) );
  AOI22_X1 U4165 ( .A1(n4664), .A2(REG2_REG_10__SCAN_IN), .B1(n3355), .B2(
        n4659), .ZN(n3356) );
  OAI211_X1 U4166 ( .C1(n3358), .C2(n4342), .A(n3357), .B(n3356), .ZN(n3359)
         );
  AOI211_X1 U4167 ( .C1(n3369), .C2(n3361), .A(n3360), .B(n3359), .ZN(n3362)
         );
  OAI21_X1 U4168 ( .B1(n3363), .B2(n4394), .A(n3362), .ZN(U3280) );
  NAND2_X1 U4169 ( .A1(n3364), .A2(n4700), .ZN(n3371) );
  NAND2_X1 U4170 ( .A1(n3962), .A2(n4440), .ZN(n3366) );
  NAND2_X1 U4171 ( .A1(n3959), .A2(n4489), .ZN(n3365) );
  OAI211_X1 U4172 ( .C1(n4409), .C2(n3367), .A(n3366), .B(n3365), .ZN(n3368)
         );
  AOI21_X1 U4173 ( .B1(n3369), .B2(n4329), .A(n3368), .ZN(n3370) );
  AND2_X1 U4174 ( .A1(n3371), .A2(n3370), .ZN(n3373) );
  MUX2_X1 U4175 ( .A(n2398), .B(n3373), .S(n4706), .Z(n3372) );
  OAI21_X1 U4176 ( .B1(n3376), .B2(n4552), .A(n3372), .ZN(U3487) );
  INV_X1 U4177 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3374) );
  MUX2_X1 U4178 ( .A(n3374), .B(n3373), .S(n4713), .Z(n3375) );
  OAI21_X1 U4179 ( .B1(n3376), .B2(n4486), .A(n3375), .ZN(U3528) );
  INV_X1 U4180 ( .A(n3377), .ZN(n3379) );
  OR2_X1 U4181 ( .A1(n3379), .A2(n3378), .ZN(n3897) );
  XNOR2_X1 U4182 ( .A(n3380), .B(n3897), .ZN(n3462) );
  INV_X1 U4183 ( .A(n3462), .ZN(n3393) );
  INV_X1 U4184 ( .A(n3381), .ZN(n3382) );
  AOI21_X1 U4185 ( .B1(n3421), .B2(n3822), .A(n3382), .ZN(n3403) );
  INV_X1 U4186 ( .A(n3395), .ZN(n3383) );
  AOI21_X1 U4187 ( .B1(n3403), .B2(n3396), .A(n3383), .ZN(n3384) );
  XNOR2_X1 U4188 ( .A(n3384), .B(n3897), .ZN(n3388) );
  OAI22_X1 U4189 ( .A1(n3562), .A2(n4444), .B1(n4409), .B2(n3385), .ZN(n3386)
         );
  AOI21_X1 U4190 ( .B1(n4440), .B2(n3574), .A(n3386), .ZN(n3387) );
  OAI21_X1 U4191 ( .B1(n3388), .B2(n4384), .A(n3387), .ZN(n3461) );
  NAND2_X1 U4192 ( .A1(n2042), .A2(n3575), .ZN(n3389) );
  NAND2_X1 U4193 ( .A1(n3438), .A2(n3389), .ZN(n3467) );
  NOR2_X1 U4194 ( .A1(n3467), .A2(n4389), .ZN(n3391) );
  OAI22_X1 U4195 ( .A1(n4566), .A2(n3325), .B1(n3578), .B2(n4634), .ZN(n3390)
         );
  AOI211_X1 U4196 ( .C1(n3461), .C2(n4566), .A(n3391), .B(n3390), .ZN(n3392)
         );
  OAI21_X1 U4197 ( .B1(n3393), .B2(n4394), .A(n3392), .ZN(U3277) );
  NAND2_X1 U4198 ( .A1(n3417), .A2(n3394), .ZN(n3397) );
  NAND2_X1 U4199 ( .A1(n3396), .A2(n3395), .ZN(n3899) );
  XNOR2_X1 U4200 ( .A(n3397), .B(n3899), .ZN(n3472) );
  NAND2_X1 U4201 ( .A1(n2065), .A2(n3487), .ZN(n3398) );
  NAND2_X1 U4202 ( .A1(n2042), .A2(n3398), .ZN(n3480) );
  INV_X1 U4203 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3399) );
  OAI22_X1 U4204 ( .A1(n4566), .A2(n3399), .B1(n3490), .B2(n4634), .ZN(n3400)
         );
  AOI21_X1 U4205 ( .B1(n4247), .B2(n3959), .A(n3400), .ZN(n3402) );
  AOI22_X1 U4206 ( .A1(n4338), .A2(n3487), .B1(n4337), .B2(n3958), .ZN(n3401)
         );
  OAI211_X1 U4207 ( .C1(n3480), .C2(n4389), .A(n3402), .B(n3401), .ZN(n3406)
         );
  XNOR2_X1 U4208 ( .A(n3403), .B(n3899), .ZN(n3404) );
  NAND2_X1 U4209 ( .A1(n3404), .A2(n4329), .ZN(n3469) );
  NOR2_X1 U4210 ( .A1(n3469), .A2(n4664), .ZN(n3405) );
  AOI211_X1 U4211 ( .C1(n4333), .C2(n3472), .A(n3406), .B(n3405), .ZN(n3407)
         );
  INV_X1 U4212 ( .A(n3407), .ZN(U3278) );
  XNOR2_X1 U4213 ( .A(n3410), .B(n3409), .ZN(n3411) );
  XNOR2_X1 U4214 ( .A(n3408), .B(n3411), .ZN(n3415) );
  AND2_X1 U4215 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4589) );
  AOI21_X1 U4216 ( .B1(n3779), .B2(n3574), .A(n4589), .ZN(n3413) );
  AOI22_X1 U4217 ( .A1(n3778), .A2(n3961), .B1(n3780), .B2(n2145), .ZN(n3412)
         );
  OAI211_X1 U4218 ( .C1(n3785), .C2(n3428), .A(n3413), .B(n3412), .ZN(n3414)
         );
  AOI21_X1 U4219 ( .B1(n3415), .B2(n3787), .A(n3414), .ZN(n3416) );
  INV_X1 U4220 ( .A(n3416), .ZN(U3233) );
  INV_X1 U4221 ( .A(n3417), .ZN(n3418) );
  AOI21_X1 U4222 ( .B1(n3420), .B2(n3419), .A(n3418), .ZN(n3552) );
  XNOR2_X1 U4223 ( .A(n3421), .B(n3879), .ZN(n3427) );
  INV_X1 U4224 ( .A(n3552), .ZN(n3425) );
  OAI22_X1 U4225 ( .A1(n3422), .A2(n4444), .B1(n4409), .B2(n3429), .ZN(n3423)
         );
  AOI21_X1 U4226 ( .B1(n3425), .B2(n3424), .A(n3423), .ZN(n3426) );
  OAI21_X1 U4227 ( .B1(n4384), .B2(n3427), .A(n3426), .ZN(n3554) );
  NAND2_X1 U4228 ( .A1(n3554), .A2(n4566), .ZN(n3434) );
  OAI22_X1 U4229 ( .A1(n4566), .A2(n3326), .B1(n3428), .B2(n4634), .ZN(n3432)
         );
  OAI21_X1 U4230 ( .B1(n3430), .B2(n3429), .A(n2065), .ZN(n3559) );
  NOR2_X1 U4231 ( .A1(n3559), .A2(n4389), .ZN(n3431) );
  AOI211_X1 U4232 ( .C1(n4247), .C2(n3961), .A(n3432), .B(n3431), .ZN(n3433)
         );
  OAI211_X1 U4233 ( .C1(n3552), .C2(n3435), .A(n3434), .B(n3433), .ZN(U3279)
         );
  XNOR2_X1 U4234 ( .A(n3913), .B(n3437), .ZN(n3510) );
  OAI21_X1 U4235 ( .B1(n2057), .B2(n3437), .A(n3436), .ZN(n3512) );
  NAND2_X1 U4236 ( .A1(n3512), .A2(n4333), .ZN(n3448) );
  INV_X1 U4237 ( .A(n3438), .ZN(n3440) );
  INV_X1 U4238 ( .A(n3499), .ZN(n3439) );
  OAI21_X1 U4239 ( .B1(n3440), .B2(n3507), .A(n3439), .ZN(n3517) );
  INV_X1 U4240 ( .A(n3517), .ZN(n3446) );
  AOI22_X1 U4241 ( .A1(n4338), .A2(n3599), .B1(n4337), .B2(n3681), .ZN(n3443)
         );
  INV_X1 U4242 ( .A(n3602), .ZN(n3441) );
  AOI22_X1 U4243 ( .A1(n4664), .A2(REG2_REG_14__SCAN_IN), .B1(n3441), .B2(
        n4659), .ZN(n3442) );
  OAI211_X1 U4244 ( .C1(n3444), .C2(n4342), .A(n3443), .B(n3442), .ZN(n3445)
         );
  AOI21_X1 U4245 ( .B1(n3446), .B2(n4651), .A(n3445), .ZN(n3447) );
  OAI211_X1 U4246 ( .C1(n3510), .C2(n3449), .A(n3448), .B(n3447), .ZN(U3276)
         );
  INV_X1 U4247 ( .A(n3451), .ZN(n3452) );
  AOI211_X1 U4248 ( .C1(n3453), .C2(n3450), .A(n3771), .B(n3452), .ZN(n3460)
         );
  NAND2_X1 U4249 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4573) );
  INV_X1 U4250 ( .A(n4573), .ZN(n3454) );
  AOI21_X1 U4251 ( .B1(n3778), .B2(n3962), .A(n3454), .ZN(n3457) );
  AOI22_X1 U4252 ( .A1(n3455), .A2(n3780), .B1(n3779), .B2(n3959), .ZN(n3456)
         );
  OAI211_X1 U4253 ( .C1(n3785), .C2(n3458), .A(n3457), .B(n3456), .ZN(n3459)
         );
  OR2_X1 U4254 ( .A1(n3460), .A2(n3459), .ZN(U3214) );
  AOI21_X1 U4255 ( .B1(n4700), .B2(n3462), .A(n3461), .ZN(n3464) );
  MUX2_X1 U4256 ( .A(n3318), .B(n3464), .S(n4713), .Z(n3463) );
  OAI21_X1 U4257 ( .B1(n4486), .B2(n3467), .A(n3463), .ZN(U3531) );
  MUX2_X1 U4258 ( .A(n3465), .B(n3464), .S(n4706), .Z(n3466) );
  OAI21_X1 U4259 ( .B1(n3467), .B2(n4552), .A(n3466), .ZN(U3493) );
  AOI22_X1 U4260 ( .A1(n3958), .A2(n4489), .B1(n4488), .B2(n3487), .ZN(n3468)
         );
  OAI211_X1 U4261 ( .C1(n3470), .C2(n4492), .A(n3469), .B(n3468), .ZN(n3471)
         );
  INV_X1 U4262 ( .A(n3471), .ZN(n3474) );
  NAND2_X1 U4263 ( .A1(n3472), .A2(n4700), .ZN(n3473) );
  AND2_X1 U4264 ( .A1(n3474), .A2(n3473), .ZN(n3477) );
  INV_X1 U4265 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3475) );
  MUX2_X1 U4266 ( .A(n3477), .B(n3475), .S(n4711), .Z(n3476) );
  OAI21_X1 U4267 ( .B1(n4486), .B2(n3480), .A(n3476), .ZN(U3530) );
  MUX2_X1 U4268 ( .A(n3478), .B(n3477), .S(n4706), .Z(n3479) );
  OAI21_X1 U4269 ( .B1(n3480), .B2(n4552), .A(n3479), .ZN(U3491) );
  INV_X1 U4270 ( .A(n3481), .ZN(n3483) );
  NAND2_X1 U4271 ( .A1(n3483), .A2(n3482), .ZN(n3484) );
  XNOR2_X1 U4272 ( .A(n3485), .B(n3484), .ZN(n3492) );
  NAND2_X1 U4273 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4595) );
  INV_X1 U4274 ( .A(n4595), .ZN(n3486) );
  AOI21_X1 U4275 ( .B1(n3778), .B2(n3959), .A(n3486), .ZN(n3489) );
  AOI22_X1 U4276 ( .A1(n3487), .A2(n3780), .B1(n3779), .B2(n3958), .ZN(n3488)
         );
  OAI211_X1 U4277 ( .C1(n3785), .C2(n3490), .A(n3489), .B(n3488), .ZN(n3491)
         );
  AOI21_X1 U4278 ( .B1(n3492), .B2(n3787), .A(n3491), .ZN(n3493) );
  INV_X1 U4279 ( .A(n3493), .ZN(U3221) );
  AOI21_X1 U4280 ( .B1(n3494), .B2(n3875), .A(n4384), .ZN(n3496) );
  NAND2_X1 U4281 ( .A1(n3496), .A2(n3495), .ZN(n3561) );
  XNOR2_X1 U4282 ( .A(n3497), .B(n3875), .ZN(n3564) );
  NAND2_X1 U4283 ( .A1(n3564), .A2(n4333), .ZN(n3506) );
  OAI21_X1 U4284 ( .B1(n3499), .B2(n3498), .A(n3544), .ZN(n3569) );
  INV_X1 U4285 ( .A(n3569), .ZN(n3504) );
  AOI22_X1 U4286 ( .A1(n4338), .A2(n3781), .B1(n4337), .B2(n3957), .ZN(n3502)
         );
  INV_X1 U4287 ( .A(n3784), .ZN(n3500) );
  AOI22_X1 U4288 ( .A1(n4664), .A2(REG2_REG_15__SCAN_IN), .B1(n3500), .B2(
        n4659), .ZN(n3501) );
  OAI211_X1 U4289 ( .C1(n3562), .C2(n4342), .A(n3502), .B(n3501), .ZN(n3503)
         );
  AOI21_X1 U4290 ( .B1(n3504), .B2(n4651), .A(n3503), .ZN(n3505) );
  OAI211_X1 U4291 ( .C1(n4664), .C2(n3561), .A(n3506), .B(n3505), .ZN(U3275)
         );
  INV_X1 U4292 ( .A(n3681), .ZN(n4493) );
  OAI22_X1 U4293 ( .A1(n4493), .A2(n4444), .B1(n4409), .B2(n3507), .ZN(n3508)
         );
  AOI21_X1 U4294 ( .B1(n4440), .B2(n3958), .A(n3508), .ZN(n3509) );
  OAI21_X1 U4295 ( .B1(n3510), .B2(n4384), .A(n3509), .ZN(n3511) );
  AOI21_X1 U4296 ( .B1(n3512), .B2(n4700), .A(n3511), .ZN(n3515) );
  INV_X1 U4297 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3988) );
  MUX2_X1 U4298 ( .A(n3515), .B(n3988), .S(n4711), .Z(n3513) );
  OAI21_X1 U4299 ( .B1(n4486), .B2(n3517), .A(n3513), .ZN(U3532) );
  MUX2_X1 U4300 ( .A(n3515), .B(n3514), .S(n2136), .Z(n3516) );
  OAI21_X1 U4301 ( .B1(n3517), .B2(n4552), .A(n3516), .ZN(U3495) );
  INV_X1 U4302 ( .A(n3534), .ZN(n3529) );
  INV_X1 U4303 ( .A(n4681), .ZN(n3521) );
  INV_X1 U4304 ( .A(n3518), .ZN(n3520) );
  NAND2_X1 U4305 ( .A1(n3521), .A2(n3522), .ZN(n3523) );
  NAND2_X1 U4306 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U4307 ( .A1(n3523), .A2(n4607), .ZN(n3526) );
  INV_X1 U4308 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U4309 ( .A1(n3534), .A2(REG1_REG_15__SCAN_IN), .ZN(n4158) );
  INV_X1 U4310 ( .A(n4158), .ZN(n3524) );
  AOI21_X1 U4311 ( .B1(n4016), .B2(n3529), .A(n3524), .ZN(n3525) );
  OAI211_X1 U4312 ( .C1(n3526), .C2(n3525), .A(n4627), .B(n4157), .ZN(n3528)
         );
  AND2_X1 U4313 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n3776) );
  AOI21_X1 U4314 ( .B1(n4626), .B2(ADDR_REG_15__SCAN_IN), .A(n3776), .ZN(n3527) );
  OAI211_X1 U4315 ( .C1(n4633), .C2(n3529), .A(n3528), .B(n3527), .ZN(n3539)
         );
  OAI22_X1 U4316 ( .A1(n3531), .A2(n3530), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4557), .ZN(n3532) );
  NOR2_X1 U4317 ( .A1(n4681), .A2(n3532), .ZN(n3533) );
  INV_X1 U4318 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U4319 ( .A1(n3534), .A2(REG2_REG_15__SCAN_IN), .ZN(n4171) );
  OR2_X1 U4320 ( .A1(n3534), .A2(REG2_REG_15__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4321 ( .A1(n4171), .A2(n3535), .ZN(n3537) );
  INV_X1 U4322 ( .A(n4172), .ZN(n3536) );
  AOI211_X1 U4323 ( .C1(n2061), .C2(n3537), .A(n3536), .B(n4620), .ZN(n3538)
         );
  OR2_X1 U4324 ( .A1(n3539), .A2(n3538), .ZN(U3255) );
  OAI21_X1 U4325 ( .B1(n3542), .B2(n3541), .A(n3540), .ZN(n4499) );
  INV_X1 U4326 ( .A(n3543), .ZN(n3588) );
  AOI21_X1 U4327 ( .B1(n4487), .B2(n3544), .A(n3588), .ZN(n4495) );
  AOI22_X1 U4328 ( .A1(n4338), .A2(n4487), .B1(n4337), .B2(n4490), .ZN(n3547)
         );
  INV_X1 U4329 ( .A(n3685), .ZN(n3545) );
  AOI22_X1 U4330 ( .A1(n4664), .A2(REG2_REG_16__SCAN_IN), .B1(n3545), .B2(
        n4659), .ZN(n3546) );
  OAI211_X1 U4331 ( .C1(n4493), .C2(n4342), .A(n3547), .B(n3546), .ZN(n3550)
         );
  OAI211_X1 U4332 ( .C1(n3548), .C2(n3878), .A(n3582), .B(n4329), .ZN(n4496)
         );
  NOR2_X1 U4333 ( .A1(n4496), .A2(n4664), .ZN(n3549) );
  AOI211_X1 U4334 ( .C1(n4495), .C2(n4651), .A(n3550), .B(n3549), .ZN(n3551)
         );
  OAI21_X1 U4335 ( .B1(n4499), .B2(n4394), .A(n3551), .ZN(U3274) );
  NOR2_X1 U4336 ( .A1(n3552), .A2(n4688), .ZN(n3553) );
  AOI211_X1 U4337 ( .C1(n4440), .C2(n3961), .A(n3554), .B(n3553), .ZN(n3556)
         );
  MUX2_X1 U4338 ( .A(n3310), .B(n3556), .S(n4713), .Z(n3555) );
  OAI21_X1 U4339 ( .B1(n4486), .B2(n3559), .A(n3555), .ZN(U3529) );
  MUX2_X1 U4340 ( .A(n3557), .B(n3556), .S(n4706), .Z(n3558) );
  OAI21_X1 U4341 ( .B1(n3559), .B2(n4552), .A(n3558), .ZN(U3489) );
  AOI22_X1 U4342 ( .A1(n3957), .A2(n4489), .B1(n4488), .B2(n3781), .ZN(n3560)
         );
  OAI211_X1 U4343 ( .C1(n3562), .C2(n4492), .A(n3561), .B(n3560), .ZN(n3563)
         );
  AOI21_X1 U4344 ( .B1(n3564), .B2(n4700), .A(n3563), .ZN(n3567) );
  MUX2_X1 U4345 ( .A(n3567), .B(n3565), .S(n2136), .Z(n3566) );
  OAI21_X1 U4346 ( .B1(n3569), .B2(n4552), .A(n3566), .ZN(U3497) );
  MUX2_X1 U4347 ( .A(n3567), .B(n4016), .S(n4711), .Z(n3568) );
  OAI21_X1 U4348 ( .B1(n4486), .B2(n3569), .A(n3568), .ZN(U3533) );
  XNOR2_X1 U4349 ( .A(n3571), .B(n3570), .ZN(n3572) );
  XNOR2_X1 U4350 ( .A(n2056), .B(n3572), .ZN(n3580) );
  AOI21_X1 U4351 ( .B1(n3778), .B2(n3574), .A(n3573), .ZN(n3577) );
  AOI22_X1 U4352 ( .A1(n3575), .A2(n3780), .B1(n3779), .B2(n3777), .ZN(n3576)
         );
  OAI211_X1 U4353 ( .C1(n3785), .C2(n3578), .A(n3577), .B(n3576), .ZN(n3579)
         );
  AOI21_X1 U4354 ( .B1(n3580), .B2(n3787), .A(n3579), .ZN(n3581) );
  INV_X1 U4355 ( .A(n3581), .ZN(U3231) );
  NAND2_X1 U4356 ( .A1(n3582), .A2(n3833), .ZN(n3583) );
  NAND2_X1 U4357 ( .A1(n3611), .A2(n3835), .ZN(n3896) );
  XNOR2_X1 U4358 ( .A(n3583), .B(n3896), .ZN(n3584) );
  NAND2_X1 U4359 ( .A1(n3584), .A2(n4329), .ZN(n4481) );
  XOR2_X1 U4360 ( .A(n3896), .B(n3585), .Z(n4484) );
  NAND2_X1 U4361 ( .A1(n4484), .A2(n4333), .ZN(n3595) );
  INV_X1 U4362 ( .A(n3610), .ZN(n3586) );
  OAI21_X1 U4363 ( .B1(n3588), .B2(n3587), .A(n3586), .ZN(n4553) );
  INV_X1 U4364 ( .A(n4553), .ZN(n3593) );
  INV_X1 U4365 ( .A(n3957), .ZN(n4482) );
  AOI22_X1 U4366 ( .A1(n4338), .A2(n4478), .B1(n4337), .B2(n4479), .ZN(n3591)
         );
  INV_X1 U4367 ( .A(n3707), .ZN(n3589) );
  AOI22_X1 U4368 ( .A1(n4664), .A2(REG2_REG_17__SCAN_IN), .B1(n3589), .B2(
        n4659), .ZN(n3590) );
  OAI211_X1 U4369 ( .C1(n4482), .C2(n4342), .A(n3591), .B(n3590), .ZN(n3592)
         );
  AOI21_X1 U4370 ( .B1(n3593), .B2(n4651), .A(n3592), .ZN(n3594) );
  OAI211_X1 U4371 ( .C1(n4664), .C2(n4481), .A(n3595), .B(n3594), .ZN(U3273)
         );
  NAND2_X1 U4372 ( .A1(n2063), .A2(n3596), .ZN(n3597) );
  XNOR2_X1 U4373 ( .A(n3598), .B(n3597), .ZN(n3604) );
  AND2_X1 U4374 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4606) );
  AOI21_X1 U4375 ( .B1(n3778), .B2(n3958), .A(n4606), .ZN(n3601) );
  AOI22_X1 U4376 ( .A1(n3599), .A2(n3780), .B1(n3779), .B2(n3681), .ZN(n3600)
         );
  OAI211_X1 U4377 ( .C1(n3785), .C2(n3602), .A(n3601), .B(n3600), .ZN(n3603)
         );
  AOI21_X1 U4378 ( .B1(n3604), .B2(n3787), .A(n3603), .ZN(n3605) );
  INV_X1 U4379 ( .A(n3605), .ZN(U3212) );
  INV_X1 U4380 ( .A(n4374), .ZN(n3607) );
  AOI21_X1 U4381 ( .B1(n3873), .B2(n3606), .A(n3607), .ZN(n4477) );
  INV_X1 U4382 ( .A(n4388), .ZN(n3608) );
  OAI211_X1 U4383 ( .C1(n3610), .C2(n3609), .A(n3608), .B(n4693), .ZN(n4475)
         );
  NAND2_X1 U4384 ( .A1(n4355), .A2(n3611), .ZN(n4379) );
  XNOR2_X1 U4385 ( .A(n4379), .B(n3873), .ZN(n3615) );
  AOI22_X1 U4386 ( .A1(n3956), .A2(n4489), .B1(n4488), .B2(n3757), .ZN(n3612)
         );
  OAI21_X1 U4387 ( .B1(n3613), .B2(n4492), .A(n3612), .ZN(n3614) );
  AOI21_X1 U4388 ( .B1(n3615), .B2(n4329), .A(n3614), .ZN(n4476) );
  OAI21_X1 U4389 ( .B1(n4190), .B2(n4475), .A(n4476), .ZN(n3617) );
  INV_X1 U4390 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4168) );
  OAI22_X1 U4391 ( .A1(n4566), .A2(n4168), .B1(n3760), .B2(n4634), .ZN(n3616)
         );
  AOI21_X1 U4392 ( .B1(n3617), .B2(n4566), .A(n3616), .ZN(n3618) );
  OAI21_X1 U4393 ( .B1(n4477), .B2(n4394), .A(n3618), .ZN(U3272) );
  INV_X1 U4394 ( .A(IR_REG_30__SCAN_IN), .ZN(n4070) );
  NAND3_X1 U4395 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4070), 
        .ZN(n3619) );
  INV_X1 U4396 ( .A(DATAI_31_), .ZN(n4083) );
  OAI22_X1 U4397 ( .A1(n3620), .A2(n3619), .B1(STATE_REG_SCAN_IN), .B2(n4083), 
        .ZN(U3321) );
  OAI22_X1 U4398 ( .A1(n4251), .A2(n3859), .B1(n3621), .B2(n4566), .ZN(n3622)
         );
  AOI21_X1 U4399 ( .B1(n4233), .B2(n4247), .A(n3622), .ZN(n3629) );
  INV_X1 U4400 ( .A(n3623), .ZN(n3627) );
  OAI22_X1 U4401 ( .A1(n3625), .A2(n4389), .B1(n3624), .B2(n4634), .ZN(n3626)
         );
  OAI21_X1 U4402 ( .B1(n3627), .B2(n3626), .A(n4566), .ZN(n3628) );
  OAI211_X1 U4403 ( .C1(n3630), .C2(n4394), .A(n3629), .B(n3628), .ZN(U3354)
         );
  NOR2_X1 U4404 ( .A1(n4228), .A2(n3785), .ZN(n3635) );
  AOI22_X1 U4405 ( .A1(n3780), .A2(n4418), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3632) );
  OAI21_X1 U4406 ( .B1(n3633), .B2(n3715), .A(n3632), .ZN(n3634) );
  AOI211_X1 U4407 ( .C1(n3779), .C2(n4233), .A(n3635), .B(n3634), .ZN(n3636)
         );
  INV_X1 U4408 ( .A(n3637), .ZN(n3743) );
  OAI21_X1 U4409 ( .B1(n3743), .B2(n3639), .A(n3638), .ZN(n3641) );
  NAND3_X1 U4410 ( .A1(n3641), .A2(n3787), .A3(n3640), .ZN(n3646) );
  OAI22_X1 U4411 ( .A1(n4263), .A2(n3717), .B1(STATE_REG_SCAN_IN), .B2(n3642), 
        .ZN(n3644) );
  OAI22_X1 U4412 ( .A1(n3088), .A2(n4304), .B1(n4298), .B2(n3715), .ZN(n3643)
         );
  NOR2_X1 U4413 ( .A1(n3644), .A2(n3643), .ZN(n3645) );
  OAI211_X1 U4414 ( .C1(n3785), .C2(n4305), .A(n3646), .B(n3645), .ZN(U3213)
         );
  NAND2_X1 U4415 ( .A1(n3649), .A2(n3648), .ZN(n3650) );
  AOI21_X1 U4416 ( .B1(n3647), .B2(n3650), .A(n3771), .ZN(n3654) );
  AND2_X1 U4417 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4194) );
  AOI21_X1 U4418 ( .B1(n3779), .B2(n3955), .A(n4194), .ZN(n3652) );
  AOI22_X1 U4419 ( .A1(n3778), .A2(n4479), .B1(n3780), .B2(n3891), .ZN(n3651)
         );
  OAI211_X1 U4420 ( .C1(n3785), .C2(n4390), .A(n3652), .B(n3651), .ZN(n3653)
         );
  OR2_X1 U4421 ( .A1(n3654), .A2(n3653), .ZN(U3216) );
  INV_X1 U4422 ( .A(n3655), .ZN(n3657) );
  NAND2_X1 U4423 ( .A1(n3657), .A2(n3656), .ZN(n3661) );
  INV_X1 U4424 ( .A(n3659), .ZN(n3736) );
  OAI211_X1 U4425 ( .C1(n3658), .C2(n3736), .A(n3733), .B(n3661), .ZN(n3660)
         );
  OAI211_X1 U4426 ( .C1(n3662), .C2(n3661), .A(n3787), .B(n3660), .ZN(n3667)
         );
  AOI22_X1 U4427 ( .A1(n4460), .A2(n3779), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3666) );
  AOI22_X1 U4428 ( .A1(n3778), .A2(n3955), .B1(n3780), .B2(n4459), .ZN(n3665)
         );
  INV_X1 U4429 ( .A(n4339), .ZN(n3663) );
  OR2_X1 U4430 ( .A1(n3785), .A2(n3663), .ZN(n3664) );
  NAND4_X1 U4431 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(U3220)
         );
  NOR2_X1 U4432 ( .A1(n3669), .A2(n2221), .ZN(n3670) );
  XNOR2_X1 U4433 ( .A(n3671), .B(n3670), .ZN(n3676) );
  NOR2_X1 U4434 ( .A1(n3785), .A2(n4270), .ZN(n3674) );
  AOI22_X1 U4435 ( .A1(n4300), .A2(n3778), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3672) );
  OAI21_X1 U4436 ( .B1(n3088), .B2(n4267), .A(n3672), .ZN(n3673) );
  AOI211_X1 U4437 ( .C1(n3779), .C2(n4419), .A(n3674), .B(n3673), .ZN(n3675)
         );
  OAI21_X1 U4438 ( .B1(n3676), .B2(n3771), .A(n3675), .ZN(U3222) );
  INV_X1 U4439 ( .A(n3773), .ZN(n3678) );
  OAI21_X1 U4440 ( .B1(n3678), .B2(n3774), .A(n3677), .ZN(n3680) );
  XNOR2_X1 U4441 ( .A(n3680), .B(n3679), .ZN(n3687) );
  AND2_X1 U4442 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4615) );
  AOI21_X1 U4443 ( .B1(n3778), .B2(n3681), .A(n4615), .ZN(n3684) );
  AOI22_X1 U4444 ( .A1(n4487), .A2(n3682), .B1(n3779), .B2(n4490), .ZN(n3683)
         );
  OAI211_X1 U4445 ( .C1(n3785), .C2(n3685), .A(n3684), .B(n3683), .ZN(n3686)
         );
  AOI21_X1 U4446 ( .B1(n3687), .B2(n3787), .A(n3686), .ZN(n3688) );
  INV_X1 U4447 ( .A(n3688), .ZN(U3223) );
  OAI211_X1 U4448 ( .C1(n3689), .C2(n3691), .A(n3690), .B(n3787), .ZN(n3699)
         );
  AOI21_X1 U4449 ( .B1(n3778), .B2(n4103), .A(n3692), .ZN(n3698) );
  AOI22_X1 U4450 ( .A1(n3694), .A2(n3780), .B1(n3779), .B2(n3693), .ZN(n3697)
         );
  OR2_X1 U4451 ( .A1(n3785), .A2(n3695), .ZN(n3696) );
  NAND4_X1 U4452 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(U3224)
         );
  INV_X1 U4453 ( .A(n3700), .ZN(n3701) );
  NOR2_X1 U4454 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  XNOR2_X1 U4455 ( .A(n3704), .B(n3703), .ZN(n3709) );
  INV_X1 U4456 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3979) );
  NOR2_X1 U4457 ( .A1(STATE_REG_SCAN_IN), .A2(n3979), .ZN(n4625) );
  AOI21_X1 U4458 ( .B1(n3779), .B2(n4479), .A(n4625), .ZN(n3706) );
  AOI22_X1 U4459 ( .A1(n3778), .A2(n3957), .B1(n3780), .B2(n4478), .ZN(n3705)
         );
  OAI211_X1 U4460 ( .C1(n3785), .C2(n3707), .A(n3706), .B(n3705), .ZN(n3708)
         );
  AOI21_X1 U4461 ( .B1(n3709), .B2(n3787), .A(n3708), .ZN(n3710) );
  INV_X1 U4462 ( .A(n3710), .ZN(U3225) );
  NAND2_X1 U4463 ( .A1(n3712), .A2(n3711), .ZN(n3713) );
  XOR2_X1 U4464 ( .A(n3714), .B(n3713), .Z(n3722) );
  INV_X1 U4465 ( .A(n3785), .ZN(n3720) );
  OAI22_X1 U4466 ( .A1(n4285), .A2(n3715), .B1(n3088), .B2(n4280), .ZN(n3719)
         );
  OAI22_X1 U4467 ( .A1(n4445), .A2(n3717), .B1(STATE_REG_SCAN_IN), .B2(n3716), 
        .ZN(n3718) );
  AOI211_X1 U4468 ( .C1(n4282), .C2(n3720), .A(n3719), .B(n3718), .ZN(n3721)
         );
  OAI21_X1 U4469 ( .B1(n3722), .B2(n3771), .A(n3721), .ZN(U3226) );
  OAI211_X1 U4470 ( .C1(n3725), .C2(n3724), .A(n3723), .B(n3787), .ZN(n3732)
         );
  NAND2_X1 U4471 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n4146) );
  INV_X1 U4472 ( .A(n4146), .ZN(n3726) );
  AOI21_X1 U4473 ( .B1(n3778), .B2(n4104), .A(n3726), .ZN(n3731) );
  AOI22_X1 U4474 ( .A1(n3727), .A2(n3780), .B1(n3779), .B2(n4102), .ZN(n3730)
         );
  OR2_X1 U4475 ( .A1(n3785), .A2(n3728), .ZN(n3729) );
  NAND4_X1 U4476 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(U3227)
         );
  INV_X1 U4477 ( .A(n3733), .ZN(n3734) );
  NOR2_X1 U4478 ( .A1(n3736), .A2(n3734), .ZN(n3735) );
  OAI22_X1 U4479 ( .A1(n3737), .A2(n3736), .B1(n3735), .B2(n3658), .ZN(n3741)
         );
  AOI22_X1 U4480 ( .A1(n3779), .A2(n4361), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3739) );
  AOI22_X1 U4481 ( .A1(n3778), .A2(n3956), .B1(n3780), .B2(n3890), .ZN(n3738)
         );
  OAI211_X1 U4482 ( .C1(n3785), .C2(n4367), .A(n3739), .B(n3738), .ZN(n3740)
         );
  AOI21_X1 U4483 ( .B1(n3741), .B2(n3787), .A(n3740), .ZN(n3742) );
  INV_X1 U4484 ( .A(n3742), .ZN(U3230) );
  AOI21_X1 U4485 ( .B1(n3745), .B2(n3744), .A(n3743), .ZN(n3751) );
  AOI22_X1 U4486 ( .A1(n4441), .A2(n3779), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n3748) );
  INV_X1 U4487 ( .A(n4318), .ZN(n3746) );
  AOI22_X1 U4488 ( .A1(n3778), .A2(n4361), .B1(n3780), .B2(n3746), .ZN(n3747)
         );
  OAI211_X1 U4489 ( .C1(n3785), .C2(n4321), .A(n3748), .B(n3747), .ZN(n3749)
         );
  INV_X1 U4490 ( .A(n3749), .ZN(n3750) );
  OAI21_X1 U4491 ( .B1(n3751), .B2(n3771), .A(n3750), .ZN(U3232) );
  XNOR2_X1 U4492 ( .A(n3753), .B(n3752), .ZN(n3754) );
  XNOR2_X1 U4493 ( .A(n3755), .B(n3754), .ZN(n3762) );
  NAND2_X1 U4494 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4165) );
  INV_X1 U4495 ( .A(n4165), .ZN(n3756) );
  AOI21_X1 U4496 ( .B1(n3779), .B2(n3956), .A(n3756), .ZN(n3759) );
  AOI22_X1 U4497 ( .A1(n3778), .A2(n4490), .B1(n3780), .B2(n3757), .ZN(n3758)
         );
  OAI211_X1 U4498 ( .C1(n3785), .C2(n3760), .A(n3759), .B(n3758), .ZN(n3761)
         );
  AOI21_X1 U4499 ( .B1(n3762), .B2(n3787), .A(n3761), .ZN(n3763) );
  INV_X1 U4500 ( .A(n3763), .ZN(U3235) );
  NAND2_X1 U4501 ( .A1(n2059), .A2(n3764), .ZN(n3765) );
  XNOR2_X1 U4502 ( .A(n3766), .B(n3765), .ZN(n3772) );
  NOR2_X1 U4503 ( .A1(n4245), .A2(n3785), .ZN(n3769) );
  AOI22_X1 U4504 ( .A1(n4427), .A2(n3778), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3767) );
  OAI21_X1 U4505 ( .B1(n3088), .B2(n4250), .A(n3767), .ZN(n3768) );
  AOI211_X1 U4506 ( .C1(n3779), .C2(n4412), .A(n3769), .B(n3768), .ZN(n3770)
         );
  OAI21_X1 U4507 ( .B1(n3772), .B2(n3771), .A(n3770), .ZN(U3237) );
  NAND2_X1 U4508 ( .A1(n3773), .A2(n3677), .ZN(n3775) );
  XNOR2_X1 U4509 ( .A(n3775), .B(n3774), .ZN(n3788) );
  AOI21_X1 U4510 ( .B1(n3778), .B2(n3777), .A(n3776), .ZN(n3783) );
  AOI22_X1 U4511 ( .A1(n3781), .A2(n3780), .B1(n3779), .B2(n3957), .ZN(n3782)
         );
  OAI211_X1 U4512 ( .C1(n3785), .C2(n3784), .A(n3783), .B(n3782), .ZN(n3786)
         );
  AOI21_X1 U4513 ( .B1(n3788), .B2(n3787), .A(n3786), .ZN(n3789) );
  INV_X1 U4514 ( .A(n3789), .ZN(U3238) );
  NOR2_X1 U4515 ( .A1(n4430), .A2(n4418), .ZN(n3848) );
  INV_X1 U4516 ( .A(n3790), .ZN(n3793) );
  OAI211_X1 U4517 ( .C1(n3793), .C2(n3941), .A(n3792), .B(n3791), .ZN(n3796)
         );
  NAND3_X1 U4518 ( .A1(n3796), .A2(n3795), .A3(n3794), .ZN(n3799) );
  NAND3_X1 U4519 ( .A1(n3799), .A2(n3798), .A3(n3797), .ZN(n3802) );
  NAND3_X1 U4520 ( .A1(n3802), .A2(n3801), .A3(n3800), .ZN(n3805) );
  NAND3_X1 U4521 ( .A1(n3805), .A2(n3804), .A3(n3803), .ZN(n3808) );
  AOI21_X1 U4522 ( .B1(n3808), .B2(n3807), .A(n3806), .ZN(n3814) );
  NAND2_X1 U4523 ( .A1(n3810), .A2(n3809), .ZN(n3813) );
  OAI211_X1 U4524 ( .C1(n3814), .C2(n3813), .A(n3812), .B(n3811), .ZN(n3817)
         );
  NAND3_X1 U4525 ( .A1(n3817), .A2(n3816), .A3(n3815), .ZN(n3820) );
  AOI21_X1 U4526 ( .B1(n3820), .B2(n3819), .A(n2121), .ZN(n3828) );
  NAND3_X1 U4527 ( .A1(n3823), .A2(n3822), .A3(n3821), .ZN(n3827) );
  NAND2_X1 U4528 ( .A1(n3824), .A2(n3831), .ZN(n3912) );
  INV_X1 U4529 ( .A(n3912), .ZN(n3826) );
  OAI211_X1 U4530 ( .C1(n3828), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3834)
         );
  INV_X1 U4531 ( .A(n3829), .ZN(n3832) );
  AOI21_X1 U4532 ( .B1(n3832), .B2(n3831), .A(n2115), .ZN(n3911) );
  NAND3_X1 U4533 ( .A1(n3834), .A2(n3911), .A3(n3833), .ZN(n3837) );
  INV_X1 U4534 ( .A(n3835), .ZN(n3836) );
  AOI21_X1 U4535 ( .B1(n3837), .B2(n3916), .A(n3836), .ZN(n3838) );
  INV_X1 U4536 ( .A(n4291), .ZN(n3867) );
  OAI211_X1 U4537 ( .C1(n3838), .C2(n3919), .A(n3918), .B(n3867), .ZN(n3839)
         );
  NAND2_X1 U4538 ( .A1(n3923), .A2(n3839), .ZN(n3841) );
  NOR2_X1 U4539 ( .A1(n3866), .A2(n3886), .ZN(n3921) );
  INV_X1 U4540 ( .A(n3921), .ZN(n3840) );
  AOI211_X1 U4541 ( .C1(n3842), .C2(n3841), .A(n3928), .B(n3840), .ZN(n3847)
         );
  AND2_X1 U4542 ( .A1(n4407), .A2(n3859), .ZN(n3843) );
  NOR2_X1 U4543 ( .A1(n3844), .A2(n3843), .ZN(n3930) );
  INV_X1 U4544 ( .A(n3930), .ZN(n3845) );
  OR4_X1 U4545 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3864) );
  OR2_X1 U4546 ( .A1(n3850), .A2(n3849), .ZN(n3926) );
  NAND2_X1 U4547 ( .A1(n3851), .A2(REG1_REG_31__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U4548 ( .A1(n2297), .A2(REG2_REG_31__SCAN_IN), .ZN(n3854) );
  INV_X1 U4549 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4500) );
  OR2_X1 U4550 ( .A1(n3852), .A2(n4500), .ZN(n3853) );
  AND3_X1 U4551 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3936) );
  INV_X1 U4552 ( .A(n3936), .ZN(n4203) );
  NAND2_X1 U4553 ( .A1(n3856), .A2(DATAI_31_), .ZN(n4204) );
  NAND2_X1 U4554 ( .A1(n4203), .A2(n4204), .ZN(n3863) );
  NOR2_X1 U4555 ( .A1(n3857), .A2(n2932), .ZN(n4400) );
  INV_X1 U4556 ( .A(n4400), .ZN(n4403) );
  OR2_X1 U4557 ( .A1(n3954), .A2(n4403), .ZN(n3858) );
  AND2_X1 U4558 ( .A1(n3863), .A2(n3858), .ZN(n3887) );
  OAI21_X1 U4559 ( .B1(n4407), .B2(n3859), .A(n3887), .ZN(n3925) );
  AOI21_X1 U4560 ( .B1(n3926), .B2(n3930), .A(n3925), .ZN(n3933) );
  NOR2_X1 U4561 ( .A1(n4203), .A2(n4204), .ZN(n3938) );
  INV_X1 U4562 ( .A(n3938), .ZN(n3861) );
  AND2_X1 U4563 ( .A1(n3954), .A2(n4403), .ZN(n3939) );
  INV_X1 U4564 ( .A(n3939), .ZN(n3860) );
  AND2_X1 U4565 ( .A1(n3861), .A2(n3860), .ZN(n3888) );
  INV_X1 U4566 ( .A(n3888), .ZN(n3862) );
  AOI22_X1 U4567 ( .A1(n3864), .A2(n3933), .B1(n3863), .B2(n3862), .ZN(n3946)
         );
  INV_X1 U4568 ( .A(n4214), .ZN(n3908) );
  XNOR2_X1 U4569 ( .A(n4419), .B(n4250), .ZN(n4243) );
  INV_X1 U4570 ( .A(n4259), .ZN(n3865) );
  NOR2_X1 U4571 ( .A1(n3866), .A2(n3865), .ZN(n4278) );
  AND2_X1 U4572 ( .A1(n3867), .A2(n4292), .ZN(n4331) );
  INV_X1 U4573 ( .A(n3868), .ZN(n3869) );
  AND4_X1 U4574 ( .A1(n2243), .A2(n3871), .A3(n3870), .A4(n3869), .ZN(n3874)
         );
  AND4_X1 U4575 ( .A1(n4331), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3882)
         );
  INV_X1 U4576 ( .A(n3875), .ZN(n3876) );
  AND4_X1 U4577 ( .A1(n4316), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3881)
         );
  NOR2_X1 U4578 ( .A1(n3879), .A2(n4660), .ZN(n3880) );
  NAND4_X1 U4579 ( .A1(n4278), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3907)
         );
  NAND2_X1 U4580 ( .A1(n4238), .A2(n3883), .ZN(n4262) );
  INV_X1 U4581 ( .A(n3884), .ZN(n3885) );
  NOR2_X1 U4582 ( .A1(n3886), .A2(n3885), .ZN(n4296) );
  NAND3_X1 U4583 ( .A1(n4296), .A2(n3888), .A3(n3887), .ZN(n3889) );
  NOR2_X1 U4584 ( .A1(n4262), .A2(n3889), .ZN(n3905) );
  XNOR2_X1 U4585 ( .A(n3955), .B(n3890), .ZN(n4357) );
  XNOR2_X1 U4586 ( .A(n3956), .B(n3891), .ZN(n4380) );
  NOR2_X1 U4587 ( .A1(n3893), .A2(n3892), .ZN(n3903) );
  NOR2_X1 U4588 ( .A1(n3895), .A2(n3894), .ZN(n3902) );
  NOR2_X1 U4589 ( .A1(n3897), .A2(n3896), .ZN(n3901) );
  NOR2_X1 U4590 ( .A1(n3899), .A2(n3898), .ZN(n3900) );
  AND4_X1 U4591 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3904)
         );
  NAND4_X1 U4592 ( .A1(n3905), .A2(n4357), .A3(n4380), .A4(n3904), .ZN(n3906)
         );
  OR4_X1 U4593 ( .A1(n3908), .A2(n4243), .A3(n3907), .A4(n3906), .ZN(n3910) );
  NOR3_X1 U4594 ( .A1(n3910), .A2(n3909), .A3(n4222), .ZN(n3943) );
  INV_X1 U4595 ( .A(n4204), .ZN(n3940) );
  OAI21_X1 U4596 ( .B1(n3913), .B2(n3912), .A(n3911), .ZN(n3917) );
  INV_X1 U4597 ( .A(n3914), .ZN(n3915) );
  AOI21_X1 U4598 ( .B1(n3917), .B2(n3916), .A(n3915), .ZN(n3920) );
  OAI21_X1 U4599 ( .B1(n3920), .B2(n3919), .A(n3918), .ZN(n3922) );
  OAI221_X1 U4600 ( .B1(n3924), .B2(n3923), .C1(n3924), .C2(n3922), .A(n3921), 
        .ZN(n3927) );
  AOI211_X1 U4601 ( .C1(n4240), .C2(n3927), .A(n3926), .B(n3925), .ZN(n3934)
         );
  NAND3_X1 U4602 ( .A1(n3931), .A2(n3930), .A3(n3929), .ZN(n3932) );
  AOI22_X1 U4603 ( .A1(n3934), .A2(n2129), .B1(n3933), .B2(n3932), .ZN(n3935)
         );
  AOI21_X1 U4604 ( .B1(n4400), .B2(n3936), .A(n3935), .ZN(n3937) );
  AOI211_X1 U4605 ( .C1(n3940), .C2(n3939), .A(n3938), .B(n3937), .ZN(n3942)
         );
  MUX2_X1 U4606 ( .A(n3943), .B(n3942), .S(n3941), .Z(n3945) );
  MUX2_X1 U4607 ( .A(n3946), .B(n3945), .S(n3944), .Z(n3947) );
  XNOR2_X1 U4608 ( .A(n3947), .B(n4190), .ZN(n3953) );
  NAND2_X1 U4609 ( .A1(n3948), .A2(n4125), .ZN(n3949) );
  OAI211_X1 U4610 ( .C1(n3950), .C2(n3952), .A(n3949), .B(B_REG_SCAN_IN), .ZN(
        n3951) );
  OAI21_X1 U4611 ( .B1(n3953), .B2(n3952), .A(n3951), .ZN(U3239) );
  MUX2_X1 U4612 ( .A(DATAO_REG_31__SCAN_IN), .B(n4203), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4613 ( .A(DATAO_REG_30__SCAN_IN), .B(n3954), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4614 ( .A(DATAO_REG_29__SCAN_IN), .B(n4407), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4615 ( .A(DATAO_REG_28__SCAN_IN), .B(n4233), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4616 ( .A(DATAO_REG_27__SCAN_IN), .B(n4412), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4617 ( .A(DATAO_REG_25__SCAN_IN), .B(n4427), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4618 ( .A(DATAO_REG_24__SCAN_IN), .B(n4300), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4619 ( .A(DATAO_REG_23__SCAN_IN), .B(n4441), .S(n3960), .Z(U3573)
         );
  MUX2_X1 U4620 ( .A(DATAO_REG_22__SCAN_IN), .B(n4460), .S(n3960), .Z(U3572)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_21__SCAN_IN), .B(n4361), .S(n3960), .Z(U3571)
         );
  MUX2_X1 U4622 ( .A(DATAO_REG_20__SCAN_IN), .B(n3955), .S(n3960), .Z(U3570)
         );
  MUX2_X1 U4623 ( .A(DATAO_REG_19__SCAN_IN), .B(n3956), .S(n3960), .Z(U3569)
         );
  MUX2_X1 U4624 ( .A(DATAO_REG_17__SCAN_IN), .B(n4490), .S(n3960), .Z(U3567)
         );
  MUX2_X1 U4625 ( .A(DATAO_REG_16__SCAN_IN), .B(n3957), .S(n3960), .Z(U3566)
         );
  MUX2_X1 U4626 ( .A(DATAO_REG_13__SCAN_IN), .B(n3958), .S(n3960), .Z(U3563)
         );
  MUX2_X1 U4627 ( .A(DATAO_REG_11__SCAN_IN), .B(n3959), .S(n3960), .Z(U3561)
         );
  MUX2_X1 U4628 ( .A(DATAO_REG_10__SCAN_IN), .B(n3961), .S(n3960), .Z(U3560)
         );
  MUX2_X1 U4629 ( .A(DATAO_REG_9__SCAN_IN), .B(n3962), .S(U4043), .Z(n4101) );
  INV_X1 U4630 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3965) );
  INV_X1 U4631 ( .A(keyinput23), .ZN(n3964) );
  OAI22_X1 U4632 ( .A1(n3965), .A2(keyinput46), .B1(n3964), .B2(
        REG1_REG_25__SCAN_IN), .ZN(n3963) );
  AOI221_X1 U4633 ( .B1(n3965), .B2(keyinput46), .C1(REG1_REG_25__SCAN_IN), 
        .C2(n3964), .A(n3963), .ZN(n3974) );
  INV_X1 U4634 ( .A(keyinput51), .ZN(n3967) );
  OAI22_X1 U4635 ( .A1(n4541), .A2(keyinput9), .B1(n3967), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n3966) );
  AOI221_X1 U4636 ( .B1(n4541), .B2(keyinput9), .C1(DATAO_REG_26__SCAN_IN), 
        .C2(n3967), .A(n3966), .ZN(n3973) );
  OAI22_X1 U4637 ( .A1(n3969), .A2(keyinput18), .B1(n3218), .B2(keyinput21), 
        .ZN(n3968) );
  AOI221_X1 U4638 ( .B1(n3969), .B2(keyinput18), .C1(keyinput21), .C2(n3218), 
        .A(n3968), .ZN(n3972) );
  INV_X1 U4639 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4406) );
  OAI22_X1 U4640 ( .A1(n4513), .A2(keyinput48), .B1(n4406), .B2(keyinput57), 
        .ZN(n3970) );
  AOI221_X1 U4641 ( .B1(n4513), .B2(keyinput48), .C1(keyinput57), .C2(n4406), 
        .A(n3970), .ZN(n3971) );
  NAND4_X1 U4642 ( .A1(n3974), .A2(n3973), .A3(n3972), .A4(n3971), .ZN(n4099)
         );
  INV_X1 U4643 ( .A(D_REG_22__SCAN_IN), .ZN(n4669) );
  INV_X1 U4644 ( .A(D_REG_28__SCAN_IN), .ZN(n4666) );
  OAI22_X1 U4645 ( .A1(n4669), .A2(keyinput37), .B1(n4666), .B2(keyinput1), 
        .ZN(n3975) );
  AOI221_X1 U4646 ( .B1(n4669), .B2(keyinput37), .C1(keyinput1), .C2(n4666), 
        .A(n3975), .ZN(n3986) );
  INV_X1 U4647 ( .A(D_REG_7__SCAN_IN), .ZN(n4672) );
  INV_X1 U4648 ( .A(D_REG_25__SCAN_IN), .ZN(n4667) );
  OAI22_X1 U4649 ( .A1(n4672), .A2(keyinput58), .B1(n4667), .B2(keyinput62), 
        .ZN(n3976) );
  AOI221_X1 U4650 ( .B1(n4672), .B2(keyinput58), .C1(keyinput62), .C2(n4667), 
        .A(n3976), .ZN(n3985) );
  INV_X1 U4651 ( .A(keyinput19), .ZN(n3978) );
  OAI22_X1 U4652 ( .A1(n3979), .A2(keyinput3), .B1(n3978), .B2(
        REG0_REG_17__SCAN_IN), .ZN(n3977) );
  AOI221_X1 U4653 ( .B1(n3979), .B2(keyinput3), .C1(REG0_REG_17__SCAN_IN), 
        .C2(n3978), .A(n3977), .ZN(n3984) );
  INV_X1 U4654 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3982) );
  INV_X1 U4655 ( .A(keyinput45), .ZN(n3981) );
  OAI22_X1 U4656 ( .A1(n3982), .A2(keyinput50), .B1(n3981), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n3980) );
  AOI221_X1 U4657 ( .B1(n3982), .B2(keyinput50), .C1(DATAO_REG_18__SCAN_IN), 
        .C2(n3981), .A(n3980), .ZN(n3983) );
  NAND4_X1 U4658 ( .A1(n3986), .A2(n3985), .A3(n3984), .A4(n3983), .ZN(n4098)
         );
  NAND2_X1 U4659 ( .A1(n2106), .A2(keyinput35), .ZN(n3987) );
  OAI221_X1 U4660 ( .B1(n3988), .B2(keyinput13), .C1(n2106), .C2(keyinput35), 
        .A(n3987), .ZN(n4000) );
  INV_X1 U4661 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3991) );
  INV_X1 U4662 ( .A(keyinput4), .ZN(n3990) );
  AOI22_X1 U4663 ( .A1(n3991), .A2(keyinput54), .B1(DATAO_REG_8__SCAN_IN), 
        .B2(n3990), .ZN(n3989) );
  OAI221_X1 U4664 ( .B1(n3991), .B2(keyinput54), .C1(n3990), .C2(
        DATAO_REG_8__SCAN_IN), .A(n3989), .ZN(n3999) );
  INV_X1 U4665 ( .A(keyinput63), .ZN(n4053) );
  INV_X1 U4666 ( .A(keyinput41), .ZN(n3993) );
  AOI22_X1 U4667 ( .A1(n4053), .A2(DATAO_REG_12__SCAN_IN), .B1(
        DATAO_REG_6__SCAN_IN), .B2(n3993), .ZN(n3992) );
  OAI221_X1 U4668 ( .B1(n4053), .B2(DATAO_REG_12__SCAN_IN), .C1(n3993), .C2(
        DATAO_REG_6__SCAN_IN), .A(n3992), .ZN(n3998) );
  INV_X1 U4669 ( .A(keyinput8), .ZN(n3996) );
  INV_X1 U4670 ( .A(keyinput20), .ZN(n3995) );
  AOI22_X1 U4671 ( .A1(n3996), .A2(DATAO_REG_2__SCAN_IN), .B1(
        DATAO_REG_15__SCAN_IN), .B2(n3995), .ZN(n3994) );
  OAI221_X1 U4672 ( .B1(n3996), .B2(DATAO_REG_2__SCAN_IN), .C1(n3995), .C2(
        DATAO_REG_15__SCAN_IN), .A(n3994), .ZN(n3997) );
  NOR4_X1 U4673 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4039)
         );
  INV_X1 U4674 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4003) );
  INV_X1 U4675 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4676 ( .A1(n4003), .A2(keyinput52), .B1(keyinput53), .B2(n4002), 
        .ZN(n4001) );
  OAI221_X1 U4677 ( .B1(n4003), .B2(keyinput52), .C1(n4002), .C2(keyinput53), 
        .A(n4001), .ZN(n4014) );
  INV_X1 U4678 ( .A(keyinput24), .ZN(n4006) );
  INV_X1 U4679 ( .A(keyinput28), .ZN(n4005) );
  AOI22_X1 U4680 ( .A1(n4006), .A2(DATAO_REG_14__SCAN_IN), .B1(
        DATAO_REG_7__SCAN_IN), .B2(n4005), .ZN(n4004) );
  OAI221_X1 U4681 ( .B1(n4006), .B2(DATAO_REG_14__SCAN_IN), .C1(n4005), .C2(
        DATAO_REG_7__SCAN_IN), .A(n4004), .ZN(n4013) );
  INV_X1 U4682 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U4683 ( .A1(n4569), .A2(keyinput38), .B1(n4008), .B2(keyinput40), 
        .ZN(n4007) );
  OAI221_X1 U4684 ( .B1(n4569), .B2(keyinput38), .C1(n4008), .C2(keyinput40), 
        .A(n4007), .ZN(n4012) );
  XNOR2_X1 U4685 ( .A(REG3_REG_2__SCAN_IN), .B(keyinput14), .ZN(n4010) );
  XNOR2_X1 U4686 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput31), .ZN(n4009) );
  NAND2_X1 U4687 ( .A1(n4010), .A2(n4009), .ZN(n4011) );
  NOR4_X1 U4688 ( .A1(n4014), .A2(n4013), .A3(n4012), .A4(n4011), .ZN(n4038)
         );
  INV_X1 U4689 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U4690 ( .A1(n4162), .A2(keyinput36), .B1(keyinput30), .B2(n4016), 
        .ZN(n4015) );
  OAI221_X1 U4691 ( .B1(n4162), .B2(keyinput36), .C1(n4016), .C2(keyinput30), 
        .A(n4015), .ZN(n4025) );
  INV_X1 U4692 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4709) );
  INV_X1 U4693 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U4694 ( .A1(n4709), .A2(keyinput39), .B1(keyinput34), .B2(n4147), 
        .ZN(n4017) );
  OAI221_X1 U4695 ( .B1(n4709), .B2(keyinput39), .C1(n4147), .C2(keyinput34), 
        .A(n4017), .ZN(n4024) );
  AOI22_X1 U4696 ( .A1(n4019), .A2(keyinput44), .B1(n2398), .B2(keyinput60), 
        .ZN(n4018) );
  OAI221_X1 U4697 ( .B1(n4019), .B2(keyinput44), .C1(n2398), .C2(keyinput60), 
        .A(n4018), .ZN(n4023) );
  XNOR2_X1 U4698 ( .A(IR_REG_6__SCAN_IN), .B(keyinput11), .ZN(n4021) );
  XNOR2_X1 U4699 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput0), .ZN(n4020) );
  NAND2_X1 U4700 ( .A1(n4021), .A2(n4020), .ZN(n4022) );
  NOR4_X1 U4701 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4037)
         );
  INV_X1 U4702 ( .A(IR_REG_1__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4703 ( .A1(n4027), .A2(keyinput55), .B1(keyinput27), .B2(n3140), 
        .ZN(n4026) );
  OAI221_X1 U4704 ( .B1(n4027), .B2(keyinput55), .C1(n3140), .C2(keyinput27), 
        .A(n4026), .ZN(n4035) );
  INV_X1 U4705 ( .A(DATAI_9_), .ZN(n4029) );
  AOI22_X1 U4706 ( .A1(n4029), .A2(keyinput7), .B1(n2585), .B2(keyinput56), 
        .ZN(n4028) );
  OAI221_X1 U4707 ( .B1(n4029), .B2(keyinput7), .C1(n2585), .C2(keyinput56), 
        .A(n4028), .ZN(n4034) );
  INV_X1 U4708 ( .A(D_REG_11__SCAN_IN), .ZN(n4671) );
  INV_X1 U4709 ( .A(D_REG_23__SCAN_IN), .ZN(n4668) );
  AOI22_X1 U4710 ( .A1(n4671), .A2(keyinput25), .B1(keyinput5), .B2(n4668), 
        .ZN(n4030) );
  OAI221_X1 U4711 ( .B1(n4671), .B2(keyinput25), .C1(n4668), .C2(keyinput5), 
        .A(n4030), .ZN(n4033) );
  INV_X1 U4712 ( .A(D_REG_21__SCAN_IN), .ZN(n4670) );
  INV_X1 U4713 ( .A(D_REG_30__SCAN_IN), .ZN(n4665) );
  AOI22_X1 U4714 ( .A1(n4670), .A2(keyinput15), .B1(keyinput43), .B2(n4665), 
        .ZN(n4031) );
  OAI221_X1 U4715 ( .B1(n4670), .B2(keyinput15), .C1(n4665), .C2(keyinput43), 
        .A(n4031), .ZN(n4032) );
  NOR4_X1 U4716 ( .A1(n4035), .A2(n4034), .A3(n4033), .A4(n4032), .ZN(n4036)
         );
  NAND4_X1 U4717 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4097)
         );
  NOR3_X1 U4718 ( .A1(keyinput43), .A2(keyinput58), .A3(keyinput37), .ZN(n4044) );
  NOR4_X1 U4719 ( .A1(keyinput45), .A2(keyinput9), .A3(keyinput23), .A4(
        keyinput51), .ZN(n4043) );
  NOR3_X1 U4720 ( .A1(keyinput50), .A2(keyinput19), .A3(keyinput3), .ZN(n4041)
         );
  NOR3_X1 U4721 ( .A1(keyinput48), .A2(keyinput18), .A3(keyinput57), .ZN(n4040) );
  AND4_X1 U4722 ( .A1(keyinput1), .A2(n4041), .A3(keyinput46), .A4(n4040), 
        .ZN(n4042) );
  NAND4_X1 U4723 ( .A1(keyinput62), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(
        n4051) );
  NAND3_X1 U4724 ( .A1(keyinput42), .A2(keyinput32), .A3(keyinput16), .ZN(
        n4050) );
  NOR2_X1 U4725 ( .A1(keyinput21), .A2(keyinput6), .ZN(n4048) );
  NAND4_X1 U4726 ( .A1(keyinput2), .A2(keyinput10), .A3(keyinput59), .A4(
        keyinput47), .ZN(n4046) );
  NAND2_X1 U4727 ( .A1(keyinput49), .A2(keyinput29), .ZN(n4045) );
  NOR4_X1 U4728 ( .A1(keyinput33), .A2(keyinput61), .A3(n4046), .A4(n4045), 
        .ZN(n4047) );
  NAND4_X1 U4729 ( .A1(keyinput22), .A2(keyinput26), .A3(n4048), .A4(n4047), 
        .ZN(n4049) );
  NOR4_X1 U4730 ( .A1(keyinput12), .A2(n4051), .A3(n4050), .A4(n4049), .ZN(
        n4068) );
  NAND2_X1 U4731 ( .A1(keyinput52), .A2(keyinput28), .ZN(n4052) );
  NOR3_X1 U4732 ( .A1(keyinput20), .A2(keyinput24), .A3(n4052), .ZN(n4058) );
  NOR3_X1 U4733 ( .A1(keyinput53), .A2(keyinput38), .A3(keyinput40), .ZN(n4057) );
  INV_X1 U4734 ( .A(keyinput35), .ZN(n4055) );
  NAND4_X1 U4735 ( .A1(keyinput4), .A2(keyinput41), .A3(keyinput8), .A4(n4053), 
        .ZN(n4054) );
  NOR4_X1 U4736 ( .A1(keyinput17), .A2(keyinput54), .A3(n4055), .A4(n4054), 
        .ZN(n4056) );
  NAND4_X1 U4737 ( .A1(n4058), .A2(keyinput31), .A3(n4057), .A4(n4056), .ZN(
        n4066) );
  NAND3_X1 U4738 ( .A1(keyinput25), .A2(keyinput5), .A3(keyinput15), .ZN(n4065) );
  NAND2_X1 U4739 ( .A1(keyinput36), .A2(keyinput34), .ZN(n4059) );
  NOR3_X1 U4740 ( .A1(keyinput14), .A2(keyinput39), .A3(n4059), .ZN(n4063) );
  NAND2_X1 U4741 ( .A1(keyinput0), .A2(keyinput30), .ZN(n4060) );
  NOR3_X1 U4742 ( .A1(keyinput60), .A2(keyinput44), .A3(n4060), .ZN(n4062) );
  NOR3_X1 U4743 ( .A1(keyinput11), .A2(keyinput55), .A3(keyinput27), .ZN(n4061) );
  NAND4_X1 U4744 ( .A1(n4063), .A2(n4062), .A3(keyinput7), .A4(n4061), .ZN(
        n4064) );
  NOR4_X1 U4745 ( .A1(keyinput56), .A2(n4066), .A3(n4065), .A4(n4064), .ZN(
        n4067) );
  AOI21_X1 U4746 ( .B1(n4068), .B2(n4067), .A(keyinput13), .ZN(n4095) );
  INV_X1 U4747 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U4748 ( .A1(n4071), .A2(keyinput49), .B1(n4070), .B2(keyinput33), 
        .ZN(n4069) );
  OAI221_X1 U4749 ( .B1(n4071), .B2(keyinput49), .C1(n4070), .C2(keyinput33), 
        .A(n4069), .ZN(n4081) );
  INV_X1 U4750 ( .A(DATAI_24_), .ZN(n4074) );
  INV_X1 U4751 ( .A(IR_REG_22__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4752 ( .A1(n4074), .A2(keyinput17), .B1(n4073), .B2(keyinput29), 
        .ZN(n4072) );
  OAI221_X1 U4753 ( .B1(n4074), .B2(keyinput17), .C1(n4073), .C2(keyinput29), 
        .A(n4072), .ZN(n4080) );
  XNOR2_X1 U4754 ( .A(IR_REG_16__SCAN_IN), .B(keyinput61), .ZN(n4078) );
  XNOR2_X1 U4755 ( .A(D_REG_0__SCAN_IN), .B(keyinput12), .ZN(n4077) );
  XNOR2_X1 U4756 ( .A(IR_REG_24__SCAN_IN), .B(keyinput32), .ZN(n4076) );
  XNOR2_X1 U4757 ( .A(IR_REG_21__SCAN_IN), .B(keyinput16), .ZN(n4075) );
  NAND4_X1 U4758 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NOR3_X1 U4759 ( .A1(n4081), .A2(n4080), .A3(n4079), .ZN(n4094) );
  AOI22_X1 U4760 ( .A1(n2484), .A2(keyinput47), .B1(keyinput42), .B2(n4083), 
        .ZN(n4082) );
  OAI221_X1 U4761 ( .B1(n2484), .B2(keyinput47), .C1(n4083), .C2(keyinput42), 
        .A(n4082), .ZN(n4092) );
  INV_X1 U4762 ( .A(DATAI_8_), .ZN(n4085) );
  AOI22_X1 U4763 ( .A1(n4085), .A2(keyinput10), .B1(keyinput59), .B2(n2292), 
        .ZN(n4084) );
  OAI221_X1 U4764 ( .B1(n4085), .B2(keyinput10), .C1(n2292), .C2(keyinput59), 
        .A(n4084), .ZN(n4091) );
  XOR2_X1 U4765 ( .A(n4500), .B(keyinput6), .Z(n4089) );
  XNOR2_X1 U4766 ( .A(IR_REG_23__SCAN_IN), .B(keyinput2), .ZN(n4088) );
  XNOR2_X1 U4767 ( .A(DATAI_12_), .B(keyinput22), .ZN(n4087) );
  XNOR2_X1 U4768 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput26), .ZN(n4086) );
  NAND4_X1 U4769 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  NOR3_X1 U4770 ( .A1(n4092), .A2(n4091), .A3(n4090), .ZN(n4093) );
  OAI211_X1 U4771 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4095), .A(n4094), .B(n4093), .ZN(n4096) );
  NOR4_X1 U4772 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4100)
         );
  XOR2_X1 U4773 ( .A(n4101), .B(n4100), .Z(U3559) );
  MUX2_X1 U4774 ( .A(DATAO_REG_5__SCAN_IN), .B(n4102), .S(n3960), .Z(U3555) );
  MUX2_X1 U4775 ( .A(DATAO_REG_4__SCAN_IN), .B(n4103), .S(n3960), .Z(U3554) );
  MUX2_X1 U4776 ( .A(DATAO_REG_3__SCAN_IN), .B(n4104), .S(n3960), .Z(U3553) );
  MUX2_X1 U4777 ( .A(DATAO_REG_1__SCAN_IN), .B(n2696), .S(n3960), .Z(U3551) );
  MUX2_X1 U4778 ( .A(DATAO_REG_0__SCAN_IN), .B(n2691), .S(n3960), .Z(U3550) );
  INV_X1 U4779 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4105) );
  NAND3_X1 U4780 ( .A1(n4627), .A2(n4105), .A3(IR_REG_0__SCAN_IN), .ZN(n4114)
         );
  AOI22_X1 U4781 ( .A1(n4626), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4113) );
  INV_X1 U4782 ( .A(n4555), .ZN(n4106) );
  AOI21_X1 U4783 ( .B1(n4106), .B2(n4105), .A(IR_REG_0__SCAN_IN), .ZN(n4111)
         );
  INV_X1 U4784 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4107) );
  AND2_X1 U4785 ( .A1(n4555), .A2(n4107), .ZN(n4108) );
  OR2_X1 U4786 ( .A1(n4108), .A2(n4564), .ZN(n4110) );
  INV_X1 U4787 ( .A(IR_REG_0__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U4788 ( .A1(n4110), .A2(n4686), .ZN(n4127) );
  OAI211_X1 U4789 ( .C1(n4111), .C2(n4110), .A(n4109), .B(n4127), .ZN(n4112)
         );
  NAND3_X1 U4790 ( .A1(n4114), .A2(n4113), .A3(n4112), .ZN(U3240) );
  NAND2_X1 U4791 ( .A1(n4180), .A2(n4563), .ZN(n4122) );
  AOI22_X1 U4792 ( .A1(n4626), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4121) );
  OAI211_X1 U4793 ( .C1(n4117), .C2(n4116), .A(n4627), .B(n4115), .ZN(n4120)
         );
  OAI211_X1 U4794 ( .C1(n4124), .C2(n4118), .A(n4593), .B(n4137), .ZN(n4119)
         );
  NAND4_X1 U4795 ( .A1(n4122), .A2(n4121), .A3(n4120), .A4(n4119), .ZN(U3241)
         );
  OR3_X1 U4796 ( .A1(n4123), .A2(n4555), .A3(n4564), .ZN(n4128) );
  NAND2_X1 U4797 ( .A1(n4125), .A2(n4124), .ZN(n4126) );
  NAND4_X1 U4798 ( .A1(n4128), .A2(U4043), .A3(n4127), .A4(n4126), .ZN(n4156)
         );
  NOR2_X1 U4799 ( .A1(n4129), .A2(STATE_REG_SCAN_IN), .ZN(n4130) );
  AOI21_X1 U4800 ( .B1(n4626), .B2(ADDR_REG_2__SCAN_IN), .A(n4130), .ZN(n4131)
         );
  OAI21_X1 U4801 ( .B1(n4633), .B2(n4133), .A(n4131), .ZN(n4132) );
  INV_X1 U4802 ( .A(n4132), .ZN(n4145) );
  MUX2_X1 U4803 ( .A(REG2_REG_2__SCAN_IN), .B(n4134), .S(n4133), .Z(n4135) );
  NAND3_X1 U4804 ( .A1(n4137), .A2(n4136), .A3(n4135), .ZN(n4138) );
  NAND3_X1 U4805 ( .A1(n4593), .A2(n4139), .A3(n4138), .ZN(n4144) );
  OAI211_X1 U4806 ( .C1(n4142), .C2(n4141), .A(n4627), .B(n4140), .ZN(n4143)
         );
  NAND4_X1 U4807 ( .A1(n4156), .A2(n4145), .A3(n4144), .A4(n4143), .ZN(U3242)
         );
  OAI21_X1 U4808 ( .B1(n4167), .B2(n4147), .A(n4146), .ZN(n4148) );
  AOI21_X1 U4809 ( .B1(n4180), .B2(n4561), .A(n4148), .ZN(n4155) );
  XOR2_X1 U4810 ( .A(REG2_REG_4__SCAN_IN), .B(n4149), .Z(n4150) );
  NAND2_X1 U4811 ( .A1(n4593), .A2(n4150), .ZN(n4154) );
  OAI211_X1 U4812 ( .C1(REG1_REG_4__SCAN_IN), .C2(n4152), .A(n4627), .B(n4151), 
        .ZN(n4153) );
  NAND4_X1 U4813 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(U3244)
         );
  NOR2_X1 U4814 ( .A1(n4175), .A2(REG1_REG_17__SCAN_IN), .ZN(n4163) );
  NOR2_X1 U4815 ( .A1(n4159), .A2(n4160), .ZN(n4161) );
  NOR2_X1 U4816 ( .A1(n4161), .A2(n4617), .ZN(n4629) );
  AOI22_X1 U4817 ( .A1(n4175), .A2(n4162), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4677), .ZN(n4628) );
  XNOR2_X1 U4818 ( .A(n4164), .B(REG1_REG_18__SCAN_IN), .ZN(n4183) );
  XNOR2_X1 U4819 ( .A(n4184), .B(n4183), .ZN(n4182) );
  INV_X1 U4820 ( .A(ADDR_REG_18__SCAN_IN), .ZN(n4166) );
  OAI21_X1 U4821 ( .B1(n4167), .B2(n4166), .A(n4165), .ZN(n4179) );
  NOR2_X1 U4822 ( .A1(n4189), .A2(n4168), .ZN(n4169) );
  AOI21_X1 U4823 ( .B1(n4189), .B2(n4168), .A(n4169), .ZN(n4177) );
  NOR2_X1 U4824 ( .A1(n4175), .A2(REG2_REG_17__SCAN_IN), .ZN(n4170) );
  AOI21_X1 U4825 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4175), .A(n4170), .ZN(n4623) );
  NAND2_X1 U4826 ( .A1(n4173), .A2(n4679), .ZN(n4174) );
  INV_X1 U4827 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4611) );
  AOI211_X1 U4828 ( .C1(n4177), .C2(n4176), .A(n4188), .B(n4620), .ZN(n4178)
         );
  AOI211_X1 U4829 ( .C1(n4180), .C2(n4189), .A(n4179), .B(n4178), .ZN(n4181)
         );
  OAI21_X1 U4830 ( .B1(n4200), .B2(n4182), .A(n4181), .ZN(U3258) );
  AOI22_X1 U4831 ( .A1(n4184), .A2(n4183), .B1(REG1_REG_18__SCAN_IN), .B2(
        n4189), .ZN(n4187) );
  INV_X1 U4832 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4185) );
  MUX2_X1 U4833 ( .A(n4185), .B(REG1_REG_19__SCAN_IN), .S(n4190), .Z(n4186) );
  XNOR2_X1 U4834 ( .A(n4187), .B(n4186), .ZN(n4201) );
  AOI21_X1 U4835 ( .B1(n4189), .B2(REG2_REG_18__SCAN_IN), .A(n4188), .ZN(n4193) );
  INV_X1 U4836 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4191) );
  MUX2_X1 U4837 ( .A(REG2_REG_19__SCAN_IN), .B(n4191), .S(n4190), .Z(n4192) );
  XNOR2_X1 U4838 ( .A(n4193), .B(n4192), .ZN(n4198) );
  AOI21_X1 U4839 ( .B1(n4626), .B2(ADDR_REG_19__SCAN_IN), .A(n4194), .ZN(n4195) );
  OAI21_X1 U4840 ( .B1(n4633), .B2(n4196), .A(n4195), .ZN(n4197) );
  AOI21_X1 U4841 ( .B1(n4198), .B2(n4593), .A(n4197), .ZN(n4199) );
  OAI21_X1 U4842 ( .B1(n4201), .B2(n4200), .A(n4199), .ZN(U3259) );
  XNOR2_X1 U4843 ( .A(n4398), .B(n4204), .ZN(n4504) );
  NAND2_X1 U4844 ( .A1(n4203), .A2(n4202), .ZN(n4402) );
  OAI21_X1 U4845 ( .B1(n4204), .B2(n4409), .A(n4402), .ZN(n4502) );
  NAND2_X1 U4846 ( .A1(n4502), .A2(n4566), .ZN(n4206) );
  NAND2_X1 U4847 ( .A1(n4664), .A2(REG2_REG_31__SCAN_IN), .ZN(n4205) );
  OAI211_X1 U4848 ( .C1(n4504), .C2(n4389), .A(n4206), .B(n4205), .ZN(U3260)
         );
  XNOR2_X1 U4849 ( .A(n4207), .B(n4214), .ZN(n4415) );
  INV_X1 U4850 ( .A(n4208), .ZN(n4209) );
  OAI21_X1 U4851 ( .B1(n4227), .B2(n4408), .A(n4209), .ZN(n4511) );
  INV_X1 U4852 ( .A(n4511), .ZN(n4219) );
  AOI22_X1 U4853 ( .A1(n4412), .A2(n4247), .B1(n4407), .B2(n4337), .ZN(n4212)
         );
  AOI22_X1 U4854 ( .A1(n4338), .A2(n4210), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4664), .ZN(n4211) );
  OAI211_X1 U4855 ( .C1(n4213), .C2(n4634), .A(n4212), .B(n4211), .ZN(n4218)
         );
  XNOR2_X1 U4856 ( .A(n4215), .B(n4214), .ZN(n4216) );
  NAND2_X1 U4857 ( .A1(n4216), .A2(n4329), .ZN(n4413) );
  NOR2_X1 U4858 ( .A1(n4413), .A2(n4664), .ZN(n4217) );
  AOI211_X1 U4859 ( .C1(n4651), .C2(n4219), .A(n4218), .B(n4217), .ZN(n4220)
         );
  OAI21_X1 U4860 ( .B1(n4415), .B2(n4394), .A(n4220), .ZN(U3262) );
  XNOR2_X1 U4861 ( .A(n4221), .B(n4222), .ZN(n4424) );
  INV_X1 U4862 ( .A(n4424), .ZN(n4237) );
  NAND2_X1 U4863 ( .A1(n4223), .A2(n4222), .ZN(n4224) );
  AOI21_X1 U4864 ( .B1(n4225), .B2(n4224), .A(n4384), .ZN(n4423) );
  NOR2_X1 U4865 ( .A1(n4252), .A2(n4231), .ZN(n4226) );
  OAI22_X1 U4866 ( .A1(n4228), .A2(n4634), .B1(n3991), .B2(n4566), .ZN(n4229)
         );
  AOI21_X1 U4867 ( .B1(n4247), .B2(n4419), .A(n4229), .ZN(n4230) );
  OAI21_X1 U4868 ( .B1(n4231), .B2(n4251), .A(n4230), .ZN(n4232) );
  AOI21_X1 U4869 ( .B1(n4337), .B2(n4233), .A(n4232), .ZN(n4234) );
  OAI21_X1 U4870 ( .B1(n4515), .B2(n4389), .A(n4234), .ZN(n4235) );
  AOI21_X1 U4871 ( .B1(n4423), .B2(n4566), .A(n4235), .ZN(n4236) );
  OAI21_X1 U4872 ( .B1(n4237), .B2(n4394), .A(n4236), .ZN(U3263) );
  INV_X1 U4873 ( .A(n4238), .ZN(n4239) );
  AOI21_X1 U4874 ( .B1(n4260), .B2(n4240), .A(n4239), .ZN(n4241) );
  XNOR2_X1 U4875 ( .A(n4241), .B(n4243), .ZN(n4242) );
  NAND2_X1 U4876 ( .A1(n4242), .A2(n4329), .ZN(n4429) );
  XNOR2_X1 U4877 ( .A(n4244), .B(n4243), .ZN(n4432) );
  NAND2_X1 U4878 ( .A1(n4432), .A2(n4333), .ZN(n4257) );
  INV_X1 U4879 ( .A(n4245), .ZN(n4246) );
  AOI22_X1 U4880 ( .A1(n4246), .A2(n4659), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4664), .ZN(n4249) );
  NAND2_X1 U4881 ( .A1(n4427), .A2(n4247), .ZN(n4248) );
  OAI211_X1 U4882 ( .C1(n4251), .C2(n4250), .A(n4249), .B(n4248), .ZN(n4255)
         );
  AND2_X1 U4883 ( .A1(n2053), .A2(n4426), .ZN(n4253) );
  OR2_X1 U4884 ( .A1(n4253), .A2(n4252), .ZN(n4519) );
  NOR2_X1 U4885 ( .A1(n4519), .A2(n4389), .ZN(n4254) );
  AOI211_X1 U4886 ( .C1(n4337), .C2(n4412), .A(n4255), .B(n4254), .ZN(n4256)
         );
  OAI211_X1 U4887 ( .C1(n4664), .C2(n4429), .A(n4257), .B(n4256), .ZN(U3264)
         );
  XNOR2_X1 U4888 ( .A(n4258), .B(n4262), .ZN(n4436) );
  INV_X1 U4889 ( .A(n4436), .ZN(n4274) );
  NAND2_X1 U4890 ( .A1(n4260), .A2(n4259), .ZN(n4261) );
  XOR2_X1 U4891 ( .A(n4262), .B(n4261), .Z(n4266) );
  OAI22_X1 U4892 ( .A1(n4263), .A2(n4492), .B1(n4267), .B2(n4409), .ZN(n4264)
         );
  AOI21_X1 U4893 ( .B1(n4419), .B2(n4489), .A(n4264), .ZN(n4265) );
  OAI21_X1 U4894 ( .B1(n4266), .B2(n4384), .A(n4265), .ZN(n4435) );
  INV_X1 U4895 ( .A(n4279), .ZN(n4268) );
  OAI21_X1 U4896 ( .B1(n4268), .B2(n4267), .A(n2053), .ZN(n4523) );
  NOR2_X1 U4897 ( .A1(n4523), .A2(n4389), .ZN(n4272) );
  INV_X1 U4898 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4269) );
  OAI22_X1 U4899 ( .A1(n4270), .A2(n4634), .B1(n4269), .B2(n4566), .ZN(n4271)
         );
  AOI211_X1 U4900 ( .C1(n4435), .C2(n4566), .A(n4272), .B(n4271), .ZN(n4273)
         );
  OAI21_X1 U4901 ( .B1(n4274), .B2(n4394), .A(n4273), .ZN(U3265) );
  XNOR2_X1 U4902 ( .A(n4275), .B(n4278), .ZN(n4276) );
  NAND2_X1 U4903 ( .A1(n4276), .A2(n4329), .ZN(n4443) );
  XOR2_X1 U4904 ( .A(n4278), .B(n4277), .Z(n4447) );
  NAND2_X1 U4905 ( .A1(n4447), .A2(n4333), .ZN(n4289) );
  INV_X1 U4906 ( .A(n4303), .ZN(n4281) );
  OAI21_X1 U4907 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(n4527) );
  INV_X1 U4908 ( .A(n4527), .ZN(n4287) );
  AOI22_X1 U4909 ( .A1(n4427), .A2(n4337), .B1(n4338), .B2(n4439), .ZN(n4284)
         );
  AOI22_X1 U4910 ( .A1(n4282), .A2(n4659), .B1(n4664), .B2(
        REG2_REG_24__SCAN_IN), .ZN(n4283) );
  OAI211_X1 U4911 ( .C1(n4285), .C2(n4342), .A(n4284), .B(n4283), .ZN(n4286)
         );
  AOI21_X1 U4912 ( .B1(n4287), .B2(n4651), .A(n4286), .ZN(n4288) );
  OAI211_X1 U4913 ( .C1(n4664), .C2(n4443), .A(n4289), .B(n4288), .ZN(U3266)
         );
  XNOR2_X1 U4914 ( .A(n4290), .B(n4296), .ZN(n4451) );
  INV_X1 U4915 ( .A(n4451), .ZN(n4310) );
  OR2_X1 U4916 ( .A1(n4328), .A2(n4291), .ZN(n4293) );
  NAND2_X1 U4917 ( .A1(n4293), .A2(n4292), .ZN(n4311) );
  INV_X1 U4918 ( .A(n4294), .ZN(n4295) );
  AOI21_X1 U4919 ( .B1(n4311), .B2(n4316), .A(n4295), .ZN(n4297) );
  XNOR2_X1 U4920 ( .A(n4297), .B(n4296), .ZN(n4302) );
  OAI22_X1 U4921 ( .A1(n4298), .A2(n4492), .B1(n4409), .B2(n4304), .ZN(n4299)
         );
  AOI21_X1 U4922 ( .B1(n4489), .B2(n4300), .A(n4299), .ZN(n4301) );
  OAI21_X1 U4923 ( .B1(n4302), .B2(n4384), .A(n4301), .ZN(n4450) );
  OAI21_X1 U4924 ( .B1(n4320), .B2(n4304), .A(n4303), .ZN(n4531) );
  NOR2_X1 U4925 ( .A1(n4531), .A2(n4389), .ZN(n4308) );
  OAI22_X1 U4926 ( .A1(n4566), .A2(n4306), .B1(n4305), .B2(n4634), .ZN(n4307)
         );
  AOI211_X1 U4927 ( .C1(n4450), .C2(n4566), .A(n4308), .B(n4307), .ZN(n4309)
         );
  OAI21_X1 U4928 ( .B1(n4310), .B2(n4394), .A(n4309), .ZN(U3267) );
  XNOR2_X1 U4929 ( .A(n4311), .B(n4316), .ZN(n4315) );
  NAND2_X1 U4930 ( .A1(n4441), .A2(n4489), .ZN(n4313) );
  NAND2_X1 U4931 ( .A1(n4361), .A2(n4440), .ZN(n4312) );
  OAI211_X1 U4932 ( .C1(n4409), .C2(n4318), .A(n4313), .B(n4312), .ZN(n4314)
         );
  AOI21_X1 U4933 ( .B1(n4315), .B2(n4329), .A(n4314), .ZN(n4455) );
  NAND2_X1 U4934 ( .A1(n4317), .A2(n4316), .ZN(n4454) );
  NAND3_X1 U4935 ( .A1(n2247), .A2(n4454), .A3(n4333), .ZN(n4326) );
  NOR2_X1 U4936 ( .A1(n4334), .A2(n4318), .ZN(n4319) );
  OR2_X1 U4937 ( .A1(n4320), .A2(n4319), .ZN(n4535) );
  INV_X1 U4938 ( .A(n4535), .ZN(n4324) );
  INV_X1 U4939 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4322) );
  OAI22_X1 U4940 ( .A1(n4566), .A2(n4322), .B1(n4321), .B2(n4634), .ZN(n4323)
         );
  AOI21_X1 U4941 ( .B1(n4324), .B2(n4651), .A(n4323), .ZN(n4325) );
  OAI211_X1 U4942 ( .C1(n4664), .C2(n4455), .A(n4326), .B(n4325), .ZN(U3268)
         );
  INV_X1 U4943 ( .A(n4331), .ZN(n4327) );
  XNOR2_X1 U4944 ( .A(n4328), .B(n4327), .ZN(n4330) );
  NAND2_X1 U4945 ( .A1(n4330), .A2(n4329), .ZN(n4462) );
  XNOR2_X1 U4946 ( .A(n4332), .B(n4331), .ZN(n4465) );
  NAND2_X1 U4947 ( .A1(n4465), .A2(n4333), .ZN(n4346) );
  INV_X1 U4948 ( .A(n4334), .ZN(n4335) );
  OAI21_X1 U4949 ( .B1(n2151), .B2(n4336), .A(n4335), .ZN(n4539) );
  INV_X1 U4950 ( .A(n4539), .ZN(n4344) );
  AOI22_X1 U4951 ( .A1(n4338), .A2(n4459), .B1(n4337), .B2(n4460), .ZN(n4341)
         );
  AOI22_X1 U4952 ( .A1(n4664), .A2(REG2_REG_21__SCAN_IN), .B1(n4339), .B2(
        n4659), .ZN(n4340) );
  OAI211_X1 U4953 ( .C1(n4463), .C2(n4342), .A(n4341), .B(n4340), .ZN(n4343)
         );
  AOI21_X1 U4954 ( .B1(n4344), .B2(n4651), .A(n4343), .ZN(n4345) );
  OAI211_X1 U4955 ( .C1(n4664), .C2(n4462), .A(n4346), .B(n4345), .ZN(U3269)
         );
  OR2_X1 U4956 ( .A1(n3606), .A2(n4347), .ZN(n4349) );
  NAND2_X1 U4957 ( .A1(n4349), .A2(n4348), .ZN(n4350) );
  XNOR2_X1 U4958 ( .A(n4350), .B(n4357), .ZN(n4364) );
  OAI22_X1 U4959 ( .A1(n4351), .A2(n4492), .B1(n4366), .B2(n4409), .ZN(n4360)
         );
  INV_X1 U4960 ( .A(n4352), .ZN(n4354) );
  OAI21_X1 U4961 ( .B1(n4355), .B2(n4354), .A(n4353), .ZN(n4356) );
  XOR2_X1 U4962 ( .A(n4357), .B(n4356), .Z(n4358) );
  NOR2_X1 U4963 ( .A1(n4358), .A2(n4384), .ZN(n4359) );
  AOI211_X1 U4964 ( .C1(n4489), .C2(n4361), .A(n4360), .B(n4359), .ZN(n4362)
         );
  OAI21_X1 U4965 ( .B1(n4364), .B2(n4363), .A(n4362), .ZN(n4468) );
  INV_X1 U4966 ( .A(n4468), .ZN(n4372) );
  INV_X1 U4967 ( .A(n4364), .ZN(n4469) );
  OAI21_X1 U4968 ( .B1(n2147), .B2(n4366), .A(n4365), .ZN(n4543) );
  INV_X1 U4969 ( .A(n4367), .ZN(n4368) );
  AOI22_X1 U4970 ( .A1(n4664), .A2(REG2_REG_20__SCAN_IN), .B1(n4368), .B2(
        n4659), .ZN(n4369) );
  OAI21_X1 U4971 ( .B1(n4543), .B2(n4389), .A(n4369), .ZN(n4370) );
  AOI21_X1 U4972 ( .B1(n4469), .B2(n4661), .A(n4370), .ZN(n4371) );
  OAI21_X1 U4973 ( .B1(n4372), .B2(n4664), .A(n4371), .ZN(U3270) );
  NAND2_X1 U4974 ( .A1(n4374), .A2(n4373), .ZN(n4375) );
  XOR2_X1 U4975 ( .A(n4380), .B(n4375), .Z(n4473) );
  INV_X1 U4976 ( .A(n4473), .ZN(n4395) );
  INV_X1 U4977 ( .A(n4376), .ZN(n4378) );
  OAI21_X1 U4978 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(n4381) );
  XNOR2_X1 U4979 ( .A(n4381), .B(n4380), .ZN(n4385) );
  OAI22_X1 U4980 ( .A1(n4463), .A2(n4444), .B1(n4409), .B2(n4387), .ZN(n4382)
         );
  AOI21_X1 U4981 ( .B1(n4440), .B2(n4479), .A(n4382), .ZN(n4383) );
  OAI21_X1 U4982 ( .B1(n4385), .B2(n4384), .A(n4383), .ZN(n4472) );
  OAI21_X1 U4983 ( .B1(n4388), .B2(n4387), .A(n4386), .ZN(n4547) );
  NOR2_X1 U4984 ( .A1(n4547), .A2(n4389), .ZN(n4392) );
  OAI22_X1 U4985 ( .A1(n4566), .A2(n4191), .B1(n4390), .B2(n4634), .ZN(n4391)
         );
  AOI211_X1 U4986 ( .C1(n4472), .C2(n4566), .A(n4392), .B(n4391), .ZN(n4393)
         );
  OAI21_X1 U4987 ( .B1(n4395), .B2(n4394), .A(n4393), .ZN(U3271) );
  NAND2_X1 U4988 ( .A1(n4502), .A2(n4713), .ZN(n4397) );
  NAND2_X1 U4989 ( .A1(n4711), .A2(REG1_REG_31__SCAN_IN), .ZN(n4396) );
  OAI211_X1 U4990 ( .C1(n4504), .C2(n4486), .A(n4397), .B(n4396), .ZN(U3549)
         );
  AOI21_X1 U4991 ( .B1(n4400), .B2(n4399), .A(n4398), .ZN(n4567) );
  NAND2_X1 U4992 ( .A1(n4567), .A2(n4401), .ZN(n4405) );
  OAI21_X1 U4993 ( .B1(n4403), .B2(n4409), .A(n4402), .ZN(n4565) );
  NAND2_X1 U4994 ( .A1(n4565), .A2(n4713), .ZN(n4404) );
  OAI211_X1 U4995 ( .C1(n4713), .C2(n4406), .A(n4405), .B(n4404), .ZN(U3548)
         );
  INV_X1 U4996 ( .A(n4407), .ZN(n4410) );
  OAI22_X1 U4997 ( .A1(n4410), .A2(n4444), .B1(n4409), .B2(n4408), .ZN(n4411)
         );
  AOI21_X1 U4998 ( .B1(n4440), .B2(n4412), .A(n4411), .ZN(n4414) );
  OAI211_X1 U4999 ( .C1(n4415), .C2(n4498), .A(n4414), .B(n4413), .ZN(n4508)
         );
  MUX2_X1 U5000 ( .A(REG1_REG_28__SCAN_IN), .B(n4508), .S(n4713), .Z(n4416) );
  INV_X1 U5001 ( .A(n4416), .ZN(n4417) );
  OAI21_X1 U5002 ( .B1(n4486), .B2(n4511), .A(n4417), .ZN(U3546) );
  AOI22_X1 U5003 ( .A1(n4419), .A2(n4440), .B1(n4418), .B2(n4488), .ZN(n4420)
         );
  OAI21_X1 U5004 ( .B1(n4421), .B2(n4444), .A(n4420), .ZN(n4422) );
  AOI211_X1 U5005 ( .C1(n4424), .C2(n4700), .A(n4423), .B(n4422), .ZN(n4512)
         );
  MUX2_X1 U5006 ( .A(n3965), .B(n4512), .S(n4713), .Z(n4425) );
  OAI21_X1 U5007 ( .B1(n4486), .B2(n4515), .A(n4425), .ZN(U3545) );
  INV_X1 U5008 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4433) );
  AOI22_X1 U5009 ( .A1(n4427), .A2(n4440), .B1(n4426), .B2(n4488), .ZN(n4428)
         );
  OAI211_X1 U5010 ( .C1(n4430), .C2(n4444), .A(n4429), .B(n4428), .ZN(n4431)
         );
  AOI21_X1 U5011 ( .B1(n4432), .B2(n4700), .A(n4431), .ZN(n4516) );
  MUX2_X1 U5012 ( .A(n4433), .B(n4516), .S(n4713), .Z(n4434) );
  OAI21_X1 U5013 ( .B1(n4486), .B2(n4519), .A(n4434), .ZN(U3544) );
  INV_X1 U5014 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4437) );
  AOI21_X1 U5015 ( .B1(n4436), .B2(n4700), .A(n4435), .ZN(n4520) );
  MUX2_X1 U5016 ( .A(n4437), .B(n4520), .S(n4713), .Z(n4438) );
  OAI21_X1 U5017 ( .B1(n4486), .B2(n4523), .A(n4438), .ZN(U3543) );
  INV_X1 U5018 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U5019 ( .A1(n4441), .A2(n4440), .B1(n4488), .B2(n4439), .ZN(n4442)
         );
  OAI211_X1 U5020 ( .C1(n4445), .C2(n4444), .A(n4443), .B(n4442), .ZN(n4446)
         );
  AOI21_X1 U5021 ( .B1(n4447), .B2(n4700), .A(n4446), .ZN(n4524) );
  MUX2_X1 U5022 ( .A(n4448), .B(n4524), .S(n4713), .Z(n4449) );
  OAI21_X1 U5023 ( .B1(n4486), .B2(n4527), .A(n4449), .ZN(U3542) );
  INV_X1 U5024 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4452) );
  AOI21_X1 U5025 ( .B1(n4451), .B2(n4700), .A(n4450), .ZN(n4528) );
  MUX2_X1 U5026 ( .A(n4452), .B(n4528), .S(n4713), .Z(n4453) );
  OAI21_X1 U5027 ( .B1(n4486), .B2(n4531), .A(n4453), .ZN(U3541) );
  NAND3_X1 U5028 ( .A1(n2247), .A2(n4454), .A3(n4700), .ZN(n4456) );
  NAND2_X1 U5029 ( .A1(n4456), .A2(n4455), .ZN(n4532) );
  MUX2_X1 U5030 ( .A(REG1_REG_22__SCAN_IN), .B(n4532), .S(n4713), .Z(n4457) );
  INV_X1 U5031 ( .A(n4457), .ZN(n4458) );
  OAI21_X1 U5032 ( .B1(n4486), .B2(n4535), .A(n4458), .ZN(U3540) );
  INV_X1 U5033 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4466) );
  AOI22_X1 U5034 ( .A1(n4460), .A2(n4489), .B1(n4488), .B2(n4459), .ZN(n4461)
         );
  OAI211_X1 U5035 ( .C1(n4463), .C2(n4492), .A(n4462), .B(n4461), .ZN(n4464)
         );
  AOI21_X1 U5036 ( .B1(n4465), .B2(n4700), .A(n4464), .ZN(n4536) );
  MUX2_X1 U5037 ( .A(n4466), .B(n4536), .S(n4713), .Z(n4467) );
  OAI21_X1 U5038 ( .B1(n4486), .B2(n4539), .A(n4467), .ZN(U3539) );
  INV_X1 U5039 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4470) );
  AOI21_X1 U5040 ( .B1(n4698), .B2(n4469), .A(n4468), .ZN(n4540) );
  MUX2_X1 U5041 ( .A(n4470), .B(n4540), .S(n4713), .Z(n4471) );
  OAI21_X1 U5042 ( .B1(n4486), .B2(n4543), .A(n4471), .ZN(U3538) );
  AOI21_X1 U5043 ( .B1(n4473), .B2(n4700), .A(n4472), .ZN(n4544) );
  MUX2_X1 U5044 ( .A(n4185), .B(n4544), .S(n4713), .Z(n4474) );
  OAI21_X1 U5045 ( .B1(n4486), .B2(n4547), .A(n4474), .ZN(U3537) );
  OAI211_X1 U5046 ( .C1(n4477), .C2(n4498), .A(n4476), .B(n4475), .ZN(n4548)
         );
  MUX2_X1 U5047 ( .A(REG1_REG_18__SCAN_IN), .B(n4548), .S(n4713), .Z(U3536) );
  AOI22_X1 U5048 ( .A1(n4479), .A2(n4489), .B1(n4478), .B2(n4488), .ZN(n4480)
         );
  OAI211_X1 U5049 ( .C1(n4482), .C2(n4492), .A(n4481), .B(n4480), .ZN(n4483)
         );
  AOI21_X1 U5050 ( .B1(n4484), .B2(n4700), .A(n4483), .ZN(n4549) );
  MUX2_X1 U5051 ( .A(n4162), .B(n4549), .S(n4713), .Z(n4485) );
  OAI21_X1 U5052 ( .B1(n4486), .B2(n4553), .A(n4485), .ZN(U3535) );
  AOI22_X1 U5053 ( .A1(n4490), .A2(n4489), .B1(n4488), .B2(n4487), .ZN(n4491)
         );
  OAI21_X1 U5054 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(n4494) );
  AOI21_X1 U5055 ( .B1(n4495), .B2(n4693), .A(n4494), .ZN(n4497) );
  OAI211_X1 U5056 ( .C1(n4499), .C2(n4498), .A(n4497), .B(n4496), .ZN(n4554)
         );
  MUX2_X1 U5057 ( .A(REG1_REG_16__SCAN_IN), .B(n4554), .S(n4713), .Z(U3534) );
  NOR2_X1 U5058 ( .A1(n4706), .A2(n4500), .ZN(n4501) );
  AOI21_X1 U5059 ( .B1(n4502), .B2(n4706), .A(n4501), .ZN(n4503) );
  OAI21_X1 U5060 ( .B1(n4504), .B2(n4552), .A(n4503), .ZN(U3517) );
  NAND2_X1 U5061 ( .A1(n4567), .A2(n4505), .ZN(n4507) );
  NAND2_X1 U5062 ( .A1(n4565), .A2(n4706), .ZN(n4506) );
  OAI211_X1 U5063 ( .C1(n4706), .C2(n2633), .A(n4507), .B(n4506), .ZN(U3516)
         );
  MUX2_X1 U5064 ( .A(REG0_REG_28__SCAN_IN), .B(n4508), .S(n4706), .Z(n4509) );
  INV_X1 U5065 ( .A(n4509), .ZN(n4510) );
  OAI21_X1 U5066 ( .B1(n4511), .B2(n4552), .A(n4510), .ZN(U3514) );
  MUX2_X1 U5067 ( .A(n4513), .B(n4512), .S(n4706), .Z(n4514) );
  OAI21_X1 U5068 ( .B1(n4515), .B2(n4552), .A(n4514), .ZN(U3513) );
  MUX2_X1 U5069 ( .A(n4517), .B(n4516), .S(n4706), .Z(n4518) );
  OAI21_X1 U5070 ( .B1(n4519), .B2(n4552), .A(n4518), .ZN(U3512) );
  MUX2_X1 U5071 ( .A(n4521), .B(n4520), .S(n4706), .Z(n4522) );
  OAI21_X1 U5072 ( .B1(n4523), .B2(n4552), .A(n4522), .ZN(U3511) );
  MUX2_X1 U5073 ( .A(n4525), .B(n4524), .S(n4706), .Z(n4526) );
  OAI21_X1 U5074 ( .B1(n4527), .B2(n4552), .A(n4526), .ZN(U3510) );
  INV_X1 U5075 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4529) );
  MUX2_X1 U5076 ( .A(n4529), .B(n4528), .S(n4706), .Z(n4530) );
  OAI21_X1 U5077 ( .B1(n4531), .B2(n4552), .A(n4530), .ZN(U3509) );
  MUX2_X1 U5078 ( .A(REG0_REG_22__SCAN_IN), .B(n4532), .S(n4706), .Z(n4533) );
  INV_X1 U5079 ( .A(n4533), .ZN(n4534) );
  OAI21_X1 U5080 ( .B1(n4535), .B2(n4552), .A(n4534), .ZN(U3508) );
  MUX2_X1 U5081 ( .A(n4537), .B(n4536), .S(n4706), .Z(n4538) );
  OAI21_X1 U5082 ( .B1(n4539), .B2(n4552), .A(n4538), .ZN(U3507) );
  MUX2_X1 U5083 ( .A(n4541), .B(n4540), .S(n4706), .Z(n4542) );
  OAI21_X1 U5084 ( .B1(n4543), .B2(n4552), .A(n4542), .ZN(U3506) );
  MUX2_X1 U5085 ( .A(n4545), .B(n4544), .S(n4706), .Z(n4546) );
  OAI21_X1 U5086 ( .B1(n4547), .B2(n4552), .A(n4546), .ZN(U3505) );
  MUX2_X1 U5087 ( .A(REG0_REG_18__SCAN_IN), .B(n4548), .S(n4706), .Z(U3503) );
  MUX2_X1 U5088 ( .A(n4550), .B(n4549), .S(n4706), .Z(n4551) );
  OAI21_X1 U5089 ( .B1(n4553), .B2(n4552), .A(n4551), .ZN(U3501) );
  MUX2_X1 U5090 ( .A(REG0_REG_16__SCAN_IN), .B(n4554), .S(n4706), .Z(U3499) );
  MUX2_X1 U5091 ( .A(DATAI_27_), .B(n4555), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5092 ( .A(DATAI_24_), .B(n4556), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5093 ( .A(n4557), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5094 ( .A(n4558), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5095 ( .A(DATAI_8_), .B(n4559), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5096 ( .A(n4560), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5097 ( .A(DATAI_4_), .B(n4561), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5098 ( .A(n4562), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5099 ( .A(n4563), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U5100 ( .A1(STATE_REG_SCAN_IN), .A2(n4564), .B1(n2576), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U5101 ( .A1(n4567), .A2(n4651), .B1(n4566), .B2(n4565), .ZN(n4568)
         );
  OAI21_X1 U5102 ( .B1(n4569), .B2(n4566), .A(n4568), .ZN(U3261) );
  OAI211_X1 U5103 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4572), .A(n4593), .B(n4571), .ZN(n4574) );
  NAND2_X1 U5104 ( .A1(n4574), .A2(n4573), .ZN(n4575) );
  AOI21_X1 U5105 ( .B1(n4626), .B2(ADDR_REG_10__SCAN_IN), .A(n4575), .ZN(n4579) );
  OAI211_X1 U5106 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4577), .A(n4627), .B(n4576), .ZN(n4578) );
  OAI211_X1 U5107 ( .C1(n4633), .C2(n2177), .A(n4579), .B(n4578), .ZN(U3250)
         );
  OAI211_X1 U5108 ( .C1(n4582), .C2(n4581), .A(n4627), .B(n4580), .ZN(n4587)
         );
  OAI211_X1 U5109 ( .C1(n4585), .C2(n4584), .A(n4593), .B(n4583), .ZN(n4586)
         );
  OAI211_X1 U5110 ( .C1(n4633), .C2(n4683), .A(n4587), .B(n4586), .ZN(n4588)
         );
  AOI211_X1 U5111 ( .C1(n4626), .C2(ADDR_REG_11__SCAN_IN), .A(n4589), .B(n4588), .ZN(n4590) );
  INV_X1 U5112 ( .A(n4590), .ZN(U3251) );
  OAI211_X1 U5113 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4594), .A(n4593), .B(n4592), .ZN(n4596) );
  NAND2_X1 U5114 ( .A1(n4596), .A2(n4595), .ZN(n4597) );
  AOI21_X1 U5115 ( .B1(n4626), .B2(ADDR_REG_12__SCAN_IN), .A(n4597), .ZN(n4601) );
  OAI211_X1 U5116 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4599), .A(n4627), .B(n4598), .ZN(n4600) );
  OAI211_X1 U5117 ( .C1(n4633), .C2(n2176), .A(n4601), .B(n4600), .ZN(U3252)
         );
  AOI211_X1 U5118 ( .C1(n4604), .C2(n4603), .A(n4602), .B(n4620), .ZN(n4605)
         );
  AOI211_X1 U5119 ( .C1(n4626), .C2(ADDR_REG_14__SCAN_IN), .A(n4606), .B(n4605), .ZN(n4610) );
  OAI211_X1 U5120 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4608), .A(n4627), .B(n4607), .ZN(n4609) );
  OAI211_X1 U5121 ( .C1(n4633), .C2(n4681), .A(n4610), .B(n4609), .ZN(U3254)
         );
  AOI221_X1 U5122 ( .B1(n4613), .B2(n4612), .C1(n4611), .C2(n4612), .A(n4620), 
        .ZN(n4614) );
  AOI211_X1 U5123 ( .C1(n4626), .C2(ADDR_REG_16__SCAN_IN), .A(n4615), .B(n4614), .ZN(n4619) );
  OAI221_X1 U5124 ( .B1(n4617), .B2(REG1_REG_16__SCAN_IN), .C1(n4617), .C2(
        n4616), .A(n4627), .ZN(n4618) );
  OAI211_X1 U5125 ( .C1(n4633), .C2(n4679), .A(n4619), .B(n4618), .ZN(U3256)
         );
  AOI221_X1 U5126 ( .B1(n4623), .B2(n4622), .C1(n4621), .C2(n4622), .A(n4620), 
        .ZN(n4624) );
  AOI211_X1 U5127 ( .C1(n4626), .C2(ADDR_REG_17__SCAN_IN), .A(n4625), .B(n4624), .ZN(n4632) );
  OAI221_X1 U5128 ( .B1(n4630), .B2(n4629), .C1(n4630), .C2(n4628), .A(n4627), 
        .ZN(n4631) );
  OAI211_X1 U5129 ( .C1(n4633), .C2(n4677), .A(n4632), .B(n4631), .ZN(U3257)
         );
  OAI22_X1 U5130 ( .A1(n4566), .A2(n2096), .B1(n4635), .B2(n4634), .ZN(n4636)
         );
  INV_X1 U5131 ( .A(n4636), .ZN(n4642) );
  INV_X1 U5132 ( .A(n4637), .ZN(n4640) );
  INV_X1 U5133 ( .A(n4638), .ZN(n4639) );
  AOI22_X1 U5134 ( .A1(n4640), .A2(n4661), .B1(n4651), .B2(n4639), .ZN(n4641)
         );
  OAI211_X1 U5135 ( .C1(n4664), .C2(n4643), .A(n4642), .B(n4641), .ZN(U3282)
         );
  AOI22_X1 U5136 ( .A1(n4664), .A2(REG2_REG_3__SCAN_IN), .B1(n4659), .B2(n4644), .ZN(n4648) );
  AOI22_X1 U5137 ( .A1(n4646), .A2(n4661), .B1(n4651), .B2(n4645), .ZN(n4647)
         );
  OAI211_X1 U5138 ( .C1(n4664), .C2(n4649), .A(n4648), .B(n4647), .ZN(U3287)
         );
  AOI22_X1 U5139 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4659), .B1(
        REG2_REG_2__SCAN_IN), .B2(n4664), .ZN(n4654) );
  AOI22_X1 U5140 ( .A1(n4652), .A2(n4661), .B1(n4651), .B2(n4650), .ZN(n4653)
         );
  OAI211_X1 U5141 ( .C1(n4664), .C2(n4655), .A(n4654), .B(n4653), .ZN(U3288)
         );
  AOI21_X1 U5142 ( .B1(n4658), .B2(n4657), .A(n4656), .ZN(n4663) );
  AOI22_X1 U5143 ( .A1(n4661), .A2(n4660), .B1(REG3_REG_0__SCAN_IN), .B2(n4659), .ZN(n4662) );
  OAI221_X1 U5144 ( .B1(n4664), .B2(n4663), .C1(n4566), .C2(n4107), .A(n4662), 
        .ZN(U3290) );
  AND2_X1 U5145 ( .A1(D_REG_31__SCAN_IN), .A2(n4674), .ZN(U3291) );
  NOR2_X1 U5146 ( .A1(n4673), .A2(n4665), .ZN(U3292) );
  AND2_X1 U5147 ( .A1(D_REG_29__SCAN_IN), .A2(n4674), .ZN(U3293) );
  NOR2_X1 U5148 ( .A1(n4673), .A2(n4666), .ZN(U3294) );
  AND2_X1 U5149 ( .A1(D_REG_27__SCAN_IN), .A2(n4674), .ZN(U3295) );
  AND2_X1 U5150 ( .A1(D_REG_26__SCAN_IN), .A2(n4674), .ZN(U3296) );
  NOR2_X1 U5151 ( .A1(n4673), .A2(n4667), .ZN(U3297) );
  AND2_X1 U5152 ( .A1(D_REG_24__SCAN_IN), .A2(n4674), .ZN(U3298) );
  NOR2_X1 U5153 ( .A1(n4673), .A2(n4668), .ZN(U3299) );
  NOR2_X1 U5154 ( .A1(n4673), .A2(n4669), .ZN(U3300) );
  NOR2_X1 U5155 ( .A1(n4673), .A2(n4670), .ZN(U3301) );
  AND2_X1 U5156 ( .A1(D_REG_20__SCAN_IN), .A2(n4674), .ZN(U3302) );
  AND2_X1 U5157 ( .A1(D_REG_19__SCAN_IN), .A2(n4674), .ZN(U3303) );
  AND2_X1 U5158 ( .A1(D_REG_18__SCAN_IN), .A2(n4674), .ZN(U3304) );
  AND2_X1 U5159 ( .A1(D_REG_17__SCAN_IN), .A2(n4674), .ZN(U3305) );
  AND2_X1 U5160 ( .A1(D_REG_16__SCAN_IN), .A2(n4674), .ZN(U3306) );
  AND2_X1 U5161 ( .A1(D_REG_15__SCAN_IN), .A2(n4674), .ZN(U3307) );
  AND2_X1 U5162 ( .A1(D_REG_14__SCAN_IN), .A2(n4674), .ZN(U3308) );
  AND2_X1 U5163 ( .A1(D_REG_13__SCAN_IN), .A2(n4674), .ZN(U3309) );
  AND2_X1 U5164 ( .A1(D_REG_12__SCAN_IN), .A2(n4674), .ZN(U3310) );
  NOR2_X1 U5165 ( .A1(n4673), .A2(n4671), .ZN(U3311) );
  AND2_X1 U5166 ( .A1(D_REG_10__SCAN_IN), .A2(n4674), .ZN(U3312) );
  AND2_X1 U5167 ( .A1(D_REG_9__SCAN_IN), .A2(n4674), .ZN(U3313) );
  AND2_X1 U5168 ( .A1(D_REG_8__SCAN_IN), .A2(n4674), .ZN(U3314) );
  NOR2_X1 U5169 ( .A1(n4673), .A2(n4672), .ZN(U3315) );
  AND2_X1 U5170 ( .A1(D_REG_6__SCAN_IN), .A2(n4674), .ZN(U3316) );
  AND2_X1 U5171 ( .A1(D_REG_5__SCAN_IN), .A2(n4674), .ZN(U3317) );
  AND2_X1 U5172 ( .A1(D_REG_4__SCAN_IN), .A2(n4674), .ZN(U3318) );
  AND2_X1 U5173 ( .A1(D_REG_3__SCAN_IN), .A2(n4674), .ZN(U3319) );
  AND2_X1 U5174 ( .A1(D_REG_2__SCAN_IN), .A2(n4674), .ZN(U3320) );
  INV_X1 U5175 ( .A(DATAI_23_), .ZN(n4676) );
  AOI21_X1 U5176 ( .B1(U3149), .B2(n4676), .A(n4675), .ZN(U3329) );
  AOI22_X1 U5177 ( .A1(STATE_REG_SCAN_IN), .A2(n4677), .B1(n2484), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5178 ( .A1(STATE_REG_SCAN_IN), .A2(n4679), .B1(n4678), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5179 ( .A1(STATE_REG_SCAN_IN), .A2(n4681), .B1(n4680), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5180 ( .A(DATAI_12_), .ZN(n4682) );
  AOI22_X1 U5181 ( .A1(STATE_REG_SCAN_IN), .A2(n2176), .B1(n4682), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5182 ( .A1(STATE_REG_SCAN_IN), .A2(n4683), .B1(n2416), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5183 ( .A(DATAI_10_), .ZN(n4684) );
  AOI22_X1 U5184 ( .A1(STATE_REG_SCAN_IN), .A2(n2177), .B1(n4684), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5185 ( .A(DATAI_0_), .ZN(n4685) );
  AOI22_X1 U5186 ( .A1(STATE_REG_SCAN_IN), .A2(n4686), .B1(n4685), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5187 ( .A1(n4706), .A2(n4687), .B1(n2293), .B2(n2136), .ZN(U3467)
         );
  NOR2_X1 U5188 ( .A1(n4689), .A2(n4688), .ZN(n4691) );
  AOI211_X1 U5189 ( .C1(n4693), .C2(n4692), .A(n4691), .B(n4690), .ZN(n4708)
         );
  AOI22_X1 U5190 ( .A1(n4706), .A2(n4708), .B1(n2286), .B2(n2136), .ZN(U3469)
         );
  INV_X1 U5191 ( .A(n4694), .ZN(n4699) );
  INV_X1 U5192 ( .A(n4695), .ZN(n4697) );
  AOI211_X1 U5193 ( .C1(n4699), .C2(n4698), .A(n4697), .B(n4696), .ZN(n4710)
         );
  AOI22_X1 U5194 ( .A1(n4706), .A2(n4710), .B1(n2321), .B2(n2136), .ZN(U3475)
         );
  NAND3_X1 U5195 ( .A1(n4702), .A2(n4701), .A3(n4700), .ZN(n4703) );
  AOI22_X1 U5196 ( .A1(n4706), .A2(n4712), .B1(n2360), .B2(n2136), .ZN(U3481)
         );
  INV_X1 U5197 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5198 ( .A1(n4713), .A2(n4708), .B1(n4707), .B2(n4711), .ZN(U3519)
         );
  AOI22_X1 U5199 ( .A1(n4713), .A2(n4710), .B1(n4709), .B2(n4711), .ZN(U3522)
         );
  AOI22_X1 U5200 ( .A1(n4713), .A2(n4712), .B1(n3016), .B2(n4711), .ZN(U3525)
         );
  CLKBUF_X3 U2276 ( .A(n2697), .Z(n2033) );
endmodule

