

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1,
         READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n11121, n11122, n11123, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11152, n11153, n11154, n11155,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313, n22314, n22315, n22316, n22317, n22318,
         n22319, n22320, n22321, n22322, n22323, n22324, n22325, n22326,
         n22327, n22328, n22329, n22330, n22331, n22332, n22333, n22334,
         n22335, n22336, n22337, n22338, n22339, n22340, n22341, n22342,
         n22343, n22344, n22345, n22346, n22347, n22348, n22349, n22350,
         n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
         n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366,
         n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374,
         n22375, n22376, n22377, n22378, n22379, n22380, n22381, n22382,
         n22383, n22384, n22385, n22386, n22387, n22388, n22389, n22390,
         n22391, n22392, n22393, n22394, n22395, n22396, n22397, n22398,
         n22399, n22400, n22401, n22402, n22403, n22404, n22405, n22406,
         n22407, n22408, n22409, n22410, n22411, n22412, n22413, n22414,
         n22415, n22416, n22417, n22418, n22419, n22420, n22421, n22422,
         n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
         n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438,
         n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446,
         n22447, n22448, n22449, n22450, n22451, n22452, n22453, n22454,
         n22455, n22456, n22457, n22458, n22459, n22460, n22461, n22462,
         n22463, n22464, n22465, n22466, n22467, n22468, n22469, n22470,
         n22471, n22472, n22473, n22474, n22475, n22476, n22477, n22478,
         n22479, n22480, n22481, n22482, n22483, n22484, n22485, n22486,
         n22487, n22488, n22489, n22490, n22491, n22492, n22493, n22494,
         n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
         n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510,
         n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518,
         n22519, n22520, n22521, n22522, n22523, n22524, n22525, n22526,
         n22527, n22528, n22529, n22530, n22531, n22532, n22533, n22534,
         n22535, n22536, n22537, n22538, n22539, n22540, n22541, n22542,
         n22543, n22544, n22545, n22546, n22547, n22548, n22549, n22550,
         n22551, n22552, n22553, n22554, n22555, n22556, n22557, n22558,
         n22559, n22560, n22561, n22562, n22563, n22564, n22565, n22566,
         n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
         n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582,
         n22583, n22584, n22585, n22586, n22587, n22588, n22589, n22590,
         n22591, n22592, n22593, n22594, n22595, n22596, n22597, n22598,
         n22599, n22600, n22601, n22602, n22603, n22604, n22605, n22606,
         n22607, n22608, n22609, n22610, n22611, n22612, n22613, n22614,
         n22615, n22616, n22617, n22618, n22619, n22620, n22621, n22622,
         n22623, n22624, n22625, n22626, n22627, n22628, n22629, n22630,
         n22631, n22632, n22633, n22634, n22635, n22636, n22637, n22638,
         n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
         n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654,
         n22655, n22656, n22657, n22658, n22659, n22660, n22661, n22662,
         n22663, n22664, n22665, n22666, n22667, n22668, n22669, n22670,
         n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
         n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
         n22687, n22688, n22689, n22690, n22691, n22692, n22693, n22694,
         n22695, n22696, n22697, n22698, n22699, n22700, n22701, n22702,
         n22703, n22704, n22705, n22706, n22707, n22708, n22709, n22710,
         n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
         n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726,
         n22727, n22728, n22729, n22730, n22731, n22732, n22733, n22734,
         n22735, n22736, n22737, n22738, n22739, n22740, n22741, n22742,
         n22743, n22744, n22745, n22746, n22747, n22748, n22749, n22750,
         n22751, n22752, n22753, n22754, n22755, n22756, n22757, n22758,
         n22759, n22760, n22761, n22762, n22763, n22764, n22765, n22766,
         n22767, n22768, n22769, n22770, n22771, n22772, n22773, n22774,
         n22775, n22776, n22777, n22778, n22779, n22780, n22781, n22782,
         n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
         n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798,
         n22799, n22800, n22801, n22802, n22803, n22804, n22805, n22806,
         n22807, n22808, n22809, n22810, n22811, n22812, n22813, n22814,
         n22815, n22816, n22817, n22818, n22819, n22820, n22821, n22822,
         n22823, n22824, n22825, n22826, n22827, n22828, n22829, n22830,
         n22831, n22832, n22833, n22834, n22835, n22836, n22837, n22838,
         n22839, n22840, n22841, n22842, n22843, n22844, n22845, n22846,
         n22847, n22848, n22849, n22850, n22851, n22852, n22853, n22854;

  INV_X1 U11228 ( .A(n11144), .ZN(n18915) );
  AND2_X1 U11229 ( .A1(n16044), .A2(n11625), .ZN(n15992) );
  CLKBUF_X2 U11230 ( .A(n18903), .Z(n11144) );
  NAND2_X1 U11231 ( .A1(n16696), .A2(n11251), .ZN(n16671) );
  NOR2_X2 U11232 ( .A1(n11183), .A2(n16705), .ZN(n16696) );
  OR2_X1 U11233 ( .A1(n21487), .A2(n21882), .ZN(n11370) );
  INV_X1 U11234 ( .A(n21885), .ZN(n21783) );
  INV_X1 U11235 ( .A(n14712), .ZN(n15910) );
  NAND2_X1 U11236 ( .A1(n12213), .A2(n15425), .ZN(n15337) );
  NAND2_X1 U11237 ( .A1(n14567), .A2(n12574), .ZN(n14648) );
  INV_X2 U11238 ( .A(n15795), .ZN(n15794) );
  CLKBUF_X2 U11240 ( .A(n13093), .Z(n13758) );
  CLKBUF_X2 U11241 ( .A(n11985), .Z(n15085) );
  BUF_X1 U11242 ( .A(n11981), .Z(n12977) );
  AND2_X1 U11243 ( .A1(n12820), .A2(n11742), .ZN(n11837) );
  CLKBUF_X2 U11244 ( .A(n11988), .Z(n12983) );
  BUF_X2 U11245 ( .A(n15715), .Z(n18379) );
  CLKBUF_X1 U11246 ( .A(n11986), .Z(n12978) );
  CLKBUF_X3 U11247 ( .A(n18153), .Z(n11128) );
  BUF_X1 U11248 ( .A(n18408), .Z(n11127) );
  CLKBUF_X2 U11249 ( .A(n15714), .Z(n11129) );
  INV_X1 U11250 ( .A(n14064), .ZN(n12393) );
  INV_X1 U11251 ( .A(n13275), .ZN(n14804) );
  AND2_X4 U11252 ( .A1(n11736), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11988) );
  AND2_X1 U11253 ( .A1(n14697), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14694) );
  CLKBUF_X1 U11254 ( .A(n19254), .Z(n11121) );
  NOR2_X1 U11255 ( .A1(n15399), .A2(n15398), .ZN(n19254) );
  NOR2_X1 U11256 ( .A1(n14840), .A2(n14825), .ZN(n11122) );
  INV_X1 U11257 ( .A(n13157), .ZN(n14825) );
  NOR2_X1 U11258 ( .A1(n14840), .A2(n14804), .ZN(n11123) );
  INV_X1 U11260 ( .A(n22854), .ZN(n11125) );
  NOR2_X1 U11261 ( .A1(n12106), .A2(n12105), .ZN(n12127) );
  AND2_X1 U11264 ( .A1(n15060), .A2(n12214), .ZN(n11134) );
  AND2_X1 U11265 ( .A1(n13037), .A2(n16572), .ZN(n13143) );
  INV_X1 U11266 ( .A(n13115), .ZN(n14537) );
  AND2_X1 U11267 ( .A1(n11745), .A2(n12820), .ZN(n12838) );
  AND2_X1 U11268 ( .A1(n12982), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12162) );
  NOR2_X1 U11269 ( .A1(n22045), .A2(n22005), .ZN(n22071) );
  NAND2_X1 U11271 ( .A1(n15604), .A2(n14470), .ZN(n15830) );
  OR2_X1 U11272 ( .A1(n16861), .A2(n11601), .ZN(n16840) );
  NAND2_X1 U11273 ( .A1(n11484), .A2(n11485), .ZN(n16899) );
  NOR2_X1 U11275 ( .A1(n20704), .A2(n18487), .ZN(n21667) );
  CLKBUF_X2 U11276 ( .A(n15714), .Z(n11130) );
  OAI21_X1 U11277 ( .B1(n20707), .B2(P3_STATE2_REG_0__SCAN_IN), .A(n21940), 
        .ZN(n18911) );
  NAND2_X1 U11278 ( .A1(n18756), .A2(n21816), .ZN(n18755) );
  INV_X2 U11279 ( .A(n21778), .ZN(n21861) );
  NOR2_X1 U11280 ( .A1(n15722), .A2(n15721), .ZN(n21434) );
  INV_X1 U11281 ( .A(n11190), .ZN(n18390) );
  NAND4_X2 U11282 ( .A1(n13155), .A2(n11193), .A3(n13154), .A4(n13153), .ZN(
        n15178) );
  INV_X2 U11284 ( .A(n12026), .ZN(n19017) );
  NOR3_X2 U11285 ( .A1(n17209), .A2(n17203), .A3(n17222), .ZN(n16924) );
  OAI211_X1 U11286 ( .C1(n15404), .C2(n15521), .A(n12234), .B(n12233), .ZN(
        n15506) );
  INV_X1 U11287 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19322) );
  NAND2_X1 U11288 ( .A1(n11370), .A2(n11368), .ZN(n21876) );
  NAND2_X1 U11289 ( .A1(n18759), .A2(n18758), .ZN(n18904) );
  NOR2_X1 U11290 ( .A1(n21487), .A2(n21450), .ZN(n21756) );
  NAND2_X1 U11291 ( .A1(n21876), .A2(n21932), .ZN(n21940) );
  AND2_X2 U11293 ( .A1(n12130), .A2(n11364), .ZN(n11363) );
  NAND2_X2 U11294 ( .A1(n20294), .A2(n12393), .ZN(n12997) );
  BUF_X1 U11295 ( .A(n12078), .Z(n12080) );
  BUF_X1 U11296 ( .A(n18408), .Z(n11126) );
  NOR2_X1 U11297 ( .A1(n21888), .A2(n21401), .ZN(n18408) );
  NAND2_X2 U11298 ( .A1(n16986), .A2(n11374), .ZN(n16861) );
  OR2_X2 U11299 ( .A1(n14213), .A2(n17853), .ZN(n11728) );
  NAND2_X4 U11300 ( .A1(n13987), .A2(n13986), .ZN(n13994) );
  OR2_X2 U11301 ( .A1(n12364), .A2(n14016), .ZN(n11696) );
  OR2_X2 U11302 ( .A1(n14213), .A2(n17351), .ZN(n11194) );
  NOR2_X4 U11303 ( .A1(n12211), .A2(n12207), .ZN(n12206) );
  NAND2_X2 U11304 ( .A1(n12220), .A2(n12212), .ZN(n12211) );
  AND2_X2 U11305 ( .A1(n11301), .A2(n21741), .ZN(n18529) );
  NOR2_X2 U11306 ( .A1(n18909), .A2(n21472), .ZN(n18908) );
  NAND2_X2 U11308 ( .A1(n11611), .A2(n13202), .ZN(n17398) );
  NAND2_X2 U11309 ( .A1(n12200), .A2(n11492), .ZN(n12426) );
  NAND2_X4 U11310 ( .A1(n13131), .A2(n11615), .ZN(n14886) );
  NAND2_X2 U11311 ( .A1(n11940), .A2(n11939), .ZN(n12005) );
  AOI211_X2 U11312 ( .C1(n20628), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n22059), .B(n20608), .ZN(n20609) );
  NAND2_X2 U11313 ( .A1(n12020), .A2(n12019), .ZN(n11689) );
  NAND2_X4 U11314 ( .A1(n11953), .A2(n11952), .ZN(n12006) );
  NOR3_X1 U11315 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21888), .A3(
        n15651), .ZN(n15714) );
  AND2_X4 U11316 ( .A1(n11308), .A2(n21398), .ZN(n18462) );
  AND2_X2 U11317 ( .A1(n21891), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n21398) );
  AND2_X4 U11318 ( .A1(n11525), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11980) );
  AND2_X4 U11319 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11525) );
  NOR3_X1 U11320 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21888), .A3(
        n15652), .ZN(n11131) );
  NOR3_X1 U11321 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21888), .A3(
        n15652), .ZN(n11132) );
  AND2_X1 U11322 ( .A1(n15060), .A2(n12214), .ZN(n11133) );
  BUF_X2 U11323 ( .A(n13102), .Z(n11136) );
  BUF_X4 U11324 ( .A(n13102), .Z(n11137) );
  INV_X1 U11325 ( .A(n13108), .ZN(n11138) );
  INV_X1 U11326 ( .A(n11138), .ZN(n11139) );
  INV_X1 U11327 ( .A(n11138), .ZN(n11140) );
  INV_X1 U11328 ( .A(n11138), .ZN(n11141) );
  INV_X1 U11329 ( .A(n11138), .ZN(n11142) );
  AND2_X1 U11330 ( .A1(n13045), .A2(n14641), .ZN(n13108) );
  NAND4_X4 U11331 ( .A1(n12033), .A2(n12032), .A3(n14174), .A4(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12527) );
  INV_X1 U11332 ( .A(n12030), .ZN(n12033) );
  NOR2_X4 U11333 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11745) );
  XNOR2_X2 U11334 ( .A(n12263), .B(n17342), .ZN(n17338) );
  NAND2_X2 U11335 ( .A1(n11686), .A2(n19045), .ZN(n12263) );
  XNOR2_X2 U11336 ( .A(n11274), .B(n12210), .ZN(n15262) );
  NAND2_X2 U11337 ( .A1(n11365), .A2(n12171), .ZN(n12210) );
  XNOR2_X2 U11338 ( .A(n16899), .B(n16898), .ZN(n16908) );
  NOR2_X1 U11339 ( .A1(n21435), .A2(n21940), .ZN(n18903) );
  OAI21_X2 U11340 ( .B1(n16860), .B2(n11708), .A(n11707), .ZN(n16834) );
  OAI21_X2 U11341 ( .B1(n16871), .B2(n16869), .A(n16867), .ZN(n16860) );
  CLKBUF_X1 U11342 ( .A(n15992), .Z(n15993) );
  NAND2_X1 U11343 ( .A1(n15617), .A2(n13527), .ZN(n15618) );
  NAND2_X1 U11344 ( .A1(n16659), .A2(n16658), .ZN(n16657) );
  OR2_X1 U11345 ( .A1(n15342), .A2(n11271), .ZN(n11270) );
  XNOR2_X1 U11346 ( .A(n12410), .B(n12409), .ZN(n15342) );
  NAND2_X1 U11347 ( .A1(n11363), .A2(n11365), .ZN(n12407) );
  CLKBUF_X2 U11348 ( .A(n13935), .Z(n13936) );
  NOR2_X1 U11349 ( .A1(n21350), .A2(n21360), .ZN(n21345) );
  INV_X1 U11350 ( .A(n16898), .ZN(n11148) );
  NAND2_X1 U11351 ( .A1(n16564), .A2(n17473), .ZN(n11284) );
  INV_X1 U11352 ( .A(n19828), .ZN(n11145) );
  AND2_X1 U11353 ( .A1(n11202), .A2(n12099), .ZN(n19878) );
  OAI22_X2 U11354 ( .A1(n21194), .A2(n21193), .B1(n21192), .B2(n21191), .ZN(
        n21379) );
  INV_X1 U11355 ( .A(n12095), .ZN(n12110) );
  CLKBUF_X2 U11356 ( .A(n12095), .Z(n12098) );
  NOR2_X1 U11357 ( .A1(n14840), .A2(n14825), .ZN(n22749) );
  NOR2_X2 U11358 ( .A1(n21687), .A2(n21849), .ZN(n21659) );
  NAND2_X1 U11359 ( .A1(n21878), .A2(n11372), .ZN(n21849) );
  NAND2_X1 U11360 ( .A1(n21886), .A2(n21861), .ZN(n21687) );
  NAND2_X1 U11361 ( .A1(n15747), .A2(n21410), .ZN(n21878) );
  INV_X4 U11362 ( .A(n20860), .ZN(n21155) );
  OAI21_X1 U11363 ( .B1(n21384), .B2(n18490), .A(n21415), .ZN(n21778) );
  NOR2_X1 U11364 ( .A1(n15798), .A2(n15797), .ZN(n15799) );
  AND2_X1 U11365 ( .A1(n12003), .A2(n14170), .ZN(n12046) );
  NAND2_X1 U11366 ( .A1(n14202), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12040) );
  NAND2_X4 U11367 ( .A1(n12997), .A2(n12031), .ZN(n14171) );
  OR3_X1 U11368 ( .A1(n15788), .A2(n11551), .A3(n11549), .ZN(n11548) );
  INV_X2 U11369 ( .A(n21434), .ZN(n21440) );
  CLKBUF_X1 U11370 ( .A(n14226), .Z(n14313) );
  NAND2_X1 U11371 ( .A1(n14797), .A2(n14886), .ZN(n21947) );
  NAND2_X2 U11372 ( .A1(n19017), .A2(n11267), .ZN(n12031) );
  INV_X1 U11373 ( .A(n11618), .ZN(n11614) );
  NAND2_X1 U11374 ( .A1(n20166), .A2(n20206), .ZN(n12030) );
  INV_X2 U11375 ( .A(n15178), .ZN(n14797) );
  NAND2_X2 U11376 ( .A1(n13922), .A2(n15178), .ZN(n14226) );
  INV_X1 U11377 ( .A(n12006), .ZN(n12011) );
  INV_X2 U11378 ( .A(n11955), .ZN(n11146) );
  NAND2_X1 U11379 ( .A1(n11592), .A2(n11591), .ZN(n12026) );
  NAND2_X1 U11380 ( .A1(n11191), .A2(n11164), .ZN(n14628) );
  OR2_X2 U11381 ( .A1(n13091), .A2(n13090), .ZN(n13156) );
  INV_X1 U11382 ( .A(n11190), .ZN(n18436) );
  INV_X4 U11383 ( .A(n18202), .ZN(n18461) );
  CLKBUF_X2 U11384 ( .A(n13231), .Z(n13832) );
  CLKBUF_X2 U11385 ( .A(n15716), .Z(n18435) );
  CLKBUF_X2 U11386 ( .A(n13238), .Z(n13805) );
  CLKBUF_X2 U11387 ( .A(n13122), .Z(n14692) );
  CLKBUF_X2 U11388 ( .A(n13237), .Z(n13806) );
  CLKBUF_X2 U11389 ( .A(n13254), .Z(n13232) );
  CLKBUF_X2 U11390 ( .A(n13203), .Z(n13833) );
  CLKBUF_X2 U11391 ( .A(n13253), .Z(n13803) );
  CLKBUF_X2 U11392 ( .A(n13208), .Z(n13804) );
  CLKBUF_X2 U11393 ( .A(n13143), .Z(n13576) );
  CLKBUF_X3 U11394 ( .A(n15713), .Z(n11152) );
  NOR2_X1 U11395 ( .A1(n15652), .A2(n15650), .ZN(n18153) );
  INV_X4 U11396 ( .A(n15724), .ZN(n18414) );
  CLKBUF_X2 U11397 ( .A(n15290), .Z(n21945) );
  AND2_X2 U11398 ( .A1(n15060), .A2(n12214), .ZN(n11986) );
  AND2_X1 U11399 ( .A1(n13305), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13046) );
  AND2_X1 U11400 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14641) );
  INV_X2 U11401 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13305) );
  NOR2_X1 U11402 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20764) );
  OAI21_X1 U11403 ( .B1(n15953), .B2(n15954), .A(n15941), .ZN(n16265) );
  AND2_X1 U11404 ( .A1(n11288), .A2(n14028), .ZN(n11287) );
  NAND2_X1 U11405 ( .A1(n11650), .A2(n16274), .ZN(n11658) );
  XNOR2_X1 U11406 ( .A(n15821), .B(n15820), .ZN(n15921) );
  OR2_X1 U11407 ( .A1(n11333), .A2(n17184), .ZN(n11330) );
  NOR3_X1 U11408 ( .A1(n15876), .A2(n15875), .A3(n15874), .ZN(n15877) );
  NAND2_X1 U11409 ( .A1(n11696), .A2(n11695), .ZN(n11694) );
  NOR2_X1 U11410 ( .A1(n15882), .A2(n19302), .ZN(n15876) );
  OR2_X1 U11411 ( .A1(n14061), .A2(n17873), .ZN(n11288) );
  OAI22_X1 U11412 ( .A1(n11358), .A2(n11357), .B1(n11362), .B2(n16900), .ZN(
        n11356) );
  AND2_X1 U11413 ( .A1(n15884), .A2(n15883), .ZN(n15885) );
  NAND2_X1 U11414 ( .A1(n17216), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17209) );
  NOR2_X1 U11415 ( .A1(n11653), .A2(n11652), .ZN(n11661) );
  NAND2_X1 U11416 ( .A1(n16275), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16274) );
  AND2_X1 U11417 ( .A1(n16929), .A2(n16927), .ZN(n16914) );
  AOI22_X1 U11418 ( .A1(n11450), .A2(n12360), .B1(n12359), .B2(n14197), .ZN(
        n12364) );
  AND2_X1 U11419 ( .A1(n14014), .A2(n16266), .ZN(n16275) );
  INV_X1 U11420 ( .A(n16266), .ZN(n11653) );
  INV_X1 U11421 ( .A(n16986), .ZN(n11147) );
  AND2_X1 U11422 ( .A1(n11570), .A2(n11379), .ZN(n11378) );
  AOI21_X1 U11423 ( .B1(n19252), .B2(n19298), .A(n11722), .ZN(n15872) );
  OAI21_X1 U11424 ( .B1(n17068), .B2(n14207), .A(n11381), .ZN(n11380) );
  AND2_X2 U11425 ( .A1(n11630), .A2(n11631), .ZN(n16069) );
  NOR2_X1 U11426 ( .A1(n16657), .A2(n11528), .ZN(n11527) );
  NAND2_X1 U11427 ( .A1(n16891), .A2(n16956), .ZN(n12324) );
  NAND2_X1 U11428 ( .A1(n11273), .A2(n11286), .ZN(n17339) );
  AND2_X1 U11429 ( .A1(n11665), .A2(n20603), .ZN(n11664) );
  AOI21_X1 U11430 ( .B1(n11667), .B2(n11428), .A(n11283), .ZN(n11427) );
  OR2_X1 U11431 ( .A1(n14009), .A2(n11666), .ZN(n11665) );
  OAI21_X1 U11432 ( .B1(n12420), .B2(n12415), .A(n12419), .ZN(n12421) );
  NAND2_X1 U11433 ( .A1(n11270), .A2(n11268), .ZN(n11337) );
  OR2_X1 U11434 ( .A1(n20619), .A2(n14008), .ZN(n11283) );
  CLKBUF_X1 U11435 ( .A(n12414), .Z(n12415) );
  NAND2_X1 U11436 ( .A1(n13362), .A2(n13361), .ZN(n15035) );
  XNOR2_X1 U11437 ( .A(n13983), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n20594) );
  NAND2_X1 U11438 ( .A1(n13982), .A2(n13981), .ZN(n13983) );
  INV_X2 U11439 ( .A(n20617), .ZN(n20603) );
  NAND2_X1 U11440 ( .A1(n11594), .A2(n12407), .ZN(n12409) );
  NAND2_X1 U11441 ( .A1(n13404), .A2(n13405), .ZN(n13965) );
  NAND2_X1 U11442 ( .A1(n19192), .A2(n19191), .ZN(n19190) );
  OR2_X1 U11443 ( .A1(n12172), .A2(n12173), .ZN(n11365) );
  XNOR2_X1 U11444 ( .A(n13335), .B(n22582), .ZN(n11649) );
  OR2_X1 U11445 ( .A1(n18791), .A2(n11302), .ZN(n11301) );
  NAND2_X2 U11446 ( .A1(n11284), .A2(n13325), .ZN(n22582) );
  AND2_X1 U11447 ( .A1(n11562), .A2(n11242), .ZN(n19161) );
  INV_X1 U11448 ( .A(n12239), .ZN(n19838) );
  NAND2_X1 U11449 ( .A1(n12096), .A2(n11202), .ZN(n19828) );
  NOR2_X2 U11450 ( .A1(n12092), .A2(n12102), .ZN(n12187) );
  NAND2_X1 U11451 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n21379), .ZN(n21369) );
  NOR2_X1 U11452 ( .A1(n14840), .A2(n14817), .ZN(n22722) );
  NOR2_X1 U11453 ( .A1(n14840), .A2(n14804), .ZN(n22776) );
  NOR2_X1 U11454 ( .A1(n14840), .A2(n14809), .ZN(n22695) );
  NOR2_X1 U11455 ( .A1(n14840), .A2(n15908), .ZN(n22839) );
  INV_X1 U11456 ( .A(n12118), .ZN(n12102) );
  AND2_X2 U11457 ( .A1(n22280), .A2(n13911), .ZN(n20628) );
  NAND2_X1 U11458 ( .A1(n12091), .A2(n12090), .ZN(n19029) );
  NAND2_X1 U11459 ( .A1(n11373), .A2(n12064), .ZN(n12436) );
  NAND2_X2 U11460 ( .A1(n20574), .A2(n14628), .ZN(n16146) );
  NOR2_X1 U11461 ( .A1(n14840), .A2(n15177), .ZN(n22608) );
  INV_X1 U11462 ( .A(n21878), .ZN(n18491) );
  NAND2_X1 U11463 ( .A1(n13268), .A2(n13267), .ZN(n13290) );
  AND2_X1 U11464 ( .A1(n12437), .A2(n12077), .ZN(n12439) );
  CLKBUF_X1 U11465 ( .A(n13292), .Z(n17438) );
  OAI211_X1 U11466 ( .C1(n13910), .C2(n22585), .A(n13201), .B(n13200), .ZN(
        n13202) );
  OR2_X1 U11467 ( .A1(n12076), .A2(n12075), .ZN(n12437) );
  INV_X2 U11468 ( .A(n16700), .ZN(n15538) );
  NOR2_X2 U11469 ( .A1(n20024), .A2(n20291), .ZN(n20025) );
  NOR2_X2 U11470 ( .A1(n20072), .A2(n20291), .ZN(n20073) );
  NOR2_X2 U11471 ( .A1(n19818), .A2(n20291), .ZN(n19819) );
  NAND2_X1 U11472 ( .A1(n13908), .A2(n13907), .ZN(n14712) );
  OR2_X1 U11473 ( .A1(n13306), .A2(n14697), .ZN(n13201) );
  OAI21_X1 U11474 ( .B1(n13306), .B2(n13179), .A(n13182), .ZN(n13252) );
  INV_X2 U11475 ( .A(n20714), .ZN(n20763) );
  NAND2_X1 U11476 ( .A1(n18866), .A2(n18474), .ZN(n18477) );
  OR2_X1 U11477 ( .A1(n12444), .A2(n12070), .ZN(n12074) );
  INV_X2 U11478 ( .A(n12444), .ZN(n15864) );
  CLKBUF_X1 U11479 ( .A(n19227), .Z(n19251) );
  OAI21_X1 U11480 ( .B1(n21874), .B2(n17408), .A(n20710), .ZN(n15749) );
  INV_X1 U11481 ( .A(n12069), .ZN(n12444) );
  AND2_X2 U11482 ( .A1(n11553), .A2(n11552), .ZN(n15795) );
  NAND2_X1 U11483 ( .A1(n12017), .A2(n12016), .ZN(n15072) );
  AND2_X1 U11484 ( .A1(n13177), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13194) );
  AND2_X1 U11485 ( .A1(n15770), .A2(n15737), .ZN(n21874) );
  AND2_X1 U11486 ( .A1(n15799), .A2(n11255), .ZN(n15377) );
  NAND3_X1 U11487 ( .A1(n18651), .A2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18698) );
  CLKBUF_X1 U11488 ( .A(n12440), .Z(n15865) );
  NAND2_X1 U11489 ( .A1(n11143), .A2(n11554), .ZN(n15798) );
  OR2_X1 U11490 ( .A1(n13023), .A2(n11295), .ZN(n12048) );
  XNOR2_X1 U11491 ( .A(n18452), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18895) );
  AND2_X1 U11492 ( .A1(n18523), .A2(n11237), .ZN(n18597) );
  OR2_X1 U11493 ( .A1(n14361), .A2(n15109), .ZN(n12441) );
  NAND2_X1 U11494 ( .A1(n13161), .A2(n14628), .ZN(n14549) );
  CLKBUF_X1 U11495 ( .A(n12386), .Z(n14029) );
  OR2_X1 U11496 ( .A1(n18495), .A2(n18450), .ZN(n18452) );
  AND2_X1 U11497 ( .A1(n11296), .A2(n11293), .ZN(n14053) );
  MUX2_X1 U11498 ( .A(n13092), .B(n14537), .S(n13156), .Z(n13114) );
  INV_X1 U11499 ( .A(n19708), .ZN(n11367) );
  OR2_X1 U11500 ( .A1(n13160), .A2(n15908), .ZN(n14686) );
  CLKBUF_X1 U11501 ( .A(n13168), .Z(n16573) );
  AND2_X1 U11502 ( .A1(n20125), .A2(n11294), .ZN(n11293) );
  BUF_X1 U11503 ( .A(n12022), .Z(n14071) );
  OR2_X2 U11504 ( .A1(n20695), .A2(n20639), .ZN(n20680) );
  NAND2_X1 U11505 ( .A1(n14809), .A2(n14839), .ZN(n14725) );
  AND2_X2 U11506 ( .A1(n19017), .A2(n19975), .ZN(n15806) );
  OR2_X1 U11507 ( .A1(n12012), .A2(n11955), .ZN(n12007) );
  INV_X1 U11508 ( .A(n14178), .ZN(n20166) );
  NAND2_X2 U11509 ( .A1(n13053), .A2(n13052), .ZN(n13157) );
  CLKBUF_X1 U11510 ( .A(n12012), .Z(n12013) );
  INV_X1 U11511 ( .A(n13922), .ZN(n14809) );
  OR2_X1 U11512 ( .A1(n15432), .A2(n19072), .ZN(n15442) );
  INV_X2 U11513 ( .A(U214), .ZN(n20695) );
  NAND2_X1 U11514 ( .A1(n11729), .A2(n11715), .ZN(n13922) );
  NAND2_X1 U11515 ( .A1(n11927), .A2(n11926), .ZN(n12012) );
  INV_X1 U11516 ( .A(n13156), .ZN(n14839) );
  AND4_X1 U11517 ( .A1(n13132), .A2(n13120), .A3(n11616), .A4(n11221), .ZN(
        n11615) );
  NAND2_X1 U11518 ( .A1(n11972), .A2(n11971), .ZN(n14178) );
  AND3_X1 U11519 ( .A1(n13044), .A2(n13043), .A3(n13042), .ZN(n13053) );
  INV_X1 U11520 ( .A(n14817), .ZN(n14548) );
  AND3_X1 U11521 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n20836), .ZN(n18807) );
  AND4_X2 U11522 ( .A1(n13081), .A2(n13080), .A3(n13079), .A4(n13078), .ZN(
        n14817) );
  AND4_X1 U11523 ( .A1(n13130), .A2(n13129), .A3(n13128), .A4(n13127), .ZN(
        n13131) );
  AND4_X1 U11524 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13155) );
  NAND2_X1 U11525 ( .A1(n11730), .A2(n11732), .ZN(n13275) );
  BUF_X2 U11526 ( .A(n11126), .Z(n18317) );
  AND4_X1 U11527 ( .A1(n13065), .A2(n13064), .A3(n13063), .A4(n13062), .ZN(
        n13081) );
  AND4_X1 U11528 ( .A1(n13031), .A2(n13030), .A3(n13029), .A4(n13028), .ZN(
        n13044) );
  AND4_X1 U11529 ( .A1(n13069), .A2(n13068), .A3(n13067), .A4(n13066), .ZN(
        n13080) );
  AND4_X1 U11530 ( .A1(n13073), .A2(n13072), .A3(n13071), .A4(n13070), .ZN(
        n13079) );
  AND4_X1 U11531 ( .A1(n13077), .A2(n13076), .A3(n13075), .A4(n13074), .ZN(
        n13078) );
  AND4_X1 U11532 ( .A1(n13119), .A2(n13118), .A3(n13117), .A4(n13116), .ZN(
        n13133) );
  BUF_X2 U11533 ( .A(n15725), .Z(n18181) );
  AND4_X1 U11534 ( .A1(n13152), .A2(n13151), .A3(n13150), .A4(n13149), .ZN(
        n13153) );
  NOR2_X1 U11535 ( .A1(n18848), .A2(n18849), .ZN(n20836) );
  AND4_X1 U11536 ( .A1(n13126), .A2(n13125), .A3(n13124), .A4(n13123), .ZN(
        n13132) );
  INV_X2 U11537 ( .A(n11746), .ZN(n12984) );
  NOR2_X1 U11538 ( .A1(n21418), .A2(n21385), .ZN(n18409) );
  AND2_X1 U11539 ( .A1(n11756), .A2(n11755), .ZN(n11376) );
  AND3_X1 U11540 ( .A1(n11759), .A2(n11758), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11762) );
  BUF_X2 U11541 ( .A(n15716), .Z(n18421) );
  INV_X2 U11542 ( .A(n20408), .ZN(n20457) );
  BUF_X4 U11543 ( .A(n18087), .Z(n11149) );
  NOR2_X1 U11544 ( .A1(n21389), .A2(n18910), .ZN(n18977) );
  NAND2_X1 U11545 ( .A1(n21398), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n21401) );
  BUF_X4 U11546 ( .A(n13144), .Z(n13835) );
  INV_X2 U11547 ( .A(n22347), .ZN(n17980) );
  INV_X1 U11548 ( .A(n11772), .ZN(n11958) );
  CLKBUF_X2 U11549 ( .A(n12979), .Z(n12973) );
  BUF_X1 U11550 ( .A(n11965), .Z(n11957) );
  AND2_X1 U11551 ( .A1(n11418), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13045) );
  AND2_X1 U11552 ( .A1(n11734), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11743) );
  NOR2_X2 U11553 ( .A1(n11646), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13047) );
  AND2_X1 U11554 ( .A1(n14641), .A2(n16572), .ZN(n13093) );
  AND2_X2 U11555 ( .A1(n13032), .A2(n14641), .ZN(n13144) );
  NOR2_X2 U11556 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13037) );
  NOR2_X1 U11557 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11736) );
  AND2_X1 U11558 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11733) );
  INV_X1 U11559 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14697) );
  NOR2_X2 U11560 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13032) );
  INV_X2 U11561 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21891) );
  NOR2_X1 U11562 ( .A1(n16840), .A2(n17091), .ZN(n16828) );
  NOR2_X4 U11563 ( .A1(n15979), .A2(n15980), .ZN(n15969) );
  NAND2_X2 U11564 ( .A1(n15992), .A2(n15994), .ZN(n15979) );
  NAND2_X2 U11565 ( .A1(n17863), .A2(n12434), .ZN(n16986) );
  OAI21_X2 U11566 ( .B1(n16338), .B2(n14012), .A(n20617), .ZN(n16307) );
  NAND2_X1 U11567 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  INV_X1 U11568 ( .A(n18779), .ZN(n18830) );
  NOR2_X4 U11569 ( .A1(n21450), .A2(n18914), .ZN(n18779) );
  OAI21_X1 U11570 ( .B1(n13306), .B2(n14727), .A(n13175), .ZN(n13178) );
  AND2_X4 U11571 ( .A1(n14886), .A2(n15178), .ZN(n14222) );
  NAND2_X2 U11572 ( .A1(n15497), .A2(n11432), .ZN(n20604) );
  NAND2_X2 U11573 ( .A1(n15499), .A2(n15498), .ZN(n15497) );
  INV_X1 U11574 ( .A(n13994), .ZN(n11153) );
  INV_X1 U11575 ( .A(n13994), .ZN(n11154) );
  OAI21_X2 U11576 ( .B1(n17039), .B2(n11341), .A(n11339), .ZN(n16891) );
  XNOR2_X1 U11577 ( .A(n13290), .B(n13289), .ZN(n16562) );
  XNOR2_X1 U11578 ( .A(n21169), .B(n18727), .ZN(n20860) );
  AOI21_X2 U11579 ( .B1(n15943), .B2(n15941), .A(n15942), .ZN(n16250) );
  AND2_X1 U11580 ( .A1(n11553), .A2(n11552), .ZN(n11157) );
  AND2_X1 U11581 ( .A1(n11553), .A2(n11552), .ZN(n11158) );
  CLKBUF_X1 U11582 ( .A(n20836), .Z(n11159) );
  NOR3_X1 U11583 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n21408), .ZN(n15713) );
  AND4_X1 U11584 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11906) );
  AND4_X1 U11585 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11904) );
  NOR2_X1 U11586 ( .A1(n11833), .A2(n11832), .ZN(n11834) );
  INV_X1 U11587 ( .A(n11831), .ZN(n11833) );
  INV_X1 U11588 ( .A(n11347), .ZN(n11346) );
  OR2_X1 U11589 ( .A1(n21943), .A2(n15169), .ZN(n16102) );
  NAND2_X1 U11590 ( .A1(n16899), .A2(n11148), .ZN(n11362) );
  OR2_X1 U11591 ( .A1(n12426), .A2(n12425), .ZN(n12430) );
  AND2_X1 U11592 ( .A1(n11241), .A2(n12129), .ZN(n11364) );
  AND3_X1 U11593 ( .A1(n20206), .A2(n14178), .A3(n12006), .ZN(n11296) );
  INV_X1 U11594 ( .A(n14725), .ZN(n14216) );
  NAND2_X1 U11595 ( .A1(n11640), .A2(n13780), .ZN(n11639) );
  NOR2_X1 U11596 ( .A1(n11641), .A2(n15943), .ZN(n11640) );
  INV_X1 U11597 ( .A(n15954), .ZN(n11641) );
  NOR2_X1 U11598 ( .A1(n11632), .A2(n11634), .ZN(n11631) );
  NAND2_X1 U11599 ( .A1(n17436), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13822) );
  NAND2_X1 U11600 ( .A1(n11170), .A2(n15372), .ZN(n11619) );
  NOR2_X2 U11601 ( .A1(n13275), .A2(n22605), .ZN(n13537) );
  AND2_X1 U11602 ( .A1(n12261), .A2(n12205), .ZN(n11458) );
  OR2_X1 U11603 ( .A1(n12298), .A2(n12308), .ZN(n12313) );
  AND3_X1 U11604 ( .A1(n12036), .A2(n11205), .A3(n12035), .ZN(n11690) );
  AOI21_X1 U11605 ( .B1(n15072), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n12018), 
        .ZN(n12019) );
  BUF_X4 U11606 ( .A(n11965), .Z(n12976) );
  NAND2_X1 U11607 ( .A1(n14053), .A2(n14479), .ZN(n14361) );
  XNOR2_X1 U11608 ( .A(n11690), .B(n11689), .ZN(n12084) );
  INV_X1 U11609 ( .A(n15830), .ZN(n15805) );
  AND2_X2 U11610 ( .A1(n14470), .A2(n14065), .ZN(n14136) );
  OAI21_X1 U11611 ( .B1(n12013), .B2(n19322), .A(n19975), .ZN(n12564) );
  AOI221_X1 U11612 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n12380), 
        .C1(n19273), .C2(n12380), .A(n12379), .ZN(n13020) );
  NOR3_X1 U11613 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n15651), .ZN(n18087) );
  OR2_X1 U11614 ( .A1(n21223), .A2(n18447), .ZN(n18446) );
  OAI211_X1 U11615 ( .C1(n15756), .C2(n15755), .A(n15764), .B(n15754), .ZN(
        n18486) );
  NOR2_X1 U11616 ( .A1(n21877), .A2(n18487), .ZN(n17985) );
  NOR2_X1 U11617 ( .A1(n14886), .A2(n15178), .ZN(n15911) );
  OR2_X1 U11618 ( .A1(n13734), .A2(n16285), .ZN(n13774) );
  INV_X1 U11619 ( .A(n11667), .ZN(n11429) );
  INV_X1 U11620 ( .A(n11432), .ZN(n11428) );
  INV_X1 U11621 ( .A(n15300), .ZN(n13430) );
  AND2_X1 U11622 ( .A1(n11658), .A2(n11656), .ZN(n15844) );
  NOR2_X1 U11623 ( .A1(n22569), .A2(n16592), .ZN(n22507) );
  INV_X1 U11624 ( .A(n14816), .ZN(n16592) );
  XNOR2_X1 U11625 ( .A(n12913), .B(n12914), .ZN(n16678) );
  NAND2_X1 U11626 ( .A1(n16678), .A2(n16677), .ZN(n16676) );
  INV_X1 U11627 ( .A(n11596), .ZN(n11595) );
  OAI21_X1 U11628 ( .B1(n17037), .B2(n11597), .A(n17864), .ZN(n11596) );
  INV_X1 U11629 ( .A(n12429), .ZN(n11597) );
  NAND2_X1 U11630 ( .A1(n12082), .A2(n12081), .ZN(n12085) );
  CLKBUF_X2 U11631 ( .A(n14085), .Z(n15828) );
  NAND2_X1 U11632 ( .A1(n11180), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11598) );
  NOR2_X1 U11633 ( .A1(n12369), .A2(n17075), .ZN(n16814) );
  AND2_X1 U11634 ( .A1(n11166), .A2(n11705), .ZN(n11704) );
  NAND2_X1 U11635 ( .A1(n11148), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11705) );
  NAND2_X1 U11636 ( .A1(n11236), .A2(n11489), .ZN(n11485) );
  NAND2_X1 U11637 ( .A1(n11336), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11335) );
  AOI21_X1 U11638 ( .B1(n14058), .B2(n14057), .A(n14056), .ZN(n14059) );
  NOR2_X1 U11639 ( .A1(n20711), .A2(n15749), .ZN(n21879) );
  NOR2_X1 U11640 ( .A1(n21666), .A2(n21703), .ZN(n21682) );
  NAND3_X1 U11641 ( .A1(n15734), .A2(n15733), .A3(n15732), .ZN(n21435) );
  AOI211_X1 U11642 ( .C1(n11131), .C2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n15731), .B(n15730), .ZN(n15732) );
  NAND2_X1 U11643 ( .A1(n15166), .A2(n15165), .ZN(n21943) );
  NOR2_X1 U11644 ( .A1(n19131), .A2(n19130), .ZN(n19129) );
  INV_X1 U11645 ( .A(n16888), .ZN(n11336) );
  OAI21_X1 U11646 ( .B1(n17656), .B2(n17657), .A(n11523), .ZN(n11522) );
  XNOR2_X1 U11647 ( .A(n17658), .B(n11524), .ZN(n11523) );
  AOI221_X1 U11648 ( .B1(DATAI_31_), .B2(keyinput_1), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_0), .A(n17655), .ZN(n17656)
         );
  XNOR2_X1 U11649 ( .A(keyinput_8), .B(DATAI_24_), .ZN(n11521) );
  OAI21_X1 U11650 ( .B1(n17500), .B2(n17501), .A(n11408), .ZN(n11407) );
  XNOR2_X1 U11651 ( .A(n17658), .B(n11409), .ZN(n11408) );
  XNOR2_X1 U11652 ( .A(n17502), .B(keyinput_136), .ZN(n11406) );
  NAND2_X1 U11653 ( .A1(n11493), .A2(n17692), .ZN(n17696) );
  OAI21_X1 U11654 ( .B1(n11496), .B2(n17688), .A(n11494), .ZN(n11493) );
  INV_X1 U11655 ( .A(keyinput_45), .ZN(n11503) );
  OAI21_X1 U11656 ( .B1(n17715), .B2(n11253), .A(n11505), .ZN(n11504) );
  INV_X1 U11657 ( .A(n17716), .ZN(n11505) );
  OAI22_X1 U11658 ( .A1(n17714), .A2(n17713), .B1(keyinput_42), .B2(
        P1_D_C_N_REG_SCAN_IN), .ZN(n17715) );
  OAI21_X1 U11659 ( .B1(n17547), .B2(n11396), .A(n11395), .ZN(n11394) );
  AND2_X1 U11660 ( .A1(n17548), .A2(keyinput_170), .ZN(n11396) );
  INV_X1 U11661 ( .A(n17549), .ZN(n11395) );
  XNOR2_X1 U11662 ( .A(n17717), .B(n11393), .ZN(n11392) );
  INV_X1 U11663 ( .A(keyinput_173), .ZN(n11393) );
  INV_X1 U11664 ( .A(n17738), .ZN(n11519) );
  INV_X1 U11665 ( .A(n17568), .ZN(n11416) );
  NAND2_X1 U11666 ( .A1(n11412), .A2(n11410), .ZN(n17583) );
  NOR2_X1 U11667 ( .A1(n17579), .A2(n11411), .ZN(n11410) );
  NAND2_X1 U11668 ( .A1(n11414), .A2(n11413), .ZN(n11412) );
  XNOR2_X1 U11669 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_199), .ZN(n11411)
         );
  CLKBUF_X1 U11670 ( .A(n11136), .Z(n13811) );
  AND2_X1 U11671 ( .A1(n14215), .A2(n14628), .ZN(n13856) );
  AOI211_X1 U11672 ( .C1(n17786), .C2(n17787), .A(n17785), .B(n17784), .ZN(
        n11512) );
  INV_X1 U11673 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11646) );
  OR2_X1 U11674 ( .A1(n12182), .A2(n12243), .ZN(n12244) );
  NAND2_X1 U11675 ( .A1(n11745), .A2(n11744), .ZN(n11772) );
  NAND2_X1 U11676 ( .A1(n11980), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11759) );
  AOI22_X1 U11677 ( .A1(n11958), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11965), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11435) );
  OR2_X1 U11678 ( .A1(n15755), .A2(n15756), .ZN(n15751) );
  NAND2_X1 U11679 ( .A1(n11624), .A2(n11622), .ZN(n13987) );
  NOR2_X1 U11680 ( .A1(n13405), .A2(n11623), .ZN(n11622) );
  INV_X1 U11681 ( .A(n13394), .ZN(n11623) );
  NAND2_X1 U11682 ( .A1(n13856), .A2(n14817), .ZN(n13183) );
  NAND2_X1 U11683 ( .A1(n13273), .A2(n13985), .ZN(n13283) );
  OAI21_X1 U11684 ( .B1(n14549), .B2(n14522), .A(n14547), .ZN(n13163) );
  OR2_X1 U11685 ( .A1(n14548), .A2(n17473), .ZN(n13314) );
  AND4_X1 U11686 ( .A1(n11847), .A2(n11846), .A3(n11845), .A4(n11844), .ZN(
        n11849) );
  NAND2_X1 U11687 ( .A1(n12128), .A2(n15109), .ZN(n12129) );
  MUX2_X1 U11688 ( .A(n11811), .B(n15410), .S(n15857), .Z(n12221) );
  AND3_X1 U11689 ( .A1(n12169), .A2(n12168), .A3(n12167), .ZN(n12399) );
  INV_X1 U11690 ( .A(n20206), .ZN(n14172) );
  NAND2_X1 U11691 ( .A1(n12001), .A2(n12000), .ZN(n11433) );
  NOR2_X1 U11692 ( .A1(n20206), .A2(n11999), .ZN(n12000) );
  AND2_X1 U11693 ( .A1(n19276), .A2(n12086), .ZN(n12118) );
  AND2_X1 U11694 ( .A1(n12116), .A2(n12117), .ZN(n12121) );
  NOR2_X1 U11695 ( .A1(n21231), .A2(n18449), .ZN(n18448) );
  INV_X1 U11696 ( .A(n11420), .ZN(n13854) );
  NOR2_X1 U11697 ( .A1(n11469), .A2(n15966), .ZN(n11468) );
  INV_X1 U11698 ( .A(n15956), .ZN(n11469) );
  AND2_X1 U11699 ( .A1(n11626), .A2(n16011), .ZN(n11625) );
  NOR2_X1 U11700 ( .A1(n16018), .A2(n11627), .ZN(n11626) );
  INV_X1 U11701 ( .A(n11628), .ZN(n11627) );
  NOR2_X1 U11702 ( .A1(n16028), .A2(n11629), .ZN(n11628) );
  INV_X1 U11703 ( .A(n16046), .ZN(n11629) );
  INV_X1 U11704 ( .A(n11283), .ZN(n14009) );
  AND2_X1 U11705 ( .A1(n11667), .A2(n14011), .ZN(n11663) );
  INV_X1 U11706 ( .A(n13822), .ZN(n13844) );
  NAND2_X1 U11707 ( .A1(n13544), .A2(n11635), .ZN(n11634) );
  INV_X1 U11708 ( .A(n16131), .ZN(n11635) );
  INV_X1 U11709 ( .A(n16137), .ZN(n13544) );
  NAND2_X1 U11710 ( .A1(n15558), .A2(n13481), .ZN(n15617) );
  INV_X1 U11711 ( .A(n15353), .ZN(n11620) );
  NOR2_X1 U11712 ( .A1(n11231), .A2(n11657), .ZN(n11656) );
  INV_X1 U11713 ( .A(n11659), .ZN(n11657) );
  NAND2_X1 U11714 ( .A1(n16037), .A2(n11481), .ZN(n11480) );
  INV_X1 U11715 ( .A(n16048), .ZN(n11481) );
  NAND2_X1 U11716 ( .A1(n11477), .A2(n14288), .ZN(n11476) );
  NOR2_X1 U11717 ( .A1(n16133), .A2(n16138), .ZN(n11477) );
  AND2_X1 U11718 ( .A1(n16390), .A2(n13993), .ZN(n11432) );
  NAND2_X1 U11719 ( .A1(n14222), .A2(n14327), .ZN(n14326) );
  AND2_X1 U11720 ( .A1(n14684), .A2(n13188), .ZN(n14544) );
  OR2_X1 U11721 ( .A1(n13244), .A2(n13243), .ZN(n13988) );
  INV_X1 U11722 ( .A(n13899), .ZN(n13891) );
  NAND2_X1 U11723 ( .A1(n11419), .A2(n13168), .ZN(n13113) );
  OR2_X1 U11724 ( .A1(n13115), .A2(n14226), .ZN(n14684) );
  AND2_X1 U11725 ( .A1(n22602), .A2(n13308), .ZN(n16585) );
  AND3_X2 U11726 ( .A1(n14886), .A2(n14548), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n13899) );
  INV_X1 U11727 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22584) );
  INV_X1 U11728 ( .A(n12304), .ZN(n11453) );
  INV_X1 U11729 ( .A(n12266), .ZN(n11457) );
  INV_X1 U11730 ( .A(n16734), .ZN(n11582) );
  NOR2_X1 U11731 ( .A1(n16757), .A2(n11580), .ZN(n11579) );
  INV_X1 U11732 ( .A(n16748), .ZN(n11580) );
  INV_X1 U11733 ( .A(n12934), .ZN(n12910) );
  AND2_X1 U11734 ( .A1(n11685), .A2(n11684), .ZN(n11683) );
  INV_X1 U11735 ( .A(n16723), .ZN(n11684) );
  AND2_X1 U11736 ( .A1(n11590), .A2(n11589), .ZN(n11588) );
  INV_X1 U11737 ( .A(n16797), .ZN(n11589) );
  AND2_X1 U11738 ( .A1(n14756), .A2(n14752), .ZN(n11585) );
  NOR2_X1 U11739 ( .A1(n12997), .A2(n12030), .ZN(n14175) );
  INV_X1 U11740 ( .A(n11975), .ZN(n14174) );
  NAND2_X1 U11741 ( .A1(n14468), .A2(n19017), .ZN(n12934) );
  INV_X1 U11742 ( .A(n14092), .ZN(n14095) );
  AOI21_X1 U11743 ( .B1(n14503), .B2(n11187), .A(n14093), .ZN(n14092) );
  AND2_X1 U11744 ( .A1(n14499), .A2(n14498), .ZN(n14088) );
  NAND2_X1 U11745 ( .A1(n11146), .A2(n12012), .ZN(n12022) );
  NAND2_X1 U11746 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11567) );
  INV_X1 U11747 ( .A(n14902), .ZN(n12461) );
  NAND2_X1 U11748 ( .A1(n12461), .A2(n11543), .ZN(n11542) );
  INV_X1 U11749 ( .A(n14910), .ZN(n11543) );
  NAND2_X1 U11750 ( .A1(n12431), .A2(n15859), .ZN(n12432) );
  NAND2_X1 U11751 ( .A1(n12074), .A2(n11204), .ZN(n12075) );
  CLKBUF_X1 U11752 ( .A(n12084), .Z(n12086) );
  OAI21_X1 U11753 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14017), .A(
        n16837), .ZN(n11450) );
  NAND2_X1 U11754 ( .A1(n16858), .A2(n12345), .ZN(n11707) );
  AND2_X1 U11755 ( .A1(n11709), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11708) );
  NAND2_X1 U11756 ( .A1(n11704), .A2(n16881), .ZN(n11443) );
  NOR2_X1 U11757 ( .A1(n11446), .A2(n11443), .ZN(n11440) );
  NAND2_X1 U11758 ( .A1(n11445), .A2(n11704), .ZN(n11444) );
  AND2_X1 U11759 ( .A1(n11703), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11447) );
  INV_X1 U11760 ( .A(n12323), .ZN(n11445) );
  INV_X1 U11761 ( .A(n16927), .ZN(n11488) );
  NOR2_X1 U11762 ( .A1(n14773), .A2(n14772), .ZN(n14771) );
  INV_X1 U11763 ( .A(n12268), .ZN(n11702) );
  OR2_X1 U11764 ( .A1(n12272), .A2(n19307), .ZN(n17868) );
  INV_X1 U11765 ( .A(n15517), .ZN(n11574) );
  NAND2_X1 U11766 ( .A1(n15342), .A2(n15521), .ZN(n12412) );
  NAND2_X1 U11767 ( .A1(n12130), .A2(n12129), .ZN(n11289) );
  NAND2_X1 U11768 ( .A1(n11192), .A2(n11767), .ZN(n11592) );
  NAND3_X1 U11769 ( .A1(n11593), .A2(n11771), .A3(n11770), .ZN(n11591) );
  AOI22_X1 U11770 ( .A1(n11958), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11767) );
  BUF_X2 U11771 ( .A(n11980), .Z(n11985) );
  OR2_X2 U11772 ( .A1(n12116), .A2(n12098), .ZN(n12092) );
  AND2_X1 U11773 ( .A1(n12116), .A2(n11449), .ZN(n12111) );
  NOR2_X1 U11774 ( .A1(n19029), .A2(n19276), .ZN(n11449) );
  AND2_X1 U11775 ( .A1(n12098), .A2(n19029), .ZN(n12096) );
  NAND2_X1 U11776 ( .A1(n11980), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11291) );
  AND2_X1 U11777 ( .A1(n11290), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11292) );
  AND2_X1 U11778 ( .A1(n11989), .A2(n11777), .ZN(n11990) );
  INV_X1 U11779 ( .A(n12023), .ZN(n11294) );
  NAND2_X1 U11780 ( .A1(n11778), .A2(n11777), .ZN(n11785) );
  INV_X1 U11781 ( .A(n12026), .ZN(n14064) );
  INV_X1 U11782 ( .A(n21409), .ZN(n15747) );
  INV_X1 U11783 ( .A(n20764), .ZN(n15652) );
  NAND2_X1 U11784 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21392), .ZN(
        n15651) );
  NOR2_X1 U11785 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11304) );
  NOR2_X1 U11786 ( .A1(n18507), .A2(n18855), .ZN(n18509) );
  NOR2_X1 U11787 ( .A1(n18879), .A2(n18501), .ZN(n18502) );
  NAND2_X1 U11788 ( .A1(n18493), .A2(n11328), .ZN(n11327) );
  NAND2_X1 U11789 ( .A1(n18495), .A2(n21375), .ZN(n11328) );
  NOR2_X1 U11790 ( .A1(n21382), .A2(n11366), .ZN(n15776) );
  NOR2_X1 U11791 ( .A1(n21440), .A2(n11367), .ZN(n11366) );
  NOR2_X1 U11792 ( .A1(n21267), .A2(n19572), .ZN(n18488) );
  NOR2_X1 U11793 ( .A1(n19490), .A2(n21440), .ZN(n21438) );
  NOR2_X1 U11794 ( .A1(n11367), .A2(n21267), .ZN(n15743) );
  NOR2_X1 U11795 ( .A1(n21433), .A2(n19490), .ZN(n21439) );
  NOR3_X1 U11796 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n21888), .A3(
        n15652), .ZN(n15715) );
  INV_X1 U11797 ( .A(n13218), .ZN(n11609) );
  NAND2_X1 U11798 ( .A1(n16102), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15196) );
  NOR3_X1 U11799 ( .A1(n15982), .A2(n11467), .A3(n11465), .ZN(n11462) );
  INV_X1 U11800 ( .A(n15916), .ZN(n11465) );
  AND2_X1 U11801 ( .A1(n11467), .A2(n14313), .ZN(n11464) );
  INV_X1 U11802 ( .A(n14226), .ZN(n14327) );
  NOR2_X1 U11803 ( .A1(n11618), .A2(n16573), .ZN(n14696) );
  AND2_X1 U11804 ( .A1(n14885), .A2(n17463), .ZN(n20463) );
  NAND2_X1 U11805 ( .A1(n22484), .A2(n14884), .ZN(n14885) );
  NOR2_X1 U11806 ( .A1(n14628), .A2(n22605), .ZN(n13293) );
  INV_X1 U11807 ( .A(n11639), .ZN(n11636) );
  OR2_X1 U11808 ( .A1(n13776), .A2(n15972), .ZN(n13799) );
  NAND2_X1 U11809 ( .A1(n13733), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13734) );
  INV_X1 U11810 ( .A(n13732), .ZN(n13733) );
  AND2_X1 U11811 ( .A1(n13737), .A2(n13736), .ZN(n15994) );
  NAND2_X1 U11812 ( .A1(n13645), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13690) );
  NOR2_X1 U11813 ( .A1(n15618), .A2(n11634), .ZN(n16217) );
  NAND2_X1 U11814 ( .A1(n11633), .A2(n13544), .ZN(n16135) );
  NAND2_X1 U11815 ( .A1(n13449), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13466) );
  INV_X1 U11816 ( .A(n15254), .ZN(n11621) );
  NAND2_X1 U11817 ( .A1(n20588), .A2(n11426), .ZN(n11424) );
  INV_X1 U11818 ( .A(n11421), .ZN(n11425) );
  AND3_X1 U11819 ( .A1(n13429), .A2(n13428), .A3(n13427), .ZN(n15300) );
  INV_X1 U11820 ( .A(n14949), .ZN(n13361) );
  INV_X1 U11821 ( .A(n14736), .ZN(n13362) );
  NAND2_X1 U11822 ( .A1(n14663), .A2(n13301), .ZN(n14738) );
  NOR2_X1 U11823 ( .A1(n11655), .A2(n11660), .ZN(n11654) );
  INV_X1 U11824 ( .A(n11656), .ZN(n11655) );
  NAND2_X1 U11825 ( .A1(n15840), .A2(n15839), .ZN(n11660) );
  NAND2_X1 U11826 ( .A1(n11651), .A2(n20617), .ZN(n11650) );
  INV_X1 U11827 ( .A(n11661), .ZN(n11651) );
  OR2_X1 U11828 ( .A1(n22289), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13914) );
  XNOR2_X1 U11829 ( .A(n13994), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16390) );
  NOR2_X1 U11830 ( .A1(n20594), .A2(n11423), .ZN(n11426) );
  INV_X1 U11831 ( .A(n13974), .ZN(n11423) );
  OR2_X1 U11832 ( .A1(n20588), .A2(n20587), .ZN(n20590) );
  AND4_X1 U11833 ( .A1(n13148), .A2(n13147), .A3(n13146), .A4(n13145), .ZN(
        n13154) );
  CLKBUF_X1 U11834 ( .A(n14672), .Z(n14673) );
  NOR2_X1 U11835 ( .A1(n22544), .A2(n16592), .ZN(n22595) );
  NOR2_X1 U11836 ( .A1(n14673), .A2(n17397), .ZN(n22604) );
  INV_X1 U11837 ( .A(n22501), .ZN(n22583) );
  AOI21_X1 U11838 ( .B1(n22571), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n16592), 
        .ZN(n22613) );
  NAND2_X1 U11839 ( .A1(n13893), .A2(n13868), .ZN(n13908) );
  NAND2_X1 U11840 ( .A1(n13906), .A2(n13905), .ZN(n13907) );
  INV_X1 U11841 ( .A(n14414), .ZN(n13868) );
  INV_X1 U11842 ( .A(n11252), .ZN(n11459) );
  NOR2_X1 U11843 ( .A1(n12301), .A2(n11455), .ZN(n11454) );
  INV_X1 U11844 ( .A(n12286), .ZN(n11455) );
  NOR2_X1 U11845 ( .A1(n14065), .A2(n12469), .ZN(n12277) );
  INV_X1 U11846 ( .A(n12031), .ZN(n15383) );
  NAND2_X1 U11847 ( .A1(n11688), .A2(n11690), .ZN(n12055) );
  INV_X1 U11848 ( .A(n11689), .ZN(n11688) );
  OR2_X1 U11849 ( .A1(n12624), .A2(n14982), .ZN(n14983) );
  AND2_X1 U11850 ( .A1(n14160), .A2(n14161), .ZN(n15808) );
  AND2_X1 U11851 ( .A1(n12916), .A2(n11674), .ZN(n11672) );
  NAND2_X1 U11852 ( .A1(n11713), .A2(n11586), .ZN(n15639) );
  AND2_X1 U11853 ( .A1(n11588), .A2(n11587), .ZN(n11586) );
  INV_X1 U11854 ( .A(n15598), .ZN(n11587) );
  NAND2_X1 U11855 ( .A1(n11713), .A2(n11588), .ZN(n16799) );
  NOR2_X1 U11856 ( .A1(n12011), .A2(n12013), .ZN(n15602) );
  NOR2_X1 U11857 ( .A1(n17299), .A2(n14746), .ZN(n15446) );
  AND2_X1 U11858 ( .A1(n14478), .A2(n22356), .ZN(n17915) );
  INV_X1 U11859 ( .A(n14371), .ZN(n15596) );
  INV_X1 U11860 ( .A(n15863), .ZN(n11528) );
  XNOR2_X1 U11861 ( .A(n12432), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17864) );
  AND2_X1 U11862 ( .A1(n12040), .A2(n12039), .ZN(n12041) );
  XNOR2_X1 U11863 ( .A(n16828), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14061) );
  AND2_X1 U11864 ( .A1(n11181), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11374) );
  AND2_X1 U11865 ( .A1(n12323), .A2(n11448), .ZN(n11446) );
  INV_X1 U11866 ( .A(n11706), .ZN(n11448) );
  NAND2_X1 U11867 ( .A1(n11362), .A2(n11360), .ZN(n11359) );
  INV_X1 U11868 ( .A(n16900), .ZN(n11360) );
  OR2_X1 U11869 ( .A1(n16652), .A2(n12203), .ZN(n16898) );
  AND2_X1 U11870 ( .A1(n19111), .A2(n12330), .ZN(n16936) );
  NAND2_X1 U11871 ( .A1(n16948), .A2(n16947), .ZN(n16949) );
  AND2_X1 U11872 ( .A1(n11713), .A2(n15001), .ZN(n16807) );
  AND3_X1 U11873 ( .A1(n14134), .A2(n14133), .A3(n14132), .ZN(n15550) );
  AND3_X1 U11874 ( .A1(n14122), .A2(n14121), .A3(n14120), .ZN(n17297) );
  AOI21_X1 U11875 ( .B1(n11697), .B2(n11701), .A(n11340), .ZN(n11339) );
  INV_X1 U11876 ( .A(n11697), .ZN(n11341) );
  INV_X1 U11877 ( .A(n17026), .ZN(n11340) );
  AOI21_X1 U11878 ( .B1(n11700), .B2(n11702), .A(n11698), .ZN(n11697) );
  INV_X1 U11879 ( .A(n17868), .ZN(n11698) );
  NAND2_X1 U11880 ( .A1(n12563), .A2(n12562), .ZN(n14473) );
  OR2_X1 U11881 ( .A1(n15076), .A2(n12560), .ZN(n12563) );
  NOR2_X1 U11882 ( .A1(n14064), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14470) );
  XNOR2_X1 U11883 ( .A(n14473), .B(n12567), .ZN(n14485) );
  AOI21_X1 U11884 ( .B1(n19029), .B2(n15124), .A(n12566), .ZN(n14484) );
  NAND2_X1 U11885 ( .A1(n14485), .A2(n14484), .ZN(n14483) );
  CLKBUF_X1 U11886 ( .A(n14041), .Z(n14042) );
  BUF_X1 U11887 ( .A(n12188), .Z(n19976) );
  AND2_X1 U11888 ( .A1(n19941), .A2(n19940), .ZN(n19998) );
  INV_X1 U11889 ( .A(n19920), .ZN(n19971) );
  AND2_X1 U11890 ( .A1(n19842), .A2(n19836), .ZN(n19942) );
  NOR2_X1 U11891 ( .A1(n12098), .A2(n17372), .ZN(n12099) );
  AND2_X1 U11892 ( .A1(n15041), .A2(n15040), .ZN(n20291) );
  INV_X1 U11893 ( .A(n15039), .ZN(n15040) );
  NAND2_X1 U11894 ( .A1(n19320), .A2(n19322), .ZN(n15041) );
  OR2_X1 U11895 ( .A1(n13020), .A2(n12382), .ZN(n15115) );
  OAI21_X1 U11896 ( .B1(n15761), .B2(n18486), .A(n15766), .ZN(n21881) );
  OR2_X1 U11897 ( .A1(n15658), .A2(n15657), .ZN(n21255) );
  INV_X1 U11898 ( .A(n11190), .ZN(n18454) );
  INV_X1 U11899 ( .A(n21398), .ZN(n15645) );
  NOR2_X1 U11900 ( .A1(n20711), .A2(n18491), .ZN(n21194) );
  OAI21_X1 U11901 ( .B1(n17985), .B2(n17984), .A(n21932), .ZN(n21191) );
  XNOR2_X1 U11902 ( .A(n18502), .B(n21506), .ZN(n18871) );
  NOR2_X1 U11903 ( .A1(n18871), .A2(n18870), .ZN(n18869) );
  OAI21_X1 U11904 ( .B1(n21682), .B2(n21885), .A(n11320), .ZN(n21705) );
  OR2_X1 U11905 ( .A1(n21683), .A2(n21784), .ZN(n11320) );
  NAND2_X1 U11906 ( .A1(n21879), .A2(n15740), .ZN(n18490) );
  AOI21_X1 U11907 ( .B1(n18518), .B2(n18517), .A(n18516), .ZN(n18820) );
  NAND2_X1 U11908 ( .A1(n11326), .A2(n18836), .ZN(n18516) );
  NAND2_X1 U11909 ( .A1(n18835), .A2(n11321), .ZN(n11326) );
  NOR2_X1 U11910 ( .A1(n18518), .A2(n11322), .ZN(n11321) );
  NAND3_X1 U11911 ( .A1(n18374), .A2(n18373), .A3(n18372), .ZN(n21450) );
  NAND2_X1 U11912 ( .A1(n18831), .A2(n18483), .ZN(n18817) );
  NAND2_X1 U11913 ( .A1(n21434), .A2(n21435), .ZN(n21432) );
  NOR2_X2 U11914 ( .A1(n21432), .A2(n21831), .ZN(n21883) );
  INV_X1 U11915 ( .A(n21255), .ZN(n21433) );
  NOR2_X1 U11916 ( .A1(n15678), .A2(n15677), .ZN(n21442) );
  CLKBUF_X1 U11917 ( .A(n14371), .Z(n15601) );
  INV_X1 U11918 ( .A(n22303), .ZN(n15163) );
  AND2_X1 U11919 ( .A1(n16102), .A2(n15174), .ZN(n22256) );
  AND2_X1 U11920 ( .A1(n16231), .A2(n14634), .ZN(n16225) );
  XNOR2_X1 U11921 ( .A(n15942), .B(n11638), .ZN(n15932) );
  NOR2_X2 U11922 ( .A1(n20628), .A2(n14579), .ZN(n20625) );
  XNOR2_X1 U11923 ( .A(n11279), .B(n16403), .ZN(n16429) );
  OAI21_X1 U11924 ( .B1(n16274), .B2(n16430), .A(n20603), .ZN(n11280) );
  NAND2_X1 U11925 ( .A1(n11282), .A2(n16414), .ZN(n11281) );
  OAI21_X1 U11926 ( .B1(n11383), .B2(n17635), .A(n17634), .ZN(n11382) );
  AOI211_X1 U11927 ( .C1(n11385), .C2(n11384), .A(n17630), .B(n17631), .ZN(
        n11383) );
  OAI211_X1 U11928 ( .C1(n15137), .C2(n13173), .A(n15132), .B(n22507), .ZN(
        n17837) );
  INV_X1 U11929 ( .A(n22669), .ZN(n22663) );
  OR2_X1 U11930 ( .A1(n14785), .A2(n11155), .ZN(n22591) );
  NOR2_X1 U11931 ( .A1(n16592), .A2(n22398), .ZN(n22669) );
  AND2_X1 U11932 ( .A1(n15399), .A2(n15591), .ZN(n19012) );
  NAND2_X1 U11933 ( .A1(n19252), .A2(n19251), .ZN(n19259) );
  AND2_X1 U11934 ( .A1(n11157), .A2(n11219), .ZN(n19131) );
  AND2_X1 U11935 ( .A1(n11227), .A2(n15365), .ZN(n11679) );
  INV_X1 U11936 ( .A(n19029), .ZN(n17372) );
  INV_X1 U11937 ( .A(n11380), .ZN(n11379) );
  NAND2_X1 U11938 ( .A1(n17064), .A2(n19292), .ZN(n11381) );
  AND2_X1 U11939 ( .A1(n11571), .A2(n11238), .ZN(n11570) );
  OR2_X1 U11940 ( .A1(n17066), .A2(n17065), .ZN(n11571) );
  XNOR2_X1 U11941 ( .A(n11436), .B(n11199), .ZN(n17071) );
  NAND2_X1 U11942 ( .A1(n11694), .A2(n11437), .ZN(n11436) );
  NOR2_X1 U11943 ( .A1(n16900), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11357) );
  INV_X1 U11944 ( .A(n11362), .ZN(n11358) );
  NOR2_X1 U11945 ( .A1(n11359), .A2(n17351), .ZN(n11354) );
  NOR2_X1 U11946 ( .A1(n11335), .A2(n19302), .ZN(n11333) );
  INV_X1 U11947 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19987) );
  INV_X1 U11948 ( .A(n19836), .ZN(n19825) );
  INV_X1 U11949 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19985) );
  INV_X1 U11950 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19871) );
  INV_X1 U11951 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19975) );
  NAND2_X1 U11952 ( .A1(n19960), .A2(n19940), .ZN(n19885) );
  INV_X1 U11953 ( .A(n21450), .ZN(n21728) );
  NOR2_X1 U11954 ( .A1(n18594), .A2(n21630), .ZN(n18667) );
  NAND3_X1 U11955 ( .A1(n22314), .A2(n18911), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n18759) );
  NOR2_X2 U11956 ( .A1(n21728), .A2(n18914), .ZN(n18812) );
  NAND2_X1 U11957 ( .A1(n21742), .A2(n21841), .ZN(n21744) );
  OAI21_X1 U11958 ( .B1(n21740), .B2(n21741), .A(n11300), .ZN(n21742) );
  OR2_X1 U11959 ( .A1(n21739), .A2(n21738), .ZN(n11300) );
  NAND2_X1 U11960 ( .A1(n21456), .A2(n21689), .ZN(n21666) );
  INV_X1 U11961 ( .A(keyinput_4), .ZN(n11524) );
  INV_X1 U11962 ( .A(keyinput_132), .ZN(n11409) );
  AOI21_X1 U11963 ( .B1(n11522), .B2(n11230), .A(n11521), .ZN(n17659) );
  NAND2_X1 U11964 ( .A1(n17684), .A2(keyinput_22), .ZN(n11499) );
  NAND2_X1 U11965 ( .A1(n17685), .A2(DATAI_10_), .ZN(n11498) );
  AOI21_X1 U11966 ( .B1(n11407), .B2(n11226), .A(n11406), .ZN(n17503) );
  AOI21_X1 U11967 ( .B1(n11501), .B2(n11500), .A(n11497), .ZN(n11496) );
  NAND2_X1 U11968 ( .A1(n11499), .A2(n11498), .ZN(n11497) );
  NOR2_X1 U11969 ( .A1(n17681), .A2(n17680), .ZN(n11500) );
  NAND2_X1 U11970 ( .A1(n17682), .A2(n17683), .ZN(n11501) );
  INV_X1 U11971 ( .A(n11495), .ZN(n11494) );
  OAI21_X1 U11972 ( .B1(n17687), .B2(keyinput_25), .A(n17686), .ZN(n11495) );
  NAND2_X1 U11973 ( .A1(n11405), .A2(n11404), .ZN(n11403) );
  NOR2_X1 U11974 ( .A1(n17518), .A2(n17517), .ZN(n11404) );
  NAND2_X1 U11975 ( .A1(n17519), .A2(n17520), .ZN(n11405) );
  AND2_X1 U11976 ( .A1(n11402), .A2(n11401), .ZN(n11400) );
  NAND2_X1 U11977 ( .A1(n17521), .A2(DATAI_10_), .ZN(n11401) );
  NAND2_X1 U11978 ( .A1(n17684), .A2(keyinput_150), .ZN(n11402) );
  INV_X1 U11979 ( .A(n17698), .ZN(n17709) );
  AOI21_X1 U11980 ( .B1(n11399), .B2(n11398), .A(n11397), .ZN(n17523) );
  XNOR2_X1 U11981 ( .A(DATAI_7_), .B(keyinput_153), .ZN(n11397) );
  INV_X1 U11982 ( .A(n17522), .ZN(n11398) );
  NAND2_X1 U11983 ( .A1(n11403), .A2(n11400), .ZN(n11399) );
  AOI211_X1 U11984 ( .C1(n11504), .C2(n11502), .A(n17722), .B(n11249), .ZN(
        n17724) );
  XNOR2_X1 U11985 ( .A(n17717), .B(n11503), .ZN(n11502) );
  AOI211_X1 U11986 ( .C1(n11394), .C2(n11392), .A(n17553), .B(n11248), .ZN(
        n17556) );
  NAND2_X1 U11987 ( .A1(n11520), .A2(n11247), .ZN(n11517) );
  NAND2_X1 U11988 ( .A1(n17740), .A2(n17741), .ZN(n11520) );
  INV_X1 U11989 ( .A(n17739), .ZN(n11518) );
  NOR2_X1 U11990 ( .A1(n17748), .A2(n17747), .ZN(n11516) );
  INV_X1 U11991 ( .A(n17569), .ZN(n11415) );
  NAND2_X1 U11992 ( .A1(n11515), .A2(n11513), .ZN(n17757) );
  NOR2_X1 U11993 ( .A1(n17752), .A2(n11514), .ZN(n11513) );
  NAND2_X1 U11994 ( .A1(n11517), .A2(n11516), .ZN(n11515) );
  XNOR2_X1 U11995 ( .A(P1_REIP_REG_12__SCAN_IN), .B(keyinput_71), .ZN(n11514)
         );
  NAND2_X1 U11996 ( .A1(n11417), .A2(n11259), .ZN(n11414) );
  NAND2_X1 U11997 ( .A1(n17570), .A2(n17571), .ZN(n11417) );
  NOR2_X1 U11998 ( .A1(n17576), .A2(n17575), .ZN(n11413) );
  NAND2_X1 U11999 ( .A1(n11391), .A2(n17592), .ZN(n11390) );
  OAI21_X1 U12000 ( .B1(n17589), .B2(n17588), .A(n17587), .ZN(n11391) );
  NOR2_X1 U12001 ( .A1(n17591), .A2(n11262), .ZN(n11389) );
  NAND2_X1 U12002 ( .A1(keyinput_100), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n11510) );
  OR2_X1 U12003 ( .A1(n13229), .A2(n13228), .ZN(n13926) );
  NAND2_X1 U12004 ( .A1(n11645), .A2(n13219), .ZN(n11644) );
  AND2_X1 U12005 ( .A1(n15210), .A2(n17473), .ZN(n11645) );
  AOI21_X1 U12006 ( .B1(n11388), .B2(n11387), .A(n11386), .ZN(n17603) );
  XNOR2_X1 U12007 ( .A(n17594), .B(keyinput_215), .ZN(n11386) );
  INV_X1 U12008 ( .A(n17593), .ZN(n11387) );
  NAND2_X1 U12009 ( .A1(n11390), .A2(n11389), .ZN(n11388) );
  NAND2_X1 U12010 ( .A1(n11511), .A2(n11508), .ZN(n11507) );
  AND2_X1 U12011 ( .A1(n17795), .A2(n11509), .ZN(n11508) );
  INV_X1 U12012 ( .A(n17791), .ZN(n11511) );
  AND2_X1 U12013 ( .A1(n17796), .A2(n11510), .ZN(n11509) );
  NAND2_X1 U12014 ( .A1(n11145), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11483) );
  NAND2_X1 U12015 ( .A1(n19878), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11482) );
  NAND2_X1 U12016 ( .A1(n11299), .A2(n11298), .ZN(n12115) );
  NAND2_X1 U12017 ( .A1(n19930), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11299) );
  NAND2_X1 U12018 ( .A1(n19950), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11298) );
  NAND2_X1 U12019 ( .A1(n12571), .A2(n12005), .ZN(n11976) );
  INV_X1 U12020 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11418) );
  CLKBUF_X1 U12021 ( .A(n13437), .Z(n13827) );
  CLKBUF_X1 U12022 ( .A(n13593), .Z(n13834) );
  OR2_X1 U12023 ( .A1(n13375), .A2(n13374), .ZN(n13967) );
  INV_X1 U12025 ( .A(n13215), .ZN(n13937) );
  NAND2_X1 U12026 ( .A1(n14804), .A2(n14817), .ZN(n11420) );
  OAI21_X1 U12027 ( .B1(n11512), .B2(n11507), .A(n17799), .ZN(n17800) );
  NAND2_X1 U12028 ( .A1(n13899), .A2(n13975), .ZN(n13901) );
  OR2_X1 U12029 ( .A1(n14886), .A2(n17473), .ZN(n13313) );
  NOR2_X1 U12030 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12820) );
  AOI22_X1 U12031 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U12032 ( .A1(n12466), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11669) );
  NAND2_X1 U12033 ( .A1(n11704), .A2(n11706), .ZN(n11703) );
  NAND2_X1 U12034 ( .A1(n12259), .A2(n12258), .ZN(n12425) );
  OR2_X1 U12035 ( .A1(n12256), .A2(n12255), .ZN(n12259) );
  XNOR2_X1 U12036 ( .A(n12426), .B(n11687), .ZN(n12414) );
  INV_X1 U12037 ( .A(n12425), .ZN(n11687) );
  INV_X1 U12038 ( .A(n12407), .ZN(n11492) );
  AND3_X1 U12039 ( .A1(n11769), .A2(n11768), .A3(n11777), .ZN(n11593) );
  NAND2_X1 U12040 ( .A1(n12121), .A2(n12110), .ZN(n12177) );
  INV_X1 U12041 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11744) );
  NAND2_X1 U12042 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U12043 ( .A1(n11377), .A2(n11434), .ZN(n11955) );
  AOI22_X1 U12044 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11918) );
  NAND2_X1 U12045 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U12046 ( .A1(n11830), .A2(n11829), .ZN(n11831) );
  XNOR2_X1 U12047 ( .A(n11777), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11832) );
  AOI21_X1 U12048 ( .B1(n21895), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n15750), .ZN(n15756) );
  NAND2_X1 U12049 ( .A1(n14825), .A2(n13275), .ZN(n14215) );
  NOR2_X1 U12050 ( .A1(n11617), .A2(n11206), .ZN(n11616) );
  AND2_X1 U12051 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11617) );
  AND2_X1 U12052 ( .A1(n15936), .A2(n15167), .ZN(n13850) );
  INV_X1 U12053 ( .A(n13995), .ZN(n11668) );
  NAND2_X1 U12054 ( .A1(n20587), .A2(n13974), .ZN(n11422) );
  AND2_X1 U12055 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13326), .ZN(
        n13353) );
  INV_X1 U12056 ( .A(n13984), .ZN(n13975) );
  NAND2_X1 U12057 ( .A1(n11479), .A2(n14307), .ZN(n11478) );
  INV_X1 U12058 ( .A(n11480), .ZN(n11479) );
  NAND2_X1 U12059 ( .A1(n20604), .A2(n13995), .ZN(n16363) );
  NOR2_X1 U12060 ( .A1(n20552), .A2(n15258), .ZN(n11472) );
  NOR2_X1 U12061 ( .A1(n13140), .A2(n11717), .ZN(n13141) );
  NAND2_X1 U12062 ( .A1(n14224), .A2(n14223), .ZN(n14229) );
  OR2_X1 U12063 ( .A1(n14797), .A2(n14825), .ZN(n13984) );
  OAI211_X1 U12064 ( .C1(n13192), .C2(n14797), .A(n13191), .B(n14541), .ZN(
        n13250) );
  AND3_X1 U12065 ( .A1(n13190), .A2(n13189), .A3(n14544), .ZN(n13191) );
  INV_X1 U12066 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14727) );
  NAND2_X1 U12067 ( .A1(n13202), .A2(n11613), .ZN(n11612) );
  AND2_X1 U12068 ( .A1(n13307), .A2(n13199), .ZN(n15135) );
  OR2_X1 U12069 ( .A1(n13324), .A2(n13323), .ZN(n13949) );
  OR2_X1 U12070 ( .A1(n13901), .A2(n14414), .ZN(n13906) );
  NAND2_X1 U12071 ( .A1(n13314), .A2(n13313), .ZN(n13893) );
  XNOR2_X1 U12072 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12999) );
  NAND2_X1 U12073 ( .A1(n12366), .A2(n12365), .ZN(n12371) );
  NOR2_X1 U12074 ( .A1(n12325), .A2(n11461), .ZN(n11460) );
  AND2_X1 U12075 ( .A1(n12206), .A2(n12205), .ZN(n12262) );
  AND2_X1 U12076 ( .A1(n12217), .A2(n12221), .ZN(n12220) );
  NAND2_X1 U12077 ( .A1(n16685), .A2(n11712), .ZN(n12913) );
  NAND2_X1 U12078 ( .A1(n11525), .A2(n11744), .ZN(n12972) );
  NAND2_X1 U12079 ( .A1(n16779), .A2(n16769), .ZN(n11575) );
  NOR2_X1 U12080 ( .A1(n15639), .A2(n15637), .ZN(n16644) );
  AND2_X1 U12081 ( .A1(n15594), .A2(n15636), .ZN(n11685) );
  NOR2_X1 U12082 ( .A1(n16872), .A2(n11556), .ZN(n11555) );
  NAND2_X1 U12083 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11551) );
  NOR2_X1 U12084 ( .A1(n15020), .A2(n11534), .ZN(n11533) );
  INV_X1 U12085 ( .A(n15203), .ZN(n11534) );
  NAND2_X1 U12086 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  NAND2_X1 U12087 ( .A1(n12010), .A2(n12048), .ZN(n12065) );
  AND2_X1 U12088 ( .A1(n11547), .A2(n11546), .ZN(n11545) );
  INV_X1 U12089 ( .A(n16682), .ZN(n11546) );
  NOR2_X1 U12090 ( .A1(n19216), .A2(n12203), .ZN(n14017) );
  AND2_X1 U12091 ( .A1(n16695), .A2(n16688), .ZN(n11547) );
  NOR2_X1 U12092 ( .A1(n11604), .A2(n17158), .ZN(n11603) );
  NOR2_X1 U12093 ( .A1(n11148), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11706) );
  INV_X1 U12094 ( .A(n16915), .ZN(n11487) );
  AND2_X1 U12095 ( .A1(n11486), .A2(n11344), .ZN(n11343) );
  NAND2_X1 U12096 ( .A1(n11347), .A2(n11345), .ZN(n11344) );
  AND2_X1 U12097 ( .A1(n11489), .A2(n16937), .ZN(n11486) );
  INV_X1 U12098 ( .A(n16947), .ZN(n11345) );
  INV_X1 U12099 ( .A(n16897), .ZN(n11489) );
  NAND2_X1 U12100 ( .A1(n11260), .A2(n11605), .ZN(n11604) );
  NOR2_X1 U12101 ( .A1(n16936), .A2(n11348), .ZN(n11347) );
  INV_X1 U12102 ( .A(n16895), .ZN(n11348) );
  NOR2_X1 U12103 ( .A1(n11532), .A2(n11531), .ZN(n11530) );
  INV_X1 U12104 ( .A(n15328), .ZN(n11531) );
  INV_X1 U12105 ( .A(n11533), .ZN(n11532) );
  AND2_X1 U12106 ( .A1(n15001), .A2(n16806), .ZN(n11590) );
  XNOR2_X1 U12107 ( .A(n12430), .B(n12203), .ZN(n12427) );
  NAND2_X1 U12108 ( .A1(n11297), .A2(n11207), .ZN(n12420) );
  INV_X1 U12109 ( .A(n12417), .ZN(n11297) );
  NAND2_X1 U12110 ( .A1(n11216), .A2(n12408), .ZN(n11594) );
  NAND4_X1 U12111 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n14089) );
  AOI21_X1 U12112 ( .B1(n14365), .B2(n14173), .A(n11266), .ZN(n14176) );
  NAND2_X1 U12113 ( .A1(n12121), .A2(n12098), .ZN(n12239) );
  INV_X1 U12114 ( .A(n19940), .ZN(n17897) );
  AND2_X1 U12115 ( .A1(n15127), .A2(n19016), .ZN(n15039) );
  INV_X1 U12116 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12214) );
  AND2_X1 U12117 ( .A1(n19987), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12381) );
  NAND2_X1 U12118 ( .A1(n21888), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15650) );
  OR2_X1 U12119 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15748), .ZN(
        n18086) );
  OR2_X1 U12120 ( .A1(n21385), .A2(n15748), .ZN(n11184) );
  NOR2_X1 U12121 ( .A1(n18714), .A2(n11314), .ZN(n11313) );
  NOR2_X1 U12122 ( .A1(n18631), .A2(n21061), .ZN(n18651) );
  OR2_X1 U12123 ( .A1(n18817), .A2(n18721), .ZN(n18550) );
  NAND2_X1 U12124 ( .A1(n18835), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18517) );
  INV_X1 U12125 ( .A(n18493), .ZN(n18494) );
  NOR2_X1 U12126 ( .A1(n21433), .A2(n21254), .ZN(n15772) );
  NOR2_X1 U12127 ( .A1(n21442), .A2(n21255), .ZN(n21396) );
  NOR2_X1 U12128 ( .A1(n21440), .A2(n15742), .ZN(n21395) );
  NAND2_X1 U12129 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21411) );
  NAND2_X1 U12130 ( .A1(n11319), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n21418) );
  INV_X1 U12131 ( .A(n15650), .ZN(n11319) );
  NAND3_X1 U12132 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15748) );
  INV_X1 U12133 ( .A(n14625), .ZN(n14883) );
  NAND2_X1 U12134 ( .A1(n13528), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13545) );
  NAND2_X1 U12135 ( .A1(n11468), .A2(n15944), .ZN(n11467) );
  INV_X1 U12136 ( .A(n11468), .ZN(n11466) );
  AOI21_X1 U12137 ( .B1(n14573), .B2(n14222), .A(n14229), .ZN(n14668) );
  INV_X1 U12138 ( .A(n16243), .ZN(n16209) );
  AND2_X1 U12139 ( .A1(n22605), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n15818) );
  NOR2_X1 U12140 ( .A1(n11639), .A2(n11638), .ZN(n11637) );
  NOR2_X1 U12141 ( .A1(n13799), .A2(n16252), .ZN(n13800) );
  AOI21_X1 U12142 ( .B1(n13798), .B2(n13797), .A(n13796), .ZN(n15954) );
  AND2_X1 U12143 ( .A1(n16254), .A2(n15167), .ZN(n13796) );
  NAND2_X1 U12144 ( .A1(n13779), .A2(n13778), .ZN(n15971) );
  OR2_X1 U12145 ( .A1(n16270), .A2(n13847), .ZN(n13778) );
  AND2_X1 U12146 ( .A1(n16298), .A2(n15167), .ZN(n13713) );
  NAND2_X1 U12147 ( .A1(n13691), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13693) );
  INV_X1 U12148 ( .A(n13690), .ZN(n13691) );
  OR2_X1 U12149 ( .A1(n16303), .A2(n13847), .ZN(n13695) );
  AND2_X1 U12150 ( .A1(n13649), .A2(n13648), .ZN(n16046) );
  AND2_X1 U12151 ( .A1(n16334), .A2(n15167), .ZN(n13626) );
  CLKBUF_X1 U12152 ( .A(n16044), .Z(n16045) );
  AND2_X1 U12153 ( .A1(n13608), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13609) );
  CLKBUF_X1 U12154 ( .A(n16070), .Z(n16123) );
  NOR2_X1 U12155 ( .A1(n13574), .A2(n22247), .ZN(n13608) );
  INV_X1 U12156 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n22247) );
  AND2_X1 U12157 ( .A1(n13496), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13528) );
  INV_X1 U12158 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13511) );
  AND2_X1 U12159 ( .A1(n16235), .A2(n16236), .ZN(n16237) );
  NOR2_X1 U12160 ( .A1(n13466), .A2(n13465), .ZN(n13467) );
  NAND2_X1 U12161 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n13467), .ZN(
        n13510) );
  CLKBUF_X1 U12162 ( .A(n15370), .Z(n15371) );
  INV_X1 U12163 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13431) );
  INV_X1 U12164 ( .A(n15036), .ZN(n13401) );
  INV_X1 U12165 ( .A(n15297), .ZN(n13402) );
  OAI21_X1 U12166 ( .B1(n13412), .B2(n13411), .A(n13410), .ZN(n13413) );
  INV_X1 U12167 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n22153) );
  NOR2_X1 U12168 ( .A1(n13396), .A2(n22153), .ZN(n13409) );
  NAND2_X1 U12169 ( .A1(n13397), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13396) );
  AOI21_X1 U12170 ( .B1(n13948), .B2(n13537), .A(n13360), .ZN(n14949) );
  NAND2_X1 U12171 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13327) );
  CLKBUF_X1 U12172 ( .A(n14736), .Z(n14950) );
  INV_X1 U12173 ( .A(n14661), .ZN(n13299) );
  INV_X1 U12174 ( .A(n14660), .ZN(n13300) );
  NAND2_X1 U12175 ( .A1(n20603), .A2(n16430), .ZN(n11659) );
  AND2_X1 U12176 ( .A1(n14320), .A2(n14319), .ZN(n15966) );
  NOR2_X1 U12177 ( .A1(n15982), .A2(n15966), .ZN(n15965) );
  NOR2_X1 U12178 ( .A1(n16062), .A2(n11480), .ZN(n16035) );
  INV_X1 U12179 ( .A(n22045), .ZN(n16532) );
  AND2_X1 U12180 ( .A1(n14297), .A2(n14296), .ZN(n16048) );
  NOR2_X1 U12181 ( .A1(n16062), .A2(n16048), .ZN(n16047) );
  NAND2_X1 U12182 ( .A1(n11474), .A2(n16125), .ZN(n11473) );
  INV_X1 U12183 ( .A(n11476), .ZN(n11474) );
  NOR2_X1 U12184 ( .A1(n16139), .A2(n11476), .ZN(n16126) );
  AND2_X1 U12185 ( .A1(n14285), .A2(n14284), .ZN(n20566) );
  NOR2_X1 U12186 ( .A1(n16139), .A2(n11475), .ZN(n20567) );
  INV_X1 U12187 ( .A(n11477), .ZN(n11475) );
  INV_X1 U12188 ( .A(n16363), .ZN(n20620) );
  NAND2_X1 U12189 ( .A1(n16345), .A2(n14006), .ZN(n20619) );
  NAND2_X1 U12190 ( .A1(n14222), .A2(n17481), .ZN(n14276) );
  OR2_X1 U12191 ( .A1(n16088), .A2(n15620), .ZN(n16139) );
  NOR2_X1 U12192 ( .A1(n20555), .A2(n20556), .ZN(n20554) );
  AND2_X1 U12193 ( .A1(n14264), .A2(n14263), .ZN(n15562) );
  OR2_X1 U12194 ( .A1(n20562), .A2(n15562), .ZN(n20555) );
  NAND2_X1 U12195 ( .A1(n20560), .A2(n20559), .ZN(n20562) );
  NAND2_X1 U12196 ( .A1(n14222), .A2(n14252), .ZN(n14253) );
  AND2_X1 U12197 ( .A1(n15357), .A2(n15356), .ZN(n20560) );
  AND2_X1 U12198 ( .A1(n15160), .A2(n11470), .ZN(n15357) );
  NOR2_X1 U12199 ( .A1(n11471), .A2(n15305), .ZN(n11470) );
  INV_X1 U12200 ( .A(n11472), .ZN(n11471) );
  NAND2_X1 U12201 ( .A1(n15160), .A2(n11472), .ZN(n15306) );
  NAND2_X1 U12202 ( .A1(n15160), .A2(n14244), .ZN(n20549) );
  NOR2_X1 U12203 ( .A1(n20570), .A2(n20571), .ZN(n20569) );
  NOR2_X1 U12204 ( .A1(n16407), .A2(n16532), .ZN(n21979) );
  INV_X1 U12205 ( .A(n22049), .ZN(n22005) );
  OR2_X1 U12206 ( .A1(n14740), .A2(n14741), .ZN(n20570) );
  AND2_X1 U12207 ( .A1(n14557), .A2(n14546), .ZN(n16550) );
  INV_X1 U12208 ( .A(n15902), .ZN(n13161) );
  NAND2_X1 U12209 ( .A1(n13292), .A2(n17473), .ZN(n13268) );
  OAI211_X1 U12210 ( .C1(n13891), .C2(n13271), .A(n13270), .B(n13269), .ZN(
        n13289) );
  CLKBUF_X1 U12211 ( .A(n14637), .Z(n14638) );
  OR2_X1 U12212 ( .A1(n13306), .A2(n13305), .ZN(n13312) );
  INV_X1 U12213 ( .A(n16573), .ZN(n17436) );
  AND2_X1 U12214 ( .A1(n14556), .A2(n14555), .ZN(n17439) );
  CLKBUF_X1 U12215 ( .A(n14619), .Z(n14688) );
  NAND2_X1 U12216 ( .A1(n13219), .A2(n13196), .ZN(n11611) );
  INV_X1 U12217 ( .A(n22528), .ZN(n16590) );
  OR2_X1 U12218 ( .A1(n14848), .A2(n22582), .ZN(n14851) );
  INV_X1 U12219 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22586) );
  NAND2_X1 U12220 ( .A1(n17626), .A2(n17627), .ZN(n11385) );
  NOR2_X1 U12221 ( .A1(n17624), .A2(n17625), .ZN(n11384) );
  NOR2_X1 U12222 ( .A1(n11648), .A2(n14638), .ZN(n14957) );
  NAND2_X1 U12223 ( .A1(n14638), .A2(n15213), .ZN(n22487) );
  INV_X1 U12224 ( .A(n14628), .ZN(n15908) );
  INV_X1 U12225 ( .A(n14838), .ZN(n14835) );
  INV_X1 U12226 ( .A(n21947), .ZN(n17464) );
  NOR2_X1 U12227 ( .A1(n14165), .A2(n14164), .ZN(n15101) );
  OR2_X1 U12228 ( .A1(n12371), .A2(n12370), .ZN(n15856) );
  AND2_X1 U12229 ( .A1(n12351), .A2(n12349), .ZN(n11913) );
  AND2_X1 U12230 ( .A1(n11913), .A2(n11912), .ZN(n12366) );
  NOR2_X1 U12231 ( .A1(n12357), .A2(n12355), .ZN(n12351) );
  OR2_X1 U12232 ( .A1(n12348), .A2(n12346), .ZN(n12357) );
  OR2_X1 U12233 ( .A1(n12343), .A2(n12341), .ZN(n12348) );
  OR2_X1 U12234 ( .A1(n16633), .A2(n11564), .ZN(n11562) );
  NAND2_X1 U12235 ( .A1(n16884), .A2(n11565), .ZN(n11564) );
  INV_X1 U12236 ( .A(n16905), .ZN(n11565) );
  NAND2_X1 U12237 ( .A1(n15794), .A2(n16884), .ZN(n11563) );
  XNOR2_X1 U12238 ( .A(n12328), .B(n11246), .ZN(n16629) );
  AND2_X1 U12239 ( .A1(n12296), .A2(n12294), .ZN(n12292) );
  NAND2_X1 U12240 ( .A1(n12287), .A2(n11174), .ZN(n12298) );
  NOR2_X1 U12241 ( .A1(n15442), .A2(n16999), .ZN(n15468) );
  NAND2_X1 U12242 ( .A1(n12287), .A2(n12286), .ZN(n12288) );
  AND2_X1 U12243 ( .A1(n11203), .A2(n12269), .ZN(n11456) );
  NOR2_X1 U12244 ( .A1(n14065), .A2(n12462), .ZN(n12273) );
  OR2_X1 U12245 ( .A1(n12274), .A2(n12273), .ZN(n12284) );
  AND2_X1 U12246 ( .A1(n12206), .A2(n11203), .ZN(n12271) );
  INV_X1 U12247 ( .A(n19253), .ZN(n19208) );
  AND4_X1 U12248 ( .A1(n12737), .A2(n12736), .A3(n12735), .A4(n12734), .ZN(
        n15572) );
  NOR2_X1 U12249 ( .A1(n11681), .A2(n12673), .ZN(n11680) );
  INV_X1 U12250 ( .A(n15024), .ZN(n11681) );
  NAND2_X1 U12251 ( .A1(n11581), .A2(n11579), .ZN(n11578) );
  NOR2_X1 U12252 ( .A1(n11583), .A2(n11582), .ZN(n11581) );
  AND3_X1 U12253 ( .A1(n11670), .A2(n12953), .A3(n16667), .ZN(n16656) );
  OAI21_X1 U12254 ( .B1(n16676), .B2(n11674), .A(n11671), .ZN(n11670) );
  INV_X1 U12255 ( .A(n11673), .ZN(n11671) );
  INV_X1 U12256 ( .A(n11579), .ZN(n11577) );
  NOR2_X1 U12257 ( .A1(n11162), .A2(n16757), .ZN(n16747) );
  XNOR2_X1 U12258 ( .A(n16692), .B(n12892), .ZN(n16687) );
  OAI21_X1 U12259 ( .B1(n16703), .B2(n16704), .A(n11711), .ZN(n16694) );
  NOR3_X1 U12260 ( .A1(n11161), .A2(n17143), .A3(n11576), .ZN(n16781) );
  NOR2_X1 U12261 ( .A1(n11161), .A2(n17143), .ZN(n16778) );
  AND2_X1 U12262 ( .A1(n15595), .A2(n11254), .ZN(n16717) );
  INV_X1 U12263 ( .A(n16718), .ZN(n11682) );
  NAND2_X1 U12264 ( .A1(n15595), .A2(n11683), .ZN(n16721) );
  AND2_X1 U12265 ( .A1(n14143), .A2(n14142), .ZN(n15598) );
  AND2_X1 U12266 ( .A1(n14141), .A2(n14140), .ZN(n16797) );
  AND2_X1 U12267 ( .A1(n15857), .A2(n12006), .ZN(n15604) );
  NAND2_X1 U12268 ( .A1(n14095), .A2(n11209), .ZN(n14761) );
  XNOR2_X1 U12269 ( .A(n14088), .B(n11569), .ZN(n14500) );
  INV_X1 U12270 ( .A(n14087), .ZN(n11569) );
  NAND2_X1 U12271 ( .A1(n14500), .A2(n14501), .ZN(n14503) );
  NAND2_X1 U12272 ( .A1(n14079), .A2(n14090), .ZN(n14499) );
  NOR2_X1 U12273 ( .A1(n14080), .A2(n14075), .ZN(n14076) );
  NAND2_X1 U12274 ( .A1(n15799), .A2(n11177), .ZN(n15802) );
  NAND2_X1 U12275 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11566) );
  AND2_X1 U12276 ( .A1(n15014), .A2(n11533), .ZN(n15329) );
  AND2_X1 U12277 ( .A1(n15014), .A2(n12478), .ZN(n15204) );
  NOR2_X1 U12278 ( .A1(n11542), .A2(n11541), .ZN(n11540) );
  INV_X1 U12279 ( .A(n14980), .ZN(n11541) );
  NAND2_X1 U12280 ( .A1(n11539), .A2(n12461), .ZN(n14911) );
  NOR2_X1 U12281 ( .A1(n14903), .A2(n11542), .ZN(n14981) );
  NAND2_X1 U12282 ( .A1(n11560), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11559) );
  NOR2_X1 U12283 ( .A1(n11188), .A2(n15809), .ZN(n15832) );
  NOR2_X1 U12284 ( .A1(n15854), .A2(n16814), .ZN(n11692) );
  INV_X1 U12285 ( .A(n16813), .ZN(n11695) );
  INV_X1 U12286 ( .A(n16814), .ZN(n11437) );
  AND2_X1 U12287 ( .A1(n19224), .A2(n15859), .ZN(n14019) );
  NAND2_X1 U12288 ( .A1(n16696), .A2(n11545), .ZN(n16680) );
  NAND2_X1 U12289 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17098), .ZN(
        n11601) );
  NOR2_X1 U12290 ( .A1(n16835), .A2(n16848), .ZN(n11451) );
  INV_X1 U12291 ( .A(n16834), .ZN(n11452) );
  CLKBUF_X1 U12292 ( .A(n16834), .Z(n16851) );
  AND2_X1 U12293 ( .A1(n16696), .A2(n16695), .ZN(n16697) );
  AOI21_X1 U12294 ( .B1(n11704), .B2(n16877), .A(n11442), .ZN(n11441) );
  AOI21_X1 U12295 ( .B1(n11214), .B2(n16877), .A(n11440), .ZN(n11439) );
  INV_X1 U12296 ( .A(n11443), .ZN(n11442) );
  OR3_X1 U12297 ( .A1(n12344), .A2(n12203), .A3(n14183), .ZN(n16867) );
  NAND2_X1 U12298 ( .A1(n11537), .A2(n11536), .ZN(n11535) );
  INV_X1 U12299 ( .A(n15567), .ZN(n11537) );
  NOR2_X1 U12300 ( .A1(n11538), .A2(n16728), .ZN(n11536) );
  NAND2_X1 U12301 ( .A1(n16896), .A2(n16937), .ZN(n16929) );
  NAND2_X1 U12302 ( .A1(n16949), .A2(n11347), .ZN(n16896) );
  OR3_X1 U12303 ( .A1(n12339), .A2(n12203), .A3(n17203), .ZN(n16927) );
  AND2_X1 U12304 ( .A1(n14771), .A2(n14135), .ZN(n11713) );
  NAND2_X1 U12305 ( .A1(n16986), .A2(n11260), .ZN(n16973) );
  AND3_X1 U12306 ( .A1(n14131), .A2(n14130), .A3(n14129), .ZN(n14772) );
  NOR2_X1 U12307 ( .A1(n11147), .A2(n11606), .ZN(n16987) );
  INV_X1 U12308 ( .A(n12435), .ZN(n11606) );
  OR2_X1 U12309 ( .A1(n17009), .A2(n16892), .ZN(n16994) );
  NAND2_X1 U12310 ( .A1(n11506), .A2(n17018), .ZN(n17009) );
  INV_X1 U12311 ( .A(n16891), .ZN(n11506) );
  NAND2_X1 U12312 ( .A1(n14751), .A2(n11232), .ZN(n17299) );
  INV_X1 U12313 ( .A(n17297), .ZN(n11584) );
  NAND2_X1 U12314 ( .A1(n17039), .A2(n17040), .ZN(n11699) );
  INV_X1 U12315 ( .A(n17352), .ZN(n17328) );
  NOR2_X1 U12316 ( .A1(n11165), .A2(n11574), .ZN(n11573) );
  NOR2_X1 U12317 ( .A1(n14096), .A2(n11165), .ZN(n15516) );
  INV_X1 U12318 ( .A(n11289), .ZN(n11274) );
  INV_X1 U12319 ( .A(n17326), .ZN(n17361) );
  INV_X1 U12320 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11741) );
  AND2_X1 U12321 ( .A1(n14483), .A2(n12569), .ZN(n14489) );
  AND2_X1 U12322 ( .A1(n12559), .A2(n12570), .ZN(n14490) );
  NAND2_X1 U12323 ( .A1(n14490), .A2(n14489), .ZN(n14488) );
  NAND2_X1 U12324 ( .A1(n14488), .A2(n12570), .ZN(n14566) );
  AND2_X1 U12325 ( .A1(n12573), .A2(n11678), .ZN(n14565) );
  INV_X1 U12326 ( .A(n12548), .ZN(n11676) );
  OR2_X1 U12327 ( .A1(n14039), .A2(n13021), .ZN(n15038) );
  INV_X1 U12328 ( .A(n19927), .ZN(n19997) );
  INV_X1 U12329 ( .A(n19878), .ZN(n19873) );
  NAND2_X1 U12330 ( .A1(n12111), .A2(n12098), .ZN(n12182) );
  OR2_X1 U12331 ( .A1(n19842), .A2(n19825), .ZN(n19920) );
  NAND2_X2 U12332 ( .A1(n11995), .A2(n11994), .ZN(n20206) );
  INV_X1 U12333 ( .A(n19942), .ZN(n19855) );
  NAND2_X1 U12334 ( .A1(n19842), .A2(n19825), .ZN(n19956) );
  INV_X1 U12335 ( .A(n19820), .ZN(n20297) );
  INV_X1 U12336 ( .A(n19821), .ZN(n20298) );
  NAND3_X1 U12337 ( .A1(n15601), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20005), 
        .ZN(n19820) );
  NAND3_X1 U12338 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n15596), .A3(n20005), 
        .ZN(n19821) );
  NAND2_X1 U12339 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20009), .ZN(n20293) );
  AND2_X1 U12340 ( .A1(n19322), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15124) );
  NOR2_X1 U12341 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20917), .ZN(n20927) );
  NAND2_X1 U12342 ( .A1(n20767), .A2(n11367), .ZN(n20770) );
  NAND2_X1 U12343 ( .A1(n21363), .A2(n21356), .ZN(n21350) );
  INV_X1 U12344 ( .A(n21414), .ZN(n11308) );
  NOR2_X1 U12345 ( .A1(n20712), .A2(n17407), .ZN(n18968) );
  OR2_X1 U12346 ( .A1(n20712), .A2(n22321), .ZN(n21193) );
  NOR2_X1 U12347 ( .A1(n20710), .A2(n20712), .ZN(n20714) );
  INV_X1 U12348 ( .A(n18740), .ZN(n18728) );
  NAND2_X1 U12349 ( .A1(n18728), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18727) );
  NAND2_X1 U12350 ( .A1(n18671), .A2(n11312), .ZN(n18740) );
  AND2_X1 U12351 ( .A1(n11313), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11312) );
  AND2_X1 U12352 ( .A1(n18687), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18671) );
  NAND3_X1 U12353 ( .A1(n18597), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18631) );
  NOR2_X1 U12354 ( .A1(n11318), .A2(n11317), .ZN(n11316) );
  INV_X1 U12355 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11317) );
  INV_X1 U12356 ( .A(n20979), .ZN(n18523) );
  NAND2_X1 U12357 ( .A1(n18523), .A2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18541) );
  NAND2_X1 U12358 ( .A1(n18782), .A2(n11173), .ZN(n18552) );
  NAND2_X1 U12359 ( .A1(n20981), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n20979) );
  INV_X1 U12360 ( .A(n18570), .ZN(n18715) );
  NAND2_X1 U12361 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21616), .ZN(
        n21604) );
  OR2_X1 U12362 ( .A1(n21562), .A2(n11257), .ZN(n21622) );
  NOR2_X1 U12363 ( .A1(n18582), .A2(n11310), .ZN(n11309) );
  NAND2_X1 U12364 ( .A1(n18782), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n20913) );
  AND3_X1 U12365 ( .A1(n18807), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18782) );
  NAND2_X1 U12366 ( .A1(n18874), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18858) );
  INV_X1 U12367 ( .A(n18911), .ZN(n18886) );
  INV_X1 U12368 ( .A(n11305), .ZN(n18679) );
  NAND2_X1 U12369 ( .A1(n21727), .A2(n21883), .ZN(n21740) );
  AND2_X1 U12370 ( .A1(n21729), .A2(n21783), .ZN(n21730) );
  OR2_X1 U12371 ( .A1(n18659), .A2(n18721), .ZN(n18705) );
  INV_X1 U12372 ( .A(n11306), .ZN(n18706) );
  AND2_X1 U12373 ( .A1(n21753), .A2(n21456), .ZN(n21758) );
  AND3_X1 U12374 ( .A1(n18643), .A2(n21753), .A3(n21643), .ZN(n18646) );
  NOR2_X1 U12375 ( .A1(n18660), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18659) );
  NOR2_X1 U12376 ( .A1(n18528), .A2(n18529), .ZN(n18756) );
  NAND2_X1 U12377 ( .A1(n18530), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n18527) );
  OR2_X1 U12378 ( .A1(n21562), .A2(n11245), .ZN(n21618) );
  INV_X1 U12379 ( .A(n21756), .ZN(n21784) );
  NOR2_X1 U12380 ( .A1(n18820), .A2(n21548), .ZN(n18819) );
  NAND2_X1 U12381 ( .A1(n18817), .A2(n18818), .ZN(n18816) );
  NAND2_X1 U12382 ( .A1(n11325), .A2(n11324), .ZN(n18835) );
  NOR2_X1 U12383 ( .A1(n18511), .A2(n18515), .ZN(n11324) );
  NAND2_X1 U12384 ( .A1(n11325), .A2(n11323), .ZN(n18514) );
  INV_X1 U12385 ( .A(n18511), .ZN(n11323) );
  XNOR2_X1 U12386 ( .A(n18548), .B(n18482), .ZN(n18832) );
  NAND2_X1 U12387 ( .A1(n18832), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18831) );
  NOR2_X1 U12388 ( .A1(n21448), .A2(n18846), .ZN(n18845) );
  NOR2_X1 U12389 ( .A1(n18869), .A2(n18504), .ZN(n18857) );
  NOR2_X1 U12390 ( .A1(n18857), .A2(n18856), .ZN(n18855) );
  XNOR2_X1 U12391 ( .A(n18477), .B(n18476), .ZN(n18854) );
  INV_X1 U12392 ( .A(n18475), .ZN(n18476) );
  INV_X1 U12393 ( .A(n21667), .ZN(n21886) );
  INV_X1 U12394 ( .A(n11327), .ZN(n18496) );
  XNOR2_X1 U12395 ( .A(n11327), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n18892) );
  NOR2_X1 U12396 ( .A1(n18892), .A2(n18891), .ZN(n18890) );
  INV_X1 U12397 ( .A(n18490), .ZN(n11372) );
  NOR2_X1 U12398 ( .A1(n18468), .A2(n18467), .ZN(n18909) );
  INV_X1 U12399 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21895) );
  INV_X1 U12400 ( .A(n21401), .ZN(n20777) );
  NAND2_X1 U12401 ( .A1(n21385), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n21414) );
  NAND2_X1 U12402 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n21408) );
  INV_X1 U12403 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21892) );
  INV_X1 U12404 ( .A(n21435), .ZN(n19657) );
  NOR2_X1 U12405 ( .A1(n15688), .A2(n15687), .ZN(n19572) );
  NOR2_X1 U12406 ( .A1(n15668), .A2(n15667), .ZN(n19490) );
  NOR2_X1 U12407 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19367), .ZN(n19705) );
  INV_X1 U12408 ( .A(n19705), .ZN(n19571) );
  AOI211_X1 U12409 ( .C1(n15777), .C2(n22370), .A(n17985), .B(n21444), .ZN(
        n21909) );
  NAND2_X1 U12410 ( .A1(n21783), .A2(n11369), .ZN(n11368) );
  INV_X1 U12411 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n22234) );
  INV_X1 U12412 ( .A(n22263), .ZN(n22246) );
  AND2_X1 U12413 ( .A1(n16102), .A2(n15185), .ZN(n22253) );
  AND2_X1 U12414 ( .A1(n16102), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22263) );
  INV_X1 U12415 ( .A(n22253), .ZN(n22267) );
  INV_X1 U12416 ( .A(n22214), .ZN(n22200) );
  INV_X1 U12417 ( .A(n16102), .ZN(n22190) );
  NOR2_X2 U12418 ( .A1(n15188), .A2(n15179), .ZN(n22255) );
  OR2_X1 U12419 ( .A1(n22256), .A2(n15176), .ZN(n22147) );
  XNOR2_X1 U12420 ( .A(n15920), .B(n15919), .ZN(n16396) );
  INV_X1 U12421 ( .A(n11463), .ZN(n15920) );
  INV_X1 U12422 ( .A(n16143), .ZN(n20572) );
  AND2_X2 U12423 ( .A1(n14220), .A2(n14219), .ZN(n20574) );
  OR2_X1 U12424 ( .A1(n15816), .A2(n15823), .ZN(n16227) );
  OR2_X1 U12425 ( .A1(n14627), .A2(n14626), .ZN(n16231) );
  INV_X1 U12426 ( .A(n16241), .ZN(n16233) );
  AND2_X1 U12427 ( .A1(n13774), .A2(n13735), .ZN(n16289) );
  AOI21_X1 U12428 ( .B1(n11632), .B2(n16218), .A(n16069), .ZN(n22257) );
  NAND2_X1 U12429 ( .A1(n11621), .A2(n13430), .ZN(n15354) );
  NAND2_X1 U12430 ( .A1(n11658), .A2(n11654), .ZN(n15841) );
  OR2_X1 U12431 ( .A1(n16463), .A2(n16460), .ZN(n16449) );
  OR2_X1 U12432 ( .A1(n13914), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22044) );
  NOR2_X1 U12433 ( .A1(n11431), .A2(n11430), .ZN(n16391) );
  INV_X1 U12434 ( .A(n13993), .ZN(n11430) );
  INV_X1 U12435 ( .A(n15497), .ZN(n11431) );
  NAND2_X1 U12436 ( .A1(n20590), .A2(n13974), .ZN(n20593) );
  AND2_X1 U12437 ( .A1(n14557), .A2(n17439), .ZN(n16548) );
  INV_X1 U12438 ( .A(n22084), .ZN(n22099) );
  INV_X1 U12439 ( .A(n11649), .ZN(n16568) );
  AOI21_X1 U12440 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n17473), .A(n17400), 
        .ZN(n22286) );
  NAND2_X1 U12441 ( .A1(n15214), .A2(n15213), .ZN(n22502) );
  INV_X1 U12442 ( .A(n22523), .ZN(n22797) );
  INV_X1 U12443 ( .A(n22795), .ZN(n16623) );
  INV_X1 U12444 ( .A(n16588), .ZN(n16621) );
  OAI21_X1 U12445 ( .B1(n22612), .B2(n22530), .A(n22613), .ZN(n14943) );
  AND2_X1 U12446 ( .A1(n14957), .A2(n11155), .ZN(n15130) );
  INV_X1 U12447 ( .A(n22540), .ZN(n22809) );
  AND2_X1 U12448 ( .A1(n22555), .A2(n22583), .ZN(n22816) );
  INV_X1 U12449 ( .A(n22642), .ZN(n22636) );
  INV_X1 U12450 ( .A(n22696), .ZN(n22690) );
  OAI211_X1 U12451 ( .C1(n22578), .C2(n22605), .A(n22595), .B(n22577), .ZN(
        n22826) );
  INV_X1 U12452 ( .A(n22820), .ZN(n22825) );
  AOI22_X1 U12453 ( .A1(n22576), .A2(n22574), .B1(n22578), .B2(n22569), .ZN(
        n22830) );
  OAI211_X1 U12454 ( .C1(n22597), .C2(n22832), .A(n22596), .B(n22595), .ZN(
        n22835) );
  INV_X1 U12455 ( .A(n22591), .ZN(n22834) );
  NOR2_X1 U12456 ( .A1(n16592), .A2(n22386), .ZN(n22609) );
  NOR2_X1 U12457 ( .A1(n16592), .A2(n22404), .ZN(n22696) );
  NOR2_X1 U12458 ( .A1(n16592), .A2(n22418), .ZN(n22750) );
  AND2_X1 U12459 ( .A1(n16181), .A2(n14816), .ZN(n22841) );
  NOR2_X1 U12460 ( .A1(n22356), .A2(n11265), .ZN(n19018) );
  NOR2_X1 U12461 ( .A1(n16633), .A2(n16905), .ZN(n16632) );
  NAND2_X1 U12462 ( .A1(n12287), .A2(n11454), .ZN(n12305) );
  NAND2_X1 U12463 ( .A1(n15871), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11552) );
  NAND2_X1 U12464 ( .A1(n15880), .A2(n19322), .ZN(n11553) );
  INV_X1 U12465 ( .A(n19215), .ZN(n19261) );
  NOR2_X1 U12466 ( .A1(n19012), .A2(n15384), .ZN(n19227) );
  OR2_X1 U12468 ( .A1(n15115), .A2(n14359), .ZN(n15591) );
  INV_X1 U12469 ( .A(n19241), .ZN(n19268) );
  INV_X1 U12470 ( .A(n19208), .ZN(n19239) );
  OR2_X1 U12471 ( .A1(n14983), .A2(n15012), .ZN(n12640) );
  AND2_X1 U12472 ( .A1(n14648), .A2(n11175), .ZN(n14907) );
  NAND2_X1 U12473 ( .A1(n14648), .A2(n11169), .ZN(n14765) );
  INV_X1 U12474 ( .A(n16732), .ZN(n16724) );
  AND2_X2 U12475 ( .A1(n13025), .A2(n19014), .ZN(n16700) );
  NAND2_X1 U12476 ( .A1(n16700), .A2(n12006), .ZN(n16732) );
  NOR2_X1 U12477 ( .A1(n16668), .A2(n11186), .ZN(n16669) );
  AND2_X1 U12478 ( .A1(n15640), .A2(n15604), .ZN(n20113) );
  AND2_X1 U12479 ( .A1(n15640), .A2(n15603), .ZN(n20114) );
  AND2_X1 U12480 ( .A1(n15640), .A2(n15597), .ZN(n20115) );
  AND2_X1 U12481 ( .A1(n14751), .A2(n14752), .ZN(n14755) );
  INV_X1 U12482 ( .A(n20117), .ZN(n16790) );
  AND2_X1 U12483 ( .A1(n15640), .A2(n14510), .ZN(n20064) );
  OR2_X1 U12484 ( .A1(n20111), .A2(n14071), .ZN(n20065) );
  INV_X1 U12485 ( .A(n20065), .ZN(n20119) );
  INV_X1 U12486 ( .A(n15640), .ZN(n20111) );
  AND2_X1 U12487 ( .A1(n15640), .A2(n12011), .ZN(n20117) );
  NAND2_X1 U12489 ( .A1(n14366), .A2(n12393), .ZN(n14477) );
  INV_X1 U12490 ( .A(n15869), .ZN(n11526) );
  OR2_X1 U12491 ( .A1(n16861), .A2(n11599), .ZN(n15861) );
  NAND2_X1 U12492 ( .A1(n11180), .A2(n11600), .ZN(n11599) );
  NOR2_X1 U12493 ( .A1(n12345), .A2(n17065), .ZN(n11600) );
  OR2_X1 U12494 ( .A1(n16908), .A2(n11359), .ZN(n11353) );
  AND2_X1 U12495 ( .A1(n11336), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11332) );
  INV_X1 U12496 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17878) );
  NAND2_X1 U12497 ( .A1(n17321), .A2(n12429), .ZN(n17865) );
  INV_X1 U12498 ( .A(n17862), .ZN(n17042) );
  OR2_X1 U12499 ( .A1(n19335), .A2(n12393), .ZN(n17853) );
  INV_X1 U12500 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15895) );
  CLKBUF_X1 U12501 ( .A(n12089), .Z(n12090) );
  INV_X1 U12502 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17049) );
  AND2_X1 U12503 ( .A1(n17877), .A2(n14425), .ZN(n17862) );
  AND2_X1 U12504 ( .A1(n17877), .A2(n17414), .ZN(n17870) );
  OR2_X1 U12505 ( .A1(n12082), .A2(n12081), .ZN(n12083) );
  INV_X1 U12506 ( .A(n17877), .ZN(n17057) );
  INV_X1 U12507 ( .A(n17853), .ZN(n17871) );
  INV_X1 U12508 ( .A(n17870), .ZN(n17852) );
  INV_X1 U12509 ( .A(n11696), .ZN(n16815) );
  NOR2_X1 U12510 ( .A1(n14207), .A2(n14206), .ZN(n14208) );
  INV_X1 U12511 ( .A(n19228), .ZN(n14206) );
  NAND2_X1 U12512 ( .A1(n11438), .A2(n11704), .ZN(n16879) );
  NAND2_X1 U12513 ( .A1(n12324), .A2(n11446), .ZN(n11438) );
  NAND2_X1 U12514 ( .A1(n16949), .A2(n16895), .ZN(n16940) );
  AND2_X1 U12515 ( .A1(n17285), .A2(n17167), .ZN(n17238) );
  NAND2_X1 U12516 ( .A1(n16891), .A2(n17027), .ZN(n17021) );
  OR2_X1 U12517 ( .A1(n17169), .A2(n14185), .ZN(n17317) );
  NAND2_X1 U12518 ( .A1(n17039), .A2(n11700), .ZN(n11338) );
  NAND2_X1 U12519 ( .A1(n17038), .A2(n17037), .ZN(n17321) );
  CLKBUF_X1 U12520 ( .A(n15507), .Z(n15514) );
  NAND2_X1 U12521 ( .A1(n11337), .A2(n12422), .ZN(n15508) );
  INV_X1 U12522 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17418) );
  NOR2_X1 U12523 ( .A1(n14473), .A2(n14472), .ZN(n19836) );
  OAI21_X1 U12524 ( .B1(n14490), .B2(n14489), .A(n14488), .ZN(n19940) );
  NAND2_X1 U12525 ( .A1(n15038), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U12526 ( .B1(n19980), .B2(n19979), .A(n20009), .ZN(n20385) );
  INV_X1 U12527 ( .A(n20381), .ZN(n20273) );
  OAI21_X1 U12528 ( .B1(n19953), .B2(n19952), .A(n19951), .ZN(n20372) );
  NAND2_X1 U12529 ( .A1(n19928), .A2(n19997), .ZN(n20232) );
  INV_X1 U12530 ( .A(n20369), .ZN(n20360) );
  AOI22_X1 U12531 ( .A1(n19906), .A2(n19905), .B1(n19904), .B2(n19903), .ZN(
        n20346) );
  INV_X1 U12532 ( .A(n20343), .ZN(n20345) );
  OAI21_X1 U12533 ( .B1(n19892), .B2(n19895), .A(n19891), .ZN(n20339) );
  OR2_X1 U12534 ( .A1(n19885), .A2(n19927), .ZN(n20343) );
  OAI21_X1 U12535 ( .B1(n19881), .B2(n19880), .A(n19879), .ZN(n20332) );
  NOR2_X2 U12536 ( .A1(n19885), .A2(n19920), .ZN(n20338) );
  AOI22_X1 U12537 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20297), .ZN(n20248) );
  AOI22_X1 U12538 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20297), .ZN(n20204) );
  INV_X1 U12539 ( .A(n20290), .ZN(n20277) );
  NOR2_X1 U12540 ( .A1(n19927), .A2(n19843), .ZN(n20312) );
  INV_X1 U12541 ( .A(n20055), .ZN(n20059) );
  AOI22_X1 U12542 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20297), .ZN(n19984) );
  INV_X1 U12543 ( .A(n20312), .ZN(n20323) );
  INV_X1 U12544 ( .A(n20280), .ZN(n20284) );
  AOI22_X1 U12545 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20297), .ZN(n20240) );
  AOI22_X1 U12546 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20297), .ZN(n20105) );
  INV_X1 U12547 ( .A(n20110), .ZN(n20102) );
  AOI21_X1 U12548 ( .B1(n20303), .B2(n20009), .A(n19830), .ZN(n20306) );
  INV_X1 U12549 ( .A(n20316), .ZN(n20304) );
  INV_X1 U12550 ( .A(n20406), .ZN(n20390) );
  AOI22_X1 U12551 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20297), .ZN(n20395) );
  INV_X1 U12552 ( .A(n20240), .ZN(n20244) );
  INV_X1 U12553 ( .A(n20248), .ZN(n20237) );
  INV_X1 U12554 ( .A(n20196), .ZN(n20200) );
  INV_X1 U12555 ( .A(n20204), .ZN(n20193) );
  AOI22_X1 U12556 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20297), .ZN(n20158) );
  INV_X1 U12557 ( .A(n20105), .ZN(n20107) );
  OR2_X1 U12558 ( .A1(n19843), .A2(n19956), .ZN(n20309) );
  INV_X1 U12559 ( .A(n20062), .ZN(n20052) );
  AOI22_X1 U12560 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20297), .ZN(n20055) );
  INV_X1 U12561 ( .A(n20405), .ZN(n20285) );
  INV_X1 U12562 ( .A(n20309), .ZN(n20299) );
  INV_X1 U12563 ( .A(n19984), .ZN(n20003) );
  INV_X1 U12564 ( .A(n17389), .ZN(n19320) );
  OR2_X1 U12565 ( .A1(n22348), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n22347) );
  NAND2_X1 U12566 ( .A1(n21026), .A2(n21155), .ZN(n21027) );
  NAND2_X1 U12567 ( .A1(n21155), .A2(n11233), .ZN(n21012) );
  NAND2_X1 U12568 ( .A1(n21012), .A2(n21013), .ZN(n21026) );
  NOR2_X1 U12569 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20968), .ZN(n20991) );
  INV_X1 U12570 ( .A(n20941), .ZN(n21102) );
  NOR2_X1 U12571 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20883), .ZN(n20905) );
  NAND2_X1 U12572 ( .A1(n21187), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21168) );
  INV_X1 U12573 ( .A(n21141), .ZN(n21183) );
  AOI211_X1 U12574 ( .C1(n11149), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n15705), .B(n15704), .ZN(n15706) );
  NOR2_X1 U12575 ( .A1(n20823), .A2(n18003), .ZN(n18014) );
  NOR2_X1 U12576 ( .A1(n20796), .A2(n17987), .ZN(n17989) );
  CLKBUF_X1 U12577 ( .A(n18350), .Z(n18315) );
  INV_X1 U12578 ( .A(n18355), .ZN(n18348) );
  NOR3_X1 U12579 ( .A1(n19657), .A2(n19708), .A3(n21191), .ZN(n18355) );
  INV_X1 U12580 ( .A(n21330), .ZN(n21295) );
  NAND2_X1 U12581 ( .A1(n21295), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n21299) );
  INV_X1 U12582 ( .A(n21341), .ZN(n21342) );
  NOR2_X1 U12583 ( .A1(n18396), .A2(n18395), .ZN(n21231) );
  INV_X1 U12584 ( .A(n21370), .ZN(n21313) );
  INV_X1 U12585 ( .A(n21236), .ZN(n21246) );
  NAND2_X1 U12586 ( .A1(n21382), .A2(n21379), .ZN(n21373) );
  NAND2_X1 U12587 ( .A1(n21294), .A2(n21379), .ZN(n21370) );
  INV_X1 U12588 ( .A(n21241), .ZN(n21377) );
  CLKBUF_X1 U12591 ( .A(n20732), .Z(n20761) );
  NAND2_X1 U12592 ( .A1(n18671), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18743) );
  NAND2_X1 U12593 ( .A1(n18680), .A2(n21747), .ZN(n21727) );
  NOR3_X1 U12594 ( .A1(n21655), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n21654), .ZN(n11371) );
  NOR2_X1 U12595 ( .A1(n21630), .A2(n21604), .ZN(n21752) );
  NOR2_X1 U12596 ( .A1(n21630), .A2(n21622), .ZN(n21456) );
  INV_X1 U12597 ( .A(n18667), .ZN(n18708) );
  NAND2_X1 U12598 ( .A1(n18523), .A2(n11316), .ZN(n18620) );
  NOR2_X1 U12599 ( .A1(n18552), .A2(n18557), .ZN(n20981) );
  NAND2_X1 U12600 ( .A1(n18861), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18848) );
  INV_X1 U12601 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18849) );
  INV_X1 U12602 ( .A(n18858), .ZN(n18861) );
  AND2_X1 U12603 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18874) );
  INV_X2 U12604 ( .A(n19703), .ZN(n19704) );
  INV_X1 U12605 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20782) );
  OAI22_X1 U12606 ( .A1(n21705), .A2(n21704), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21707) );
  NOR2_X1 U12607 ( .A1(n21596), .A2(n18769), .ZN(n21616) );
  NOR2_X2 U12608 ( .A1(n21728), .A2(n21547), .ZN(n21865) );
  NOR2_X2 U12609 ( .A1(n21447), .A2(n21937), .ZN(n21841) );
  NOR4_X1 U12610 ( .A1(n21446), .A2(n21445), .A3(n21444), .A4(n21443), .ZN(
        n21447) );
  NAND2_X1 U12611 ( .A1(n21841), .A2(n21883), .ZN(n21547) );
  INV_X1 U12612 ( .A(n21849), .ZN(n21859) );
  INV_X1 U12613 ( .A(n21761), .ZN(n21754) );
  INV_X1 U12614 ( .A(n21841), .ZN(n21808) );
  NOR2_X1 U12615 ( .A1(n19571), .A2(n19389), .ZN(n18917) );
  INV_X1 U12616 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21904) );
  INV_X1 U12617 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19698) );
  INV_X1 U12618 ( .A(n21937), .ZN(n21932) );
  NOR2_X1 U12619 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n21936), .ZN(n21917) );
  CLKBUF_X1 U12620 ( .A(n19360), .Z(n19699) );
  OAI21_X1 U12621 ( .B1(n16429), .B2(n22280), .A(n14015), .ZN(P1_U2969) );
  AOI21_X1 U12622 ( .B1(n11382), .B2(n17830), .A(n17829), .ZN(n17839) );
  OAI21_X1 U12623 ( .B1(n17067), .B2(n19302), .A(n11378), .ZN(n17069) );
  AOI21_X1 U12624 ( .B1(n16908), .B2(n11352), .A(n11361), .ZN(n11349) );
  NAND2_X1 U12625 ( .A1(n11354), .A2(n11351), .ZN(n11350) );
  AND2_X1 U12626 ( .A1(n11172), .A2(n19299), .ZN(n11352) );
  AND2_X1 U12627 ( .A1(n11336), .A2(n11224), .ZN(n11334) );
  AOI22_X1 U12628 ( .A1(n18667), .A2(n11371), .B1(n21661), .B2(n18812), .ZN(
        n18709) );
  NAND2_X1 U12629 ( .A1(n11558), .A2(n11560), .ZN(n15436) );
  AND2_X1 U12630 ( .A1(n11621), .A2(n11170), .ZN(n11160) );
  OR2_X1 U12631 ( .A1(n16626), .A2(n16627), .ZN(n11161) );
  OR3_X1 U12632 ( .A1(n11161), .A2(n11575), .A3(n11250), .ZN(n11162) );
  NOR2_X1 U12633 ( .A1(n17849), .A2(n11561), .ZN(n11560) );
  NAND2_X1 U12634 ( .A1(n16044), .A2(n11628), .ZN(n11163) );
  NOR2_X1 U12635 ( .A1(n15275), .A2(n11559), .ZN(n15437) );
  AND4_X1 U12636 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        n11164) );
  NAND2_X1 U12637 ( .A1(n14972), .A2(n14889), .ZN(n11165) );
  INV_X1 U12638 ( .A(n12441), .ZN(n12466) );
  NOR2_X2 U12639 ( .A1(n15698), .A2(n15697), .ZN(n19708) );
  INV_X1 U12640 ( .A(n12413), .ZN(n11269) );
  AND4_X1 U12641 ( .A1(n16889), .A2(n12340), .A3(n16915), .A4(n16927), .ZN(
        n11166) );
  NAND2_X1 U12642 ( .A1(n16986), .A2(n11603), .ZN(n16880) );
  AND2_X1 U12643 ( .A1(n11530), .A2(n11529), .ZN(n11167) );
  AND2_X1 U12644 ( .A1(n11560), .A2(n11557), .ZN(n11168) );
  NOR2_X1 U12645 ( .A1(n11548), .A2(n16902), .ZN(n15783) );
  NAND2_X1 U12646 ( .A1(n15595), .A2(n11685), .ZN(n15635) );
  NOR2_X1 U12647 ( .A1(n15434), .A2(n17878), .ZN(n15435) );
  NOR2_X1 U12648 ( .A1(n15788), .A2(n12538), .ZN(n15787) );
  NOR3_X1 U12649 ( .A1(n15788), .A2(n11551), .A3(n12538), .ZN(n15786) );
  AND2_X1 U12650 ( .A1(n15025), .A2(n11227), .ZN(n15332) );
  NAND2_X1 U12651 ( .A1(n11143), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15782) );
  NOR3_X1 U12652 ( .A1(n15442), .A2(n11566), .A3(n11567), .ZN(n15464) );
  AND2_X1 U12653 ( .A1(n14647), .A2(n11724), .ZN(n11169) );
  AND2_X1 U12654 ( .A1(n13430), .A2(n11620), .ZN(n11170) );
  AND2_X1 U12655 ( .A1(n11454), .A2(n11453), .ZN(n11171) );
  AND2_X1 U12656 ( .A1(n16900), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11172) );
  AND2_X1 U12657 ( .A1(n11309), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11173) );
  AND2_X1 U12658 ( .A1(n11171), .A2(n12299), .ZN(n11174) );
  INV_X1 U12659 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16966) );
  AND2_X1 U12660 ( .A1(n11169), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11175) );
  NAND2_X1 U12661 ( .A1(n14751), .A2(n11223), .ZN(n15456) );
  AND2_X1 U12662 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11176) );
  AND2_X1 U12663 ( .A1(n11176), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11177) );
  AND2_X1 U12664 ( .A1(n11555), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11178) );
  AND2_X1 U12665 ( .A1(n11460), .A2(n11246), .ZN(n11179) );
  INV_X1 U12666 ( .A(n17157), .ZN(n11605) );
  AND2_X1 U12667 ( .A1(n11602), .A2(n17098), .ZN(n11180) );
  AND2_X1 U12668 ( .A1(n11603), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11181) );
  AND2_X2 U12669 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11735), .ZN(
        n11813) );
  OR2_X1 U12670 ( .A1(n15568), .A2(n11535), .ZN(n11182) );
  OR2_X1 U12671 ( .A1(n16710), .A2(n16709), .ZN(n11183) );
  NAND2_X1 U12672 ( .A1(n12206), .A2(n11458), .ZN(n12260) );
  OR2_X1 U12673 ( .A1(n16139), .A2(n11473), .ZN(n11185) );
  AND2_X1 U12674 ( .A1(n11675), .A2(n12950), .ZN(n11186) );
  OR2_X1 U12675 ( .A1(n14088), .A2(n14087), .ZN(n11187) );
  INV_X1 U12676 ( .A(n18409), .ZN(n20786) );
  INV_X2 U12677 ( .A(n20786), .ZN(n18456) );
  OR2_X1 U12678 ( .A1(n11162), .A2(n11578), .ZN(n11188) );
  NAND2_X2 U12679 ( .A1(n12979), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12150) );
  NAND2_X1 U12680 ( .A1(n16044), .A2(n16046), .ZN(n16027) );
  OR3_X1 U12681 ( .A1(n16062), .A2(n11478), .A3(n16002), .ZN(n11189) );
  NOR2_X1 U12682 ( .A1(n15275), .A2(n17849), .ZN(n15375) );
  AND2_X1 U12683 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15274) );
  AND2_X1 U12684 ( .A1(n16044), .A2(n11626), .ZN(n16009) );
  INV_X1 U12685 ( .A(n11295), .ZN(n14479) );
  OR2_X1 U12686 ( .A1(n15651), .A2(n21411), .ZN(n11190) );
  AND4_X1 U12687 ( .A1(n13097), .A2(n13096), .A3(n13095), .A4(n13094), .ZN(
        n11191) );
  AND4_X1 U12688 ( .A1(n11766), .A2(n11765), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(n11764), .ZN(n11192) );
  AND2_X1 U12689 ( .A1(n13142), .A2(n13141), .ZN(n11193) );
  INV_X1 U12690 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17860) );
  NAND2_X1 U12691 ( .A1(n11699), .A2(n12268), .ZN(n17866) );
  XNOR2_X1 U12692 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15860), .ZN(
        n11195) );
  INV_X2 U12693 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11777) );
  AND2_X1 U12694 ( .A1(n12292), .A2(n11179), .ZN(n11196) );
  NOR2_X1 U12695 ( .A1(n16861), .A2(n12345), .ZN(n11197) );
  AND2_X1 U12696 ( .A1(n12287), .A2(n11171), .ZN(n11198) );
  AND2_X1 U12697 ( .A1(n12375), .A2(n15855), .ZN(n11199) );
  NAND2_X1 U12698 ( .A1(n13304), .A2(n13303), .ZN(n13335) );
  NOR2_X1 U12699 ( .A1(n16861), .A2(n11598), .ZN(n11200) );
  AND4_X1 U12700 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n11201) );
  AND2_X1 U12701 ( .A1(n12116), .A2(n15076), .ZN(n11202) );
  NOR2_X1 U12702 ( .A1(n11604), .A2(n11147), .ZN(n16888) );
  NAND2_X1 U12703 ( .A1(n15952), .A2(n15954), .ZN(n15941) );
  AND2_X1 U12704 ( .A1(n11457), .A2(n11458), .ZN(n11203) );
  XNOR2_X1 U12705 ( .A(n11527), .B(n11526), .ZN(n19252) );
  AND3_X1 U12706 ( .A1(n12072), .A2(n11669), .A3(n12073), .ZN(n11204) );
  INV_X2 U12707 ( .A(n21294), .ZN(n21267) );
  OR2_X1 U12708 ( .A1(n12441), .A2(n17053), .ZN(n11205) );
  AND2_X1 U12709 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U12710 ( .A1(n12085), .A2(n12083), .ZN(n15076) );
  NAND2_X1 U12711 ( .A1(n12413), .A2(n15522), .ZN(n11207) );
  OR3_X1 U12712 ( .A1(n11161), .A2(n11575), .A3(n17143), .ZN(n11208) );
  NAND3_X1 U12713 ( .A1(n14503), .A2(n11187), .A3(n14093), .ZN(n11209) );
  AND2_X1 U12714 ( .A1(n20590), .A2(n11426), .ZN(n11210) );
  NAND2_X1 U12715 ( .A1(n12111), .A2(n12110), .ZN(n12181) );
  INV_X1 U12716 ( .A(n12181), .ZN(n19902) );
  AND2_X1 U12717 ( .A1(n12116), .A2(n12118), .ZN(n11211) );
  NAND2_X1 U12718 ( .A1(n15274), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15275) );
  INV_X1 U12719 ( .A(n15275), .ZN(n11558) );
  NOR2_X1 U12720 ( .A1(n21562), .A2(n18520), .ZN(n11212) );
  INV_X1 U12721 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n21392) );
  AND2_X1 U12722 ( .A1(n11296), .A2(n20125), .ZN(n11213) );
  OAI21_X1 U12723 ( .B1(n17166), .B2(n19302), .A(n17165), .ZN(n11361) );
  NAND2_X1 U12724 ( .A1(n11447), .A2(n11444), .ZN(n11214) );
  AND2_X1 U12725 ( .A1(n16986), .A2(n11181), .ZN(n11215) );
  NAND2_X1 U12726 ( .A1(n16696), .A2(n11547), .ZN(n16679) );
  OR2_X1 U12727 ( .A1(n12210), .A2(n11289), .ZN(n11216) );
  AND3_X1 U12728 ( .A1(n11982), .A2(n11292), .A3(n11291), .ZN(n11217) );
  INV_X1 U12729 ( .A(n13196), .ZN(n11613) );
  AND2_X1 U12730 ( .A1(n12005), .A2(n11955), .ZN(n11218) );
  NAND2_X1 U12731 ( .A1(n19112), .A2(n19123), .ZN(n11219) );
  OR2_X1 U12732 ( .A1(n15982), .A2(n11467), .ZN(n11220) );
  AND2_X1 U12733 ( .A1(n13133), .A2(n13121), .ZN(n11221) );
  NAND2_X1 U12734 ( .A1(n14804), .A2(n13157), .ZN(n13184) );
  NAND2_X1 U12735 ( .A1(n13983), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11222) );
  NAND2_X1 U12736 ( .A1(n14648), .A2(n14647), .ZN(n14646) );
  NOR2_X1 U12737 ( .A1(n11182), .A2(n16641), .ZN(n16624) );
  NAND2_X1 U12738 ( .A1(n11558), .A2(n11168), .ZN(n15434) );
  AND2_X1 U12739 ( .A1(n15595), .A2(n15594), .ZN(n15592) );
  NAND2_X1 U12740 ( .A1(n15025), .A2(n15024), .ZN(n15023) );
  AND2_X1 U12741 ( .A1(n15025), .A2(n11680), .ZN(n15200) );
  NAND2_X1 U12742 ( .A1(n15014), .A2(n11530), .ZN(n15327) );
  INV_X1 U12743 ( .A(n12203), .ZN(n15859) );
  NAND2_X1 U12744 ( .A1(n14839), .A2(n13922), .ZN(n11618) );
  AND2_X1 U12745 ( .A1(n11585), .A2(n15457), .ZN(n11223) );
  NOR2_X2 U12746 ( .A1(n18446), .A2(n21728), .ZN(n18721) );
  NAND2_X1 U12747 ( .A1(n11713), .A2(n11590), .ZN(n16796) );
  INV_X1 U12748 ( .A(n15817), .ZN(n11638) );
  NAND2_X1 U12749 ( .A1(n11338), .A2(n11697), .ZN(n17028) );
  INV_X1 U12750 ( .A(n11648), .ZN(n22555) );
  NOR3_X1 U12751 ( .A1(n15442), .A2(n11568), .A3(n16999), .ZN(n15465) );
  AND2_X1 U12752 ( .A1(n15435), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15431) );
  AND2_X1 U12753 ( .A1(n17377), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11224) );
  OR3_X1 U12754 ( .A1(n15442), .A2(n11567), .A3(n11568), .ZN(n11225) );
  XNOR2_X1 U12755 ( .A(DATAI_27_), .B(keyinput_133), .ZN(n11226) );
  INV_X1 U12756 ( .A(n13936), .ZN(n11647) );
  AND2_X1 U12757 ( .A1(n11680), .A2(n15334), .ZN(n11227) );
  OR3_X1 U12758 ( .A1(n15568), .A2(n15567), .A3(n11538), .ZN(n11228) );
  OR2_X1 U12759 ( .A1(n16062), .A2(n11478), .ZN(n11229) );
  XOR2_X1 U12760 ( .A(DATAI_27_), .B(keyinput_5), .Z(n11230) );
  INV_X1 U12761 ( .A(n15020), .ZN(n12478) );
  NOR2_X1 U12762 ( .A1(n15015), .A2(n15016), .ZN(n15014) );
  INV_X1 U12763 ( .A(n11701), .ZN(n11700) );
  OAI21_X1 U12764 ( .B1(n17040), .B2(n11702), .A(n17867), .ZN(n11701) );
  AND2_X1 U12765 ( .A1(n20603), .A2(n16414), .ZN(n11231) );
  AND2_X1 U12766 ( .A1(n11223), .A2(n11584), .ZN(n11232) );
  INV_X1 U12767 ( .A(n15618), .ZN(n11633) );
  OR2_X1 U12768 ( .A1(n21011), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11233) );
  NAND2_X1 U12769 ( .A1(n13696), .A2(n13695), .ZN(n16018) );
  AND2_X1 U12770 ( .A1(n13389), .A2(n13388), .ZN(n13405) );
  INV_X1 U12771 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16999) );
  OR2_X1 U12772 ( .A1(n16139), .A2(n16138), .ZN(n11234) );
  OR3_X1 U12773 ( .A1(n15788), .A2(n12538), .A3(n11550), .ZN(n11235) );
  INV_X1 U12774 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11568) );
  OR2_X1 U12775 ( .A1(n11488), .A2(n11487), .ZN(n11236) );
  INV_X1 U12776 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16919) );
  INV_X1 U12777 ( .A(n17351), .ZN(n19299) );
  AND2_X1 U12778 ( .A1(n11316), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11237) );
  NOR2_X1 U12779 ( .A1(n17062), .A2(n17063), .ZN(n11238) );
  NOR2_X1 U12780 ( .A1(n16632), .A2(n15794), .ZN(n11239) );
  NOR2_X1 U12781 ( .A1(n12549), .A2(n11676), .ZN(n11240) );
  AND2_X1 U12782 ( .A1(n12171), .A2(n14066), .ZN(n11241) );
  AND2_X1 U12783 ( .A1(n11563), .A2(n11158), .ZN(n11242) );
  NAND2_X1 U12784 ( .A1(n11572), .A2(n14889), .ZN(n14890) );
  NAND2_X1 U12785 ( .A1(n11143), .A2(n11178), .ZN(n15780) );
  NOR2_X1 U12786 ( .A1(n14650), .A2(n14656), .ZN(n14655) );
  AND2_X1 U12787 ( .A1(n14751), .A2(n11585), .ZN(n14754) );
  AND2_X1 U12788 ( .A1(n11143), .A2(n11555), .ZN(n11243) );
  AND2_X1 U12789 ( .A1(n15799), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14024) );
  AND2_X1 U12790 ( .A1(n18671), .A2(n11313), .ZN(n11244) );
  INV_X1 U12791 ( .A(n15366), .ZN(n11529) );
  OR2_X1 U12792 ( .A1(n18520), .A2(n21596), .ZN(n11245) );
  NAND2_X1 U12793 ( .A1(n14112), .A2(n14111), .ZN(n14751) );
  OR2_X1 U12794 ( .A1(n14065), .A2(n11909), .ZN(n11246) );
  AND3_X1 U12795 ( .A1(n11519), .A2(n17749), .A3(n11518), .ZN(n11247) );
  XNOR2_X1 U12796 ( .A(n13178), .B(n13194), .ZN(n14919) );
  INV_X1 U12797 ( .A(n12291), .ZN(n11461) );
  OR2_X1 U12798 ( .A1(n17555), .A2(n17554), .ZN(n11248) );
  OR2_X1 U12799 ( .A1(n17721), .A2(n17723), .ZN(n11249) );
  INV_X1 U12800 ( .A(n12012), .ZN(n12571) );
  OR2_X1 U12801 ( .A1(n17143), .A2(n16763), .ZN(n11250) );
  OR2_X2 U12802 ( .A1(n17449), .A2(n22303), .ZN(n22280) );
  INV_X1 U12803 ( .A(n22280), .ZN(n20595) );
  AND2_X1 U12804 ( .A1(n11545), .A2(n11544), .ZN(n11251) );
  AND2_X1 U12805 ( .A1(n15857), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n11252) );
  AND2_X1 U12806 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_42), .ZN(n11253) );
  AND2_X1 U12807 ( .A1(n11683), .A2(n11682), .ZN(n11254) );
  AND2_X1 U12808 ( .A1(n11177), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11255) );
  AND2_X1 U12809 ( .A1(n11179), .A2(n11459), .ZN(n11256) );
  OR2_X1 U12810 ( .A1(n11245), .A2(n11303), .ZN(n11257) );
  INV_X1 U12811 ( .A(n21877), .ZN(n11369) );
  INV_X1 U12812 ( .A(n16216), .ZN(n11632) );
  NAND2_X1 U12813 ( .A1(n15799), .A2(n11176), .ZN(n14023) );
  AND2_X1 U12814 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15060) );
  AND2_X1 U12815 ( .A1(n18782), .A2(n11309), .ZN(n11258) );
  AND3_X1 U12816 ( .A1(n11416), .A2(n17577), .A3(n11415), .ZN(n11259) );
  INV_X1 U12817 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11556) );
  INV_X1 U12818 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11322) );
  AND2_X1 U12819 ( .A1(n12435), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11260) );
  OR2_X1 U12820 ( .A1(n18711), .A2(n21654), .ZN(n11261) );
  INV_X1 U12821 ( .A(n17076), .ZN(n11602) );
  INV_X1 U12822 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11303) );
  AND2_X1 U12823 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_212), .ZN(n11262)
         );
  INV_X1 U12824 ( .A(n14011), .ZN(n11666) );
  INV_X1 U12825 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11314) );
  INV_X1 U12826 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11310) );
  INV_X1 U12827 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11550) );
  INV_X1 U12828 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11311) );
  NOR2_X1 U12829 ( .A1(n14840), .A2(n14797), .ZN(n11263) );
  OR3_X1 U12830 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14792), .A3(n13173), 
        .ZN(n14840) );
  CLKBUF_X1 U12831 ( .A(n21148), .Z(n11264) );
  NOR4_X1 U12832 ( .A1(n21389), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n21148)
         );
  NOR2_X1 U12833 ( .A1(n12023), .A2(n11267), .ZN(n12024) );
  NAND2_X1 U12834 ( .A1(n11267), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11295) );
  AND2_X1 U12835 ( .A1(n12393), .A2(n11267), .ZN(n15390) );
  NAND2_X1 U12836 ( .A1(n20294), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11265) );
  INV_X2 U12837 ( .A(n11267), .ZN(n20294) );
  AND2_X1 U12838 ( .A1(n14053), .A2(n11267), .ZN(n15122) );
  NOR2_X1 U12839 ( .A1(n11433), .A2(n11267), .ZN(n14041) );
  AND2_X1 U12840 ( .A1(n14172), .A2(n11267), .ZN(n11266) );
  OAI21_X1 U12841 ( .B1(n14039), .B2(n11267), .A(n11954), .ZN(n14040) );
  NAND2_X4 U12842 ( .A1(n11785), .A2(n11784), .ZN(n11267) );
  AOI21_X1 U12843 ( .B1(n12411), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n11269), .ZN(n11268) );
  INV_X1 U12844 ( .A(n12411), .ZN(n11271) );
  NAND2_X1 U12845 ( .A1(n12412), .A2(n12411), .ZN(n12417) );
  NAND2_X2 U12846 ( .A1(n11272), .A2(n12409), .ZN(n12411) );
  INV_X1 U12847 ( .A(n12410), .ZN(n11272) );
  NAND2_X2 U12848 ( .A1(n17856), .A2(n12424), .ZN(n17038) );
  NAND2_X2 U12849 ( .A1(n17339), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17856) );
  NAND2_X1 U12850 ( .A1(n15507), .A2(n12416), .ZN(n11273) );
  NOR2_X2 U12851 ( .A1(n16973), .A2(n17240), .ZN(n17216) );
  NAND2_X1 U12852 ( .A1(n11278), .A2(n11275), .ZN(P2_U2994) );
  AOI21_X1 U12853 ( .B1(n11276), .B2(n17843), .A(n16912), .ZN(n11275) );
  NAND2_X1 U12854 ( .A1(n11277), .A2(n11335), .ZN(n11276) );
  NAND2_X1 U12855 ( .A1(n16924), .A2(n11332), .ZN(n11277) );
  OR2_X1 U12856 ( .A1(n17185), .A2(n17853), .ZN(n11278) );
  NAND3_X1 U12857 ( .A1(n12025), .A2(n14171), .A3(n14047), .ZN(n13022) );
  AND4_X2 U12858 ( .A1(n12025), .A2(n12033), .A3(n14171), .A4(n14047), .ZN(
        n14202) );
  NAND3_X1 U12859 ( .A1(n11281), .A2(n16246), .A3(n11280), .ZN(n11279) );
  NAND2_X1 U12860 ( .A1(n16274), .A2(n11661), .ZN(n11282) );
  INV_X1 U12861 ( .A(n13363), .ZN(n13365) );
  NAND3_X1 U12862 ( .A1(n13304), .A2(n13303), .A3(n22582), .ZN(n13363) );
  NAND2_X2 U12863 ( .A1(n11285), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13306) );
  NAND3_X1 U12864 ( .A1(n13172), .A2(n13176), .A3(n13171), .ZN(n11285) );
  INV_X2 U12865 ( .A(n13994), .ZN(n20617) );
  AND2_X2 U12866 ( .A1(n13046), .A2(n16572), .ZN(n13122) );
  AND2_X2 U12867 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16572) );
  INV_X1 U12868 ( .A(n12421), .ZN(n11286) );
  NAND2_X1 U12869 ( .A1(n11728), .A2(n11287), .ZN(P2_U2986) );
  INV_X2 U12870 ( .A(n12972), .ZN(n12982) );
  NAND3_X1 U12871 ( .A1(n11525), .A2(n11744), .A3(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11290) );
  NOR2_X2 U12872 ( .A1(n12109), .A2(n12107), .ZN(n19950) );
  NOR2_X2 U12873 ( .A1(n12109), .A2(n12108), .ZN(n19930) );
  OR2_X2 U12874 ( .A1(n12110), .A2(n12116), .ZN(n12109) );
  NAND2_X1 U12875 ( .A1(n18685), .A2(n21748), .ZN(n18680) );
  NAND3_X1 U12876 ( .A1(n18588), .A2(n11304), .A3(n11303), .ZN(n11302) );
  OAI211_X2 U12877 ( .C1(n11306), .C2(n11261), .A(n18678), .B(n18705), .ZN(
        n11305) );
  OR2_X2 U12878 ( .A1(n18659), .A2(n11307), .ZN(n11306) );
  OR2_X2 U12879 ( .A1(n18647), .A2(n21768), .ZN(n11307) );
  INV_X2 U12880 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21385) );
  INV_X1 U12881 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11315) );
  INV_X1 U12882 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11318) );
  INV_X2 U12883 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21888) );
  INV_X1 U12884 ( .A(n18845), .ZN(n11325) );
  NAND2_X1 U12886 ( .A1(n11331), .A2(n11329), .ZN(P2_U3026) );
  AOI21_X1 U12887 ( .B1(n11334), .B2(n16924), .A(n11330), .ZN(n11329) );
  OR2_X1 U12888 ( .A1(n17185), .A2(n17351), .ZN(n11331) );
  NAND3_X1 U12889 ( .A1(n11337), .A2(n12422), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15507) );
  OR2_X1 U12890 ( .A1(n16948), .A2(n11346), .ZN(n11342) );
  NAND2_X1 U12891 ( .A1(n11342), .A2(n11343), .ZN(n11484) );
  INV_X1 U12892 ( .A(n16908), .ZN(n11351) );
  OAI211_X1 U12893 ( .C1(n11356), .C2(n17351), .A(n11350), .B(n11349), .ZN(
        P2_U3025) );
  NAND2_X1 U12894 ( .A1(n16908), .A2(n11172), .ZN(n11355) );
  NAND3_X1 U12895 ( .A1(n11355), .A2(n11356), .A3(n11353), .ZN(n17154) );
  NOR2_X2 U12896 ( .A1(n21255), .A2(n19490), .ZN(n21382) );
  OR2_X2 U12897 ( .A1(n21831), .A2(n21435), .ZN(n21885) );
  XNOR2_X2 U12898 ( .A(n12436), .B(n12439), .ZN(n12116) );
  NAND2_X1 U12899 ( .A1(n12078), .A2(n12079), .ZN(n11373) );
  NAND3_X1 U12900 ( .A1(n11376), .A2(n11375), .A3(n11753), .ZN(n11377) );
  AND2_X1 U12901 ( .A1(n11754), .A2(n11777), .ZN(n11375) );
  NAND3_X1 U12902 ( .A1(n12412), .A2(n12411), .A3(n11269), .ZN(n12422) );
  NAND4_X1 U12903 ( .A1(n14804), .A2(n13157), .A3(n14548), .A4(n14628), .ZN(
        n13168) );
  NAND3_X1 U12904 ( .A1(n14809), .A2(n14628), .A3(n11420), .ZN(n11419) );
  OAI21_X1 U12905 ( .B1(n16562), .B2(n13984), .A(n13924), .ZN(n14514) );
  OAI21_X2 U12906 ( .B1(n16255), .B2(n16258), .A(n20617), .ZN(n16266) );
  NAND2_X2 U12907 ( .A1(n16307), .A2(n14013), .ZN(n16255) );
  OAI21_X1 U12908 ( .B1(n20594), .B2(n11422), .A(n11222), .ZN(n11421) );
  NAND2_X1 U12909 ( .A1(n11424), .A2(n11425), .ZN(n15499) );
  OAI21_X1 U12910 ( .B1(n15497), .B2(n11429), .A(n11427), .ZN(n16338) );
  NAND2_X1 U12911 ( .A1(n12002), .A2(n11433), .ZN(n14170) );
  NAND4_X1 U12912 ( .A1(n11762), .A2(n11760), .A3(n11435), .A4(n11761), .ZN(
        n11434) );
  NAND2_X2 U12913 ( .A1(n12265), .A2(n12264), .ZN(n17039) );
  OAI21_X2 U12914 ( .B1(n12324), .B2(n11441), .A(n11439), .ZN(n16871) );
  AND2_X2 U12915 ( .A1(n11452), .A2(n11451), .ZN(n16837) );
  NAND2_X1 U12916 ( .A1(n12206), .A2(n11456), .ZN(n12274) );
  NAND2_X1 U12917 ( .A1(n12292), .A2(n11256), .ZN(n12343) );
  NAND2_X1 U12918 ( .A1(n12292), .A2(n11460), .ZN(n12328) );
  NAND2_X1 U12919 ( .A1(n12292), .A2(n12291), .ZN(n12326) );
  NAND2_X2 U12920 ( .A1(n14226), .A2(n14222), .ZN(n14321) );
  AND2_X2 U12921 ( .A1(n14694), .A2(n13047), .ZN(n13254) );
  AOI211_X1 U12922 ( .C1(n15982), .C2(n14226), .A(n11462), .B(n11464), .ZN(
        n11463) );
  NOR2_X1 U12923 ( .A1(n15982), .A2(n11466), .ZN(n15945) );
  NAND4_X1 U12924 ( .A1(n12103), .A2(n12104), .A3(n11483), .A4(n11482), .ZN(
        n12105) );
  NAND2_X1 U12925 ( .A1(n11492), .A2(n12200), .ZN(n11491) );
  NAND2_X1 U12926 ( .A1(n11490), .A2(n19034), .ZN(n12235) );
  NAND3_X1 U12927 ( .A1(n11491), .A2(n12203), .A3(n12202), .ZN(n11490) );
  NAND2_X1 U12928 ( .A1(n12426), .A2(n12202), .ZN(n12413) );
  NAND3_X1 U12929 ( .A1(n12011), .A2(n12571), .A3(n11218), .ZN(n11975) );
  NOR2_X1 U12930 ( .A1(n11525), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15089) );
  AND2_X2 U12931 ( .A1(n11525), .A2(n11757), .ZN(n11964) );
  AND2_X1 U12932 ( .A1(n12820), .A2(n11525), .ZN(n12795) );
  NOR2_X1 U12933 ( .A1(n11745), .A2(n11525), .ZN(n15069) );
  NAND3_X1 U12934 ( .A1(n12032), .A2(n14174), .A3(n12033), .ZN(n15061) );
  NAND2_X1 U12935 ( .A1(n15014), .A2(n11167), .ZN(n15539) );
  NOR2_X1 U12936 ( .A1(n15568), .A2(n15567), .ZN(n15611) );
  INV_X1 U12937 ( .A(n15610), .ZN(n11538) );
  INV_X1 U12938 ( .A(n14903), .ZN(n11539) );
  NAND2_X1 U12939 ( .A1(n11539), .A2(n11540), .ZN(n15015) );
  AOI21_X2 U12940 ( .B1(n12436), .B2(n12439), .A(n12438), .ZN(n14652) );
  INV_X1 U12941 ( .A(n16673), .ZN(n11544) );
  NAND2_X1 U12942 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11549) );
  AND2_X1 U12943 ( .A1(n11178), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11554) );
  INV_X1 U12944 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11561) );
  AND2_X1 U12945 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U12946 ( .A1(n11562), .A2(n11563), .ZN(n19153) );
  INV_X1 U12947 ( .A(n14096), .ZN(n11572) );
  NAND2_X1 U12948 ( .A1(n11572), .A2(n11573), .ZN(n14109) );
  INV_X1 U12949 ( .A(n16779), .ZN(n11576) );
  NOR2_X1 U12950 ( .A1(n11162), .A2(n11577), .ZN(n14160) );
  INV_X1 U12951 ( .A(n14161), .ZN(n11583) );
  OAI21_X2 U12952 ( .B1(n17038), .B2(n11597), .A(n11595), .ZN(n17863) );
  INV_X1 U12953 ( .A(n14919), .ZN(n11610) );
  INV_X1 U12954 ( .A(n13202), .ZN(n11608) );
  OAI211_X1 U12955 ( .C1(n11608), .C2(n13219), .A(n11612), .B(n11607), .ZN(
        n14672) );
  NAND3_X1 U12956 ( .A1(n11608), .A2(n13219), .A3(n13196), .ZN(n11607) );
  NAND2_X2 U12957 ( .A1(n11610), .A2(n11609), .ZN(n13219) );
  NAND3_X1 U12958 ( .A1(n11614), .A2(n14825), .A3(n13854), .ZN(n13160) );
  NAND4_X1 U12959 ( .A1(n11614), .A2(n14825), .A3(n13854), .A4(n14886), .ZN(
        n15902) );
  INV_X1 U12960 ( .A(n14886), .ZN(n15177) );
  NOR2_X2 U12961 ( .A1(n15254), .A2(n11619), .ZN(n15370) );
  INV_X1 U12962 ( .A(n13395), .ZN(n11624) );
  NAND2_X1 U12963 ( .A1(n11624), .A2(n13394), .ZN(n13404) );
  INV_X1 U12964 ( .A(n15618), .ZN(n11630) );
  AND2_X2 U12965 ( .A1(n15969), .A2(n13780), .ZN(n15952) );
  AND2_X1 U12966 ( .A1(n15969), .A2(n11636), .ZN(n15942) );
  NAND2_X1 U12967 ( .A1(n15969), .A2(n11637), .ZN(n15821) );
  NAND2_X1 U12968 ( .A1(n13249), .A2(n13274), .ZN(n13282) );
  NAND2_X1 U12969 ( .A1(n11644), .A2(n11642), .ZN(n13274) );
  NAND2_X1 U12970 ( .A1(n13219), .A2(n15210), .ZN(n14636) );
  NAND2_X1 U12971 ( .A1(n11644), .A2(n13230), .ZN(n13925) );
  NOR2_X1 U12972 ( .A1(n13248), .A2(n11643), .ZN(n11642) );
  INV_X1 U12973 ( .A(n13230), .ZN(n11643) );
  NAND2_X1 U12974 ( .A1(n11649), .A2(n13975), .ZN(n13921) );
  NAND2_X1 U12975 ( .A1(n11649), .A2(n13537), .ZN(n13334) );
  NAND2_X1 U12976 ( .A1(n16568), .A2(n11647), .ZN(n22512) );
  NAND2_X1 U12977 ( .A1(n11649), .A2(n11647), .ZN(n11648) );
  NAND2_X1 U12978 ( .A1(n11658), .A2(n11659), .ZN(n16245) );
  INV_X1 U12979 ( .A(n16441), .ZN(n11652) );
  NAND2_X1 U12980 ( .A1(n20604), .A2(n11663), .ZN(n11662) );
  NAND2_X1 U12981 ( .A1(n11662), .A2(n11664), .ZN(n16309) );
  NOR2_X2 U12982 ( .A1(n14010), .A2(n11668), .ZN(n11667) );
  INV_X2 U12983 ( .A(n12466), .ZN(n15868) );
  NAND2_X1 U12984 ( .A1(n11672), .A2(n16676), .ZN(n16667) );
  NAND2_X1 U12985 ( .A1(n16676), .A2(n12916), .ZN(n11675) );
  OAI21_X1 U12986 ( .B1(n12916), .B2(n11674), .A(n16670), .ZN(n11673) );
  INV_X1 U12987 ( .A(n12950), .ZN(n11674) );
  NAND2_X1 U12988 ( .A1(n12116), .A2(n15124), .ZN(n11677) );
  NAND2_X1 U12989 ( .A1(n11677), .A2(n12548), .ZN(n12550) );
  NAND2_X1 U12990 ( .A1(n11677), .A2(n11240), .ZN(n11678) );
  NAND2_X1 U12991 ( .A1(n15025), .A2(n11679), .ZN(n15364) );
  NAND2_X1 U12992 ( .A1(n12414), .A2(n12203), .ZN(n11686) );
  XNOR2_X1 U12993 ( .A(n11691), .B(n11195), .ZN(n15886) );
  OAI21_X2 U12994 ( .B1(n11694), .B2(n11693), .A(n11692), .ZN(n11691) );
  INV_X1 U12995 ( .A(n15855), .ZN(n11693) );
  INV_X1 U12996 ( .A(n16858), .ZN(n11709) );
  NAND2_X1 U12997 ( .A1(n16069), .A2(n11726), .ZN(n16070) );
  NAND2_X1 U12998 ( .A1(n12407), .A2(n12201), .ZN(n12202) );
  NOR2_X1 U12999 ( .A1(n12092), .A2(n12101), .ZN(n12188) );
  OR2_X1 U13000 ( .A1(n14566), .A2(n14565), .ZN(n14568) );
  NOR2_X1 U13001 ( .A1(n14840), .A2(n14839), .ZN(n22668) );
  AOI21_X1 U13002 ( .B1(n15921), .B2(n20614), .A(n15847), .ZN(n15848) );
  INV_X1 U13003 ( .A(n15932), .ZN(n16150) );
  NAND2_X1 U13004 ( .A1(n15932), .A2(n14221), .ZN(n14334) );
  NOR2_X1 U13005 ( .A1(n22542), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11710) );
  INV_X1 U13006 ( .A(n15200), .ZN(n15331) );
  INV_X1 U13007 ( .A(n22456), .ZN(n22414) );
  OR2_X1 U13008 ( .A1(n12858), .A2(n19017), .ZN(n11711) );
  OR2_X1 U13009 ( .A1(n12895), .A2(n16692), .ZN(n11712) );
  INV_X1 U13010 ( .A(n16146), .ZN(n14221) );
  INV_X1 U13011 ( .A(n11143), .ZN(n15785) );
  AND2_X1 U13012 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11714) );
  AND4_X1 U13013 ( .A1(n13106), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n11715) );
  NAND2_X1 U13014 ( .A1(n14046), .A2(n12006), .ZN(n14045) );
  AND2_X1 U13015 ( .A1(n16578), .A2(n14694), .ZN(n11716) );
  AND2_X1 U13016 ( .A1(n13253), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11717) );
  INV_X1 U13017 ( .A(n22559), .ZN(n22607) );
  INV_X1 U13018 ( .A(n11958), .ZN(n11746) );
  OR4_X1 U13019 ( .A1(n17079), .A2(n17076), .A3(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A4(n17065), .ZN(n11718) );
  INV_X1 U13020 ( .A(n18917), .ZN(n19703) );
  OR2_X1 U13021 ( .A1(n13115), .A2(n14886), .ZN(n11719) );
  OR2_X1 U13022 ( .A1(n19256), .A2(n19255), .ZN(n11720) );
  AND2_X1 U13023 ( .A1(n15602), .A2(n15857), .ZN(n11721) );
  NOR2_X1 U13024 ( .A1(n17066), .A2(n15871), .ZN(n11722) );
  AND2_X1 U13025 ( .A1(n14211), .A2(n14210), .ZN(n11723) );
  OR2_X1 U13026 ( .A1(n22369), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19006) );
  AND2_X1 U13027 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11724) );
  AND2_X1 U13028 ( .A1(n13027), .A2(n13026), .ZN(n11725) );
  INV_X1 U13029 ( .A(n17873), .ZN(n17843) );
  INV_X1 U13030 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n15308) );
  AND2_X1 U13031 ( .A1(n14212), .A2(n14205), .ZN(n19298) );
  INV_X1 U13032 ( .A(n19298), .ZN(n14207) );
  INV_X1 U13033 ( .A(n12143), .ZN(n11860) );
  AND2_X2 U13034 ( .A1(n14694), .A2(n13032), .ZN(n13231) );
  INV_X1 U13035 ( .A(n14388), .ZN(n14442) );
  INV_X1 U13036 ( .A(n18697), .ZN(n18758) );
  NAND2_X1 U13037 ( .A1(n12012), .A2(n11955), .ZN(n12023) );
  AND2_X1 U13038 ( .A1(n13592), .A2(n13591), .ZN(n11726) );
  OR2_X1 U13039 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13847) );
  AND4_X1 U13040 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n11727) );
  INV_X1 U13041 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17416) );
  AND2_X2 U13042 ( .A1(n13047), .A2(n13046), .ZN(n13238) );
  AND4_X1 U13043 ( .A1(n13112), .A2(n13111), .A3(n13110), .A4(n13109), .ZN(
        n11729) );
  AND4_X1 U13044 ( .A1(n13057), .A2(n13056), .A3(n13055), .A4(n13054), .ZN(
        n11730) );
  AND2_X2 U13045 ( .A1(n14694), .A2(n16572), .ZN(n13253) );
  AND2_X1 U13046 ( .A1(n14696), .A2(n15914), .ZN(n11731) );
  AND2_X2 U13047 ( .A1(n13045), .A2(n14694), .ZN(n13237) );
  AND4_X1 U13048 ( .A1(n13061), .A2(n13060), .A3(n13059), .A4(n13058), .ZN(
        n11732) );
  INV_X1 U13049 ( .A(n13170), .ZN(n14556) );
  OAI22_X1 U13050 ( .A1(n17690), .A2(keyinput_26), .B1(n17689), .B2(DATAI_6_), 
        .ZN(n17691) );
  INV_X1 U13051 ( .A(n17691), .ZN(n17692) );
  XNOR2_X1 U13052 ( .A(READY1), .B(keyinput_36), .ZN(n17707) );
  AOI21_X1 U13053 ( .B1(n17709), .B2(n17708), .A(n17707), .ZN(n17710) );
  XNOR2_X1 U13054 ( .A(keyinput_84), .B(P1_EBX_REG_31__SCAN_IN), .ZN(n17765)
         );
  AOI21_X1 U13055 ( .B1(n17767), .B2(n17766), .A(n17765), .ZN(n17768) );
  INV_X1 U13056 ( .A(n17768), .ZN(n17769) );
  OAI211_X1 U13057 ( .C1(n17780), .C2(n17779), .A(n17778), .B(n17777), .ZN(
        n17786) );
  OR2_X1 U13058 ( .A1(n12182), .A2(n12940), .ZN(n12183) );
  OAI22_X1 U13059 ( .A1(n15312), .A2(keyinput_107), .B1(n17797), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n17798) );
  INV_X1 U13060 ( .A(n17798), .ZN(n17799) );
  OR2_X1 U13061 ( .A1(n13874), .A2(n13878), .ZN(n13860) );
  NAND2_X1 U13062 ( .A1(n12189), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12104) );
  AND2_X1 U13063 ( .A1(n14071), .A2(n12393), .ZN(n11974) );
  NAND2_X1 U13064 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11758) );
  OAI22_X1 U13065 ( .A1(n12239), .A2(n12120), .B1(n12174), .B2(n12119), .ZN(
        n12124) );
  AOI22_X1 U13066 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11959) );
  AND2_X1 U13067 ( .A1(n13864), .A2(n13863), .ZN(n13871) );
  OR2_X1 U13068 ( .A1(n13345), .A2(n13344), .ZN(n13957) );
  NAND2_X1 U13069 ( .A1(n12006), .A2(n11954), .ZN(n11977) );
  INV_X1 U13070 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11757) );
  INV_X1 U13071 ( .A(n12005), .ZN(n11954) );
  AND2_X1 U13072 ( .A1(n11921), .A2(n11920), .ZN(n11925) );
  AND2_X1 U13073 ( .A1(n13526), .A2(n15616), .ZN(n13527) );
  OR2_X1 U13074 ( .A1(n13387), .A2(n13386), .ZN(n13978) );
  OR2_X1 U13075 ( .A1(n13214), .A2(n13213), .ZN(n13215) );
  AND4_X1 U13076 ( .A1(n13036), .A2(n13035), .A3(n13034), .A4(n13033), .ZN(
        n13043) );
  INV_X1 U13077 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12538) );
  INV_X1 U13078 ( .A(n12160), .ZN(n12584) );
  AND3_X1 U13079 ( .A1(n11934), .A2(n11933), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11938) );
  INV_X1 U13080 ( .A(n18452), .ZN(n18451) );
  NAND2_X1 U13081 ( .A1(n13867), .A2(n13869), .ZN(n14414) );
  INV_X1 U13082 ( .A(n13914), .ZN(n13310) );
  INV_X1 U13083 ( .A(n15971), .ZN(n13780) );
  INV_X1 U13084 ( .A(n13643), .ZN(n13644) );
  INV_X1 U13085 ( .A(n13413), .ZN(n13414) );
  INV_X1 U13086 ( .A(n13293), .ZN(n13412) );
  AND2_X1 U13087 ( .A1(n14279), .A2(n14278), .ZN(n16138) );
  INV_X1 U13088 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13179) );
  OR2_X1 U13089 ( .A1(n13264), .A2(n13263), .ZN(n13927) );
  AND4_X1 U13090 ( .A1(n13051), .A2(n13050), .A3(n13049), .A4(n13048), .ZN(
        n13052) );
  NAND2_X1 U13091 ( .A1(n18721), .A2(n21833), .ZN(n18526) );
  AND2_X1 U13092 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18505), .ZN(
        n18507) );
  OR2_X1 U13093 ( .A1(n15168), .A2(n22108), .ZN(n15169) );
  AND3_X1 U13094 ( .A1(n13462), .A2(n13461), .A3(n13460), .ZN(n13463) );
  NAND2_X1 U13095 ( .A1(n13835), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13120) );
  NAND2_X1 U13096 ( .A1(n13800), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15170) );
  INV_X1 U13097 ( .A(n13412), .ZN(n13849) );
  AND2_X1 U13098 ( .A1(n13644), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13645) );
  INV_X1 U13099 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13465) );
  XNOR2_X1 U13100 ( .A(n13282), .B(n13283), .ZN(n14637) );
  AND2_X1 U13101 ( .A1(n14250), .A2(n14249), .ZN(n15258) );
  OAI21_X1 U13102 ( .B1(n16594), .B2(n16593), .A(n22595), .ZN(n16616) );
  OR2_X1 U13103 ( .A1(n14848), .A2(n22486), .ZN(n14785) );
  INV_X1 U13104 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22585) );
  AOI21_X1 U13105 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19898), .A(
        n11834), .ZN(n12380) );
  AND2_X1 U13106 ( .A1(n14150), .A2(n14149), .ZN(n17143) );
  AND2_X1 U13107 ( .A1(n14145), .A2(n14144), .ZN(n15637) );
  INV_X1 U13108 ( .A(n15550), .ZN(n14135) );
  OAI21_X1 U13109 ( .B1(n14761), .B2(n14760), .A(n14095), .ZN(n14096) );
  AND2_X1 U13110 ( .A1(n12361), .A2(n17111), .ZN(n16848) );
  AND2_X1 U13111 ( .A1(n17006), .A2(n17008), .ZN(n16993) );
  INV_X1 U13112 ( .A(n12399), .ZN(n14077) );
  AND2_X1 U13113 ( .A1(n13020), .A2(n14479), .ZN(n13021) );
  AND2_X1 U13114 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12551) );
  CLKBUF_X3 U13115 ( .A(n15725), .Z(n18455) );
  NAND2_X1 U13116 ( .A1(n18527), .A2(n18526), .ZN(n18528) );
  NOR2_X1 U13117 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18550), .ZN(
        n18802) );
  OR2_X1 U13118 ( .A1(n17409), .A2(n21197), .ZN(n15774) );
  INV_X1 U13119 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17392) );
  AND2_X1 U13120 ( .A1(n16021), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n16012) );
  NOR2_X1 U13121 ( .A1(n13545), .A2(n22234), .ZN(n13561) );
  NAND2_X1 U13122 ( .A1(n13312), .A2(n13311), .ZN(n14849) );
  INV_X1 U13123 ( .A(n22272), .ZN(n22249) );
  XNOR2_X1 U13124 ( .A(n13252), .B(n13251), .ZN(n13292) );
  NAND2_X1 U13125 ( .A1(n15910), .A2(n15163), .ZN(n14625) );
  AND2_X1 U13126 ( .A1(n16231), .A2(n14635), .ZN(n15824) );
  OR2_X1 U13127 ( .A1(n13693), .A2(n13692), .ZN(n13732) );
  NAND2_X1 U13128 ( .A1(n13561), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13574) );
  NOR2_X1 U13129 ( .A1(n13510), .A2(n13511), .ZN(n13496) );
  NOR2_X1 U13130 ( .A1(n13432), .A2(n13431), .ZN(n13449) );
  AND3_X1 U13131 ( .A1(n14540), .A2(n11614), .A3(n13857), .ZN(n14533) );
  INV_X1 U13132 ( .A(n20628), .ZN(n16384) );
  INV_X1 U13133 ( .A(n16318), .ZN(n16327) );
  NAND2_X1 U13134 ( .A1(n14557), .A2(n15904), .ZN(n22049) );
  INV_X1 U13135 ( .A(n14638), .ZN(n14778) );
  NOR2_X1 U13136 ( .A1(n22512), .A2(n14638), .ZN(n15214) );
  NOR3_X1 U13137 ( .A1(n14916), .A2(n22607), .A3(n22560), .ZN(n22612) );
  AND2_X1 U13138 ( .A1(n13936), .A2(n22486), .ZN(n14917) );
  INV_X1 U13139 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n22571) );
  AOI21_X1 U13140 ( .B1(n14640), .B2(n16559), .A(n22298), .ZN(n14792) );
  OR2_X1 U13141 ( .A1(n14785), .A2(n15213), .ZN(n22823) );
  NOR2_X1 U13142 ( .A1(n15794), .A2(n19140), .ZN(n16638) );
  INV_X1 U13143 ( .A(n11121), .ZN(n19210) );
  INV_X1 U13144 ( .A(n19237), .ZN(n19256) );
  INV_X1 U13145 ( .A(n16663), .ZN(n12953) );
  INV_X1 U13146 ( .A(n16667), .ZN(n16668) );
  AND4_X1 U13147 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n16718) );
  AND3_X1 U13148 ( .A1(n14126), .A2(n14125), .A3(n14124), .ZN(n14746) );
  NAND2_X1 U13149 ( .A1(n14109), .A2(n14108), .ZN(n14749) );
  INV_X1 U13150 ( .A(n12540), .ZN(n12541) );
  INV_X1 U13151 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19072) );
  AND2_X1 U13152 ( .A1(n16993), .A2(n16995), .ZN(n16956) );
  NOR2_X1 U13153 ( .A1(n17378), .A2(n19279), .ZN(n17295) );
  INV_X1 U13154 ( .A(n19292), .ZN(n17371) );
  INV_X1 U13155 ( .A(n14038), .ZN(n14060) );
  INV_X1 U13156 ( .A(n19928), .ZN(n19929) );
  NOR2_X1 U13157 ( .A1(n20291), .A2(n15037), .ZN(n20005) );
  INV_X1 U13158 ( .A(n20291), .ZN(n20009) );
  INV_X1 U13159 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19903) );
  INV_X1 U13160 ( .A(n21881), .ZN(n18484) );
  NOR2_X1 U13161 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n21022), .ZN(n21037) );
  NAND2_X1 U13162 ( .A1(n20941), .A2(n20912), .ZN(n21046) );
  NOR2_X1 U13163 ( .A1(n21432), .A2(n15737), .ZN(n20711) );
  INV_X1 U13164 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18619) );
  INV_X1 U13165 ( .A(n18721), .ZN(n21741) );
  INV_X1 U13166 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21743) );
  NAND2_X1 U13167 ( .A1(n18686), .A2(n18721), .ZN(n18685) );
  NOR2_X1 U13168 ( .A1(n18490), .A2(n18489), .ZN(n21410) );
  INV_X1 U13169 ( .A(n21815), .ZN(n21814) );
  OR2_X1 U13170 ( .A1(n21563), .A2(n18520), .ZN(n18769) );
  INV_X1 U13171 ( .A(n18481), .ZN(n18482) );
  INV_X1 U13172 ( .A(n21883), .ZN(n21487) );
  AOI21_X1 U13173 ( .B1(n21927), .B2(n18359), .A(n21428), .ZN(n19367) );
  NOR2_X1 U13174 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22559) );
  OR2_X1 U13175 ( .A1(n22214), .A2(n22190), .ZN(n22273) );
  INV_X1 U13176 ( .A(n22264), .ZN(n22251) );
  NOR2_X2 U13177 ( .A1(n15188), .A2(n15187), .ZN(n22214) );
  INV_X1 U13178 ( .A(n16227), .ZN(n16211) );
  AND2_X1 U13179 ( .A1(n15824), .A2(n15823), .ZN(n16229) );
  INV_X1 U13180 ( .A(n16231), .ZN(n16240) );
  OR2_X1 U13181 ( .A1(n16225), .A2(n15824), .ZN(n16241) );
  INV_X1 U13182 ( .A(n22414), .ZN(n22479) );
  NAND2_X1 U13183 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n13609), .ZN(
        n13643) );
  AOI21_X1 U13184 ( .B1(n16239), .B2(n16238), .A(n16237), .ZN(n22220) );
  NAND2_X1 U13185 ( .A1(n13409), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13432) );
  AND2_X1 U13186 ( .A1(n13353), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13397) );
  AND2_X1 U13187 ( .A1(n13853), .A2(n22559), .ZN(n20614) );
  NAND2_X1 U13188 ( .A1(n14531), .A2(n14530), .ZN(n14557) );
  NAND2_X1 U13189 ( .A1(n21956), .A2(n21955), .ZN(n22060) );
  INV_X1 U13190 ( .A(n22067), .ZN(n22098) );
  OR2_X1 U13191 ( .A1(n16550), .A2(n16548), .ZN(n22045) );
  INV_X1 U13192 ( .A(n14636), .ZN(n22593) );
  NOR2_X1 U13193 ( .A1(n14712), .A2(n13173), .ZN(n22298) );
  INV_X1 U13194 ( .A(n22490), .ZN(n22783) );
  INV_X1 U13195 ( .A(n22502), .ZN(n22789) );
  NOR2_X2 U13196 ( .A1(n22512), .A2(n22501), .ZN(n22796) );
  NOR2_X1 U13197 ( .A1(n22512), .A2(n22487), .ZN(n22795) );
  OAI211_X1 U13198 ( .C1(n22563), .C2(n14854), .A(n14850), .B(n22613), .ZN(
        n14877) );
  INV_X1 U13199 ( .A(n22526), .ZN(n22802) );
  AND2_X1 U13200 ( .A1(n14917), .A2(n22583), .ZN(n22803) );
  AND2_X1 U13201 ( .A1(n14917), .A2(n22554), .ZN(n15157) );
  INV_X1 U13202 ( .A(n11155), .ZN(n15213) );
  AND2_X1 U13203 ( .A1(n22556), .A2(n22593), .ZN(n22550) );
  NOR2_X1 U13204 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14792), .ZN(n14816) );
  INV_X1 U13205 ( .A(n22823), .ZN(n14828) );
  INV_X1 U13206 ( .A(n22646), .ZN(n22637) );
  INV_X1 U13207 ( .A(n22781), .ZN(n22772) );
  NOR2_X1 U13208 ( .A1(n16592), .A2(n22392), .ZN(n22642) );
  AND2_X1 U13209 ( .A1(n13936), .A2(n22488), .ZN(n22844) );
  AND2_X1 U13210 ( .A1(n15308), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13910) );
  INV_X1 U13211 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n17473) );
  INV_X1 U13212 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n22343) );
  INV_X1 U13213 ( .A(n20520), .ZN(n20515) );
  NAND2_X1 U13214 ( .A1(n19259), .A2(n19258), .ZN(n19260) );
  NOR2_X1 U13215 ( .A1(n15794), .A2(n19160), .ZN(n19179) );
  NOR2_X1 U13216 ( .A1(n19975), .A2(n19237), .ZN(n19253) );
  NOR2_X1 U13217 ( .A1(n15794), .A2(n19316), .ZN(n19265) );
  AND2_X1 U13218 ( .A1(n19012), .A2(n15393), .ZN(n19237) );
  INV_X1 U13219 ( .A(n19332), .ZN(n19014) );
  INV_X1 U13220 ( .A(n14477), .ZN(n14463) );
  AOI21_X1 U13221 ( .B1(n19252), .B2(n17870), .A(n15881), .ZN(n15884) );
  INV_X1 U13222 ( .A(n19294), .ZN(n19124) );
  OAI211_X1 U13223 ( .C1(n19269), .C2(n17371), .A(n15873), .B(n11718), .ZN(
        n15874) );
  AND2_X1 U13224 ( .A1(n14212), .A2(n14063), .ZN(n19292) );
  NOR2_X1 U13225 ( .A1(n11147), .A2(n17282), .ZN(n17030) );
  INV_X1 U13226 ( .A(n19302), .ZN(n17377) );
  AOI21_X1 U13227 ( .B1(n14060), .B2(n14059), .A(n19332), .ZN(n14212) );
  INV_X1 U13228 ( .A(n19941), .ZN(n19960) );
  OAI21_X1 U13229 ( .B1(n14485), .B2(n14484), .A(n14483), .ZN(n19842) );
  OAI21_X1 U13230 ( .B1(n20397), .B2(n20010), .A(n20009), .ZN(n20402) );
  INV_X1 U13231 ( .A(n20289), .ZN(n20398) );
  AND2_X1 U13232 ( .A1(n19998), .A2(n19957), .ZN(n20384) );
  INV_X1 U13233 ( .A(n20232), .ZN(n20371) );
  OR2_X1 U13234 ( .A1(n19924), .A2(n19923), .ZN(n20359) );
  NOR2_X1 U13235 ( .A1(n19956), .A2(n19929), .ZN(n20352) );
  AND2_X1 U13236 ( .A1(n19941), .A2(n17897), .ZN(n19928) );
  OR2_X1 U13237 ( .A1(n19842), .A2(n19836), .ZN(n19927) );
  NOR2_X2 U13238 ( .A1(n19885), .A2(n19956), .ZN(n20331) );
  NOR2_X1 U13239 ( .A1(n19885), .A2(n19855), .ZN(n20319) );
  INV_X1 U13240 ( .A(n20158), .ZN(n20160) );
  INV_X1 U13241 ( .A(n20164), .ZN(n20155) );
  NAND2_X1 U13242 ( .A1(n19960), .A2(n17897), .ZN(n19843) );
  INV_X1 U13243 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n22354) );
  NAND2_X1 U13244 ( .A1(n21932), .A2(n18484), .ZN(n20712) );
  NOR2_X1 U13245 ( .A1(n21116), .A2(n21115), .ZN(n21156) );
  INV_X1 U13246 ( .A(n21046), .ZN(n21076) );
  NOR2_X1 U13247 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20999), .ZN(n21015) );
  NOR2_X1 U13248 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20944), .ZN(n20959) );
  NOR2_X1 U13249 ( .A1(n20769), .A2(n20770), .ZN(n20941) );
  INV_X1 U13250 ( .A(n21168), .ZN(n21159) );
  INV_X1 U13251 ( .A(n20802), .ZN(n21179) );
  NOR2_X1 U13252 ( .A1(n18314), .A2(n18313), .ZN(n18329) );
  INV_X1 U13253 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20823) );
  NOR2_X1 U13254 ( .A1(n21299), .A2(n21300), .ZN(n21326) );
  NOR4_X1 U13255 ( .A1(n21344), .A2(n21293), .A3(n21292), .A4(n21291), .ZN(
        n21337) );
  NAND2_X1 U13256 ( .A1(n21345), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n21344) );
  NOR2_X1 U13257 ( .A1(n21369), .A2(n21249), .ZN(n21363) );
  NOR2_X1 U13258 ( .A1(n21244), .A2(n21243), .ZN(n21236) );
  INV_X1 U13259 ( .A(n21373), .ZN(n21376) );
  NOR2_X1 U13260 ( .A1(n20750), .A2(n20714), .ZN(n20732) );
  NOR2_X1 U13261 ( .A1(n18910), .A2(n18886), .ZN(n18697) );
  INV_X1 U13262 ( .A(n21817), .ZN(n21458) );
  NAND2_X1 U13263 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18550), .ZN(
        n21563) );
  NOR2_X1 U13264 ( .A1(n18519), .A2(n18819), .ZN(n21562) );
  NAND2_X1 U13265 ( .A1(n21744), .A2(n21743), .ZN(n21745) );
  INV_X2 U13266 ( .A(n21659), .ZN(n21831) );
  NOR2_X1 U13267 ( .A1(n21559), .A2(n21558), .ZN(n21614) );
  INV_X1 U13268 ( .A(n21617), .ZN(n21722) );
  NAND2_X1 U13269 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n21917), .ZN(n21937) );
  INV_X1 U13270 ( .A(n21926), .ZN(n21428) );
  INV_X1 U13271 ( .A(n19772), .ZN(n19782) );
  INV_X1 U13272 ( .A(n19629), .ZN(n19752) );
  AND2_X1 U13273 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19704), .ZN(n19485) );
  INV_X1 U13274 ( .A(n19712), .ZN(n19797) );
  INV_X1 U13275 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n21389) );
  AND2_X1 U13276 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22323), .ZN(n18997) );
  NAND2_X2 U13277 ( .A1(n14346), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n16158)
         );
  NOR2_X1 U13278 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14358), .ZN(n19360)
         );
  NAND2_X1 U13279 ( .A1(n15912), .A2(n14883), .ZN(n15165) );
  INV_X1 U13280 ( .A(n22255), .ZN(n22278) );
  INV_X1 U13281 ( .A(n22256), .ZN(n22268) );
  NAND2_X1 U13282 ( .A1(n20574), .A2(n15908), .ZN(n16143) );
  NAND2_X1 U13283 ( .A1(n15921), .A2(n15822), .ZN(n15826) );
  OAI21_X1 U13284 ( .B1(n16237), .B2(n16085), .A(n16084), .ZN(n16385) );
  INV_X1 U13285 ( .A(n20463), .ZN(n20481) );
  OR2_X1 U13286 ( .A1(n15165), .A2(n14493), .ZN(n22478) );
  INV_X1 U13287 ( .A(n20625), .ZN(n20634) );
  NAND2_X1 U13288 ( .A1(n14557), .A2(n14550), .ZN(n22067) );
  NAND2_X1 U13289 ( .A1(n14557), .A2(n14536), .ZN(n22084) );
  INV_X1 U13290 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U13291 ( .A1(n22491), .A2(n22497), .B1(n22493), .B2(n22544), .ZN(
        n22787) );
  AOI211_X2 U13292 ( .C1(n22607), .C2(n22492), .A(n15212), .B(n15211), .ZN(
        n15253) );
  AOI22_X1 U13293 ( .A1(n22504), .A2(n22508), .B1(n22544), .B2(n11710), .ZN(
        n22793) );
  AOI22_X1 U13294 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22519), .B1(n22521), 
        .B2(n22518), .ZN(n22800) );
  OR2_X1 U13295 ( .A1(n14851), .A2(n11155), .ZN(n22526) );
  OR2_X1 U13296 ( .A1(n14851), .A2(n15213), .ZN(n16588) );
  AOI22_X1 U13297 ( .A1(n22529), .A2(n22536), .B1(n11710), .B2(n22569), .ZN(
        n22807) );
  INV_X1 U13298 ( .A(n15157), .ZN(n17833) );
  INV_X1 U13299 ( .A(n15130), .ZN(n17834) );
  NAND2_X1 U13300 ( .A1(n14957), .A2(n15213), .ZN(n22540) );
  AOI22_X1 U13301 ( .A1(n22545), .A2(n22550), .B1(n22544), .B2(n22543), .ZN(
        n22813) );
  NAND2_X1 U13302 ( .A1(n22555), .A2(n22554), .ZN(n22820) );
  INV_X1 U13303 ( .A(n22609), .ZN(n22581) );
  INV_X1 U13304 ( .A(n22750), .ZN(n22744) );
  INV_X1 U13305 ( .A(n14784), .ZN(n14847) );
  NAND3_X1 U13306 ( .A1(n13936), .A2(n22583), .A3(n22582), .ZN(n22848) );
  NAND2_X1 U13307 ( .A1(n13910), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n22303) );
  INV_X1 U13308 ( .A(n22308), .ZN(n17432) );
  AND2_X1 U13309 ( .A1(n22343), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22853) );
  INV_X1 U13310 ( .A(n20510), .ZN(n22331) );
  OR2_X1 U13311 ( .A1(n15115), .A2(n14368), .ZN(n15399) );
  NAND2_X1 U13312 ( .A1(n15111), .A2(n19014), .ZN(n19335) );
  NAND2_X1 U13313 ( .A1(n15804), .A2(n15803), .ZN(n15814) );
  NAND2_X1 U13314 ( .A1(n15388), .A2(n15387), .ZN(n19215) );
  NAND2_X1 U13315 ( .A1(n14568), .A2(n14567), .ZN(n19941) );
  AND2_X1 U13316 ( .A1(n14509), .A2(n19014), .ZN(n15640) );
  NOR2_X1 U13317 ( .A1(n20119), .A2(n20117), .ZN(n20071) );
  INV_X1 U13318 ( .A(n20064), .ZN(n15004) );
  INV_X1 U13319 ( .A(n17915), .ZN(n17949) );
  OAI21_X1 U13320 ( .B1(n14367), .B2(n14368), .A(n14477), .ZN(n14388) );
  INV_X1 U13321 ( .A(n14442), .ZN(n14467) );
  NOR2_X1 U13322 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  OR2_X1 U13323 ( .A1(n19335), .A2(n19017), .ZN(n17873) );
  NAND2_X1 U13324 ( .A1(n19335), .A2(n12536), .ZN(n17877) );
  NAND2_X1 U13325 ( .A1(n14212), .A2(n15097), .ZN(n17351) );
  NAND2_X1 U13326 ( .A1(n14212), .A2(n15102), .ZN(n19302) );
  INV_X1 U13327 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19898) );
  INV_X1 U13328 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19273) );
  NAND2_X1 U13329 ( .A1(n19998), .A2(n19997), .ZN(n20289) );
  NAND2_X1 U13330 ( .A1(n19998), .A2(n19971), .ZN(n20394) );
  INV_X1 U13331 ( .A(n20384), .ZN(n20276) );
  NAND2_X1 U13332 ( .A1(n19998), .A2(n19942), .ZN(n20381) );
  NAND2_X1 U13333 ( .A1(n19928), .A2(n19971), .ZN(n20369) );
  INV_X1 U13334 ( .A(n20352), .ZN(n20363) );
  NAND2_X1 U13335 ( .A1(n19942), .A2(n19928), .ZN(n20356) );
  INV_X1 U13336 ( .A(n20338), .ZN(n20262) );
  AOI22_X1 U13337 ( .A1(n19877), .A2(n19880), .B1(n19876), .B2(n19875), .ZN(
        n20336) );
  INV_X1 U13338 ( .A(n20319), .ZN(n20329) );
  AOI22_X1 U13339 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20297), .ZN(n20062) );
  AOI22_X1 U13340 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20297), .ZN(n20290) );
  OR2_X1 U13341 ( .A1(n19843), .A2(n19920), .ZN(n20316) );
  OR2_X1 U13342 ( .A1(n19843), .A2(n19855), .ZN(n20405) );
  INV_X1 U13343 ( .A(n20300), .ZN(n20210) );
  INV_X1 U13344 ( .A(n22312), .ZN(n17413) );
  CLKBUF_X1 U13345 ( .A(n17975), .Z(n22351) );
  AOI21_X1 U13346 ( .B1(n21879), .B2(n21878), .A(n20712), .ZN(n20767) );
  OR2_X1 U13347 ( .A1(n21087), .A2(n21086), .ZN(n21116) );
  INV_X1 U13348 ( .A(n21161), .ZN(n21184) );
  OR3_X1 U13349 ( .A1(n21102), .A2(n20887), .A3(P3_REIP_REG_9__SCAN_IN), .ZN(
        n20895) );
  INV_X1 U13350 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20800) );
  AND2_X1 U13351 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18124), .ZN(n18111) );
  NOR2_X1 U13352 ( .A1(n18348), .A2(n21267), .ZN(n18352) );
  NAND2_X1 U13353 ( .A1(n21255), .A2(n21313), .ZN(n21341) );
  NOR2_X1 U13354 ( .A1(n21213), .A2(n21362), .ZN(n21217) );
  NOR2_X1 U13355 ( .A1(n18385), .A2(n18384), .ZN(n21223) );
  NOR2_X1 U13356 ( .A1(n18406), .A2(n18405), .ZN(n21248) );
  NOR2_X1 U13357 ( .A1(n21871), .A2(n18968), .ZN(n18979) );
  INV_X1 U13358 ( .A(n18968), .ZN(n18967) );
  INV_X1 U13359 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n21850) );
  INV_X1 U13360 ( .A(n18812), .ZN(n18829) );
  INV_X1 U13361 ( .A(n18904), .ZN(n18896) );
  INV_X1 U13362 ( .A(n21865), .ZN(n21790) );
  INV_X1 U13363 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21869) );
  NAND2_X1 U13364 ( .A1(n21822), .A2(n21808), .ZN(n21761) );
  INV_X1 U13365 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21903) );
  INV_X1 U13366 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19447) );
  INV_X1 U13367 ( .A(n19768), .ZN(n19679) );
  INV_X1 U13368 ( .A(n19746), .ZN(n19738) );
  INV_X1 U13369 ( .A(n19607), .ZN(n19602) );
  INV_X1 U13370 ( .A(n19484), .ZN(n19481) );
  INV_X1 U13371 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n21936) );
  INV_X1 U13372 ( .A(n22317), .ZN(n17404) );
  INV_X1 U13373 ( .A(n16158), .ZN(n15823) );
  NAND2_X1 U13374 ( .A1(n14334), .A2(n14333), .ZN(P1_U2842) );
  OAI21_X1 U13375 ( .B1(n17071), .B2(n17853), .A(n12545), .ZN(P2_U2984) );
  NAND2_X1 U13376 ( .A1(n11723), .A2(n11194), .ZN(P2_U3018) );
  AND2_X4 U13377 ( .A1(n11745), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11965) );
  AND2_X2 U13378 ( .A1(n12976), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12160) );
  NAND2_X1 U13379 ( .A1(n12976), .A2(n11777), .ZN(n11862) );
  INV_X2 U13380 ( .A(n11862), .ZN(n12782) );
  AOI22_X1 U13381 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11740) );
  AND2_X4 U13382 ( .A1(n11733), .A2(n11741), .ZN(n12979) );
  INV_X1 U13383 ( .A(n12150), .ZN(n12648) );
  INV_X1 U13384 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11734) );
  AND2_X4 U13385 ( .A1(n11743), .A2(n11757), .ZN(n11981) );
  AND2_X2 U13386 ( .A1(n12977), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12615) );
  AOI22_X1 U13387 ( .A1(n12648), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11739) );
  NAND3_X1 U13388 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12376) );
  INV_X1 U13389 ( .A(n12376), .ZN(n11735) );
  AOI22_X1 U13390 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11813), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11738) );
  AND2_X2 U13391 ( .A1(n12983), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12159) );
  NOR2_X1 U13392 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12376), .ZN(
        n12152) );
  AOI22_X1 U13393 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11737) );
  NAND4_X1 U13394 ( .A1(n11740), .A2(n11739), .A3(n11738), .A4(n11737), .ZN(
        n11752) );
  NOR2_X1 U13395 ( .A1(n11741), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11742) );
  AOI22_X1 U13396 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11837), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11750) );
  AND2_X1 U13397 ( .A1(n11743), .A2(n12820), .ZN(n11788) );
  AOI22_X1 U13398 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11749) );
  AND2_X2 U13399 ( .A1(n12973), .A2(n11777), .ZN(n12846) );
  AND2_X2 U13400 ( .A1(n12984), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12161) );
  AOI22_X1 U13401 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12161), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11748) );
  NAND2_X2 U13402 ( .A1(n12978), .A2(n11777), .ZN(n12837) );
  INV_X1 U13403 ( .A(n12837), .ZN(n12686) );
  AND2_X2 U13404 ( .A1(n15085), .A2(n11777), .ZN(n12143) );
  AOI22_X1 U13405 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11747) );
  NAND4_X1 U13406 ( .A1(n11750), .A2(n11749), .A3(n11748), .A4(n11747), .ZN(
        n11751) );
  NOR2_X1 U13407 ( .A1(n11752), .A2(n11751), .ZN(n12400) );
  AOI22_X1 U13408 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U13409 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U13410 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11133), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U13411 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U13412 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U13413 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11760) );
  INV_X2 U13414 ( .A(n11146), .ZN(n15857) );
  OR2_X1 U13415 ( .A1(n12400), .A2(n15857), .ZN(n14070) );
  INV_X1 U13416 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14486) );
  INV_X1 U13417 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14474) );
  NAND3_X1 U13418 ( .A1(n15857), .A2(n14486), .A3(n14474), .ZN(n11763) );
  NAND2_X1 U13419 ( .A1(n14070), .A2(n11763), .ZN(n12217) );
  AOI22_X1 U13420 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11964), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11766) );
  AOI22_X1 U13421 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U13422 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11133), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U13423 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11133), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11769) );
  AOI22_X1 U13424 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11768) );
  AOI22_X1 U13425 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11771) );
  AOI22_X1 U13426 ( .A1(n11958), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11964), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11770) );
  INV_X2 U13427 ( .A(n11772), .ZN(n11987) );
  AOI22_X1 U13428 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11776) );
  AOI22_X1 U13429 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U13430 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U13431 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11773) );
  NAND4_X1 U13432 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11778) );
  AOI22_X1 U13433 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11782) );
  AOI22_X1 U13434 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11781) );
  AOI22_X1 U13435 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11780) );
  AOI22_X1 U13436 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11779) );
  NAND4_X1 U13437 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  NAND2_X1 U13438 ( .A1(n11783), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11784) );
  INV_X1 U13439 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11787) );
  INV_X1 U13440 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11786) );
  OAI22_X1 U13441 ( .A1(n12150), .A2(n11787), .B1(n12837), .B2(n11786), .ZN(
        n11794) );
  NAND2_X1 U13442 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11792) );
  NAND2_X1 U13443 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U13444 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11790) );
  AOI22_X1 U13445 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U13446 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  NOR2_X1 U13447 ( .A1(n11794), .A2(n11793), .ZN(n11802) );
  AOI22_X1 U13448 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U13449 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11798) );
  NAND2_X1 U13450 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11797) );
  NAND2_X1 U13451 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U13452 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n11795) );
  AND4_X1 U13453 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11800) );
  AOI22_X1 U13454 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U13455 ( .A1(n15383), .A2(n14089), .ZN(n11810) );
  NAND2_X1 U13456 ( .A1(n12999), .A2(n12381), .ZN(n11804) );
  NAND2_X1 U13457 ( .A1(n19985), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U13458 ( .A1(n11804), .A2(n11803), .ZN(n11808) );
  INV_X1 U13459 ( .A(n11808), .ZN(n11806) );
  XNOR2_X1 U13460 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11807) );
  INV_X1 U13461 ( .A(n11807), .ZN(n11805) );
  NAND2_X1 U13462 ( .A1(n11806), .A2(n11805), .ZN(n11809) );
  NAND2_X1 U13463 ( .A1(n11808), .A2(n11807), .ZN(n11830) );
  AND2_X1 U13464 ( .A1(n11809), .A2(n11830), .ZN(n12998) );
  NAND2_X1 U13465 ( .A1(n12031), .A2(n12998), .ZN(n13009) );
  NAND2_X1 U13466 ( .A1(n11810), .A2(n13009), .ZN(n11811) );
  INV_X1 U13467 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n15410) );
  INV_X1 U13468 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12097) );
  INV_X1 U13469 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11812) );
  OAI22_X1 U13470 ( .A1(n12150), .A2(n12097), .B1(n12837), .B2(n11812), .ZN(
        n11819) );
  NAND2_X1 U13471 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U13472 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U13473 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11815) );
  AOI22_X1 U13474 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11814) );
  NAND4_X1 U13475 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11818) );
  NOR2_X1 U13476 ( .A1(n11819), .A2(n11818), .ZN(n11828) );
  AOI22_X1 U13477 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11827) );
  INV_X1 U13478 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12120) );
  INV_X1 U13479 ( .A(n12162), .ZN(n11878) );
  INV_X1 U13480 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11820) );
  OAI22_X1 U13481 ( .A1(n12584), .A2(n12120), .B1(n11878), .B2(n11820), .ZN(
        n11824) );
  INV_X1 U13482 ( .A(n12161), .ZN(n11881) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12754) );
  NAND2_X1 U13484 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U13485 ( .A1(n12795), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11821) );
  OAI211_X1 U13486 ( .C1(n11881), .C2(n12754), .A(n11822), .B(n11821), .ZN(
        n11823) );
  NOR2_X1 U13487 ( .A1(n11824), .A2(n11823), .ZN(n11826) );
  AOI22_X1 U13488 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U13489 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n14100) );
  NAND2_X1 U13490 ( .A1(n19871), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11829) );
  XNOR2_X1 U13491 ( .A(n11831), .B(n11832), .ZN(n13011) );
  MUX2_X1 U13492 ( .A(n14100), .B(n13011), .S(n12031), .Z(n12387) );
  INV_X1 U13493 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12071) );
  MUX2_X1 U13494 ( .A(n12387), .B(n12071), .S(n15857), .Z(n12212) );
  NAND3_X1 U13495 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12380), .A3(
        n19273), .ZN(n12995) );
  INV_X1 U13496 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11836) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11835) );
  OAI22_X1 U13498 ( .A1(n12150), .A2(n11836), .B1(n12837), .B2(n11835), .ZN(
        n11843) );
  NAND2_X1 U13499 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U13500 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U13501 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11839) );
  AOI22_X1 U13502 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11838) );
  NAND4_X1 U13503 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n11842) );
  NOR2_X1 U13504 ( .A1(n11843), .A2(n11842), .ZN(n11851) );
  AOI22_X1 U13505 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U13506 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11847) );
  NAND2_X1 U13507 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U13508 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U13509 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11844) );
  AOI22_X1 U13510 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11848) );
  NAND4_X1 U13511 ( .A1(n11851), .A2(n11850), .A3(n11849), .A4(n11848), .ZN(
        n14066) );
  MUX2_X1 U13512 ( .A(n12995), .B(n14066), .S(n15383), .Z(n12388) );
  INV_X1 U13513 ( .A(n12388), .ZN(n11852) );
  MUX2_X1 U13514 ( .A(n11852), .B(P2_EBX_REG_4__SCAN_IN), .S(n15857), .Z(
        n12207) );
  INV_X1 U13515 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n12445) );
  INV_X1 U13516 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12190) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11853) );
  OAI22_X1 U13518 ( .A1(n12150), .A2(n12190), .B1(n12837), .B2(n11853), .ZN(
        n11859) );
  NAND2_X1 U13519 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U13520 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U13521 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11855) );
  AOI22_X1 U13522 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11854) );
  NAND4_X1 U13523 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11858) );
  NOR2_X1 U13524 ( .A1(n11859), .A2(n11858), .ZN(n11870) );
  AOI22_X1 U13525 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11869) );
  INV_X1 U13526 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11861) );
  INV_X1 U13527 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12657) );
  OAI22_X1 U13528 ( .A1(n11862), .A2(n11861), .B1(n11860), .B2(n12657), .ZN(
        n11866) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U13530 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U13531 ( .A1(n12795), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11863) );
  OAI211_X1 U13532 ( .C1(n12584), .C2(n12176), .A(n11864), .B(n11863), .ZN(
        n11865) );
  NOR2_X1 U13533 ( .A1(n11866), .A2(n11865), .ZN(n11868) );
  AOI22_X1 U13534 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12162), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11867) );
  NAND4_X1 U13535 ( .A1(n11870), .A2(n11869), .A3(n11868), .A4(n11867), .ZN(
        n14103) );
  MUX2_X1 U13536 ( .A(n12445), .B(n14103), .S(n14065), .Z(n12205) );
  INV_X1 U13537 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19044) );
  INV_X1 U13538 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12248) );
  INV_X1 U13539 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11871) );
  OAI22_X1 U13540 ( .A1(n12150), .A2(n12248), .B1(n12837), .B2(n11871), .ZN(
        n11877) );
  NAND2_X1 U13541 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11875) );
  NAND2_X1 U13542 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11874) );
  NAND2_X1 U13543 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11873) );
  AOI22_X1 U13544 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U13545 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  NOR2_X1 U13546 ( .A1(n11877), .A2(n11876), .ZN(n11887) );
  AOI22_X1 U13547 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11886) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12240) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12243) );
  OAI22_X1 U13550 ( .A1(n12584), .A2(n12240), .B1(n11878), .B2(n12243), .ZN(
        n11883) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12804) );
  NAND2_X1 U13552 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11880) );
  NAND2_X1 U13553 ( .A1(n12795), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11879) );
  OAI211_X1 U13554 ( .C1(n11881), .C2(n12804), .A(n11880), .B(n11879), .ZN(
        n11882) );
  NOR2_X1 U13555 ( .A1(n11883), .A2(n11882), .ZN(n11885) );
  AOI22_X1 U13556 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11884) );
  NAND4_X1 U13557 ( .A1(n11887), .A2(n11886), .A3(n11885), .A4(n11884), .ZN(
        n14107) );
  MUX2_X1 U13558 ( .A(n19044), .B(n14107), .S(n14065), .Z(n12261) );
  NAND2_X1 U13559 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11891) );
  NAND2_X1 U13560 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11890) );
  NAND2_X1 U13561 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11889) );
  NAND2_X1 U13562 ( .A1(n12143), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11888) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11893) );
  INV_X1 U13564 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11892) );
  OAI22_X1 U13565 ( .A1(n12150), .A2(n11893), .B1(n12837), .B2(n11892), .ZN(
        n11899) );
  NAND2_X1 U13566 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11897) );
  NAND2_X1 U13567 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11896) );
  NAND2_X1 U13568 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11895) );
  AOI22_X1 U13569 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11894) );
  NAND4_X1 U13570 ( .A1(n11897), .A2(n11896), .A3(n11895), .A4(n11894), .ZN(
        n11898) );
  NOR2_X1 U13571 ( .A1(n11899), .A2(n11898), .ZN(n11905) );
  AOI22_X1 U13572 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11903) );
  NAND2_X1 U13573 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11902) );
  NAND2_X1 U13574 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11901) );
  NAND2_X1 U13575 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11900) );
  AND3_X2 U13576 ( .A1(n11906), .A2(n11905), .A3(n11904), .ZN(n12203) );
  MUX2_X1 U13577 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12203), .S(n14065), .Z(
        n12266) );
  NAND2_X1 U13578 ( .A1(n15857), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12269) );
  INV_X1 U13579 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12462) );
  INV_X1 U13580 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n11907) );
  NOR2_X1 U13581 ( .A1(n14065), .A2(n11907), .ZN(n12282) );
  OR2_X2 U13582 ( .A1(n12284), .A2(n12282), .ZN(n12278) );
  INV_X1 U13583 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12469) );
  NOR2_X4 U13584 ( .A1(n12278), .A2(n12277), .ZN(n12287) );
  NAND2_X1 U13585 ( .A1(n15857), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12286) );
  INV_X1 U13586 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11908) );
  NOR2_X1 U13587 ( .A1(n14065), .A2(n11908), .ZN(n12301) );
  INV_X1 U13588 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n15549) );
  NOR2_X1 U13589 ( .A1(n14065), .A2(n15549), .ZN(n12304) );
  NAND2_X1 U13590 ( .A1(n15857), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12299) );
  INV_X1 U13591 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12487) );
  NOR2_X1 U13592 ( .A1(n14065), .A2(n12487), .ZN(n12308) );
  INV_X1 U13593 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12491) );
  NOR2_X1 U13594 ( .A1(n14065), .A2(n12491), .ZN(n12311) );
  NOR2_X2 U13595 ( .A1(n12313), .A2(n12311), .ZN(n12296) );
  NAND2_X1 U13596 ( .A1(n15857), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U13597 ( .A1(n15857), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12291) );
  INV_X1 U13598 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16646) );
  NOR2_X1 U13599 ( .A1(n14065), .A2(n16646), .ZN(n12325) );
  INV_X1 U13600 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n11909) );
  INV_X1 U13601 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12510) );
  NOR2_X1 U13602 ( .A1(n14065), .A2(n12510), .ZN(n12341) );
  INV_X1 U13603 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n11910) );
  NOR2_X1 U13604 ( .A1(n14065), .A2(n11910), .ZN(n12346) );
  INV_X1 U13605 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n11911) );
  NOR2_X1 U13606 ( .A1(n14065), .A2(n11911), .ZN(n12355) );
  NAND2_X1 U13607 ( .A1(n15857), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U13608 ( .A1(n15857), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11912) );
  NOR2_X1 U13609 ( .A1(n11913), .A2(n11912), .ZN(n11914) );
  OR2_X1 U13610 ( .A1(n12366), .A2(n11914), .ZN(n19216) );
  AOI22_X1 U13611 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U13612 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11915) );
  AND3_X1 U13613 ( .A1(n11916), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11915), .ZN(n11919) );
  AOI22_X1 U13614 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11917) );
  NAND3_X1 U13615 ( .A1(n11919), .A2(n11918), .A3(n11917), .ZN(n11927) );
  AOI21_X1 U13616 ( .B1(n11980), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U13617 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U13618 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U13619 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11922) );
  NAND4_X1 U13620 ( .A1(n11925), .A2(n11924), .A3(n11923), .A4(n11922), .ZN(
        n11926) );
  AOI22_X1 U13621 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11928) );
  AND2_X1 U13622 ( .A1(n11928), .A2(n11777), .ZN(n11932) );
  AOI22_X1 U13623 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U13624 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U13625 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11929) );
  NAND4_X1 U13626 ( .A1(n11932), .A2(n11931), .A3(n11930), .A4(n11929), .ZN(
        n11940) );
  NAND2_X1 U13627 ( .A1(n11980), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11934) );
  AOI22_X1 U13628 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U13629 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U13630 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U13631 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  AOI22_X1 U13632 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U13633 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11942) );
  AND2_X1 U13634 ( .A1(n11942), .A2(n11941), .ZN(n11944) );
  AOI22_X1 U13635 ( .A1(n11957), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11943) );
  NAND3_X1 U13636 ( .A1(n11945), .A2(n11944), .A3(n11943), .ZN(n11946) );
  NAND2_X1 U13637 ( .A1(n11946), .A2(n11777), .ZN(n11953) );
  AOI22_X1 U13638 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n11965), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U13639 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U13640 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U13641 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11980), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U13642 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NAND2_X1 U13643 ( .A1(n11951), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11952) );
  NAND2_X1 U13644 ( .A1(n12007), .A2(n12023), .ZN(n14046) );
  NAND2_X1 U13645 ( .A1(n11954), .A2(n12022), .ZN(n14043) );
  INV_X1 U13646 ( .A(n14043), .ZN(n11956) );
  AOI21_X1 U13647 ( .B1(n14045), .B2(n11977), .A(n11956), .ZN(n11973) );
  AOI22_X1 U13648 ( .A1(n11957), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11958), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U13649 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U13650 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11986), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U13651 ( .A1(n11962), .A2(n11961), .A3(n11960), .A4(n11959), .ZN(
        n11963) );
  NAND2_X1 U13652 ( .A1(n11963), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11972) );
  AOI22_X1 U13653 ( .A1(n11964), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U13654 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U13655 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U13656 ( .A1(n11965), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11966) );
  NAND4_X1 U13657 ( .A1(n11969), .A2(n11968), .A3(n11967), .A4(n11966), .ZN(
        n11970) );
  NAND2_X1 U13658 ( .A1(n11970), .A2(n11777), .ZN(n11971) );
  MUX2_X2 U13659 ( .A(n14174), .B(n11973), .S(n14178), .Z(n12043) );
  NAND2_X1 U13660 ( .A1(n11975), .A2(n11974), .ZN(n12044) );
  NAND2_X1 U13661 ( .A1(n12044), .A2(n20294), .ZN(n12003) );
  NAND2_X1 U13662 ( .A1(n11977), .A2(n11976), .ZN(n11979) );
  NAND2_X1 U13663 ( .A1(n12022), .A2(n14178), .ZN(n11978) );
  NAND2_X1 U13664 ( .A1(n11979), .A2(n11978), .ZN(n11998) );
  AOI22_X1 U13665 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U13666 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U13667 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11983) );
  NAND3_X1 U13668 ( .A1(n11217), .A2(n11984), .A3(n11983), .ZN(n11995) );
  AOI22_X1 U13669 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11985), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U13670 ( .A1(n11981), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11134), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U13671 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11987), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U13672 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11988), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11989) );
  NAND4_X1 U13673 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  NAND2_X1 U13674 ( .A1(n12007), .A2(n20206), .ZN(n11996) );
  OAI21_X1 U13675 ( .B1(n11998), .B2(n11996), .A(n20294), .ZN(n11997) );
  INV_X1 U13676 ( .A(n11997), .ZN(n12002) );
  INV_X1 U13677 ( .A(n11998), .ZN(n12001) );
  NAND3_X1 U13678 ( .A1(n12005), .A2(n12006), .A3(n11146), .ZN(n11999) );
  OAI21_X1 U13679 ( .B1(n12043), .B2(n12031), .A(n12046), .ZN(n12004) );
  NAND2_X1 U13680 ( .A1(n12004), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12010) );
  INV_X1 U13681 ( .A(n14053), .ZN(n14031) );
  INV_X1 U13682 ( .A(n12007), .ZN(n12008) );
  NAND2_X1 U13683 ( .A1(n11213), .A2(n12008), .ZN(n12386) );
  NAND3_X1 U13684 ( .A1(n12386), .A2(n20206), .A3(n19017), .ZN(n12009) );
  NAND2_X1 U13685 ( .A1(n14031), .A2(n12009), .ZN(n13023) );
  NAND2_X1 U13686 ( .A1(n12065), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12020) );
  INV_X1 U13687 ( .A(n14041), .ZN(n12015) );
  NAND2_X1 U13688 ( .A1(n14175), .A2(n11721), .ZN(n12014) );
  NAND2_X1 U13689 ( .A1(n12015), .A2(n12014), .ZN(n12021) );
  INV_X1 U13690 ( .A(n12021), .ZN(n12017) );
  INV_X1 U13691 ( .A(n15122), .ZN(n12016) );
  NAND2_X1 U13692 ( .A1(n19322), .A2(n17416), .ZN(n19309) );
  NOR2_X1 U13693 ( .A1(n19309), .A2(n19985), .ZN(n12018) );
  NAND2_X1 U13694 ( .A1(n12021), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12029) );
  INV_X1 U13695 ( .A(n12022), .ZN(n14078) );
  MUX2_X1 U13696 ( .A(n14078), .B(n12024), .S(n20166), .Z(n12025) );
  INV_X1 U13697 ( .A(n11977), .ZN(n14047) );
  INV_X1 U13698 ( .A(n14361), .ZN(n12027) );
  NAND3_X2 U13699 ( .A1(n12029), .A2(n12040), .A3(n12028), .ZN(n12069) );
  NAND2_X1 U13700 ( .A1(n12069), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12036) );
  INV_X1 U13701 ( .A(n12031), .ZN(n12032) );
  INV_X1 U13702 ( .A(n12527), .ZN(n12034) );
  AOI22_X1 U13703 ( .A1(n12034), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12035) );
  INV_X1 U13704 ( .A(n14064), .ZN(n15109) );
  INV_X1 U13705 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17053) );
  NAND2_X1 U13706 ( .A1(n15383), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12037) );
  NOR2_X1 U13707 ( .A1(n12037), .A2(n12030), .ZN(n12038) );
  INV_X1 U13708 ( .A(n12527), .ZN(n12440) );
  OAI22_X1 U13709 ( .A1(n12065), .A2(n12038), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n12440), .ZN(n12042) );
  INV_X1 U13710 ( .A(n19309), .ZN(n12066) );
  NAND2_X1 U13711 ( .A1(n12066), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U13712 ( .A1(n12042), .A2(n12041), .ZN(n12082) );
  NAND2_X1 U13713 ( .A1(n12069), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12054) );
  INV_X1 U13714 ( .A(n12043), .ZN(n12045) );
  NAND2_X1 U13715 ( .A1(n12045), .A2(n12044), .ZN(n14166) );
  NAND2_X1 U13716 ( .A1(n14166), .A2(n12046), .ZN(n12047) );
  NAND2_X1 U13717 ( .A1(n12047), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12053) );
  INV_X1 U13718 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n14423) );
  OAI21_X1 U13719 ( .B1(n12441), .B2(n14423), .A(n12048), .ZN(n12051) );
  NAND2_X1 U13720 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12049) );
  OAI211_X1 U13721 ( .C1(n12527), .C2(n14474), .A(n19309), .B(n12049), .ZN(
        n12050) );
  NOR2_X1 U13722 ( .A1(n12051), .A2(n12050), .ZN(n12052) );
  NAND3_X1 U13723 ( .A1(n12054), .A2(n12053), .A3(n12052), .ZN(n12081) );
  NAND2_X1 U13724 ( .A1(n12084), .A2(n12085), .ZN(n12089) );
  NAND2_X1 U13725 ( .A1(n12089), .A2(n12055), .ZN(n12078) );
  NAND2_X1 U13726 ( .A1(n12065), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12057) );
  AOI21_X1 U13727 ( .B1(n19322), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U13728 ( .A1(n12057), .A2(n12056), .ZN(n12062) );
  INV_X1 U13729 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U13730 ( .A1(n12069), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12059) );
  AOI22_X1 U13731 ( .A1(n12440), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12058) );
  OAI211_X1 U13732 ( .C1(n12441), .C2(n12060), .A(n12059), .B(n12058), .ZN(
        n12061) );
  OR2_X2 U13733 ( .A1(n12062), .A2(n12061), .ZN(n12064) );
  NAND2_X1 U13734 ( .A1(n12062), .A2(n12061), .ZN(n12063) );
  AND2_X2 U13735 ( .A1(n12064), .A2(n12063), .ZN(n12079) );
  NAND2_X1 U13736 ( .A1(n12065), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12068) );
  NAND2_X1 U13737 ( .A1(n12066), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12067) );
  NAND2_X1 U13738 ( .A1(n12068), .A2(n12067), .ZN(n12076) );
  INV_X1 U13739 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12070) );
  INV_X1 U13740 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n15268) );
  NAND2_X1 U13741 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12073) );
  OR2_X1 U13742 ( .A1(n12527), .A2(n12071), .ZN(n12072) );
  NAND2_X1 U13743 ( .A1(n12076), .A2(n12075), .ZN(n12077) );
  XNOR2_X2 U13744 ( .A(n12080), .B(n12079), .ZN(n12095) );
  NOR2_X1 U13745 ( .A1(n15076), .A2(n12086), .ZN(n12117) );
  INV_X1 U13746 ( .A(n12117), .ZN(n12108) );
  NOR2_X2 U13747 ( .A1(n12092), .A2(n12108), .ZN(n19993) );
  INV_X1 U13748 ( .A(n12085), .ZN(n12088) );
  INV_X1 U13749 ( .A(n12086), .ZN(n12087) );
  NAND2_X1 U13750 ( .A1(n12088), .A2(n12087), .ZN(n12091) );
  NAND2_X1 U13751 ( .A1(n19029), .A2(n15076), .ZN(n12101) );
  AOI22_X1 U13752 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19993), .B1(
        n12188), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12094) );
  INV_X1 U13753 ( .A(n15076), .ZN(n19276) );
  OR2_X1 U13754 ( .A1(n19029), .A2(n19276), .ZN(n12107) );
  NOR2_X2 U13755 ( .A1(n12092), .A2(n12107), .ZN(n20012) );
  AOI22_X1 U13756 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20012), .B1(
        n12187), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U13757 ( .A1(n12094), .A2(n12093), .ZN(n12106) );
  INV_X1 U13758 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12100) );
  NOR2_X2 U13759 ( .A1(n12109), .A2(n12101), .ZN(n12189) );
  NOR2_X2 U13760 ( .A1(n12109), .A2(n12102), .ZN(n19911) );
  NAND2_X1 U13761 ( .A1(n19911), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U13762 ( .A1(n19852), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12113) );
  NAND2_X1 U13763 ( .A1(n19902), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12112) );
  NAND3_X1 U13764 ( .A1(n12113), .A2(n12112), .A3(n19017), .ZN(n12114) );
  NOR2_X1 U13765 ( .A1(n12115), .A2(n12114), .ZN(n12126) );
  NAND2_X1 U13766 ( .A1(n11211), .A2(n12110), .ZN(n12174) );
  INV_X1 U13767 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12119) );
  NAND2_X1 U13768 ( .A1(n11211), .A2(n12098), .ZN(n12178) );
  INV_X1 U13769 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12122) );
  OAI22_X1 U13770 ( .A1(n12754), .A2(n12177), .B1(n12178), .B2(n12122), .ZN(
        n12123) );
  NOR2_X1 U13771 ( .A1(n12124), .A2(n12123), .ZN(n12125) );
  NAND3_X1 U13772 ( .A1(n12127), .A2(n12126), .A3(n12125), .ZN(n12130) );
  INV_X1 U13773 ( .A(n14100), .ZN(n12128) );
  INV_X1 U13774 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12722) );
  INV_X1 U13775 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12131) );
  OAI22_X1 U13776 ( .A1(n12722), .A2(n12177), .B1(n12174), .B2(n12131), .ZN(
        n12134) );
  INV_X1 U13777 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12132) );
  INV_X1 U13778 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15052) );
  OAI22_X1 U13779 ( .A1(n12132), .A2(n19828), .B1(n12178), .B2(n15052), .ZN(
        n12133) );
  NOR2_X1 U13780 ( .A1(n12134), .A2(n12133), .ZN(n12138) );
  AOI21_X1 U13781 ( .B1(n19838), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n15109), .ZN(n12137) );
  INV_X1 U13782 ( .A(n12182), .ZN(n19852) );
  AOI22_X1 U13783 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19852), .B1(
        n19902), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12136) );
  NAND2_X1 U13784 ( .A1(n19930), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12135) );
  NAND4_X1 U13785 ( .A1(n12138), .A2(n12137), .A3(n12136), .A4(n12135), .ZN(
        n12173) );
  AOI22_X1 U13786 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19993), .B1(
        n12187), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U13787 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19950), .B1(
        n19911), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U13788 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12188), .B1(
        n12189), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U13789 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20012), .B1(
        n19878), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12139) );
  NAND4_X1 U13790 ( .A1(n12142), .A2(n12141), .A3(n12140), .A4(n12139), .ZN(
        n12172) );
  NAND2_X1 U13791 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12147) );
  NAND2_X1 U13792 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12146) );
  NAND2_X1 U13793 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12145) );
  NAND2_X1 U13794 ( .A1(n12143), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12144) );
  AND4_X1 U13795 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12169) );
  INV_X1 U13796 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12149) );
  INV_X1 U13797 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12148) );
  OAI22_X1 U13798 ( .A1(n12150), .A2(n12149), .B1(n12837), .B2(n12148), .ZN(
        n12158) );
  NAND2_X1 U13799 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12156) );
  NAND2_X1 U13800 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12155) );
  NAND2_X1 U13801 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12154) );
  INV_X1 U13802 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U13803 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12152), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12153) );
  NAND4_X1 U13804 ( .A1(n12156), .A2(n12155), .A3(n12154), .A4(n12153), .ZN(
        n12157) );
  NOR2_X1 U13805 ( .A1(n12158), .A2(n12157), .ZN(n12168) );
  AOI22_X1 U13806 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U13807 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12165) );
  NAND2_X1 U13808 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12164) );
  NAND2_X1 U13809 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12163) );
  AND4_X1 U13810 ( .A1(n12166), .A2(n12165), .A3(n12164), .A4(n12163), .ZN(
        n12167) );
  NAND2_X1 U13811 ( .A1(n14077), .A2(n15109), .ZN(n14420) );
  OR2_X1 U13812 ( .A1(n12400), .A2(n14420), .ZN(n12397) );
  INV_X1 U13813 ( .A(n14089), .ZN(n12170) );
  NAND2_X1 U13814 ( .A1(n12397), .A2(n12170), .ZN(n12171) );
  INV_X1 U13815 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12175) );
  OAI22_X1 U13816 ( .A1(n12176), .A2(n12239), .B1(n12174), .B2(n12175), .ZN(
        n12180) );
  INV_X1 U13817 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12787) );
  INV_X1 U13818 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12658) );
  OAI22_X1 U13819 ( .A1(n12787), .A2(n12177), .B1(n12178), .B2(n12658), .ZN(
        n12179) );
  NOR2_X1 U13820 ( .A1(n12180), .A2(n12179), .ZN(n12186) );
  AOI22_X1 U13821 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19930), .B1(
        n19950), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12185) );
  OR2_X1 U13822 ( .A1(n12181), .A2(n12657), .ZN(n12184) );
  INV_X1 U13823 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U13824 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12187), .B1(
        n20012), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U13825 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19976), .B1(
        n19993), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U13826 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12189), .B1(
        n19911), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12194) );
  INV_X1 U13827 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12191) );
  OAI22_X1 U13828 ( .A1(n12191), .A2(n19873), .B1(n19828), .B2(n12190), .ZN(
        n12192) );
  INV_X1 U13829 ( .A(n12192), .ZN(n12193) );
  NAND2_X1 U13830 ( .A1(n11727), .A2(n11201), .ZN(n12199) );
  INV_X1 U13831 ( .A(n14103), .ZN(n12197) );
  NAND2_X1 U13832 ( .A1(n12197), .A2(n15109), .ZN(n12198) );
  NAND2_X1 U13833 ( .A1(n12199), .A2(n12198), .ZN(n12201) );
  INV_X1 U13834 ( .A(n12201), .ZN(n12200) );
  INV_X1 U13835 ( .A(n12262), .ZN(n12204) );
  OAI21_X1 U13836 ( .B1(n12206), .B2(n12205), .A(n12204), .ZN(n19034) );
  INV_X1 U13837 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15522) );
  XNOR2_X1 U13838 ( .A(n12235), .B(n15522), .ZN(n15505) );
  INV_X1 U13839 ( .A(n12206), .ZN(n12209) );
  NAND2_X1 U13840 ( .A1(n12207), .A2(n12211), .ZN(n12208) );
  NAND2_X1 U13841 ( .A1(n12209), .A2(n12208), .ZN(n15404) );
  INV_X1 U13842 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15521) );
  NAND2_X1 U13843 ( .A1(n15262), .A2(n12203), .ZN(n12213) );
  OAI21_X1 U13844 ( .B1(n12220), .B2(n12212), .A(n12211), .ZN(n15425) );
  INV_X1 U13845 ( .A(n12381), .ZN(n12216) );
  NAND2_X1 U13846 ( .A1(n12214), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12215) );
  NAND2_X1 U13847 ( .A1(n12216), .A2(n12215), .ZN(n13002) );
  INV_X1 U13848 ( .A(n13002), .ZN(n13000) );
  MUX2_X1 U13849 ( .A(n13000), .B(n14077), .S(n15383), .Z(n12390) );
  MUX2_X1 U13850 ( .A(n12390), .B(P2_EBX_REG_0__SCAN_IN), .S(n15857), .Z(
        n15582) );
  NAND2_X1 U13851 ( .A1(n15582), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14417) );
  INV_X1 U13852 ( .A(n12217), .ZN(n12223) );
  NAND3_X1 U13853 ( .A1(n15857), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n12218) );
  NAND2_X1 U13854 ( .A1(n12223), .A2(n12218), .ZN(n19025) );
  AND2_X1 U13855 ( .A1(n14417), .A2(n19025), .ZN(n17054) );
  NOR2_X1 U13856 ( .A1(n14417), .A2(n19025), .ZN(n17055) );
  NOR2_X1 U13857 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17055), .ZN(
        n12219) );
  NOR2_X1 U13858 ( .A1(n17054), .A2(n12219), .ZN(n15887) );
  INV_X1 U13859 ( .A(n12220), .ZN(n12225) );
  INV_X1 U13860 ( .A(n12221), .ZN(n12222) );
  NAND2_X1 U13861 ( .A1(n12223), .A2(n12222), .ZN(n12224) );
  NAND2_X1 U13862 ( .A1(n12225), .A2(n12224), .ZN(n12226) );
  XNOR2_X1 U13863 ( .A(n12226), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n15888) );
  NAND2_X1 U13864 ( .A1(n15887), .A2(n15888), .ZN(n12228) );
  INV_X1 U13865 ( .A(n12226), .ZN(n15413) );
  NAND2_X1 U13866 ( .A1(n15413), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12227) );
  AND2_X1 U13867 ( .A1(n12228), .A2(n12227), .ZN(n12230) );
  AND2_X1 U13868 ( .A1(n15404), .A2(n15521), .ZN(n12231) );
  AOI21_X1 U13869 ( .B1(n12230), .B2(n12070), .A(n12231), .ZN(n12229) );
  NAND2_X1 U13870 ( .A1(n15337), .A2(n12229), .ZN(n12234) );
  INV_X1 U13871 ( .A(n12230), .ZN(n15338) );
  INV_X1 U13872 ( .A(n12231), .ZN(n12232) );
  NAND3_X1 U13873 ( .A1(n15338), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n12232), .ZN(n12233) );
  NAND2_X1 U13874 ( .A1(n15505), .A2(n15506), .ZN(n12237) );
  NAND2_X1 U13875 ( .A1(n12235), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12236) );
  NAND2_X1 U13876 ( .A1(n12237), .A2(n12236), .ZN(n17337) );
  INV_X1 U13877 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12238) );
  OAI22_X1 U13878 ( .A1(n12804), .A2(n12177), .B1(n12174), .B2(n12238), .ZN(
        n12242) );
  INV_X1 U13879 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12680) );
  OAI22_X1 U13880 ( .A1(n12240), .A2(n12239), .B1(n12178), .B2(n12680), .ZN(
        n12241) );
  NOR2_X1 U13881 ( .A1(n12242), .A2(n12241), .ZN(n12247) );
  AOI22_X1 U13882 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19950), .B1(
        n19930), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12246) );
  NAND2_X1 U13883 ( .A1(n19902), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12245) );
  NAND4_X1 U13884 ( .A1(n12247), .A2(n12246), .A3(n12245), .A4(n12244), .ZN(
        n12256) );
  AOI22_X1 U13885 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20012), .B1(
        n12187), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U13886 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19993), .B1(
        n19976), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U13887 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19911), .B1(
        n12189), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12252) );
  INV_X1 U13888 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12249) );
  OAI22_X1 U13889 ( .A1(n12249), .A2(n19873), .B1(n19828), .B2(n12248), .ZN(
        n12250) );
  INV_X1 U13890 ( .A(n12250), .ZN(n12251) );
  NAND4_X1 U13891 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12255) );
  INV_X1 U13892 ( .A(n14107), .ZN(n12257) );
  NAND2_X1 U13893 ( .A1(n12257), .A2(n15109), .ZN(n12258) );
  OAI21_X1 U13894 ( .B1(n12262), .B2(n12261), .A(n12260), .ZN(n19045) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17342) );
  NAND2_X1 U13896 ( .A1(n17337), .A2(n17338), .ZN(n12265) );
  NAND2_X1 U13897 ( .A1(n12263), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12264) );
  XNOR2_X1 U13898 ( .A(n12260), .B(n12266), .ZN(n12267) );
  XNOR2_X1 U13899 ( .A(n12267), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17040) );
  INV_X1 U13900 ( .A(n12267), .ZN(n15492) );
  NAND2_X1 U13901 ( .A1(n15492), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12268) );
  INV_X1 U13902 ( .A(n12269), .ZN(n12270) );
  XNOR2_X1 U13903 ( .A(n12271), .B(n12270), .ZN(n15482) );
  NAND2_X1 U13904 ( .A1(n15482), .A2(n15859), .ZN(n12272) );
  INV_X1 U13905 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n19307) );
  NAND2_X1 U13906 ( .A1(n12272), .A2(n19307), .ZN(n17867) );
  NAND2_X1 U13907 ( .A1(n12274), .A2(n12273), .ZN(n12275) );
  NAND2_X1 U13908 ( .A1(n12284), .A2(n12275), .ZN(n15463) );
  OR2_X1 U13909 ( .A1(n15463), .A2(n12203), .ZN(n12276) );
  INV_X1 U13910 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17282) );
  NAND2_X1 U13911 ( .A1(n12276), .A2(n17282), .ZN(n17026) );
  AND2_X1 U13912 ( .A1(n12278), .A2(n12277), .ZN(n12279) );
  NOR2_X1 U13913 ( .A1(n12287), .A2(n12279), .ZN(n19078) );
  INV_X1 U13914 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17283) );
  NOR2_X1 U13915 ( .A1(n12203), .A2(n17283), .ZN(n12280) );
  NAND2_X1 U13916 ( .A1(n19078), .A2(n12280), .ZN(n17006) );
  INV_X1 U13917 ( .A(n15463), .ZN(n12281) );
  NAND3_X1 U13918 ( .A1(n12281), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n15859), .ZN(n17027) );
  INV_X1 U13919 ( .A(n12282), .ZN(n12283) );
  XNOR2_X1 U13920 ( .A(n12284), .B(n12283), .ZN(n19066) );
  NAND2_X1 U13921 ( .A1(n19066), .A2(n15859), .ZN(n12316) );
  INV_X1 U13922 ( .A(n12316), .ZN(n12285) );
  NAND2_X1 U13923 ( .A1(n12285), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17019) );
  AND2_X1 U13924 ( .A1(n17027), .A2(n17019), .ZN(n17008) );
  OR2_X1 U13925 ( .A1(n12287), .A2(n12286), .ZN(n12289) );
  AND2_X1 U13926 ( .A1(n12289), .A2(n12288), .ZN(n12307) );
  INV_X1 U13927 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17269) );
  NOR2_X1 U13928 ( .A1(n12203), .A2(n17269), .ZN(n12290) );
  NAND2_X1 U13929 ( .A1(n12307), .A2(n12290), .ZN(n16995) );
  XNOR2_X1 U13930 ( .A(n12292), .B(n11461), .ZN(n19148) );
  NAND2_X1 U13931 ( .A1(n19148), .A2(n15859), .ZN(n12293) );
  INV_X1 U13932 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17188) );
  NAND2_X1 U13933 ( .A1(n12293), .A2(n17188), .ZN(n16916) );
  INV_X1 U13934 ( .A(n12294), .ZN(n12295) );
  XNOR2_X1 U13935 ( .A(n12296), .B(n12295), .ZN(n19134) );
  NAND2_X1 U13936 ( .A1(n19134), .A2(n15859), .ZN(n12297) );
  INV_X1 U13937 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17203) );
  NAND2_X1 U13938 ( .A1(n12297), .A2(n17203), .ZN(n16928) );
  NAND2_X1 U13939 ( .A1(n16916), .A2(n16928), .ZN(n16897) );
  OR2_X1 U13940 ( .A1(n11198), .A2(n12299), .ZN(n12300) );
  NAND2_X1 U13941 ( .A1(n12298), .A2(n12300), .ZN(n15477) );
  INV_X1 U13942 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17240) );
  OAI21_X1 U13943 ( .B1(n15477), .B2(n12203), .A(n17240), .ZN(n16963) );
  INV_X1 U13944 ( .A(n12301), .ZN(n12302) );
  XNOR2_X1 U13945 ( .A(n12288), .B(n12302), .ZN(n19088) );
  NAND2_X1 U13946 ( .A1(n19088), .A2(n15859), .ZN(n12303) );
  INV_X1 U13947 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17258) );
  NAND2_X1 U13948 ( .A1(n12303), .A2(n17258), .ZN(n16958) );
  AND2_X1 U13949 ( .A1(n12305), .A2(n12304), .ZN(n12306) );
  OR2_X1 U13950 ( .A1(n12306), .A2(n11198), .ZN(n15557) );
  INV_X1 U13951 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14186) );
  OAI21_X1 U13952 ( .B1(n15557), .B2(n12203), .A(n14186), .ZN(n16961) );
  INV_X1 U13953 ( .A(n12307), .ZN(n15452) );
  OAI21_X1 U13954 ( .B1(n15452), .B2(n12203), .A(n17269), .ZN(n16996) );
  NAND4_X1 U13955 ( .A1(n16963), .A2(n16958), .A3(n16961), .A4(n16996), .ZN(
        n16894) );
  INV_X1 U13956 ( .A(n16894), .ZN(n12319) );
  INV_X1 U13957 ( .A(n12308), .ZN(n12309) );
  XNOR2_X1 U13958 ( .A(n12298), .B(n12309), .ZN(n19108) );
  NAND2_X1 U13959 ( .A1(n19108), .A2(n15859), .ZN(n12310) );
  XNOR2_X1 U13960 ( .A(n12310), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16947) );
  INV_X1 U13961 ( .A(n12311), .ZN(n12312) );
  XNOR2_X1 U13962 ( .A(n12313), .B(n12312), .ZN(n19111) );
  NAND2_X1 U13963 ( .A1(n19111), .A2(n15859), .ZN(n12314) );
  INV_X1 U13964 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17222) );
  NAND2_X1 U13965 ( .A1(n12314), .A2(n17222), .ZN(n16937) );
  NAND2_X1 U13966 ( .A1(n19078), .A2(n15859), .ZN(n12315) );
  NAND2_X1 U13967 ( .A1(n12315), .A2(n17283), .ZN(n17007) );
  INV_X1 U13968 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17294) );
  NAND2_X1 U13969 ( .A1(n12316), .A2(n17294), .ZN(n17018) );
  NAND2_X1 U13970 ( .A1(n17007), .A2(n17018), .ZN(n12317) );
  NAND2_X1 U13971 ( .A1(n16993), .A2(n12317), .ZN(n12318) );
  NAND4_X1 U13972 ( .A1(n12319), .A2(n16947), .A3(n16937), .A4(n12318), .ZN(
        n12320) );
  NOR2_X1 U13973 ( .A1(n16897), .A2(n12320), .ZN(n12322) );
  NAND2_X1 U13974 ( .A1(n16629), .A2(n15859), .ZN(n12321) );
  INV_X1 U13975 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17158) );
  NAND2_X1 U13976 ( .A1(n12321), .A2(n17158), .ZN(n16890) );
  AND2_X1 U13977 ( .A1(n12322), .A2(n16890), .ZN(n12323) );
  INV_X1 U13978 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17183) );
  NAND2_X1 U13979 ( .A1(n12326), .A2(n12325), .ZN(n12327) );
  NAND2_X1 U13980 ( .A1(n12328), .A2(n12327), .ZN(n16652) );
  NOR2_X1 U13981 ( .A1(n12203), .A2(n17158), .ZN(n12329) );
  NAND2_X1 U13982 ( .A1(n16629), .A2(n12329), .ZN(n16889) );
  NOR2_X1 U13983 ( .A1(n12203), .A2(n17222), .ZN(n12330) );
  INV_X1 U13984 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17217) );
  NOR2_X1 U13985 ( .A1(n12203), .A2(n17217), .ZN(n12331) );
  NAND2_X1 U13986 ( .A1(n19108), .A2(n12331), .ZN(n16895) );
  NOR2_X1 U13987 ( .A1(n12203), .A2(n17258), .ZN(n12332) );
  NAND2_X1 U13988 ( .A1(n19088), .A2(n12332), .ZN(n16957) );
  INV_X1 U13989 ( .A(n15477), .ZN(n12334) );
  NOR2_X1 U13990 ( .A1(n12203), .A2(n17240), .ZN(n12333) );
  NAND2_X1 U13991 ( .A1(n12334), .A2(n12333), .ZN(n16962) );
  INV_X1 U13992 ( .A(n15557), .ZN(n12336) );
  NOR2_X1 U13993 ( .A1(n12203), .A2(n14186), .ZN(n12335) );
  NAND2_X1 U13994 ( .A1(n12336), .A2(n12335), .ZN(n16960) );
  NAND4_X1 U13995 ( .A1(n16895), .A2(n16957), .A3(n16962), .A4(n16960), .ZN(
        n12337) );
  NOR2_X1 U13996 ( .A1(n16936), .A2(n12337), .ZN(n12340) );
  NOR2_X1 U13997 ( .A1(n12203), .A2(n17188), .ZN(n12338) );
  NAND2_X1 U13998 ( .A1(n19148), .A2(n12338), .ZN(n16915) );
  INV_X1 U13999 ( .A(n19134), .ZN(n12339) );
  XNOR2_X1 U14000 ( .A(n11196), .B(n11252), .ZN(n19151) );
  NAND2_X1 U14001 ( .A1(n19151), .A2(n15859), .ZN(n16877) );
  INV_X1 U14002 ( .A(n12341), .ZN(n12342) );
  XNOR2_X1 U14003 ( .A(n12343), .B(n12342), .ZN(n19164) );
  AOI21_X1 U14004 ( .B1(n19164), .B2(n15859), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16869) );
  INV_X1 U14005 ( .A(n19164), .ZN(n12344) );
  INV_X1 U14006 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14183) );
  INV_X1 U14007 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12345) );
  INV_X1 U14008 ( .A(n12346), .ZN(n12347) );
  XNOR2_X1 U14009 ( .A(n12348), .B(n12347), .ZN(n19173) );
  NAND2_X1 U14010 ( .A1(n19173), .A2(n15859), .ZN(n16858) );
  INV_X1 U14011 ( .A(n12349), .ZN(n12350) );
  XNOR2_X1 U14012 ( .A(n12351), .B(n12350), .ZN(n19197) );
  NAND2_X1 U14013 ( .A1(n19197), .A2(n15859), .ZN(n12352) );
  INV_X1 U14014 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17100) );
  NAND2_X1 U14015 ( .A1(n12352), .A2(n17100), .ZN(n12354) );
  NOR2_X1 U14016 ( .A1(n12203), .A2(n17100), .ZN(n12353) );
  NAND2_X1 U14017 ( .A1(n19197), .A2(n12353), .ZN(n12363) );
  NAND2_X1 U14018 ( .A1(n12354), .A2(n12363), .ZN(n16835) );
  INV_X1 U14019 ( .A(n12355), .ZN(n12356) );
  XNOR2_X1 U14020 ( .A(n12357), .B(n12356), .ZN(n19185) );
  NAND2_X1 U14021 ( .A1(n19185), .A2(n15859), .ZN(n12361) );
  INV_X1 U14022 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17111) );
  NAND2_X1 U14023 ( .A1(n15857), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12365) );
  INV_X1 U14024 ( .A(n12365), .ZN(n12358) );
  XNOR2_X1 U14025 ( .A(n12366), .B(n12358), .ZN(n19224) );
  OAI21_X1 U14026 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n14019), .ZN(n12360) );
  INV_X1 U14027 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14197) );
  INV_X1 U14028 ( .A(n14019), .ZN(n12359) );
  INV_X1 U14029 ( .A(n12361), .ZN(n12362) );
  NAND2_X1 U14030 ( .A1(n12362), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16847) );
  NAND2_X1 U14031 ( .A1(n12363), .A2(n16847), .ZN(n14016) );
  INV_X1 U14032 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n12367) );
  NOR2_X1 U14033 ( .A1(n14065), .A2(n12367), .ZN(n12370) );
  XNOR2_X1 U14034 ( .A(n12371), .B(n12370), .ZN(n19236) );
  NOR2_X1 U14035 ( .A1(n19236), .A2(n12203), .ZN(n12368) );
  NOR2_X1 U14036 ( .A1(n12368), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16813) );
  INV_X1 U14037 ( .A(n12368), .ZN(n12369) );
  INV_X1 U14038 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17075) );
  INV_X1 U14039 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12372) );
  NOR2_X1 U14040 ( .A1(n14065), .A2(n12372), .ZN(n12373) );
  XNOR2_X1 U14041 ( .A(n15856), .B(n12373), .ZN(n15815) );
  INV_X1 U14042 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17065) );
  OR2_X1 U14043 ( .A1(n12203), .A2(n17065), .ZN(n12374) );
  NOR2_X1 U14044 ( .A1(n15815), .A2(n12374), .ZN(n15854) );
  INV_X1 U14045 ( .A(n15854), .ZN(n12375) );
  OAI21_X1 U14046 ( .B1(n15815), .B2(n12203), .A(n17065), .ZN(n15855) );
  AND2_X1 U14047 ( .A1(n12376), .A2(n19273), .ZN(n15107) );
  NAND2_X1 U14048 ( .A1(n12150), .A2(n15107), .ZN(n12378) );
  INV_X1 U14049 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12377) );
  NAND2_X1 U14050 ( .A1(n12378), .A2(n12377), .ZN(n17880) );
  NOR2_X1 U14051 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n17418), .ZN(
        n12379) );
  NAND3_X1 U14052 ( .A1(n12995), .A2(n13011), .A3(n12998), .ZN(n12383) );
  XNOR2_X1 U14053 ( .A(n12999), .B(n12381), .ZN(n13003) );
  NOR2_X1 U14054 ( .A1(n12383), .A2(n13003), .ZN(n12382) );
  NOR2_X1 U14055 ( .A1(n12383), .A2(n13002), .ZN(n12384) );
  NOR2_X1 U14056 ( .A1(n15115), .A2(n12384), .ZN(n12385) );
  MUX2_X1 U14057 ( .A(n17880), .B(n12385), .S(n17416), .Z(n19318) );
  NOR2_X1 U14058 ( .A1(n14029), .A2(n12031), .ZN(n15097) );
  NAND2_X1 U14059 ( .A1(n19318), .A2(n15097), .ZN(n12396) );
  NAND2_X1 U14060 ( .A1(n12388), .A2(n12387), .ZN(n13016) );
  INV_X1 U14061 ( .A(n13009), .ZN(n12389) );
  AOI21_X1 U14062 ( .B1(n12390), .B2(n12999), .A(n12389), .ZN(n12391) );
  NOR2_X1 U14063 ( .A1(n13016), .A2(n12391), .ZN(n12392) );
  OR2_X1 U14064 ( .A1(n12392), .A2(n13020), .ZN(n15103) );
  INV_X1 U14065 ( .A(n15103), .ZN(n12395) );
  INV_X1 U14066 ( .A(n15390), .ZN(n12394) );
  NOR2_X1 U14067 ( .A1(n14029), .A2(n12394), .ZN(n15102) );
  NAND2_X1 U14068 ( .A1(n12395), .A2(n15102), .ZN(n14055) );
  NAND2_X1 U14069 ( .A1(n12396), .A2(n14055), .ZN(n15111) );
  NAND3_X1 U14070 ( .A1(n17416), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n19332) );
  INV_X1 U14071 ( .A(n12397), .ZN(n12398) );
  XOR2_X1 U14072 ( .A(n14089), .B(n12398), .Z(n15891) );
  XNOR2_X1 U14073 ( .A(n12400), .B(n12399), .ZN(n12401) );
  NAND2_X1 U14074 ( .A1(n14420), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14422) );
  NOR2_X1 U14075 ( .A1(n12401), .A2(n14422), .ZN(n12402) );
  INV_X1 U14076 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17052) );
  XNOR2_X1 U14077 ( .A(n12401), .B(n14422), .ZN(n17051) );
  NOR2_X1 U14078 ( .A1(n17052), .A2(n17051), .ZN(n17050) );
  NOR2_X1 U14079 ( .A1(n12402), .A2(n17050), .ZN(n12403) );
  XOR2_X1 U14080 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12403), .Z(
        n15890) );
  NOR2_X1 U14081 ( .A1(n15891), .A2(n15890), .ZN(n15889) );
  INV_X1 U14082 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17362) );
  NOR2_X1 U14083 ( .A1(n12403), .A2(n17362), .ZN(n12404) );
  OR2_X1 U14084 ( .A1(n15889), .A2(n12404), .ZN(n12405) );
  XNOR2_X1 U14085 ( .A(n12405), .B(n12070), .ZN(n15261) );
  NAND2_X1 U14086 ( .A1(n12405), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12406) );
  INV_X1 U14087 ( .A(n14066), .ZN(n12408) );
  AND2_X1 U14088 ( .A1(n12417), .A2(n12415), .ZN(n12416) );
  MUX2_X1 U14089 ( .A(n12425), .B(n15522), .S(n12413), .Z(n12418) );
  OAI21_X1 U14090 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12415), .A(
        n12418), .ZN(n12419) );
  NAND2_X1 U14091 ( .A1(n15507), .A2(n12422), .ZN(n12423) );
  NAND2_X1 U14092 ( .A1(n12423), .A2(n12415), .ZN(n12424) );
  XNOR2_X1 U14093 ( .A(n12427), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17037) );
  INV_X1 U14094 ( .A(n12427), .ZN(n12428) );
  NAND2_X1 U14095 ( .A1(n12428), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12429) );
  INV_X1 U14096 ( .A(n12430), .ZN(n12431) );
  INV_X1 U14097 ( .A(n12432), .ZN(n12433) );
  NAND2_X1 U14098 ( .A1(n12433), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12434) );
  AND2_X1 U14099 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17284) );
  NAND2_X1 U14100 ( .A1(n17284), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17247) );
  NAND2_X1 U14101 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14187) );
  NOR2_X1 U14102 ( .A1(n17247), .A2(n14187), .ZN(n12435) );
  AND3_X1 U14103 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17171) );
  NAND4_X1 U14104 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A4(n17171), .ZN(n17157) );
  INV_X1 U14105 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16881) );
  AND2_X1 U14106 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17098) );
  AND2_X1 U14107 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17077) );
  NAND2_X1 U14108 ( .A1(n17077), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17076) );
  XNOR2_X1 U14109 ( .A(n11200), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17067) );
  NOR2_X1 U14110 ( .A1(n17067), .A2(n17873), .ZN(n12544) );
  INV_X1 U14111 ( .A(n12437), .ZN(n12438) );
  AOI22_X1 U14112 ( .A1(n15865), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12443) );
  NAND2_X1 U14113 ( .A1(n12466), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12442) );
  OAI211_X1 U14114 ( .C1(n12444), .C2(n15521), .A(n12443), .B(n12442), .ZN(
        n14651) );
  NAND2_X1 U14115 ( .A1(n14652), .A2(n14651), .ZN(n14650) );
  INV_X1 U14116 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14106) );
  NAND2_X1 U14117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12447) );
  OR2_X1 U14118 ( .A1(n12527), .A2(n12445), .ZN(n12446) );
  OAI211_X1 U14119 ( .C1(n15868), .C2(n14106), .A(n12447), .B(n12446), .ZN(
        n12448) );
  AOI21_X1 U14120 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n12448), .ZN(n14656) );
  AOI22_X1 U14121 ( .A1(n15865), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12450) );
  NAND2_X1 U14122 ( .A1(n12466), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12449) );
  OAI211_X1 U14123 ( .C1(n12444), .C2(n17342), .A(n12450), .B(n12449), .ZN(
        n14680) );
  NAND2_X1 U14124 ( .A1(n14655), .A2(n14680), .ZN(n14679) );
  INV_X1 U14125 ( .A(n14679), .ZN(n14766) );
  NAND2_X1 U14126 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12456) );
  INV_X1 U14127 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n17044) );
  NAND2_X1 U14128 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12453) );
  INV_X1 U14129 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n12451) );
  OR2_X1 U14130 ( .A1(n12527), .A2(n12451), .ZN(n12452) );
  OAI211_X1 U14131 ( .C1(n15868), .C2(n17044), .A(n12453), .B(n12452), .ZN(
        n12454) );
  INV_X1 U14132 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U14133 ( .A1(n12456), .A2(n12455), .ZN(n14767) );
  NAND2_X1 U14134 ( .A1(n14766), .A2(n14767), .ZN(n14903) );
  INV_X1 U14135 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U14136 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12459) );
  INV_X1 U14137 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n12457) );
  OR2_X1 U14138 ( .A1(n12527), .A2(n12457), .ZN(n12458) );
  OAI211_X1 U14139 ( .C1(n15868), .C2(n14116), .A(n12459), .B(n12458), .ZN(
        n12460) );
  AOI21_X1 U14140 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n12460), .ZN(n14902) );
  INV_X1 U14141 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n17961) );
  NAND2_X1 U14142 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12464) );
  OR2_X1 U14143 ( .A1(n12527), .A2(n12462), .ZN(n12463) );
  OAI211_X1 U14144 ( .C1(n15868), .C2(n17961), .A(n12464), .B(n12463), .ZN(
        n12465) );
  AOI21_X1 U14145 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n12465), .ZN(n14910) );
  INV_X1 U14146 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n17962) );
  NAND2_X1 U14147 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12468) );
  AOI22_X1 U14148 ( .A1(n15865), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12467) );
  OAI211_X1 U14149 ( .C1(n15868), .C2(n17962), .A(n12468), .B(n12467), .ZN(
        n14980) );
  INV_X1 U14150 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12472) );
  NAND2_X1 U14151 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12471) );
  OR2_X1 U14152 ( .A1(n12527), .A2(n12469), .ZN(n12470) );
  OAI211_X1 U14153 ( .C1(n15868), .C2(n12472), .A(n12471), .B(n12470), .ZN(
        n12473) );
  AOI21_X1 U14154 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n12473), .ZN(n15016) );
  INV_X1 U14155 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n17963) );
  NAND2_X1 U14156 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12476) );
  INV_X1 U14157 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12474) );
  OR2_X1 U14158 ( .A1(n12527), .A2(n12474), .ZN(n12475) );
  OAI211_X1 U14159 ( .C1(n15868), .C2(n17963), .A(n12476), .B(n12475), .ZN(
        n12477) );
  AOI21_X1 U14160 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n12477), .ZN(n15020) );
  INV_X1 U14161 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19084) );
  NAND2_X1 U14162 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12480) );
  AOI22_X1 U14163 ( .A1(n15865), .A2(P2_EBX_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12479) );
  OAI211_X1 U14164 ( .C1(n15868), .C2(n19084), .A(n12480), .B(n12479), .ZN(
        n15203) );
  INV_X1 U14165 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n17964) );
  NAND2_X1 U14166 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12482) );
  AOI22_X1 U14167 ( .A1(n15865), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12481) );
  OAI211_X1 U14168 ( .C1(n15868), .C2(n17964), .A(n12482), .B(n12481), .ZN(
        n15328) );
  INV_X1 U14169 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n17965) );
  NAND2_X1 U14170 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12485) );
  INV_X1 U14171 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12483) );
  OR2_X1 U14172 ( .A1(n12527), .A2(n12483), .ZN(n12484) );
  OAI211_X1 U14173 ( .C1(n15868), .C2(n17965), .A(n12485), .B(n12484), .ZN(
        n12486) );
  AOI21_X1 U14174 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12486), .ZN(n15366) );
  INV_X1 U14175 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n17966) );
  NAND2_X1 U14176 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12489) );
  OR2_X1 U14177 ( .A1(n12527), .A2(n12487), .ZN(n12488) );
  OAI211_X1 U14178 ( .C1(n15868), .C2(n17966), .A(n12489), .B(n12488), .ZN(
        n12490) );
  AOI21_X1 U14179 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n12490), .ZN(n15540) );
  OR2_X2 U14180 ( .A1(n15539), .A2(n15540), .ZN(n15568) );
  INV_X1 U14181 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n17967) );
  NAND2_X1 U14182 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12493) );
  OR2_X1 U14183 ( .A1(n12527), .A2(n12491), .ZN(n12492) );
  OAI211_X1 U14184 ( .C1(n15868), .C2(n17967), .A(n12493), .B(n12492), .ZN(
        n12494) );
  AOI21_X1 U14185 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12494), .ZN(n15567) );
  INV_X1 U14186 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n17968) );
  NAND2_X1 U14187 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12496) );
  AOI22_X1 U14188 ( .A1(n15865), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12495) );
  OAI211_X1 U14189 ( .C1(n15868), .C2(n17968), .A(n12496), .B(n12495), .ZN(
        n15610) );
  INV_X1 U14190 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n17969) );
  NAND2_X1 U14191 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12499) );
  INV_X1 U14192 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12497) );
  OR2_X1 U14193 ( .A1(n12527), .A2(n12497), .ZN(n12498) );
  OAI211_X1 U14194 ( .C1(n15868), .C2(n17969), .A(n12499), .B(n12498), .ZN(
        n12500) );
  AOI21_X1 U14195 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n12500), .ZN(n16728) );
  INV_X1 U14196 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n17970) );
  NAND2_X1 U14197 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12502) );
  OR2_X1 U14198 ( .A1(n12527), .A2(n16646), .ZN(n12501) );
  OAI211_X1 U14199 ( .C1(n15868), .C2(n17970), .A(n12502), .B(n12501), .ZN(
        n12503) );
  AOI21_X1 U14200 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n12503), .ZN(n16641) );
  INV_X1 U14201 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n16901) );
  NAND2_X1 U14202 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12505) );
  AOI22_X1 U14203 ( .A1(n15865), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n12504) );
  OAI211_X1 U14204 ( .C1(n15868), .C2(n16901), .A(n12505), .B(n12504), .ZN(
        n16625) );
  NAND2_X1 U14205 ( .A1(n16624), .A2(n16625), .ZN(n16710) );
  INV_X1 U14206 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16882) );
  NAND2_X1 U14207 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12508) );
  INV_X1 U14208 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n12506) );
  OR2_X1 U14209 ( .A1(n12527), .A2(n12506), .ZN(n12507) );
  OAI211_X1 U14210 ( .C1(n15868), .C2(n16882), .A(n12508), .B(n12507), .ZN(
        n12509) );
  AOI21_X1 U14211 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n12509), .ZN(n16709) );
  INV_X1 U14212 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n17971) );
  NAND2_X1 U14213 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12512) );
  OR2_X1 U14214 ( .A1(n12527), .A2(n12510), .ZN(n12511) );
  OAI211_X1 U14215 ( .C1(n15868), .C2(n17971), .A(n12512), .B(n12511), .ZN(
        n12513) );
  AOI21_X1 U14216 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n12513), .ZN(n16705) );
  INV_X1 U14217 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16862) );
  NAND2_X1 U14218 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12515) );
  AOI22_X1 U14219 ( .A1(n15865), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12514) );
  OAI211_X1 U14220 ( .C1(n15868), .C2(n16862), .A(n12515), .B(n12514), .ZN(
        n16695) );
  INV_X1 U14221 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17972) );
  NAND2_X1 U14222 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12517) );
  AOI22_X1 U14223 ( .A1(n15865), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12516) );
  OAI211_X1 U14224 ( .C1(n15868), .C2(n17972), .A(n12517), .B(n12516), .ZN(
        n16688) );
  INV_X1 U14225 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17973) );
  NAND2_X1 U14226 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12520) );
  INV_X1 U14227 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n12518) );
  OR2_X1 U14228 ( .A1(n12527), .A2(n12518), .ZN(n12519) );
  OAI211_X1 U14229 ( .C1(n15868), .C2(n17973), .A(n12520), .B(n12519), .ZN(
        n12521) );
  AOI21_X1 U14230 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12521), .ZN(n16682) );
  INV_X1 U14231 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19207) );
  NAND2_X1 U14232 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12524) );
  INV_X1 U14233 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n12522) );
  OR2_X1 U14234 ( .A1(n12527), .A2(n12522), .ZN(n12523) );
  OAI211_X1 U14235 ( .C1(n15868), .C2(n19207), .A(n12524), .B(n12523), .ZN(
        n12525) );
  AOI21_X1 U14236 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12525), .ZN(n16673) );
  INV_X1 U14237 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n14159) );
  NAND2_X1 U14238 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12529) );
  INV_X1 U14239 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n12526) );
  OR2_X1 U14240 ( .A1(n12527), .A2(n12526), .ZN(n12528) );
  OAI211_X1 U14241 ( .C1(n15868), .C2(n14159), .A(n12529), .B(n12528), .ZN(
        n12530) );
  AOI21_X1 U14242 ( .B1(n15864), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12530), .ZN(n14022) );
  INV_X1 U14244 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17974) );
  NAND2_X1 U14245 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12532) );
  AOI22_X1 U14246 ( .A1(n15865), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12531) );
  OAI211_X1 U14247 ( .C1(n15868), .C2(n17974), .A(n12532), .B(n12531), .ZN(
        n16658) );
  INV_X1 U14248 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17976) );
  NAND2_X1 U14249 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12534) );
  AOI22_X1 U14250 ( .A1(n15865), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12533) );
  OAI211_X1 U14251 ( .C1(n15868), .C2(n17976), .A(n12534), .B(n12533), .ZN(
        n15863) );
  XNOR2_X1 U14252 ( .A(n16657), .B(n15863), .ZN(n17061) );
  NAND2_X1 U14253 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n15127) );
  INV_X1 U14254 ( .A(n15127), .ZN(n12535) );
  NOR2_X1 U14255 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n12535), .ZN(n17879) );
  NAND2_X1 U14256 ( .A1(n17879), .A2(n19322), .ZN(n12536) );
  AND2_X1 U14257 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17414) );
  NAND2_X1 U14258 ( .A1(n17061), .A2(n17870), .ZN(n12542) );
  INV_X1 U14259 ( .A(n15124), .ZN(n12560) );
  INV_X1 U14260 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19841) );
  NAND2_X1 U14261 ( .A1(n19841), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U14262 ( .A1(n12560), .A2(n12537), .ZN(n14425) );
  INV_X1 U14263 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17849) );
  NAND2_X1 U14264 ( .A1(n15431), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15432) );
  NAND2_X1 U14265 ( .A1(n15464), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15788) );
  INV_X1 U14266 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16902) );
  INV_X1 U14267 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16872) );
  INV_X1 U14268 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16852) );
  INV_X1 U14269 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15797) );
  INV_X1 U14270 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16818) );
  INV_X1 U14271 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n15376) );
  XNOR2_X1 U14272 ( .A(n15802), .B(n15376), .ZN(n19264) );
  NAND2_X1 U14273 ( .A1(n17416), .A2(n19975), .ZN(n19311) );
  NOR2_X1 U14274 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19311), .ZN(n17840) );
  NAND2_X2 U14275 ( .A1(n17840), .A2(n19322), .ZN(n19294) );
  NOR2_X1 U14276 ( .A1(n19294), .A2(n17976), .ZN(n17063) );
  AOI21_X1 U14277 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17063), .ZN(n12539) );
  OAI21_X1 U14278 ( .B1(n17042), .B2(n19264), .A(n12539), .ZN(n12540) );
  NAND2_X1 U14279 ( .A1(n12542), .A2(n12541), .ZN(n12543) );
  NAND2_X1 U14280 ( .A1(n12551), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12553) );
  NAND2_X1 U14281 ( .A1(n19903), .A2(n19975), .ZN(n15037) );
  AOI21_X1 U14282 ( .B1(n19898), .B2(n12553), .A(n15037), .ZN(n12547) );
  INV_X1 U14283 ( .A(n12553), .ZN(n12546) );
  NAND2_X1 U14284 ( .A1(n12546), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20008) );
  AND2_X1 U14285 ( .A1(n12547), .A2(n20008), .ZN(n19848) );
  AOI21_X1 U14286 ( .B1(n12564), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19848), .ZN(n12548) );
  AND2_X1 U14287 ( .A1(n12013), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14468) );
  INV_X1 U14288 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12755) );
  NOR2_X1 U14289 ( .A1(n12934), .A2(n12755), .ZN(n12549) );
  NAND2_X1 U14290 ( .A1(n12550), .A2(n12549), .ZN(n12573) );
  NAND2_X1 U14291 ( .A1(n12095), .A2(n15124), .ZN(n12556) );
  INV_X1 U14292 ( .A(n12551), .ZN(n19958) );
  NAND2_X1 U14293 ( .A1(n19958), .A2(n19871), .ZN(n12552) );
  NAND2_X1 U14294 ( .A1(n12553), .A2(n12552), .ZN(n19849) );
  NOR2_X1 U14295 ( .A1(n19849), .A2(n15037), .ZN(n12554) );
  AOI21_X1 U14296 ( .B1(n12564), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12554), .ZN(n12555) );
  NAND2_X1 U14297 ( .A1(n12556), .A2(n12555), .ZN(n12558) );
  INV_X1 U14298 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12739) );
  NOR2_X1 U14299 ( .A1(n12934), .A2(n12739), .ZN(n12557) );
  OR2_X1 U14300 ( .A1(n12558), .A2(n12557), .ZN(n12559) );
  NAND2_X1 U14301 ( .A1(n12558), .A2(n12557), .ZN(n12570) );
  NOR2_X1 U14302 ( .A1(n15037), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12561) );
  AOI21_X1 U14303 ( .B1(n12564), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12561), .ZN(n12562) );
  NAND2_X1 U14304 ( .A1(n12910), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12567) );
  OAI21_X1 U14305 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19958), .ZN(n19972) );
  NAND2_X1 U14306 ( .A1(n12564), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12565) );
  OAI21_X1 U14307 ( .B1(n19972), .B2(n15037), .A(n12565), .ZN(n12566) );
  INV_X1 U14308 ( .A(n14473), .ZN(n12568) );
  NAND2_X1 U14309 ( .A1(n12568), .A2(n12567), .ZN(n12569) );
  NAND2_X1 U14310 ( .A1(n14565), .A2(n14566), .ZN(n14567) );
  NAND2_X1 U14311 ( .A1(n12571), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12572) );
  AND2_X1 U14312 ( .A1(n12573), .A2(n12572), .ZN(n12574) );
  INV_X1 U14313 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12771) );
  NOR2_X1 U14314 ( .A1(n12934), .A2(n12771), .ZN(n14647) );
  INV_X1 U14315 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12575) );
  INV_X1 U14316 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12582) );
  NAND2_X1 U14317 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12579) );
  NAND2_X1 U14318 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12578) );
  NAND2_X1 U14319 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12577) );
  AOI22_X1 U14320 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12576) );
  AND4_X1 U14321 ( .A1(n12579), .A2(n12578), .A3(n12577), .A4(n12576), .ZN(
        n12581) );
  NAND2_X1 U14322 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12580) );
  OAI211_X1 U14323 ( .C1(n12582), .C2(n12150), .A(n12581), .B(n12580), .ZN(
        n12583) );
  INV_X1 U14324 ( .A(n12583), .ZN(n12592) );
  AOI22_X1 U14325 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12588) );
  NAND2_X1 U14326 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U14327 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12586) );
  NAND2_X1 U14328 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12585) );
  AND4_X1 U14329 ( .A1(n12588), .A2(n12587), .A3(n12586), .A4(n12585), .ZN(
        n12591) );
  AOI22_X1 U14330 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U14331 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U14332 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n14906) );
  NAND2_X1 U14333 ( .A1(n14907), .A2(n14906), .ZN(n14905) );
  NAND2_X1 U14334 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U14335 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12596) );
  NAND2_X1 U14336 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12595) );
  NAND2_X1 U14337 ( .A1(n12795), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12594) );
  AOI22_X1 U14338 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12593) );
  AND4_X1 U14339 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12597) );
  OAI211_X1 U14340 ( .C1(n20209), .C2(n12150), .A(n12598), .B(n12597), .ZN(
        n12599) );
  INV_X1 U14341 ( .A(n12599), .ZN(n12607) );
  AOI22_X1 U14342 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U14343 ( .A1(n12143), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12602) );
  NAND2_X1 U14344 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12601) );
  NAND2_X1 U14345 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12600) );
  AND4_X1 U14346 ( .A1(n12603), .A2(n12602), .A3(n12601), .A4(n12600), .ZN(
        n12606) );
  AOI22_X1 U14347 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12605) );
  AOI22_X1 U14348 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12604) );
  NAND4_X1 U14349 ( .A1(n12607), .A2(n12606), .A3(n12605), .A4(n12604), .ZN(
        n14984) );
  INV_X1 U14350 ( .A(n14984), .ZN(n12624) );
  INV_X1 U14351 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12608) );
  OAI22_X1 U14352 ( .A1(n12150), .A2(n15052), .B1(n12837), .B2(n12608), .ZN(
        n12614) );
  NAND2_X1 U14353 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12612) );
  NAND2_X1 U14354 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U14355 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12610) );
  AOI22_X1 U14356 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12609) );
  NAND4_X1 U14357 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        n12613) );
  NOR2_X1 U14358 ( .A1(n12614), .A2(n12613), .ZN(n12623) );
  AOI22_X1 U14359 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U14360 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U14361 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12618) );
  NAND2_X1 U14362 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U14363 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12616) );
  AND4_X1 U14364 ( .A1(n12619), .A2(n12618), .A3(n12617), .A4(n12616), .ZN(
        n12621) );
  AOI22_X1 U14365 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12620) );
  NAND4_X1 U14366 ( .A1(n12623), .A2(n12622), .A3(n12621), .A4(n12620), .ZN(
        n14117) );
  INV_X1 U14367 ( .A(n14117), .ZN(n14982) );
  INV_X1 U14368 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12625) );
  OAI22_X1 U14369 ( .A1(n12150), .A2(n12122), .B1(n12837), .B2(n12625), .ZN(
        n12631) );
  NAND2_X1 U14370 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12629) );
  NAND2_X1 U14371 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12628) );
  NAND2_X1 U14372 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12627) );
  AOI22_X1 U14373 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12626) );
  NAND4_X1 U14374 ( .A1(n12629), .A2(n12628), .A3(n12627), .A4(n12626), .ZN(
        n12630) );
  NOR2_X1 U14375 ( .A1(n12631), .A2(n12630), .ZN(n12639) );
  AOI22_X1 U14376 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U14377 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12635) );
  NAND2_X1 U14378 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12634) );
  NAND2_X1 U14379 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12633) );
  NAND2_X1 U14380 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12632) );
  AND4_X1 U14381 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12637) );
  AOI22_X1 U14382 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12636) );
  NAND4_X1 U14383 ( .A1(n12639), .A2(n12638), .A3(n12637), .A4(n12636), .ZN(
        n14123) );
  INV_X1 U14384 ( .A(n14123), .ZN(n15012) );
  NOR2_X2 U14385 ( .A1(n14905), .A2(n12640), .ZN(n15025) );
  NAND2_X1 U14386 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12647) );
  AOI22_X1 U14387 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11837), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U14388 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n12642) );
  NAND2_X1 U14389 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12839), .ZN(
        n12641) );
  NAND2_X1 U14390 ( .A1(n12642), .A2(n12641), .ZN(n12643) );
  AOI21_X1 U14391 ( .B1(n12838), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n12643), .ZN(n12645) );
  NAND2_X1 U14392 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12644) );
  AND4_X1 U14393 ( .A1(n12647), .A2(n12646), .A3(n12645), .A4(n12644), .ZN(
        n12656) );
  AOI22_X1 U14394 ( .A1(n12648), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12615), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U14395 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U14396 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12651) );
  NAND2_X1 U14397 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12650) );
  NAND2_X1 U14398 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12649) );
  AND4_X1 U14399 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        n12654) );
  AOI22_X1 U14400 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12653) );
  NAND4_X1 U14401 ( .A1(n12656), .A2(n12655), .A3(n12654), .A4(n12653), .ZN(
        n15024) );
  OAI22_X1 U14402 ( .A1(n12150), .A2(n12658), .B1(n12837), .B2(n12657), .ZN(
        n12664) );
  NAND2_X1 U14403 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12662) );
  NAND2_X1 U14404 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12661) );
  NAND2_X1 U14405 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12660) );
  AOI22_X1 U14406 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12659) );
  NAND4_X1 U14407 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n12659), .ZN(
        n12663) );
  NOR2_X1 U14408 ( .A1(n12664), .A2(n12663), .ZN(n12672) );
  AOI22_X1 U14409 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U14410 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U14411 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12667) );
  NAND2_X1 U14412 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12666) );
  NAND2_X1 U14413 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12665) );
  AND4_X1 U14414 ( .A1(n12668), .A2(n12667), .A3(n12666), .A4(n12665), .ZN(
        n12670) );
  AOI22_X1 U14415 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12669) );
  NAND4_X1 U14416 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n15201) );
  INV_X1 U14417 ( .A(n15201), .ZN(n12673) );
  NAND2_X1 U14418 ( .A1(n12846), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U14419 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U14420 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12676) );
  NAND2_X1 U14421 ( .A1(n12795), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12675) );
  AOI22_X1 U14422 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12674) );
  AND4_X1 U14423 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12678) );
  OAI211_X1 U14424 ( .C1(n12680), .C2(n12150), .A(n12679), .B(n12678), .ZN(
        n12681) );
  INV_X1 U14425 ( .A(n12681), .ZN(n12690) );
  AOI22_X1 U14426 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U14427 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12684) );
  NAND2_X1 U14428 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12683) );
  NAND2_X1 U14429 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12682) );
  AND4_X1 U14430 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12689) );
  AOI22_X1 U14431 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U14432 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12687) );
  NAND4_X1 U14433 ( .A1(n12690), .A2(n12689), .A3(n12688), .A4(n12687), .ZN(
        n15334) );
  INV_X1 U14434 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19824) );
  INV_X1 U14435 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12691) );
  OAI22_X1 U14436 ( .A1(n12150), .A2(n19824), .B1(n12837), .B2(n12691), .ZN(
        n12697) );
  NAND2_X1 U14437 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12695) );
  NAND2_X1 U14438 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12694) );
  NAND2_X1 U14439 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12693) );
  AOI22_X1 U14440 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12692) );
  NAND4_X1 U14441 ( .A1(n12695), .A2(n12694), .A3(n12693), .A4(n12692), .ZN(
        n12696) );
  NOR2_X1 U14442 ( .A1(n12697), .A2(n12696), .ZN(n12705) );
  AOI22_X1 U14443 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n12615), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12704) );
  AOI22_X1 U14444 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12701) );
  NAND2_X1 U14445 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12700) );
  NAND2_X1 U14446 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12699) );
  NAND2_X1 U14447 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12698) );
  AND4_X1 U14448 ( .A1(n12701), .A2(n12700), .A3(n12699), .A4(n12698), .ZN(
        n12703) );
  AOI22_X1 U14449 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U14450 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n15365) );
  INV_X1 U14451 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12706) );
  OAI22_X1 U14452 ( .A1(n12150), .A2(n12151), .B1(n12837), .B2(n12706), .ZN(
        n12712) );
  NAND2_X1 U14453 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12710) );
  NAND2_X1 U14454 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12709) );
  NAND2_X1 U14455 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12708) );
  AOI22_X1 U14456 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12707) );
  NAND4_X1 U14457 ( .A1(n12710), .A2(n12709), .A3(n12708), .A4(n12707), .ZN(
        n12711) );
  NOR2_X1 U14458 ( .A1(n12712), .A2(n12711), .ZN(n12720) );
  AOI22_X1 U14459 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U14460 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12716) );
  NAND2_X1 U14461 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12715) );
  NAND2_X1 U14462 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12714) );
  NAND2_X1 U14463 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12713) );
  AND4_X1 U14464 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12718) );
  AOI22_X1 U14465 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12717) );
  NAND4_X1 U14466 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        n15536) );
  INV_X1 U14467 ( .A(n15536), .ZN(n12721) );
  OR2_X2 U14468 ( .A1(n15364), .A2(n12721), .ZN(n15571) );
  INV_X1 U14469 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12723) );
  OAI22_X1 U14470 ( .A1(n12150), .A2(n12723), .B1(n12837), .B2(n12722), .ZN(
        n12729) );
  NAND2_X1 U14471 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12727) );
  NAND2_X1 U14472 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U14473 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12725) );
  AOI22_X1 U14474 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12724) );
  NAND4_X1 U14475 ( .A1(n12727), .A2(n12726), .A3(n12725), .A4(n12724), .ZN(
        n12728) );
  NOR2_X1 U14476 ( .A1(n12729), .A2(n12728), .ZN(n12737) );
  AOI22_X1 U14477 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12736) );
  AOI22_X1 U14478 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12733) );
  NAND2_X1 U14479 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12732) );
  NAND2_X1 U14480 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12731) );
  NAND2_X1 U14481 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12730) );
  AND4_X1 U14482 ( .A1(n12733), .A2(n12732), .A3(n12731), .A4(n12730), .ZN(
        n12735) );
  AOI22_X1 U14483 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12734) );
  NOR2_X4 U14484 ( .A1(n15571), .A2(n15572), .ZN(n15595) );
  INV_X1 U14485 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12738) );
  OAI22_X1 U14486 ( .A1(n12150), .A2(n12739), .B1(n12837), .B2(n12738), .ZN(
        n12745) );
  NAND2_X1 U14487 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12743) );
  NAND2_X1 U14488 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12742) );
  NAND2_X1 U14489 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12741) );
  AOI22_X1 U14490 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12740) );
  NAND4_X1 U14491 ( .A1(n12743), .A2(n12742), .A3(n12741), .A4(n12740), .ZN(
        n12744) );
  NOR2_X1 U14492 ( .A1(n12745), .A2(n12744), .ZN(n12753) );
  AOI22_X1 U14493 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12752) );
  AOI22_X1 U14494 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U14495 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12748) );
  NAND2_X1 U14496 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12747) );
  NAND2_X1 U14497 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12746) );
  AND4_X1 U14498 ( .A1(n12749), .A2(n12748), .A3(n12747), .A4(n12746), .ZN(
        n12751) );
  AOI22_X1 U14499 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12750) );
  NAND4_X1 U14500 ( .A1(n12753), .A2(n12752), .A3(n12751), .A4(n12750), .ZN(
        n15594) );
  OAI22_X1 U14501 ( .A1(n12150), .A2(n12755), .B1(n12837), .B2(n12754), .ZN(
        n12761) );
  NAND2_X1 U14502 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U14503 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12758) );
  NAND2_X1 U14504 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12757) );
  AOI22_X1 U14505 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12756) );
  NAND4_X1 U14506 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n12756), .ZN(
        n12760) );
  NOR2_X1 U14507 ( .A1(n12761), .A2(n12760), .ZN(n12769) );
  AOI22_X1 U14508 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U14509 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U14510 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12764) );
  NAND2_X1 U14511 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12763) );
  NAND2_X1 U14512 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12762) );
  AND4_X1 U14513 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12767) );
  AOI22_X1 U14514 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12766) );
  NAND4_X1 U14515 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n15636) );
  INV_X1 U14516 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12770) );
  OAI22_X1 U14517 ( .A1(n12150), .A2(n12771), .B1(n12837), .B2(n12770), .ZN(
        n12777) );
  NAND2_X1 U14518 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12775) );
  NAND2_X1 U14519 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12774) );
  NAND2_X1 U14520 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12773) );
  AOI22_X1 U14521 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12772) );
  NAND4_X1 U14522 ( .A1(n12775), .A2(n12774), .A3(n12773), .A4(n12772), .ZN(
        n12776) );
  NOR2_X1 U14523 ( .A1(n12777), .A2(n12776), .ZN(n12786) );
  AOI22_X1 U14524 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U14525 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U14526 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12780) );
  NAND2_X1 U14527 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12779) );
  NAND2_X1 U14528 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12778) );
  AND4_X1 U14529 ( .A1(n12781), .A2(n12780), .A3(n12779), .A4(n12778), .ZN(
        n12784) );
  AOI22_X1 U14530 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12783) );
  AND4_X1 U14531 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n16723) );
  INV_X1 U14532 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12788) );
  OAI22_X1 U14533 ( .A1(n12150), .A2(n12788), .B1(n12837), .B2(n12787), .ZN(
        n12794) );
  NAND2_X1 U14534 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12792) );
  NAND2_X1 U14535 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12791) );
  NAND2_X1 U14536 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12790) );
  AOI22_X1 U14537 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U14538 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12793) );
  NOR2_X1 U14539 ( .A1(n12794), .A2(n12793), .ZN(n12803) );
  AOI22_X1 U14540 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U14541 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U14542 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U14543 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12797) );
  NAND2_X1 U14544 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12796) );
  AND4_X1 U14545 ( .A1(n12799), .A2(n12798), .A3(n12797), .A4(n12796), .ZN(
        n12801) );
  AOI22_X1 U14546 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12800) );
  INV_X1 U14547 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12805) );
  OAI22_X1 U14548 ( .A1(n12150), .A2(n12805), .B1(n12837), .B2(n12804), .ZN(
        n12811) );
  NAND2_X1 U14549 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12809) );
  NAND2_X1 U14550 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12808) );
  NAND2_X1 U14551 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12807) );
  AOI22_X1 U14552 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12839), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12806) );
  NAND4_X1 U14553 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n12810) );
  NOR2_X1 U14554 ( .A1(n12811), .A2(n12810), .ZN(n12819) );
  AOI22_X1 U14555 ( .A1(n12615), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U14556 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U14557 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12814) );
  NAND2_X1 U14558 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12813) );
  NAND2_X1 U14559 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12812) );
  AND4_X1 U14560 ( .A1(n12815), .A2(n12814), .A3(n12813), .A4(n12812), .ZN(
        n12817) );
  AOI22_X1 U14561 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12816) );
  NAND4_X1 U14562 ( .A1(n12819), .A2(n12818), .A3(n12817), .A4(n12816), .ZN(
        n16712) );
  NAND2_X1 U14563 ( .A1(n16717), .A2(n16712), .ZN(n16703) );
  AOI22_X1 U14564 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12827) );
  AOI22_X1 U14565 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U14566 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12825) );
  NAND2_X1 U14567 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12823) );
  AND2_X1 U14568 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12821) );
  OR2_X1 U14569 ( .A1(n12821), .A2(n12820), .ZN(n12985) );
  NAND2_X1 U14570 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12822) );
  AND3_X1 U14571 ( .A1(n12823), .A2(n12985), .A3(n12822), .ZN(n12824) );
  NAND4_X1 U14572 ( .A1(n12827), .A2(n12826), .A3(n12825), .A4(n12824), .ZN(
        n12835) );
  AOI22_X1 U14573 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U14574 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U14575 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12831) );
  NAND2_X1 U14576 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12829) );
  INV_X1 U14577 ( .A(n12985), .ZN(n12957) );
  NAND2_X1 U14578 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12828) );
  AND3_X1 U14579 ( .A1(n12829), .A2(n12957), .A3(n12828), .ZN(n12830) );
  NAND4_X1 U14580 ( .A1(n12833), .A2(n12832), .A3(n12831), .A4(n12830), .ZN(
        n12834) );
  NAND2_X1 U14581 ( .A1(n12835), .A2(n12834), .ZN(n12855) );
  INV_X1 U14582 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12836) );
  OAI22_X1 U14583 ( .A1(n12150), .A2(n12575), .B1(n12837), .B2(n12836), .ZN(
        n12845) );
  NAND2_X1 U14584 ( .A1(n11788), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12843) );
  NAND2_X1 U14585 ( .A1(n12838), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12842) );
  NAND2_X1 U14586 ( .A1(n11837), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12841) );
  AOI22_X1 U14587 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12839), .ZN(n12840) );
  NAND4_X1 U14588 ( .A1(n12843), .A2(n12842), .A3(n12841), .A4(n12840), .ZN(
        n12844) );
  NOR2_X1 U14589 ( .A1(n12845), .A2(n12844), .ZN(n12854) );
  AOI22_X1 U14590 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12615), .B1(
        n12846), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12853) );
  AOI22_X1 U14591 ( .A1(n12159), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12795), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U14592 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12849) );
  NAND2_X1 U14593 ( .A1(n12161), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n12848) );
  NAND2_X1 U14594 ( .A1(n12162), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12847) );
  AND4_X1 U14595 ( .A1(n12850), .A2(n12849), .A3(n12848), .A4(n12847), .ZN(
        n12852) );
  AOI22_X1 U14596 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12143), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U14597 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12857) );
  XOR2_X1 U14598 ( .A(n12855), .B(n12857), .Z(n16704) );
  INV_X1 U14599 ( .A(n12855), .ZN(n12856) );
  NAND2_X1 U14600 ( .A1(n12857), .A2(n12856), .ZN(n12858) );
  INV_X1 U14601 ( .A(n12858), .ZN(n12874) );
  NAND2_X1 U14602 ( .A1(n12910), .A2(n12874), .ZN(n12876) );
  AOI22_X1 U14603 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12984), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12864) );
  NAND2_X1 U14604 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12860) );
  NAND2_X1 U14605 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12859) );
  AND3_X1 U14606 ( .A1(n12957), .A2(n12860), .A3(n12859), .ZN(n12863) );
  AOI22_X1 U14607 ( .A1(n12977), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12862) );
  AOI22_X1 U14608 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12861) );
  NAND4_X1 U14609 ( .A1(n12864), .A2(n12863), .A3(n12862), .A4(n12861), .ZN(
        n12872) );
  AOI22_X1 U14610 ( .A1(n12977), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12976), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12870) );
  NAND2_X1 U14611 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12866) );
  NAND2_X1 U14612 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12865) );
  AND3_X1 U14613 ( .A1(n12866), .A2(n12985), .A3(n12865), .ZN(n12869) );
  AOI22_X1 U14614 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U14615 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12867) );
  NAND4_X1 U14616 ( .A1(n12870), .A2(n12869), .A3(n12868), .A4(n12867), .ZN(
        n12871) );
  AND2_X1 U14617 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  INV_X1 U14618 ( .A(n12873), .ZN(n12875) );
  AND2_X1 U14619 ( .A1(n12874), .A2(n12873), .ZN(n12891) );
  AOI22_X1 U14620 ( .A1(n12876), .A2(n12875), .B1(n12891), .B2(n19017), .ZN(
        n16693) );
  NAND2_X1 U14621 ( .A1(n16694), .A2(n16693), .ZN(n16692) );
  AOI22_X1 U14622 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12882) );
  AOI22_X1 U14623 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U14624 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12880) );
  NAND2_X1 U14625 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n12878) );
  NAND2_X1 U14626 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12877) );
  AND3_X1 U14627 ( .A1(n12878), .A2(n12985), .A3(n12877), .ZN(n12879) );
  NAND4_X1 U14628 ( .A1(n12882), .A2(n12881), .A3(n12880), .A4(n12879), .ZN(
        n12890) );
  AOI22_X1 U14629 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U14630 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U14631 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12886) );
  NAND2_X1 U14632 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12884) );
  NAND2_X1 U14633 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12883) );
  AND3_X1 U14634 ( .A1(n12884), .A2(n12957), .A3(n12883), .ZN(n12885) );
  NAND4_X1 U14635 ( .A1(n12888), .A2(n12887), .A3(n12886), .A4(n12885), .ZN(
        n12889) );
  AND2_X1 U14636 ( .A1(n12890), .A2(n12889), .ZN(n12893) );
  NAND2_X1 U14637 ( .A1(n12891), .A2(n12893), .ZN(n12931) );
  OAI211_X1 U14638 ( .C1(n12891), .C2(n12893), .A(n12910), .B(n12931), .ZN(
        n12895) );
  INV_X1 U14639 ( .A(n12895), .ZN(n12892) );
  INV_X1 U14640 ( .A(n12893), .ZN(n12894) );
  NOR2_X1 U14641 ( .A1(n14064), .A2(n12894), .ZN(n16686) );
  NAND2_X1 U14642 ( .A1(n16687), .A2(n16686), .ZN(n16685) );
  AOI22_X1 U14643 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U14644 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U14645 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12899) );
  NAND2_X1 U14646 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12897) );
  NAND2_X1 U14647 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12896) );
  AND3_X1 U14648 ( .A1(n12897), .A2(n12985), .A3(n12896), .ZN(n12898) );
  NAND4_X1 U14649 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        n12909) );
  AOI22_X1 U14650 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U14651 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U14652 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12905) );
  NAND2_X1 U14653 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12903) );
  NAND2_X1 U14654 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12902) );
  AND3_X1 U14655 ( .A1(n12903), .A2(n12957), .A3(n12902), .ZN(n12904) );
  NAND4_X1 U14656 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12908) );
  AND2_X1 U14657 ( .A1(n12909), .A2(n12908), .ZN(n12932) );
  XNOR2_X1 U14658 ( .A(n12931), .B(n12932), .ZN(n12911) );
  NAND2_X1 U14659 ( .A1(n12911), .A2(n12910), .ZN(n12914) );
  INV_X1 U14660 ( .A(n12932), .ZN(n12912) );
  NOR2_X1 U14661 ( .A1(n19017), .A2(n12912), .ZN(n16677) );
  INV_X1 U14662 ( .A(n12914), .ZN(n12915) );
  NAND2_X1 U14663 ( .A1(n12913), .A2(n12915), .ZN(n12916) );
  AOI22_X1 U14664 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U14665 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U14666 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12920) );
  NAND2_X1 U14667 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n12918) );
  NAND2_X1 U14668 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12917) );
  AND3_X1 U14669 ( .A1(n12918), .A2(n12985), .A3(n12917), .ZN(n12919) );
  NAND4_X1 U14670 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12930) );
  AOI22_X1 U14671 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U14672 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U14673 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12926) );
  NAND2_X1 U14674 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12924) );
  NAND2_X1 U14675 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12923) );
  AND3_X1 U14676 ( .A1(n12924), .A2(n12957), .A3(n12923), .ZN(n12925) );
  NAND4_X1 U14677 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n12929) );
  NAND2_X1 U14678 ( .A1(n12930), .A2(n12929), .ZN(n12951) );
  INV_X1 U14679 ( .A(n12931), .ZN(n12933) );
  NAND2_X1 U14680 ( .A1(n12933), .A2(n12932), .ZN(n12935) );
  NOR2_X1 U14681 ( .A1(n12935), .A2(n12951), .ZN(n16662) );
  AOI211_X1 U14682 ( .C1(n12951), .C2(n12935), .A(n12934), .B(n16662), .ZN(
        n12950) );
  AOI22_X1 U14683 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U14684 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12936) );
  NAND2_X1 U14685 ( .A1(n12937), .A2(n12936), .ZN(n12949) );
  AOI22_X1 U14686 ( .A1(n15085), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12976), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12939) );
  AOI21_X1 U14687 ( .B1(n12983), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n12985), .ZN(n12938) );
  OAI211_X1 U14688 ( .C1(n11746), .C2(n12940), .A(n12939), .B(n12938), .ZN(
        n12948) );
  AOI22_X1 U14689 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12977), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14690 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12941) );
  NAND2_X1 U14691 ( .A1(n12942), .A2(n12941), .ZN(n12947) );
  AOI22_X1 U14692 ( .A1(n15085), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12976), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12945) );
  NAND2_X1 U14693 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12944) );
  NAND2_X1 U14694 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12943) );
  NAND4_X1 U14695 ( .A1(n12945), .A2(n12985), .A3(n12944), .A4(n12943), .ZN(
        n12946) );
  OAI22_X1 U14696 ( .A1(n12949), .A2(n12948), .B1(n12947), .B2(n12946), .ZN(
        n16663) );
  INV_X1 U14697 ( .A(n12951), .ZN(n12952) );
  NAND2_X1 U14698 ( .A1(n15109), .A2(n12952), .ZN(n16670) );
  INV_X1 U14699 ( .A(n16662), .ZN(n12954) );
  NOR3_X1 U14700 ( .A1(n12954), .A2(n12393), .A3(n16663), .ZN(n16653) );
  AOI22_X1 U14701 ( .A1(n12976), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12984), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12961) );
  NAND2_X1 U14702 ( .A1(n15085), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n12956) );
  NAND2_X1 U14703 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12955) );
  AND3_X1 U14704 ( .A1(n12957), .A2(n12956), .A3(n12955), .ZN(n12960) );
  AOI22_X1 U14705 ( .A1(n12973), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U14706 ( .A1(n12977), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12958) );
  NAND4_X1 U14707 ( .A1(n12961), .A2(n12960), .A3(n12959), .A4(n12958), .ZN(
        n12969) );
  AOI22_X1 U14708 ( .A1(n12977), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12984), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U14709 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U14710 ( .A1(n11957), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12982), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12965) );
  NAND2_X1 U14711 ( .A1(n15085), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12963) );
  NAND2_X1 U14712 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12962) );
  AND3_X1 U14713 ( .A1(n12963), .A2(n12962), .A3(n12985), .ZN(n12964) );
  NAND4_X1 U14714 ( .A1(n12967), .A2(n12966), .A3(n12965), .A4(n12964), .ZN(
        n12968) );
  AND2_X1 U14715 ( .A1(n12969), .A2(n12968), .ZN(n16654) );
  OAI21_X1 U14716 ( .B1(n16656), .B2(n16653), .A(n16654), .ZN(n12994) );
  AOI22_X1 U14717 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n12984), .B1(
        n12976), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12971) );
  AOI21_X1 U14718 ( .B1(n12983), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A(
        n12985), .ZN(n12970) );
  OAI211_X1 U14719 ( .C1(n12972), .C2(n19824), .A(n12971), .B(n12970), .ZN(
        n12992) );
  AOI22_X1 U14720 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n12977), .B1(
        n12973), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U14721 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n15085), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12974) );
  NAND2_X1 U14722 ( .A1(n12975), .A2(n12974), .ZN(n12991) );
  AOI22_X1 U14723 ( .A1(n12977), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12976), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12981) );
  AOI22_X1 U14724 ( .A1(n12979), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12978), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U14725 ( .A1(n12981), .A2(n12980), .ZN(n12990) );
  AOI22_X1 U14726 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15085), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12988) );
  NAND2_X1 U14727 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12987) );
  NAND2_X1 U14728 ( .A1(n12984), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12986) );
  NAND4_X1 U14729 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12989) );
  OAI22_X1 U14730 ( .A1(n12992), .A2(n12991), .B1(n12990), .B2(n12989), .ZN(
        n12993) );
  XNOR2_X1 U14731 ( .A(n12994), .B(n12993), .ZN(n15853) );
  NOR2_X1 U14732 ( .A1(n12995), .A2(n12031), .ZN(n12996) );
  OR2_X1 U14733 ( .A1(n13020), .A2(n12996), .ZN(n13018) );
  INV_X1 U14734 ( .A(n12998), .ZN(n13008) );
  NAND2_X1 U14735 ( .A1(n13000), .A2(n12999), .ZN(n13001) );
  NAND2_X1 U14736 ( .A1(n15383), .A2(n13001), .ZN(n13007) );
  NAND2_X1 U14737 ( .A1(n15109), .A2(n13002), .ZN(n13005) );
  INV_X1 U14738 ( .A(n13003), .ZN(n13004) );
  NAND3_X1 U14739 ( .A1(n13005), .A2(n20294), .A3(n13004), .ZN(n13006) );
  OAI211_X1 U14740 ( .C1(n12997), .C2(n13008), .A(n13007), .B(n13006), .ZN(
        n13014) );
  OAI21_X1 U14741 ( .B1(n14479), .B2(n15109), .A(n13008), .ZN(n13010) );
  NAND2_X1 U14742 ( .A1(n13010), .A2(n13009), .ZN(n13013) );
  INV_X1 U14743 ( .A(n13011), .ZN(n13012) );
  AOI21_X1 U14744 ( .B1(n13014), .B2(n13013), .A(n13012), .ZN(n13015) );
  AOI21_X1 U14745 ( .B1(n13016), .B2(n12031), .A(n13015), .ZN(n13017) );
  NOR2_X1 U14746 ( .A1(n13018), .A2(n13017), .ZN(n13019) );
  MUX2_X1 U14747 ( .A(n19273), .B(n13019), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n14039) );
  INV_X1 U14748 ( .A(n15038), .ZN(n15100) );
  INV_X1 U14749 ( .A(n13022), .ZN(n13024) );
  AND2_X1 U14750 ( .A1(n13024), .A2(n13023), .ZN(n15059) );
  NAND2_X1 U14751 ( .A1(n15100), .A2(n15059), .ZN(n15055) );
  NAND2_X1 U14752 ( .A1(n15055), .A2(n15061), .ZN(n13025) );
  NAND2_X1 U14753 ( .A1(n17061), .A2(n16700), .ZN(n13027) );
  NAND2_X1 U14754 ( .A1(n15538), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13026) );
  OAI21_X1 U14755 ( .B1(n15853), .B2(n16732), .A(n11725), .ZN(P2_U2857) );
  AND2_X2 U14756 ( .A1(n13045), .A2(n13046), .ZN(n13102) );
  NAND2_X1 U14757 ( .A1(n11135), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13031) );
  AND2_X2 U14758 ( .A1(n13045), .A2(n13037), .ZN(n13437) );
  NAND2_X1 U14759 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n13030) );
  AND2_X2 U14760 ( .A1(n13046), .A2(n13032), .ZN(n13203) );
  NAND2_X1 U14761 ( .A1(n13203), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n13029) );
  NAND2_X1 U14762 ( .A1(n13093), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13028) );
  NAND2_X1 U14763 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n13036) );
  NAND2_X1 U14764 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n13035) );
  NAND2_X1 U14765 ( .A1(n13143), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n13034) );
  AND2_X2 U14766 ( .A1(n13037), .A2(n13032), .ZN(n13208) );
  NAND2_X1 U14767 ( .A1(n13208), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13033) );
  AND2_X2 U14768 ( .A1(n13047), .A2(n13037), .ZN(n13107) );
  NAND2_X1 U14769 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n13040) );
  NAND2_X1 U14770 ( .A1(n13253), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13039) );
  NAND2_X1 U14771 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13038) );
  NAND3_X1 U14772 ( .A1(n13040), .A2(n13039), .A3(n13038), .ZN(n13041) );
  NOR2_X1 U14773 ( .A1(n11714), .A2(n13041), .ZN(n13042) );
  NAND2_X1 U14774 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13051) );
  AND2_X2 U14775 ( .A1(n13047), .A2(n14641), .ZN(n13593) );
  NAND2_X1 U14776 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13050) );
  NAND2_X1 U14777 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13049) );
  NAND2_X1 U14778 ( .A1(n13144), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13048) );
  AOI22_X1 U14779 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13208), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U14780 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13056) );
  AOI22_X1 U14781 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13143), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13055) );
  AOI22_X1 U14782 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13144), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13054) );
  AOI22_X1 U14783 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13061) );
  AOI22_X1 U14784 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13253), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U14785 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13203), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U14786 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13093), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13058) );
  NAND2_X1 U14787 ( .A1(n13157), .A2(n13275), .ZN(n13092) );
  NAND2_X1 U14788 ( .A1(n11135), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13065) );
  NAND2_X1 U14789 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n13064) );
  NAND2_X1 U14790 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13063) );
  NAND2_X1 U14791 ( .A1(n13093), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13062) );
  NAND2_X1 U14792 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13069) );
  NAND2_X1 U14793 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n13068) );
  NAND2_X1 U14794 ( .A1(n13253), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13067) );
  NAND2_X1 U14795 ( .A1(n13203), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13066) );
  NAND2_X1 U14796 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13073) );
  NAND2_X1 U14797 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n13072) );
  NAND2_X1 U14798 ( .A1(n13208), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13071) );
  NAND2_X1 U14799 ( .A1(n13143), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n13070) );
  NAND2_X1 U14800 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13077) );
  NAND2_X1 U14801 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13076) );
  NAND2_X1 U14802 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n13075) );
  NAND2_X1 U14803 ( .A1(n13144), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13074) );
  NAND2_X2 U14804 ( .A1(n13157), .A2(n14817), .ZN(n13115) );
  AOI22_X1 U14805 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13253), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14806 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13231), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14807 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13203), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13083) );
  AOI22_X1 U14808 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13208), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13082) );
  NAND4_X1 U14809 ( .A1(n13085), .A2(n13084), .A3(n13083), .A4(n13082), .ZN(
        n13091) );
  AOI22_X1 U14810 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13089) );
  AOI22_X1 U14811 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13088) );
  AOI22_X1 U14812 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13093), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13087) );
  AOI22_X1 U14813 ( .A1(n13143), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13144), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13086) );
  NAND4_X1 U14814 ( .A1(n13089), .A2(n13088), .A3(n13087), .A4(n13086), .ZN(
        n13090) );
  AOI22_X1 U14815 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U14816 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13253), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13096) );
  AOI22_X1 U14817 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13203), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U14818 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13093), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U14819 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U14820 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13208), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U14821 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13143), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U14822 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13144), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U14823 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13106) );
  AOI22_X1 U14824 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13253), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U14825 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13203), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U14826 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13093), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U14827 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13238), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13112) );
  AOI22_X1 U14828 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13208), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U14829 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13143), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13110) );
  AOI22_X1 U14830 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13144), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13109) );
  NAND2_X1 U14831 ( .A1(n13114), .A2(n13113), .ZN(n13170) );
  NAND2_X1 U14832 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13119) );
  NAND2_X1 U14833 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13118) );
  NAND2_X1 U14834 ( .A1(n13253), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13117) );
  NAND2_X1 U14835 ( .A1(n13203), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13116) );
  NAND2_X1 U14836 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13121) );
  NAND2_X1 U14837 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13126) );
  NAND2_X1 U14838 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13125) );
  NAND2_X1 U14839 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13124) );
  NAND2_X1 U14840 ( .A1(n13093), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13123) );
  NAND2_X1 U14841 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13130) );
  NAND2_X1 U14842 ( .A1(n11140), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13129) );
  NAND2_X1 U14843 ( .A1(n13208), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13128) );
  NAND2_X1 U14844 ( .A1(n13143), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13127) );
  NOR2_X2 U14845 ( .A1(n13170), .A2(n11719), .ZN(n14409) );
  NAND2_X1 U14846 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13137) );
  NAND2_X1 U14847 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13136) );
  NAND2_X1 U14848 ( .A1(n13254), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13135) );
  NAND2_X1 U14849 ( .A1(n13108), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n13134) );
  NAND2_X1 U14850 ( .A1(n13203), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13142) );
  NAND2_X1 U14851 ( .A1(n11137), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13139) );
  NAND2_X1 U14852 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13138) );
  NAND2_X1 U14853 ( .A1(n13139), .A2(n13138), .ZN(n13140) );
  NAND2_X1 U14854 ( .A1(n13238), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13148) );
  NAND2_X1 U14855 ( .A1(n13231), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13147) );
  NAND2_X1 U14856 ( .A1(n13143), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13146) );
  NAND2_X1 U14857 ( .A1(n13144), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U14858 ( .A1(n13237), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13152) );
  NAND2_X1 U14859 ( .A1(n13122), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13151) );
  NAND2_X1 U14860 ( .A1(n13208), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13150) );
  NAND2_X1 U14861 ( .A1(n13093), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13149) );
  NAND2_X1 U14862 ( .A1(n14409), .A2(n14797), .ZN(n14619) );
  INV_X1 U14863 ( .A(n14686), .ZN(n13158) );
  NAND2_X1 U14864 ( .A1(n13158), .A2(n14222), .ZN(n13159) );
  NAND2_X1 U14865 ( .A1(n14619), .A2(n13159), .ZN(n14532) );
  XNOR2_X1 U14866 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n14522) );
  AND2_X1 U14867 ( .A1(n15911), .A2(n14825), .ZN(n14683) );
  NAND2_X1 U14868 ( .A1(n13275), .A2(n14628), .ZN(n14629) );
  NOR2_X1 U14869 ( .A1(n14725), .A2(n14629), .ZN(n13162) );
  NAND2_X1 U14870 ( .A1(n14683), .A2(n13162), .ZN(n14547) );
  NOR2_X1 U14871 ( .A1(n14532), .A2(n13163), .ZN(n13176) );
  INV_X1 U14872 ( .A(n13183), .ZN(n13164) );
  INV_X1 U14873 ( .A(n13184), .ZN(n13165) );
  NAND2_X1 U14874 ( .A1(n13164), .A2(n13184), .ZN(n13169) );
  NAND2_X1 U14875 ( .A1(n13165), .A2(n21947), .ZN(n13166) );
  NAND2_X1 U14876 ( .A1(n13169), .A2(n13166), .ZN(n14519) );
  NAND2_X1 U14877 ( .A1(n14519), .A2(n11614), .ZN(n13167) );
  NAND2_X1 U14878 ( .A1(n13167), .A2(n14886), .ZN(n14542) );
  NAND2_X1 U14879 ( .A1(n13169), .A2(n16573), .ZN(n13192) );
  NAND2_X1 U14880 ( .A1(n15177), .A2(n15178), .ZN(n15195) );
  AND4_X2 U14881 ( .A1(n14542), .A2(n13192), .A3(n15195), .A4(n14684), .ZN(
        n13172) );
  OAI21_X1 U14882 ( .B1(n13170), .B2(n14216), .A(n15177), .ZN(n13171) );
  INV_X1 U14883 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U14884 ( .A1(n13173), .A2(n15308), .ZN(n22289) );
  NAND2_X1 U14885 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13198) );
  OAI21_X1 U14886 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n13198), .ZN(n22542) );
  INV_X1 U14887 ( .A(n13910), .ZN(n13180) );
  NAND2_X1 U14888 ( .A1(n13180), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13193) );
  OAI21_X1 U14889 ( .B1(n13914), .B2(n22542), .A(n13193), .ZN(n13174) );
  INV_X1 U14890 ( .A(n13174), .ZN(n13175) );
  INV_X1 U14891 ( .A(n13176), .ZN(n13177) );
  MUX2_X1 U14892 ( .A(n13180), .B(n13310), .S(n22571), .Z(n13181) );
  INV_X1 U14893 ( .A(n13181), .ZN(n13182) );
  NAND2_X1 U14894 ( .A1(n13183), .A2(n17464), .ZN(n13190) );
  INV_X1 U14895 ( .A(n15911), .ZN(n15175) );
  AND2_X1 U14896 ( .A1(n15175), .A2(n14226), .ZN(n15899) );
  NAND2_X1 U14897 ( .A1(n13184), .A2(n13922), .ZN(n13187) );
  OR2_X1 U14898 ( .A1(n22289), .A2(n17473), .ZN(n20637) );
  AOI21_X1 U14899 ( .B1(n13156), .B2(n14886), .A(n20637), .ZN(n13185) );
  NAND2_X1 U14900 ( .A1(n15195), .A2(n13185), .ZN(n13186) );
  AOI21_X1 U14901 ( .B1(n15899), .B2(n13187), .A(n13186), .ZN(n13189) );
  NAND2_X1 U14902 ( .A1(n14216), .A2(n14804), .ZN(n13188) );
  NAND2_X1 U14903 ( .A1(n13170), .A2(n15911), .ZN(n14541) );
  NAND2_X1 U14904 ( .A1(n13252), .A2(n13250), .ZN(n13218) );
  INV_X1 U14905 ( .A(n13193), .ZN(n13195) );
  OAI21_X1 U14906 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n13195), .A(
        n13194), .ZN(n13196) );
  INV_X1 U14907 ( .A(n13198), .ZN(n13197) );
  NAND2_X1 U14908 ( .A1(n13197), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13307) );
  NAND2_X1 U14909 ( .A1(n13198), .A2(n22585), .ZN(n13199) );
  NAND2_X1 U14910 ( .A1(n13310), .A2(n15135), .ZN(n13200) );
  AOI22_X1 U14911 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U14912 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U14913 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U14914 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13204) );
  NAND4_X1 U14915 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        n13214) );
  AOI22_X1 U14916 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13212) );
  AOI22_X1 U14917 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U14918 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U14919 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13209) );
  NAND4_X1 U14920 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13213) );
  OAI22_X2 U14921 ( .A1(n14672), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13937), 
        .B2(n13314), .ZN(n13217) );
  INV_X1 U14922 ( .A(n13313), .ZN(n13245) );
  AOI22_X1 U14923 ( .A1(n13899), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13245), .B2(n13215), .ZN(n13216) );
  XNOR2_X2 U14924 ( .A(n13217), .B(n13216), .ZN(n13303) );
  NAND2_X1 U14925 ( .A1(n14919), .A2(n13218), .ZN(n15210) );
  INV_X1 U14926 ( .A(n13314), .ZN(n13272) );
  AOI22_X1 U14927 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13122), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U14928 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U14929 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U14930 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13220) );
  NAND4_X1 U14931 ( .A1(n13223), .A2(n13222), .A3(n13221), .A4(n13220), .ZN(
        n13229) );
  AOI22_X1 U14932 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U14933 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13143), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13226) );
  AOI22_X1 U14934 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13144), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U14935 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13224) );
  NAND4_X1 U14936 ( .A1(n13227), .A2(n13226), .A3(n13225), .A4(n13224), .ZN(
        n13228) );
  NAND2_X1 U14937 ( .A1(n13272), .A2(n13926), .ZN(n13230) );
  AOI22_X1 U14938 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U14939 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U14940 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13122), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U14941 ( .A1(n11142), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13233) );
  NAND4_X1 U14942 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13244) );
  AOI22_X1 U14943 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U14944 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13241) );
  AOI22_X1 U14945 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13240) );
  AOI22_X1 U14946 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13239) );
  NAND4_X1 U14947 ( .A1(n13242), .A2(n13241), .A3(n13240), .A4(n13239), .ZN(
        n13243) );
  NAND2_X1 U14948 ( .A1(n13899), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13247) );
  NAND2_X1 U14949 ( .A1(n13245), .A2(n13926), .ZN(n13246) );
  OAI211_X1 U14950 ( .C1(n13314), .C2(n13988), .A(n13247), .B(n13246), .ZN(
        n13248) );
  NAND2_X1 U14951 ( .A1(n13925), .A2(n13248), .ZN(n13249) );
  INV_X1 U14952 ( .A(n13250), .ZN(n13251) );
  INV_X1 U14953 ( .A(n13988), .ZN(n13265) );
  AOI22_X1 U14954 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U14955 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13232), .B1(
        n11139), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U14956 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13122), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13256) );
  AOI22_X1 U14957 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13255) );
  NAND4_X1 U14958 ( .A1(n13258), .A2(n13257), .A3(n13256), .A4(n13255), .ZN(
        n13264) );
  AOI22_X1 U14959 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n13763), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U14960 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U14961 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13260) );
  AOI22_X1 U14962 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13259) );
  NAND4_X1 U14963 ( .A1(n13262), .A2(n13261), .A3(n13260), .A4(n13259), .ZN(
        n13263) );
  XNOR2_X1 U14964 ( .A(n13265), .B(n13927), .ZN(n13266) );
  NAND2_X1 U14965 ( .A1(n13266), .A2(n13272), .ZN(n13267) );
  INV_X1 U14966 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13271) );
  AOI21_X1 U14967 ( .B1(n14817), .B2(n13988), .A(n17473), .ZN(n13270) );
  NAND2_X1 U14968 ( .A1(n15177), .A2(n13927), .ZN(n13269) );
  NAND2_X1 U14969 ( .A1(n13290), .A2(n13289), .ZN(n13273) );
  NAND2_X1 U14970 ( .A1(n13272), .A2(n13988), .ZN(n13985) );
  OAI21_X2 U14971 ( .B1(n13282), .B2(n13283), .A(n13274), .ZN(n13302) );
  XNOR2_X1 U14972 ( .A(n13303), .B(n13302), .ZN(n13935) );
  INV_X2 U14973 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n22605) );
  NAND2_X1 U14974 ( .A1(n13935), .A2(n13537), .ZN(n13280) );
  INV_X1 U14975 ( .A(n14629), .ZN(n14635) );
  NAND2_X1 U14976 ( .A1(n14635), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13351) );
  INV_X2 U14977 ( .A(n13847), .ZN(n15167) );
  XNOR2_X1 U14978 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n22113) );
  AOI21_X1 U14979 ( .B1(n15167), .B2(n22113), .A(n15818), .ZN(n13277) );
  NAND2_X1 U14980 ( .A1(n13293), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n13276) );
  OAI211_X1 U14981 ( .C1(n13351), .C2(n14697), .A(n13277), .B(n13276), .ZN(
        n13278) );
  INV_X1 U14982 ( .A(n13278), .ZN(n13279) );
  NAND2_X1 U14983 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  NAND2_X1 U14984 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13301) );
  NAND2_X1 U14985 ( .A1(n13281), .A2(n13301), .ZN(n14660) );
  NAND2_X1 U14986 ( .A1(n14637), .A2(n13537), .ZN(n13288) );
  AOI22_X1 U14987 ( .A1(n13293), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n22605), .ZN(n13286) );
  INV_X1 U14988 ( .A(n13351), .ZN(n13284) );
  NAND2_X1 U14989 ( .A1(n13284), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13285) );
  AND2_X1 U14990 ( .A1(n13286), .A2(n13285), .ZN(n13287) );
  NAND2_X1 U14991 ( .A1(n13288), .A2(n13287), .ZN(n14572) );
  NAND2_X1 U14992 ( .A1(n11155), .A2(n14804), .ZN(n13291) );
  NAND2_X1 U14993 ( .A1(n13291), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14574) );
  NAND2_X1 U14994 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13295) );
  NAND2_X1 U14995 ( .A1(n13293), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n13294) );
  OAI211_X1 U14996 ( .C1(n13351), .C2(n13179), .A(n13295), .B(n13294), .ZN(
        n13296) );
  AOI21_X1 U14997 ( .B1(n17438), .B2(n13537), .A(n13296), .ZN(n13297) );
  OR2_X1 U14998 ( .A1(n14574), .A2(n13297), .ZN(n14575) );
  INV_X1 U14999 ( .A(n13297), .ZN(n14576) );
  OR2_X1 U15000 ( .A1(n14576), .A2(n13847), .ZN(n13298) );
  NAND2_X1 U15001 ( .A1(n14575), .A2(n13298), .ZN(n14571) );
  NAND2_X1 U15002 ( .A1(n14572), .A2(n14571), .ZN(n14661) );
  NAND2_X1 U15003 ( .A1(n13300), .A2(n13299), .ZN(n14663) );
  INV_X1 U15004 ( .A(n13302), .ZN(n13304) );
  INV_X1 U15005 ( .A(n13307), .ZN(n14918) );
  NAND2_X1 U15006 ( .A1(n14918), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n22602) );
  NAND2_X1 U15007 ( .A1(n13307), .A2(n22586), .ZN(n13308) );
  NOR2_X1 U15008 ( .A1(n13910), .A2(n22586), .ZN(n13309) );
  AOI21_X1 U15009 ( .B1(n16585), .B2(n13310), .A(n13309), .ZN(n13311) );
  XNOR2_X2 U15010 ( .A(n17398), .B(n14849), .ZN(n16564) );
  AOI22_X1 U15011 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13318) );
  AOI22_X1 U15012 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13317) );
  AOI22_X1 U15013 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U15014 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13315) );
  NAND4_X1 U15015 ( .A1(n13318), .A2(n13317), .A3(n13316), .A4(n13315), .ZN(
        n13324) );
  AOI22_X1 U15016 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13322) );
  AOI22_X1 U15017 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U15018 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13320) );
  AOI22_X1 U15019 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13319) );
  NAND4_X1 U15020 ( .A1(n13322), .A2(n13321), .A3(n13320), .A4(n13319), .ZN(
        n13323) );
  AOI22_X1 U15021 ( .A1(n13893), .A2(n13949), .B1(n13899), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13325) );
  INV_X1 U15022 ( .A(n13327), .ZN(n13326) );
  INV_X1 U15023 ( .A(n13353), .ZN(n13355) );
  INV_X1 U15024 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13328) );
  NAND2_X1 U15025 ( .A1(n13328), .A2(n13327), .ZN(n13329) );
  NAND2_X1 U15026 ( .A1(n13355), .A2(n13329), .ZN(n15186) );
  AOI22_X1 U15027 ( .A1(n15186), .A2(n15167), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13331) );
  NAND2_X1 U15028 ( .A1(n13849), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n13330) );
  OAI211_X1 U15029 ( .C1(n13351), .C2(n13305), .A(n13331), .B(n13330), .ZN(
        n13332) );
  INV_X1 U15030 ( .A(n13332), .ZN(n13333) );
  NAND2_X1 U15031 ( .A1(n13334), .A2(n13333), .ZN(n14737) );
  NAND2_X1 U15032 ( .A1(n14738), .A2(n14737), .ZN(n14736) );
  AOI22_X1 U15033 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13339) );
  AOI22_X1 U15034 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13338) );
  AOI22_X1 U15035 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13337) );
  AOI22_X1 U15036 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13336) );
  NAND4_X1 U15037 ( .A1(n13339), .A2(n13338), .A3(n13337), .A4(n13336), .ZN(
        n13345) );
  AOI22_X1 U15038 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13343) );
  AOI22_X1 U15039 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13342) );
  AOI22_X1 U15040 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13341) );
  AOI22_X1 U15041 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13340) );
  NAND4_X1 U15042 ( .A1(n13343), .A2(n13342), .A3(n13341), .A4(n13340), .ZN(
        n13344) );
  NAND2_X1 U15043 ( .A1(n13893), .A2(n13957), .ZN(n13347) );
  NAND2_X1 U15044 ( .A1(n13899), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13346) );
  NAND2_X1 U15045 ( .A1(n13347), .A2(n13346), .ZN(n13364) );
  XNOR2_X1 U15046 ( .A(n13363), .B(n13364), .ZN(n13948) );
  INV_X1 U15047 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13350) );
  NAND2_X1 U15048 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13349) );
  NAND2_X1 U15049 ( .A1(n13849), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n13348) );
  OAI211_X1 U15050 ( .C1(n13351), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        n13352) );
  NAND2_X1 U15051 ( .A1(n13352), .A2(n13847), .ZN(n13359) );
  INV_X1 U15052 ( .A(n13397), .ZN(n13357) );
  INV_X1 U15053 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U15054 ( .A1(n13355), .A2(n13354), .ZN(n13356) );
  NAND2_X1 U15055 ( .A1(n13357), .A2(n13356), .ZN(n22138) );
  NAND2_X1 U15056 ( .A1(n22138), .A2(n15167), .ZN(n13358) );
  NAND2_X1 U15057 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  NAND2_X1 U15058 ( .A1(n13365), .A2(n13364), .ZN(n13395) );
  AOI22_X1 U15059 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13369) );
  AOI22_X1 U15060 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13368) );
  AOI22_X1 U15061 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13367) );
  AOI22_X1 U15062 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13366) );
  NAND4_X1 U15063 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n13366), .ZN(
        n13375) );
  AOI22_X1 U15064 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U15065 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13372) );
  AOI22_X1 U15066 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13371) );
  AOI22_X1 U15067 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13370) );
  NAND4_X1 U15068 ( .A1(n13373), .A2(n13372), .A3(n13371), .A4(n13370), .ZN(
        n13374) );
  NAND2_X1 U15069 ( .A1(n13893), .A2(n13967), .ZN(n13377) );
  NAND2_X1 U15070 ( .A1(n13899), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n13376) );
  NAND2_X1 U15071 ( .A1(n13377), .A2(n13376), .ZN(n13394) );
  AOI22_X1 U15072 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13381) );
  AOI22_X1 U15073 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13380) );
  AOI22_X1 U15074 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13379) );
  AOI22_X1 U15075 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13378) );
  NAND4_X1 U15076 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n13378), .ZN(
        n13387) );
  AOI22_X1 U15077 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13385) );
  AOI22_X1 U15078 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13384) );
  AOI22_X1 U15079 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U15080 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13382) );
  NAND4_X1 U15081 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13386) );
  NAND2_X1 U15082 ( .A1(n13893), .A2(n13978), .ZN(n13389) );
  NAND2_X1 U15083 ( .A1(n13899), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n13388) );
  INV_X1 U15084 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n15299) );
  NAND2_X1 U15085 ( .A1(n13396), .A2(n22153), .ZN(n13391) );
  INV_X1 U15086 ( .A(n13409), .ZN(n13390) );
  NAND2_X1 U15087 ( .A1(n13391), .A2(n13390), .ZN(n22157) );
  AOI22_X1 U15088 ( .A1(n22157), .A2(n15167), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13392) );
  OAI21_X1 U15089 ( .B1(n13412), .B2(n15299), .A(n13392), .ZN(n13393) );
  AOI21_X1 U15090 ( .B1(n13965), .B2(n13537), .A(n13393), .ZN(n15297) );
  XNOR2_X1 U15091 ( .A(n13395), .B(n13394), .ZN(n13956) );
  INV_X1 U15092 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13399) );
  OAI21_X1 U15093 ( .B1(n13397), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n13396), .ZN(n22141) );
  AOI22_X1 U15094 ( .A1(n22141), .A2(n15167), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n13398) );
  OAI21_X1 U15095 ( .B1(n13412), .B2(n13399), .A(n13398), .ZN(n13400) );
  AOI21_X1 U15096 ( .B1(n13956), .B2(n13537), .A(n13400), .ZN(n15036) );
  NAND2_X1 U15097 ( .A1(n13402), .A2(n13401), .ZN(n13403) );
  NOR2_X2 U15098 ( .A1(n15035), .A2(n13403), .ZN(n15256) );
  INV_X1 U15099 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13407) );
  NAND2_X1 U15100 ( .A1(n13893), .A2(n13988), .ZN(n13406) );
  OAI21_X1 U15101 ( .B1(n13407), .B2(n13891), .A(n13406), .ZN(n13408) );
  XNOR2_X1 U15102 ( .A(n13987), .B(n13408), .ZN(n13976) );
  NAND2_X1 U15103 ( .A1(n13976), .A2(n13537), .ZN(n13415) );
  INV_X1 U15104 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13411) );
  OAI21_X1 U15105 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13409), .A(
        n13432), .ZN(n22165) );
  AOI22_X1 U15106 ( .A1(n15167), .A2(n22165), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U15107 ( .A1(n13415), .A2(n13414), .ZN(n15255) );
  NAND2_X1 U15108 ( .A1(n15256), .A2(n15255), .ZN(n15254) );
  AOI22_X1 U15109 ( .A1(n13437), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U15110 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13803), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U15111 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n11141), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15112 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13416) );
  NAND4_X1 U15113 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        n13425) );
  AOI22_X1 U15114 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n13834), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U15115 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13232), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U15116 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15117 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13832), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13420) );
  NAND4_X1 U15118 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n13420), .ZN(
        n13424) );
  OAI21_X1 U15119 ( .B1(n13425), .B2(n13424), .A(n13537), .ZN(n13429) );
  NAND2_X1 U15120 ( .A1(n13849), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n13428) );
  INV_X1 U15121 ( .A(n13432), .ZN(n13426) );
  XNOR2_X1 U15122 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n13426), .ZN(
        n15501) );
  AOI22_X1 U15123 ( .A1(n15167), .A2(n15501), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13427) );
  XOR2_X1 U15124 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n13449), .Z(n22183) );
  INV_X1 U15125 ( .A(n22183), .ZN(n13448) );
  AOI22_X1 U15126 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13436) );
  AOI22_X1 U15127 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13435) );
  AOI22_X1 U15128 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15129 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13433) );
  NAND4_X1 U15130 ( .A1(n13436), .A2(n13435), .A3(n13434), .A4(n13433), .ZN(
        n13443) );
  AOI22_X1 U15131 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13441) );
  AOI22_X1 U15132 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U15133 ( .A1(n13576), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U15134 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13438) );
  NAND4_X1 U15135 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13442) );
  OAI21_X1 U15136 ( .B1(n13443), .B2(n13442), .A(n13537), .ZN(n13446) );
  NAND2_X1 U15137 ( .A1(n13849), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n13445) );
  NAND2_X1 U15138 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13444) );
  NAND3_X1 U15139 ( .A1(n13446), .A2(n13445), .A3(n13444), .ZN(n13447) );
  AOI21_X1 U15140 ( .B1(n13448), .B2(n15167), .A(n13447), .ZN(n15353) );
  XNOR2_X1 U15141 ( .A(n13466), .B(n13465), .ZN(n22194) );
  NAND2_X1 U15142 ( .A1(n22194), .A2(n15167), .ZN(n13464) );
  AOI22_X1 U15143 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U15144 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13452) );
  AOI22_X1 U15145 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U15146 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13450) );
  NAND4_X1 U15147 ( .A1(n13453), .A2(n13452), .A3(n13451), .A4(n13450), .ZN(
        n13459) );
  AOI22_X1 U15148 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U15149 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U15150 ( .A1(n13593), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15151 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13454) );
  NAND4_X1 U15152 ( .A1(n13457), .A2(n13456), .A3(n13455), .A4(n13454), .ZN(
        n13458) );
  OAI21_X1 U15153 ( .B1(n13459), .B2(n13458), .A(n13537), .ZN(n13462) );
  NAND2_X1 U15154 ( .A1(n13849), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U15155 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13460) );
  NAND2_X1 U15156 ( .A1(n13464), .A2(n13463), .ZN(n15372) );
  NAND2_X1 U15157 ( .A1(n13849), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n13469) );
  OAI21_X1 U15158 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n13467), .A(
        n13510), .ZN(n22206) );
  AOI22_X1 U15159 ( .A1(n15167), .A2(n22206), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U15160 ( .A1(n13469), .A2(n13468), .ZN(n15559) );
  NAND2_X1 U15161 ( .A1(n15370), .A2(n15559), .ZN(n15558) );
  AOI22_X1 U15162 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13473) );
  AOI22_X1 U15163 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15164 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U15165 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13470) );
  NAND4_X1 U15166 ( .A1(n13473), .A2(n13472), .A3(n13471), .A4(n13470), .ZN(
        n13479) );
  AOI22_X1 U15167 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13477) );
  AOI22_X1 U15168 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13476) );
  AOI22_X1 U15169 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13475) );
  AOI22_X1 U15170 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13474) );
  NAND4_X1 U15171 ( .A1(n13477), .A2(n13476), .A3(n13475), .A4(n13474), .ZN(
        n13478) );
  OR2_X1 U15172 ( .A1(n13479), .A2(n13478), .ZN(n13480) );
  AND2_X1 U15173 ( .A1(n13537), .A2(n13480), .ZN(n15560) );
  NAND2_X1 U15174 ( .A1(n15370), .A2(n15560), .ZN(n13481) );
  XNOR2_X1 U15175 ( .A(n13528), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16371) );
  AOI22_X1 U15176 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U15177 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13484) );
  AOI22_X1 U15178 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15179 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13482) );
  NAND4_X1 U15180 ( .A1(n13485), .A2(n13484), .A3(n13483), .A4(n13482), .ZN(
        n13491) );
  AOI22_X1 U15181 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13489) );
  AOI22_X1 U15182 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13488) );
  AOI22_X1 U15183 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U15184 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13486) );
  NAND4_X1 U15185 ( .A1(n13489), .A2(n13488), .A3(n13487), .A4(n13486), .ZN(
        n13490) );
  OAI21_X1 U15186 ( .B1(n13491), .B2(n13490), .A(n13537), .ZN(n13494) );
  NAND2_X1 U15187 ( .A1(n13849), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n13493) );
  NAND2_X1 U15188 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13492) );
  NAND3_X1 U15189 ( .A1(n13494), .A2(n13493), .A3(n13492), .ZN(n13495) );
  AOI21_X1 U15190 ( .B1(n16371), .B2(n15167), .A(n13495), .ZN(n15619) );
  INV_X1 U15191 ( .A(n15619), .ZN(n13526) );
  XOR2_X1 U15192 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n13496), .Z(
        n16388) );
  AOI22_X1 U15193 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13500) );
  AOI22_X1 U15194 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13499) );
  AOI22_X1 U15195 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13498) );
  AOI22_X1 U15196 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13497) );
  NAND4_X1 U15197 ( .A1(n13500), .A2(n13499), .A3(n13498), .A4(n13497), .ZN(
        n13506) );
  AOI22_X1 U15198 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13504) );
  AOI22_X1 U15199 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13503) );
  AOI22_X1 U15200 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13502) );
  AOI22_X1 U15201 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13501) );
  NAND4_X1 U15202 ( .A1(n13504), .A2(n13503), .A3(n13502), .A4(n13501), .ZN(
        n13505) );
  OR2_X1 U15203 ( .A1(n13506), .A2(n13505), .ZN(n13507) );
  AOI22_X1 U15204 ( .A1(n13537), .A2(n13507), .B1(n15818), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n13509) );
  NAND2_X1 U15205 ( .A1(n13849), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n13508) );
  OAI211_X1 U15206 ( .C1(n16388), .C2(n13847), .A(n13509), .B(n13508), .ZN(
        n16085) );
  XOR2_X1 U15207 ( .A(n13511), .B(n13510), .Z(n22221) );
  AOI22_X1 U15208 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U15209 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13514) );
  AOI22_X1 U15210 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13513) );
  AOI22_X1 U15211 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13512) );
  NAND4_X1 U15212 ( .A1(n13515), .A2(n13514), .A3(n13513), .A4(n13512), .ZN(
        n13521) );
  AOI22_X1 U15213 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13519) );
  AOI22_X1 U15214 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13518) );
  AOI22_X1 U15215 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13517) );
  AOI22_X1 U15216 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13516) );
  NAND4_X1 U15217 ( .A1(n13519), .A2(n13518), .A3(n13517), .A4(n13516), .ZN(
        n13520) );
  OAI21_X1 U15218 ( .B1(n13521), .B2(n13520), .A(n13537), .ZN(n13524) );
  NAND2_X1 U15219 ( .A1(n13849), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n13523) );
  NAND2_X1 U15220 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13522) );
  AND3_X1 U15221 ( .A1(n13524), .A2(n13523), .A3(n13522), .ZN(n13525) );
  OAI21_X1 U15222 ( .B1(n22221), .B2(n13847), .A(n13525), .ZN(n16236) );
  AND2_X1 U15223 ( .A1(n16085), .A2(n16236), .ZN(n15616) );
  XOR2_X1 U15224 ( .A(n22234), .B(n13545), .Z(n22231) );
  INV_X1 U15225 ( .A(n22231), .ZN(n16359) );
  AOI22_X1 U15226 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13532) );
  AOI22_X1 U15227 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13531) );
  AOI22_X1 U15228 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13530) );
  AOI22_X1 U15229 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13529) );
  NAND4_X1 U15230 ( .A1(n13532), .A2(n13531), .A3(n13530), .A4(n13529), .ZN(
        n13539) );
  AOI22_X1 U15231 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13536) );
  AOI22_X1 U15232 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13535) );
  AOI22_X1 U15233 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13534) );
  AOI22_X1 U15234 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13533) );
  NAND4_X1 U15235 ( .A1(n13536), .A2(n13535), .A3(n13534), .A4(n13533), .ZN(
        n13538) );
  OAI21_X1 U15236 ( .B1(n13539), .B2(n13538), .A(n13537), .ZN(n13542) );
  NAND2_X1 U15237 ( .A1(n13849), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13541) );
  NAND2_X1 U15238 ( .A1(n15818), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13540) );
  NAND3_X1 U15239 ( .A1(n13542), .A2(n13541), .A3(n13540), .ZN(n13543) );
  AOI21_X1 U15240 ( .B1(n16359), .B2(n15167), .A(n13543), .ZN(n16137) );
  INV_X1 U15241 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n22236) );
  XNOR2_X1 U15242 ( .A(n13561), .B(n22236), .ZN(n22239) );
  NAND2_X1 U15243 ( .A1(n22239), .A2(n15167), .ZN(n13560) );
  AOI22_X1 U15244 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13549) );
  AOI22_X1 U15245 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13548) );
  AOI22_X1 U15246 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13547) );
  AOI22_X1 U15247 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13546) );
  NAND4_X1 U15248 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13555) );
  AOI22_X1 U15249 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13232), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13553) );
  AOI22_X1 U15250 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n13763), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U15251 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n11141), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13551) );
  AOI22_X1 U15252 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n13832), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13550) );
  NAND4_X1 U15253 ( .A1(n13553), .A2(n13552), .A3(n13551), .A4(n13550), .ZN(
        n13554) );
  NOR2_X1 U15254 ( .A1(n13555), .A2(n13554), .ZN(n13558) );
  AOI21_X1 U15255 ( .B1(n22236), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13556) );
  AOI21_X1 U15256 ( .B1(n13849), .B2(P1_EAX_REG_16__SCAN_IN), .A(n13556), .ZN(
        n13557) );
  OAI21_X1 U15257 ( .B1(n13822), .B2(n13558), .A(n13557), .ZN(n13559) );
  NAND2_X1 U15258 ( .A1(n13560), .A2(n13559), .ZN(n16131) );
  XOR2_X1 U15259 ( .A(n22247), .B(n13574), .Z(n22252) );
  AOI22_X1 U15260 ( .A1(n13293), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n15818), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13573) );
  AOI22_X1 U15261 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13565) );
  AOI22_X1 U15262 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13564) );
  AOI22_X1 U15263 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13563) );
  AOI22_X1 U15264 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13562) );
  NAND4_X1 U15265 ( .A1(n13565), .A2(n13564), .A3(n13563), .A4(n13562), .ZN(
        n13571) );
  AOI22_X1 U15266 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13569) );
  AOI22_X1 U15267 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13568) );
  AOI22_X1 U15268 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15269 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13566) );
  NAND4_X1 U15270 ( .A1(n13569), .A2(n13568), .A3(n13567), .A4(n13566), .ZN(
        n13570) );
  OAI21_X1 U15271 ( .B1(n13571), .B2(n13570), .A(n13844), .ZN(n13572) );
  OAI211_X1 U15272 ( .C1(n22252), .C2(n13847), .A(n13573), .B(n13572), .ZN(
        n16216) );
  INV_X1 U15273 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13575) );
  XNOR2_X1 U15274 ( .A(n13608), .B(n13575), .ZN(n16339) );
  NAND2_X1 U15275 ( .A1(n16339), .A2(n15167), .ZN(n13592) );
  AOI22_X1 U15276 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13580) );
  AOI22_X1 U15277 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13579) );
  AOI22_X1 U15278 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13578) );
  AOI22_X1 U15279 ( .A1(n13804), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13577) );
  NAND4_X1 U15280 ( .A1(n13580), .A2(n13579), .A3(n13578), .A4(n13577), .ZN(
        n13588) );
  NAND2_X1 U15281 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13582) );
  NAND2_X1 U15282 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13581) );
  AND3_X1 U15283 ( .A1(n13582), .A2(n13581), .A3(n13847), .ZN(n13586) );
  AOI22_X1 U15284 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13585) );
  AOI22_X1 U15285 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13584) );
  AOI22_X1 U15286 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11139), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13583) );
  NAND4_X1 U15287 ( .A1(n13586), .A2(n13585), .A3(n13584), .A4(n13583), .ZN(
        n13587) );
  NAND2_X1 U15288 ( .A1(n13822), .A2(n13847), .ZN(n13660) );
  OAI21_X1 U15289 ( .B1(n13588), .B2(n13587), .A(n13660), .ZN(n13590) );
  AOI22_X1 U15290 ( .A1(n13293), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n22605), .ZN(n13589) );
  NAND2_X1 U15291 ( .A1(n13590), .A2(n13589), .ZN(n13591) );
  AOI22_X1 U15292 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13597) );
  AOI22_X1 U15293 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13593), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U15294 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13595) );
  AOI22_X1 U15295 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13594) );
  NAND4_X1 U15296 ( .A1(n13597), .A2(n13596), .A3(n13595), .A4(n13594), .ZN(
        n13603) );
  AOI22_X1 U15297 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13601) );
  AOI22_X1 U15298 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U15299 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13599) );
  AOI22_X1 U15300 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13598) );
  NAND4_X1 U15301 ( .A1(n13601), .A2(n13600), .A3(n13599), .A4(n13598), .ZN(
        n13602) );
  NOR2_X1 U15302 ( .A1(n13603), .A2(n13602), .ZN(n13607) );
  NAND2_X1 U15303 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13604) );
  NAND2_X1 U15304 ( .A1(n13847), .A2(n13604), .ZN(n13605) );
  AOI21_X1 U15305 ( .B1(n13849), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13605), .ZN(
        n13606) );
  OAI21_X1 U15306 ( .B1(n13822), .B2(n13607), .A(n13606), .ZN(n13612) );
  OAI21_X1 U15307 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n13609), .A(
        n13643), .ZN(n22266) );
  INV_X1 U15308 ( .A(n22266), .ZN(n13610) );
  NAND2_X1 U15309 ( .A1(n13610), .A2(n15167), .ZN(n13611) );
  NAND2_X1 U15310 ( .A1(n13612), .A2(n13611), .ZN(n16122) );
  NOR2_X2 U15311 ( .A1(n16070), .A2(n16122), .ZN(n16057) );
  AOI22_X1 U15312 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13827), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13618) );
  AOI22_X1 U15313 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13617) );
  AOI22_X1 U15314 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13616) );
  AOI21_X1 U15315 ( .B1(n13758), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n15167), .ZN(n13614) );
  NAND2_X1 U15316 ( .A1(n13835), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13613) );
  AND2_X1 U15317 ( .A1(n13614), .A2(n13613), .ZN(n13615) );
  NAND4_X1 U15318 ( .A1(n13618), .A2(n13617), .A3(n13616), .A4(n13615), .ZN(
        n13624) );
  AOI22_X1 U15319 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11142), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13622) );
  AOI22_X1 U15320 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U15321 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13620) );
  AOI22_X1 U15322 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13619) );
  NAND4_X1 U15323 ( .A1(n13622), .A2(n13621), .A3(n13620), .A4(n13619), .ZN(
        n13623) );
  OR2_X1 U15324 ( .A1(n13624), .A2(n13623), .ZN(n13625) );
  NAND2_X1 U15325 ( .A1(n13660), .A2(n13625), .ZN(n13628) );
  AOI22_X1 U15326 ( .A1(n13293), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n22605), .ZN(n13627) );
  XNOR2_X1 U15327 ( .A(n13643), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16334) );
  AOI21_X1 U15328 ( .B1(n13628), .B2(n13627), .A(n13626), .ZN(n16059) );
  AND2_X2 U15329 ( .A1(n16057), .A2(n16059), .ZN(n16044) );
  AOI22_X1 U15330 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13632) );
  AOI22_X1 U15331 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13631) );
  AOI22_X1 U15332 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13630) );
  AOI22_X1 U15333 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13629) );
  NAND4_X1 U15334 ( .A1(n13632), .A2(n13631), .A3(n13630), .A4(n13629), .ZN(
        n13638) );
  AOI22_X1 U15335 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13636) );
  AOI22_X1 U15336 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13635) );
  AOI22_X1 U15337 ( .A1(n11142), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13634) );
  AOI22_X1 U15338 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13633) );
  NAND4_X1 U15339 ( .A1(n13636), .A2(n13635), .A3(n13634), .A4(n13633), .ZN(
        n13637) );
  NOR2_X1 U15340 ( .A1(n13638), .A2(n13637), .ZN(n13642) );
  NAND2_X1 U15341 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13639) );
  NAND2_X1 U15342 ( .A1(n13847), .A2(n13639), .ZN(n13640) );
  AOI21_X1 U15343 ( .B1(n13849), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13640), .ZN(
        n13641) );
  OAI21_X1 U15344 ( .B1(n13822), .B2(n13642), .A(n13641), .ZN(n13649) );
  INV_X1 U15345 ( .A(n13645), .ZN(n13646) );
  INV_X1 U15346 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16321) );
  NAND2_X1 U15347 ( .A1(n13646), .A2(n16321), .ZN(n13647) );
  AND2_X1 U15348 ( .A1(n13690), .A2(n13647), .ZN(n16325) );
  NAND2_X1 U15349 ( .A1(n16325), .A2(n15167), .ZN(n13648) );
  AOI22_X1 U15350 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13653) );
  AOI22_X1 U15351 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U15352 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13651) );
  AOI22_X1 U15353 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13650) );
  NAND4_X1 U15354 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13662) );
  NAND2_X1 U15355 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13655) );
  NAND2_X1 U15356 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13654) );
  AND3_X1 U15357 ( .A1(n13655), .A2(n13654), .A3(n13847), .ZN(n13659) );
  AOI22_X1 U15358 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13827), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U15359 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13657) );
  AOI22_X1 U15360 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13656) );
  NAND4_X1 U15361 ( .A1(n13659), .A2(n13658), .A3(n13657), .A4(n13656), .ZN(
        n13661) );
  OAI21_X1 U15362 ( .B1(n13662), .B2(n13661), .A(n13660), .ZN(n13664) );
  AOI22_X1 U15363 ( .A1(n13293), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n22605), .ZN(n13663) );
  NAND2_X1 U15364 ( .A1(n13664), .A2(n13663), .ZN(n13666) );
  XNOR2_X1 U15365 ( .A(n13690), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16311) );
  NAND2_X1 U15366 ( .A1(n16311), .A2(n15167), .ZN(n13665) );
  NAND2_X1 U15367 ( .A1(n13666), .A2(n13665), .ZN(n16028) );
  AOI22_X1 U15368 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n13827), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U15369 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n13232), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U15370 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U15371 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13667) );
  NAND4_X1 U15372 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13676) );
  AOI22_X1 U15373 ( .A1(n13107), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U15374 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n11141), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U15375 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U15376 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U15377 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13675) );
  NOR2_X1 U15378 ( .A1(n13676), .A2(n13675), .ZN(n13698) );
  AOI22_X1 U15379 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13827), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U15380 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13679) );
  AOI22_X1 U15381 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13678) );
  AOI22_X1 U15382 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13677) );
  NAND4_X1 U15383 ( .A1(n13680), .A2(n13679), .A3(n13678), .A4(n13677), .ZN(
        n13686) );
  AOI22_X1 U15384 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11139), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13684) );
  AOI22_X1 U15385 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13683) );
  AOI22_X1 U15386 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13682) );
  AOI22_X1 U15387 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13681) );
  NAND4_X1 U15388 ( .A1(n13684), .A2(n13683), .A3(n13682), .A4(n13681), .ZN(
        n13685) );
  NOR2_X1 U15389 ( .A1(n13686), .A2(n13685), .ZN(n13697) );
  XNOR2_X1 U15390 ( .A(n13698), .B(n13697), .ZN(n13689) );
  INV_X1 U15391 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13692) );
  AOI21_X1 U15392 ( .B1(n13692), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13687) );
  AOI21_X1 U15393 ( .B1(n13849), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13687), .ZN(
        n13688) );
  OAI21_X1 U15394 ( .B1(n13822), .B2(n13689), .A(n13688), .ZN(n13696) );
  NAND2_X1 U15395 ( .A1(n13693), .A2(n13692), .ZN(n13694) );
  NAND2_X1 U15396 ( .A1(n13732), .A2(n13694), .ZN(n16303) );
  NOR2_X1 U15397 ( .A1(n13698), .A2(n13697), .ZN(n13717) );
  AOI22_X1 U15398 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U15399 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U15400 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U15401 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U15402 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13708) );
  AOI22_X1 U15403 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U15404 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U15405 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U15406 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13703) );
  NAND4_X1 U15407 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13707) );
  OR2_X1 U15408 ( .A1(n13708), .A2(n13707), .ZN(n13716) );
  INV_X1 U15409 ( .A(n13716), .ZN(n13709) );
  XNOR2_X1 U15410 ( .A(n13717), .B(n13709), .ZN(n13710) );
  NAND2_X1 U15411 ( .A1(n13710), .A2(n13844), .ZN(n13715) );
  NAND2_X1 U15412 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13711) );
  NAND2_X1 U15413 ( .A1(n13847), .A2(n13711), .ZN(n13712) );
  AOI21_X1 U15414 ( .B1(n13849), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13712), .ZN(
        n13714) );
  XNOR2_X1 U15415 ( .A(n13732), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16298) );
  AOI21_X1 U15416 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n16011) );
  NAND2_X1 U15417 ( .A1(n13717), .A2(n13716), .ZN(n13738) );
  AOI22_X1 U15418 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13721) );
  AOI22_X1 U15419 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U15420 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13719) );
  AOI22_X1 U15421 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13718) );
  NAND4_X1 U15422 ( .A1(n13721), .A2(n13720), .A3(n13719), .A4(n13718), .ZN(
        n13727) );
  AOI22_X1 U15423 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13811), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13725) );
  AOI22_X1 U15424 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13724) );
  AOI22_X1 U15425 ( .A1(n13833), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13723) );
  AOI22_X1 U15426 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13722) );
  NAND4_X1 U15427 ( .A1(n13725), .A2(n13724), .A3(n13723), .A4(n13722), .ZN(
        n13726) );
  NOR2_X1 U15428 ( .A1(n13727), .A2(n13726), .ZN(n13739) );
  XNOR2_X1 U15429 ( .A(n13738), .B(n13739), .ZN(n13731) );
  NAND2_X1 U15430 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13728) );
  NAND2_X1 U15431 ( .A1(n13847), .A2(n13728), .ZN(n13729) );
  AOI21_X1 U15432 ( .B1(n13849), .B2(P1_EAX_REG_25__SCAN_IN), .A(n13729), .ZN(
        n13730) );
  OAI21_X1 U15433 ( .B1(n13731), .B2(n13822), .A(n13730), .ZN(n13737) );
  INV_X1 U15434 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16285) );
  NAND2_X1 U15435 ( .A1(n13734), .A2(n16285), .ZN(n13735) );
  NAND2_X1 U15436 ( .A1(n16289), .A2(n15167), .ZN(n13736) );
  NOR2_X1 U15437 ( .A1(n13739), .A2(n13738), .ZN(n13757) );
  AOI22_X1 U15438 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13743) );
  AOI22_X1 U15439 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13742) );
  AOI22_X1 U15440 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13741) );
  AOI22_X1 U15441 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13740) );
  NAND4_X1 U15442 ( .A1(n13743), .A2(n13742), .A3(n13741), .A4(n13740), .ZN(
        n13749) );
  AOI22_X1 U15443 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13747) );
  AOI22_X1 U15444 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U15445 ( .A1(n11142), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13745) );
  AOI22_X1 U15446 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13744) );
  NAND4_X1 U15447 ( .A1(n13747), .A2(n13746), .A3(n13745), .A4(n13744), .ZN(
        n13748) );
  OR2_X1 U15448 ( .A1(n13749), .A2(n13748), .ZN(n13756) );
  XNOR2_X1 U15449 ( .A(n13757), .B(n13756), .ZN(n13753) );
  NAND2_X1 U15450 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13750) );
  NAND2_X1 U15451 ( .A1(n13847), .A2(n13750), .ZN(n13751) );
  AOI21_X1 U15452 ( .B1(n13849), .B2(P1_EAX_REG_26__SCAN_IN), .A(n13751), .ZN(
        n13752) );
  OAI21_X1 U15453 ( .B1(n13753), .B2(n13822), .A(n13752), .ZN(n13755) );
  XNOR2_X1 U15454 ( .A(n13774), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16276) );
  NAND2_X1 U15455 ( .A1(n16276), .A2(n15167), .ZN(n13754) );
  NAND2_X1 U15456 ( .A1(n13755), .A2(n13754), .ZN(n15980) );
  NAND2_X1 U15457 ( .A1(n13757), .A2(n13756), .ZN(n13781) );
  AOI22_X1 U15458 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U15459 ( .A1(n13803), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U15460 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13760) );
  AOI22_X1 U15461 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13759) );
  NAND4_X1 U15462 ( .A1(n13762), .A2(n13761), .A3(n13760), .A4(n13759), .ZN(
        n13769) );
  AOI22_X1 U15463 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13763), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13767) );
  AOI22_X1 U15464 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13766) );
  AOI22_X1 U15465 ( .A1(n11139), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13765) );
  AOI22_X1 U15466 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13764) );
  NAND4_X1 U15467 ( .A1(n13767), .A2(n13766), .A3(n13765), .A4(n13764), .ZN(
        n13768) );
  NOR2_X1 U15468 ( .A1(n13769), .A2(n13768), .ZN(n13782) );
  XNOR2_X1 U15469 ( .A(n13781), .B(n13782), .ZN(n13773) );
  NAND2_X1 U15470 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13770) );
  NAND2_X1 U15471 ( .A1(n13847), .A2(n13770), .ZN(n13771) );
  AOI21_X1 U15472 ( .B1(n13849), .B2(P1_EAX_REG_27__SCAN_IN), .A(n13771), .ZN(
        n13772) );
  OAI21_X1 U15473 ( .B1(n13773), .B2(n13822), .A(n13772), .ZN(n13779) );
  INV_X1 U15474 ( .A(n13774), .ZN(n13775) );
  NAND2_X1 U15475 ( .A1(n13775), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13776) );
  INV_X1 U15476 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15972) );
  NAND2_X1 U15477 ( .A1(n13776), .A2(n15972), .ZN(n13777) );
  NAND2_X1 U15478 ( .A1(n13799), .A2(n13777), .ZN(n16270) );
  NOR2_X1 U15479 ( .A1(n13782), .A2(n13781), .ZN(n13819) );
  AOI22_X1 U15480 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11137), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13786) );
  AOI22_X1 U15481 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13785) );
  AOI22_X1 U15482 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13784) );
  AOI22_X1 U15483 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13783) );
  NAND4_X1 U15484 ( .A1(n13786), .A2(n13785), .A3(n13784), .A4(n13783), .ZN(
        n13792) );
  AOI22_X1 U15485 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13805), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13790) );
  AOI22_X1 U15486 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13789) );
  AOI22_X1 U15487 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13788) );
  AOI22_X1 U15488 ( .A1(n13832), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13787) );
  NAND4_X1 U15489 ( .A1(n13790), .A2(n13789), .A3(n13788), .A4(n13787), .ZN(
        n13791) );
  OR2_X1 U15490 ( .A1(n13792), .A2(n13791), .ZN(n13818) );
  INV_X1 U15491 ( .A(n13818), .ZN(n13793) );
  XNOR2_X1 U15492 ( .A(n13819), .B(n13793), .ZN(n13794) );
  NAND2_X1 U15493 ( .A1(n13794), .A2(n13844), .ZN(n13798) );
  INV_X1 U15494 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16252) );
  AOI21_X1 U15495 ( .B1(n16252), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13795) );
  AOI21_X1 U15496 ( .B1(n13849), .B2(P1_EAX_REG_28__SCAN_IN), .A(n13795), .ZN(
        n13797) );
  XNOR2_X1 U15497 ( .A(n13799), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16254) );
  INV_X1 U15498 ( .A(n13800), .ZN(n13801) );
  INV_X1 U15499 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15946) );
  NAND2_X1 U15500 ( .A1(n13801), .A2(n15946), .ZN(n13802) );
  NAND2_X1 U15501 ( .A1(n15170), .A2(n13802), .ZN(n16248) );
  AOI22_X1 U15502 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U15503 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13809) );
  AOI22_X1 U15504 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13808) );
  AOI22_X1 U15505 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13807) );
  NAND4_X1 U15506 ( .A1(n13810), .A2(n13809), .A3(n13808), .A4(n13807), .ZN(
        n13817) );
  AOI22_X1 U15507 ( .A1(n13811), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14692), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13815) );
  AOI22_X1 U15508 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13814) );
  AOI22_X1 U15509 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13813) );
  AOI22_X1 U15510 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13812) );
  NAND4_X1 U15511 ( .A1(n13815), .A2(n13814), .A3(n13813), .A4(n13812), .ZN(
        n13816) );
  NOR2_X1 U15512 ( .A1(n13817), .A2(n13816), .ZN(n13826) );
  NAND2_X1 U15513 ( .A1(n13819), .A2(n13818), .ZN(n13825) );
  XNOR2_X1 U15514 ( .A(n13826), .B(n13825), .ZN(n13823) );
  AOI21_X1 U15515 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n22605), .A(
        n15167), .ZN(n13821) );
  NAND2_X1 U15516 ( .A1(n13293), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n13820) );
  OAI211_X1 U15517 ( .C1(n13823), .C2(n13822), .A(n13821), .B(n13820), .ZN(
        n13824) );
  OAI21_X1 U15518 ( .B1(n13847), .B2(n16248), .A(n13824), .ZN(n15943) );
  NOR2_X1 U15519 ( .A1(n13826), .A2(n13825), .ZN(n13843) );
  AOI22_X1 U15520 ( .A1(n13806), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11136), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U15521 ( .A1(n13827), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13803), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13830) );
  AOI22_X1 U15522 ( .A1(n14692), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13758), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13829) );
  AOI22_X1 U15523 ( .A1(n13232), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13804), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13828) );
  NAND4_X1 U15524 ( .A1(n13831), .A2(n13830), .A3(n13829), .A4(n13828), .ZN(
        n13841) );
  AOI22_X1 U15525 ( .A1(n11141), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n13832), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13839) );
  AOI22_X1 U15526 ( .A1(n13834), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13833), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13838) );
  AOI22_X1 U15527 ( .A1(n13763), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13576), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13837) );
  AOI22_X1 U15528 ( .A1(n13805), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13835), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13836) );
  NAND4_X1 U15529 ( .A1(n13839), .A2(n13838), .A3(n13837), .A4(n13836), .ZN(
        n13840) );
  NOR2_X1 U15530 ( .A1(n13841), .A2(n13840), .ZN(n13842) );
  XNOR2_X1 U15531 ( .A(n13843), .B(n13842), .ZN(n13845) );
  NAND2_X1 U15532 ( .A1(n13845), .A2(n13844), .ZN(n13852) );
  NAND2_X1 U15533 ( .A1(n22605), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13846) );
  NAND2_X1 U15534 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  AOI21_X1 U15535 ( .B1(n13849), .B2(P1_EAX_REG_30__SCAN_IN), .A(n13848), .ZN(
        n13851) );
  XNOR2_X1 U15536 ( .A(n15170), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15936) );
  AOI21_X1 U15537 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(n15817) );
  NAND3_X1 U15538 ( .A1(n17473), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n22290) );
  INV_X1 U15539 ( .A(n22290), .ZN(n13853) );
  INV_X1 U15540 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13916) );
  NAND2_X1 U15541 ( .A1(n13854), .A2(n13157), .ZN(n13855) );
  AND2_X1 U15542 ( .A1(n13856), .A2(n13855), .ZN(n14540) );
  NAND2_X1 U15543 ( .A1(n16573), .A2(n15177), .ZN(n13857) );
  NAND2_X1 U15544 ( .A1(n22584), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13859) );
  NAND2_X1 U15545 ( .A1(n14727), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n13858) );
  NAND2_X1 U15546 ( .A1(n13859), .A2(n13858), .ZN(n13874) );
  NAND2_X1 U15547 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n22571), .ZN(
        n13878) );
  NAND2_X1 U15548 ( .A1(n13860), .A2(n13859), .ZN(n13890) );
  XNOR2_X1 U15549 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13888) );
  NAND2_X1 U15550 ( .A1(n13890), .A2(n13888), .ZN(n13862) );
  NAND2_X1 U15551 ( .A1(n22585), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13861) );
  NAND2_X1 U15552 ( .A1(n13862), .A2(n13861), .ZN(n13872) );
  NAND2_X1 U15553 ( .A1(n22586), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13864) );
  NAND2_X1 U15554 ( .A1(n13305), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13863) );
  NAND2_X1 U15555 ( .A1(n13872), .A2(n13871), .ZN(n13866) );
  INV_X1 U15556 ( .A(n13864), .ZN(n13870) );
  AOI21_X1 U15557 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17477), .A(
        n13870), .ZN(n13865) );
  NAND2_X1 U15558 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  NAND2_X1 U15559 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13350), .ZN(
        n13869) );
  OAI22_X1 U15560 ( .A1(n13872), .A2(n13871), .B1(n13870), .B2(n13869), .ZN(
        n14413) );
  INV_X1 U15561 ( .A(n14413), .ZN(n13902) );
  INV_X1 U15562 ( .A(n13893), .ZN(n13876) );
  INV_X1 U15563 ( .A(n13878), .ZN(n13873) );
  XNOR2_X1 U15564 ( .A(n13874), .B(n13873), .ZN(n14411) );
  OAI22_X1 U15565 ( .A1(n17473), .A2(n13157), .B1(n13891), .B2(n14411), .ZN(
        n13881) );
  INV_X1 U15566 ( .A(n13881), .ZN(n13875) );
  OAI21_X1 U15567 ( .B1(n13876), .B2(n14797), .A(n13875), .ZN(n13887) );
  INV_X1 U15568 ( .A(n14411), .ZN(n13877) );
  OAI21_X1 U15569 ( .B1(n13893), .B2(n13984), .A(n13877), .ZN(n13886) );
  OAI21_X1 U15570 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n22571), .A(
        n13878), .ZN(n13880) );
  INV_X1 U15571 ( .A(n13880), .ZN(n13879) );
  NAND2_X1 U15572 ( .A1(n13893), .A2(n13879), .ZN(n13884) );
  AOI21_X1 U15573 ( .B1(n14825), .B2(n14886), .A(n15178), .ZN(n13894) );
  AOI211_X1 U15574 ( .C1(n14537), .C2(n14886), .A(n13880), .B(n13894), .ZN(
        n13883) );
  NOR3_X1 U15575 ( .A1(n15178), .A2(n14411), .A3(n13881), .ZN(n13882) );
  AOI211_X1 U15576 ( .C1(n13901), .C2(n13884), .A(n13883), .B(n13882), .ZN(
        n13885) );
  AOI21_X1 U15577 ( .B1(n13887), .B2(n13886), .A(n13885), .ZN(n13897) );
  INV_X1 U15578 ( .A(n13888), .ZN(n13889) );
  XNOR2_X1 U15579 ( .A(n13890), .B(n13889), .ZN(n14410) );
  NOR2_X1 U15580 ( .A1(n14410), .A2(n13891), .ZN(n13892) );
  AOI211_X1 U15581 ( .C1(n14410), .C2(n13893), .A(n13892), .B(n13894), .ZN(
        n13896) );
  NAND3_X1 U15582 ( .A1(n14410), .A2(n13894), .A3(n13893), .ZN(n13895) );
  OAI21_X1 U15583 ( .B1(n13897), .B2(n13896), .A(n13895), .ZN(n13898) );
  OAI21_X1 U15584 ( .B1(n13899), .B2(n13902), .A(n13898), .ZN(n13900) );
  OAI21_X1 U15585 ( .B1(n13902), .B2(n13901), .A(n13900), .ZN(n13903) );
  AOI21_X1 U15586 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n17473), .A(
        n13903), .ZN(n13904) );
  INV_X1 U15587 ( .A(n13904), .ZN(n13905) );
  NOR2_X1 U15588 ( .A1(n14712), .A2(n13115), .ZN(n13909) );
  NAND2_X1 U15589 ( .A1(n14533), .A2(n13909), .ZN(n17449) );
  NAND2_X1 U15590 ( .A1(n22607), .A2(n13914), .ZN(n21944) );
  NAND2_X1 U15591 ( .A1(n21944), .A2(n17473), .ZN(n13911) );
  NAND2_X1 U15592 ( .A1(n17473), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13913) );
  INV_X1 U15593 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n22590) );
  NAND2_X1 U15594 ( .A1(n22590), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13912) );
  AND2_X1 U15595 ( .A1(n13913), .A2(n13912), .ZN(n14579) );
  NAND2_X1 U15596 ( .A1(n20625), .A2(n15936), .ZN(n13915) );
  INV_X2 U15597 ( .A(n22044), .ZN(n22108) );
  NAND2_X1 U15598 ( .A1(n22108), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n16423) );
  OAI211_X1 U15599 ( .C1(n13916), .C2(n16384), .A(n13915), .B(n16423), .ZN(
        n13917) );
  AOI21_X1 U15600 ( .B1(n15932), .B2(n20614), .A(n13917), .ZN(n14015) );
  NAND2_X1 U15601 ( .A1(n13926), .A2(n13927), .ZN(n13938) );
  NAND2_X1 U15602 ( .A1(n13938), .A2(n13937), .ZN(n13950) );
  INV_X1 U15603 ( .A(n13949), .ZN(n13918) );
  XNOR2_X1 U15604 ( .A(n13950), .B(n13918), .ZN(n13919) );
  NAND2_X1 U15605 ( .A1(n13919), .A2(n17464), .ZN(n13920) );
  NAND2_X1 U15606 ( .A1(n13921), .A2(n13920), .ZN(n13946) );
  INV_X1 U15607 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21992) );
  XNOR2_X1 U15608 ( .A(n13946), .B(n21992), .ZN(n14990) );
  NAND2_X1 U15609 ( .A1(n15177), .A2(n13922), .ZN(n13939) );
  OAI21_X1 U15610 ( .B1(n21947), .B2(n13927), .A(n13939), .ZN(n13923) );
  INV_X1 U15611 ( .A(n13923), .ZN(n13924) );
  NAND2_X1 U15612 ( .A1(n14514), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14515) );
  OR2_X1 U15613 ( .A1(n13925), .A2(n13984), .ZN(n13931) );
  OAI21_X1 U15614 ( .B1(n13927), .B2(n13926), .A(n13938), .ZN(n13928) );
  OAI211_X1 U15615 ( .C1(n13928), .C2(n21947), .A(n11614), .B(n13157), .ZN(
        n13929) );
  INV_X1 U15616 ( .A(n13929), .ZN(n13930) );
  NAND2_X1 U15617 ( .A1(n13931), .A2(n13930), .ZN(n13932) );
  XNOR2_X1 U15618 ( .A(n14515), .B(n13932), .ZN(n14616) );
  NAND2_X1 U15619 ( .A1(n14616), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15030) );
  INV_X1 U15620 ( .A(n13932), .ZN(n13933) );
  OR2_X1 U15621 ( .A1(n14515), .A2(n13933), .ZN(n13934) );
  NAND2_X1 U15622 ( .A1(n15030), .A2(n13934), .ZN(n13944) );
  INV_X1 U15623 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21974) );
  XNOR2_X1 U15624 ( .A(n13944), .B(n21974), .ZN(n14997) );
  NAND2_X1 U15625 ( .A1(n13936), .A2(n13975), .ZN(n13943) );
  XNOR2_X1 U15626 ( .A(n13938), .B(n13937), .ZN(n13941) );
  INV_X1 U15627 ( .A(n13939), .ZN(n13940) );
  AOI21_X1 U15628 ( .B1(n13941), .B2(n17464), .A(n13940), .ZN(n13942) );
  NAND2_X1 U15629 ( .A1(n13943), .A2(n13942), .ZN(n14996) );
  NAND2_X1 U15630 ( .A1(n14997), .A2(n14996), .ZN(n14995) );
  NAND2_X1 U15631 ( .A1(n13944), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13945) );
  NAND2_X1 U15632 ( .A1(n14995), .A2(n13945), .ZN(n14989) );
  NAND2_X1 U15633 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  NAND2_X1 U15634 ( .A1(n13946), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13947) );
  NAND2_X1 U15635 ( .A1(n14988), .A2(n13947), .ZN(n20577) );
  NAND2_X1 U15636 ( .A1(n13948), .A2(n13975), .ZN(n13953) );
  NAND2_X1 U15637 ( .A1(n13950), .A2(n13949), .ZN(n13959) );
  XNOR2_X1 U15638 ( .A(n13959), .B(n13957), .ZN(n13951) );
  NAND2_X1 U15639 ( .A1(n13951), .A2(n17464), .ZN(n13952) );
  NAND2_X1 U15640 ( .A1(n13953), .A2(n13952), .ZN(n13954) );
  INV_X1 U15641 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21986) );
  XNOR2_X1 U15642 ( .A(n13954), .B(n21986), .ZN(n20576) );
  NAND2_X1 U15643 ( .A1(n20577), .A2(n20576), .ZN(n20575) );
  NAND2_X1 U15644 ( .A1(n13954), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13955) );
  NAND2_X1 U15645 ( .A1(n20575), .A2(n13955), .ZN(n20583) );
  NAND2_X1 U15646 ( .A1(n13956), .A2(n13975), .ZN(n13962) );
  INV_X1 U15647 ( .A(n13957), .ZN(n13958) );
  OR2_X1 U15648 ( .A1(n13959), .A2(n13958), .ZN(n13966) );
  XNOR2_X1 U15649 ( .A(n13966), .B(n13967), .ZN(n13960) );
  NAND2_X1 U15650 ( .A1(n13960), .A2(n17464), .ZN(n13961) );
  NAND2_X1 U15651 ( .A1(n13962), .A2(n13961), .ZN(n13963) );
  INV_X1 U15652 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21954) );
  XNOR2_X1 U15653 ( .A(n13963), .B(n21954), .ZN(n20582) );
  NAND2_X1 U15654 ( .A1(n20583), .A2(n20582), .ZN(n20581) );
  NAND2_X1 U15655 ( .A1(n13963), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13964) );
  NAND2_X1 U15656 ( .A1(n20581), .A2(n13964), .ZN(n20588) );
  NAND3_X1 U15657 ( .A1(n13987), .A2(n13975), .A3(n13965), .ZN(n13971) );
  INV_X1 U15658 ( .A(n13966), .ZN(n13968) );
  NAND2_X1 U15659 ( .A1(n13968), .A2(n13967), .ZN(n13977) );
  XNOR2_X1 U15660 ( .A(n13977), .B(n13978), .ZN(n13969) );
  NAND2_X1 U15661 ( .A1(n13969), .A2(n17464), .ZN(n13970) );
  NAND2_X1 U15662 ( .A1(n13971), .A2(n13970), .ZN(n13972) );
  XNOR2_X1 U15663 ( .A(n13972), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20587) );
  INV_X1 U15664 ( .A(n13972), .ZN(n13973) );
  INV_X1 U15665 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21999) );
  NAND2_X1 U15666 ( .A1(n13973), .A2(n21999), .ZN(n13974) );
  NAND2_X1 U15667 ( .A1(n13976), .A2(n13975), .ZN(n13982) );
  INV_X1 U15668 ( .A(n13977), .ZN(n13979) );
  NAND2_X1 U15669 ( .A1(n13979), .A2(n13978), .ZN(n13990) );
  XNOR2_X1 U15670 ( .A(n13990), .B(n13988), .ZN(n13980) );
  NAND2_X1 U15671 ( .A1(n13980), .A2(n17464), .ZN(n13981) );
  NOR2_X1 U15672 ( .A1(n13985), .A2(n13984), .ZN(n13986) );
  NAND2_X1 U15673 ( .A1(n17464), .A2(n13988), .ZN(n13989) );
  OR2_X1 U15674 ( .A1(n13990), .A2(n13989), .ZN(n13991) );
  NAND2_X1 U15675 ( .A1(n13994), .A2(n13991), .ZN(n13992) );
  INV_X1 U15676 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n22030) );
  XNOR2_X1 U15677 ( .A(n13992), .B(n22030), .ZN(n15498) );
  NAND2_X1 U15678 ( .A1(n13992), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13993) );
  INV_X1 U15679 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n22038) );
  NAND2_X1 U15680 ( .A1(n20603), .A2(n22038), .ZN(n13995) );
  NAND2_X1 U15681 ( .A1(n11153), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16366) );
  INV_X1 U15682 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U15683 ( .A1(n13994), .A2(n14268), .ZN(n13996) );
  NAND2_X1 U15684 ( .A1(n16366), .A2(n13996), .ZN(n16381) );
  INV_X1 U15685 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n22053) );
  NAND2_X1 U15686 ( .A1(n13994), .A2(n22053), .ZN(n16380) );
  NAND2_X1 U15687 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13997) );
  NAND2_X1 U15688 ( .A1(n13994), .A2(n13997), .ZN(n16378) );
  NAND2_X1 U15689 ( .A1(n16380), .A2(n16378), .ZN(n13998) );
  NOR2_X1 U15690 ( .A1(n16381), .A2(n13998), .ZN(n16364) );
  INV_X1 U15691 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21957) );
  NAND2_X1 U15692 ( .A1(n13994), .A2(n21957), .ZN(n13999) );
  NAND2_X1 U15693 ( .A1(n16364), .A2(n13999), .ZN(n16346) );
  NAND2_X1 U15694 ( .A1(n16346), .A2(n20603), .ZN(n20618) );
  INV_X1 U15695 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14281) );
  NAND2_X1 U15696 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22078) );
  INV_X1 U15697 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14000) );
  NAND2_X1 U15698 ( .A1(n20617), .A2(n14000), .ZN(n16348) );
  OAI21_X1 U15699 ( .B1(n14281), .B2(n22078), .A(n16348), .ZN(n14001) );
  NAND2_X1 U15700 ( .A1(n20618), .A2(n14001), .ZN(n14010) );
  INV_X1 U15701 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14259) );
  INV_X1 U15702 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14002) );
  NAND2_X1 U15703 ( .A1(n14259), .A2(n14002), .ZN(n14003) );
  NAND2_X1 U15704 ( .A1(n11154), .A2(n14003), .ZN(n16376) );
  NAND2_X1 U15705 ( .A1(n11154), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16379) );
  NAND2_X1 U15706 ( .A1(n16376), .A2(n16379), .ZN(n16365) );
  NAND2_X1 U15707 ( .A1(n11154), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14004) );
  NAND2_X1 U15708 ( .A1(n16366), .A2(n14004), .ZN(n14005) );
  NOR2_X1 U15709 ( .A1(n16365), .A2(n14005), .ZN(n16345) );
  NAND2_X1 U15710 ( .A1(n20617), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14006) );
  NOR2_X1 U15711 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14007) );
  NOR2_X1 U15712 ( .A1(n13994), .A2(n14007), .ZN(n14008) );
  NAND3_X1 U15713 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n22104) );
  INV_X1 U15714 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n22072) );
  NOR2_X1 U15715 ( .A1(n22104), .A2(n22072), .ZN(n14011) );
  NAND2_X1 U15716 ( .A1(n16309), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14013) );
  INV_X1 U15717 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16328) );
  INV_X1 U15718 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16529) );
  INV_X1 U15719 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16510) );
  NAND4_X1 U15720 ( .A1(n16328), .A2(n16529), .A3(n22072), .A4(n16510), .ZN(
        n14012) );
  INV_X1 U15721 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16483) );
  INV_X1 U15722 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16471) );
  INV_X1 U15723 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16479) );
  NAND3_X1 U15724 ( .A1(n16483), .A2(n16471), .A3(n16479), .ZN(n16258) );
  NAND2_X1 U15725 ( .A1(n14013), .A2(n20603), .ZN(n16282) );
  AND2_X1 U15726 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16459) );
  NAND2_X1 U15727 ( .A1(n16459), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16412) );
  NAND2_X1 U15728 ( .A1(n20603), .A2(n16412), .ZN(n16256) );
  AND2_X1 U15729 ( .A1(n16282), .A2(n16256), .ZN(n14014) );
  NOR2_X1 U15730 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16441) );
  XNOR2_X1 U15731 ( .A(n20603), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16246) );
  NAND2_X1 U15732 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16430) );
  INV_X1 U15733 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16403) );
  OR2_X2 U15734 ( .A1(n16837), .A2(n14016), .ZN(n14018) );
  NOR2_X2 U15735 ( .A1(n14018), .A2(n14017), .ZN(n16826) );
  INV_X1 U15736 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17091) );
  NAND2_X1 U15737 ( .A1(n14018), .A2(n14017), .ZN(n16824) );
  OAI21_X1 U15738 ( .B1(n16826), .B2(n17091), .A(n16824), .ZN(n14021) );
  XNOR2_X1 U15739 ( .A(n14019), .B(n14197), .ZN(n14020) );
  XNOR2_X1 U15740 ( .A(n14021), .B(n14020), .ZN(n14213) );
  AOI21_X1 U15741 ( .B1(n14022), .B2(n16671), .A(n16659), .ZN(n19228) );
  OR2_X1 U15742 ( .A1(n14024), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14025) );
  NAND2_X1 U15743 ( .A1(n14023), .A2(n14025), .ZN(n19231) );
  NOR2_X1 U15744 ( .A1(n19294), .A2(n14159), .ZN(n14198) );
  AOI21_X1 U15745 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14198), .ZN(n14026) );
  OAI21_X1 U15746 ( .B1(n17042), .B2(n19231), .A(n14026), .ZN(n14027) );
  AOI21_X1 U15747 ( .B1(n19228), .B2(n17870), .A(n14027), .ZN(n14028) );
  INV_X1 U15748 ( .A(n14029), .ZN(n14033) );
  INV_X1 U15749 ( .A(n15115), .ZN(n14030) );
  NAND2_X1 U15750 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n22349) );
  NAND2_X1 U15751 ( .A1(n14030), .A2(n22349), .ZN(n14367) );
  NOR2_X1 U15752 ( .A1(n14367), .A2(n14031), .ZN(n14032) );
  AOI21_X1 U15753 ( .B1(n19318), .B2(n14033), .A(n14032), .ZN(n14035) );
  INV_X1 U15754 ( .A(n22349), .ZN(n22359) );
  INV_X1 U15755 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n22348) );
  INV_X1 U15756 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n22366) );
  NAND2_X1 U15757 ( .A1(n22348), .A2(n22366), .ZN(n22350) );
  NAND2_X2 U15758 ( .A1(n22354), .A2(n17980), .ZN(n17977) );
  OAI21_X1 U15759 ( .B1(n22354), .B2(n22350), .A(n17977), .ZN(n22356) );
  INV_X1 U15760 ( .A(n22356), .ZN(n14051) );
  NOR2_X1 U15761 ( .A1(n22359), .A2(n14051), .ZN(n15395) );
  NAND3_X1 U15762 ( .A1(n15038), .A2(n15395), .A3(n14172), .ZN(n14034) );
  NAND2_X1 U15763 ( .A1(n14035), .A2(n14034), .ZN(n14037) );
  NOR2_X1 U15764 ( .A1(n14367), .A2(n20206), .ZN(n14036) );
  MUX2_X1 U15765 ( .A(n14037), .B(n14036), .S(n15109), .Z(n14038) );
  INV_X1 U15766 ( .A(n14040), .ZN(n14058) );
  NAND2_X1 U15767 ( .A1(n15038), .A2(n19017), .ZN(n14057) );
  AND2_X1 U15768 ( .A1(n14043), .A2(n20206), .ZN(n14044) );
  OR2_X1 U15769 ( .A1(n14042), .A2(n14044), .ZN(n14050) );
  NAND2_X1 U15770 ( .A1(n14045), .A2(n15390), .ZN(n14169) );
  OR2_X1 U15771 ( .A1(n14046), .A2(n11954), .ZN(n14167) );
  NAND2_X1 U15772 ( .A1(n14047), .A2(n15109), .ZN(n14164) );
  OAI211_X1 U15773 ( .C1(n20294), .C2(n12011), .A(n14164), .B(n20206), .ZN(
        n14048) );
  AND4_X1 U15774 ( .A1(n14169), .A2(n12030), .A3(n14167), .A4(n14048), .ZN(
        n14049) );
  NAND2_X1 U15775 ( .A1(n14050), .A2(n14049), .ZN(n14165) );
  NOR2_X1 U15776 ( .A1(n14367), .A2(n14051), .ZN(n14052) );
  AND2_X1 U15777 ( .A1(n14053), .A2(n14052), .ZN(n14054) );
  NOR2_X1 U15778 ( .A1(n14165), .A2(n14054), .ZN(n15057) );
  NAND2_X1 U15779 ( .A1(n14055), .A2(n15057), .ZN(n14056) );
  OR2_X1 U15780 ( .A1(n14061), .A2(n19302), .ZN(n14211) );
  INV_X1 U15781 ( .A(n15059), .ZN(n15098) );
  OR2_X1 U15782 ( .A1(n14042), .A2(n15122), .ZN(n15112) );
  NAND2_X1 U15783 ( .A1(n15112), .A2(n19017), .ZN(n14062) );
  NAND2_X1 U15784 ( .A1(n15098), .A2(n14062), .ZN(n14063) );
  INV_X1 U15785 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n14069) );
  NOR2_X1 U15786 ( .A1(n12006), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U15787 ( .A1(n15828), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14068) );
  NAND2_X1 U15788 ( .A1(n14136), .A2(n14066), .ZN(n14067) );
  OAI211_X1 U15789 ( .C1(n15830), .C2(n14069), .A(n14068), .B(n14067), .ZN(
        n14972) );
  INV_X1 U15790 ( .A(n14070), .ZN(n14074) );
  AND2_X1 U15791 ( .A1(n12006), .A2(n19975), .ZN(n14080) );
  NAND2_X1 U15792 ( .A1(n14071), .A2(n14080), .ZN(n14072) );
  OAI21_X1 U15793 ( .B1(n19975), .B2(n19985), .A(n14072), .ZN(n14073) );
  AOI21_X1 U15794 ( .B1(n14074), .B2(n14470), .A(n14073), .ZN(n14501) );
  AND2_X1 U15795 ( .A1(n19987), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14075) );
  AOI21_X1 U15796 ( .B1(n14136), .B2(n14077), .A(n14076), .ZN(n14079) );
  NAND2_X1 U15797 ( .A1(n14078), .A2(n15806), .ZN(n14090) );
  INV_X1 U15798 ( .A(n14080), .ZN(n14083) );
  INV_X1 U15799 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n14081) );
  NAND2_X1 U15800 ( .A1(n19975), .A2(n14081), .ZN(n14082) );
  AOI22_X1 U15801 ( .A1(n19017), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n14083), .B2(n14082), .ZN(n14084) );
  OAI21_X1 U15802 ( .B1(n15830), .B2(n14423), .A(n14084), .ZN(n14498) );
  AOI22_X1 U15803 ( .A1(n14085), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14086) );
  OAI21_X1 U15804 ( .B1(n15830), .B2(n17053), .A(n14086), .ZN(n14087) );
  NAND2_X1 U15805 ( .A1(n14136), .A2(n14089), .ZN(n14091) );
  OAI211_X1 U15806 ( .C1(n19975), .C2(n19871), .A(n14091), .B(n14090), .ZN(
        n14093) );
  AOI22_X1 U15807 ( .A1(n15828), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14094) );
  OAI21_X1 U15808 ( .B1(n15830), .B2(n12060), .A(n14094), .ZN(n14760) );
  NAND2_X1 U15809 ( .A1(n15828), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n14098) );
  NAND2_X1 U15810 ( .A1(n15806), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14097) );
  OAI211_X1 U15811 ( .C1(n19898), .C2(n19975), .A(n14098), .B(n14097), .ZN(
        n14099) );
  INV_X1 U15812 ( .A(n14099), .ZN(n14102) );
  NAND2_X1 U15813 ( .A1(n14136), .A2(n14100), .ZN(n14101) );
  OAI211_X1 U15814 ( .C1(n15830), .C2(n15268), .A(n14102), .B(n14101), .ZN(
        n14889) );
  AOI22_X1 U15815 ( .A1(n15828), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14105) );
  NAND2_X1 U15816 ( .A1(n14136), .A2(n14103), .ZN(n14104) );
  OAI211_X1 U15817 ( .C1(n15830), .C2(n14106), .A(n14105), .B(n14104), .ZN(
        n15517) );
  NAND2_X1 U15818 ( .A1(n14136), .A2(n14107), .ZN(n14108) );
  INV_X1 U15819 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19046) );
  AOI22_X1 U15820 ( .A1(n15828), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14110) );
  OAI21_X1 U15821 ( .B1(n15830), .B2(n19046), .A(n14110), .ZN(n14750) );
  NAND2_X1 U15822 ( .A1(n14749), .A2(n14750), .ZN(n14112) );
  NAND2_X1 U15823 ( .A1(n14136), .A2(n15859), .ZN(n14111) );
  AOI22_X1 U15824 ( .A1(n15828), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14113) );
  OAI21_X1 U15825 ( .B1(n15830), .B2(n17044), .A(n14113), .ZN(n14752) );
  AOI22_X1 U15826 ( .A1(n15828), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14115) );
  NAND2_X1 U15827 ( .A1(n14136), .A2(n14906), .ZN(n14114) );
  OAI211_X1 U15828 ( .C1(n15830), .C2(n14116), .A(n14115), .B(n14114), .ZN(
        n14756) );
  AOI22_X1 U15829 ( .A1(n15828), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n15806), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U15830 ( .A1(n14136), .A2(n14117), .ZN(n14118) );
  OAI211_X1 U15831 ( .C1(n15830), .C2(n17961), .A(n14119), .B(n14118), .ZN(
        n15457) );
  NAND2_X1 U15832 ( .A1(n15805), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U15833 ( .A1(n15828), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14121) );
  NAND2_X1 U15834 ( .A1(n14136), .A2(n14984), .ZN(n14120) );
  NAND2_X1 U15835 ( .A1(n15805), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U15836 ( .A1(n15828), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U15837 ( .A1(n14136), .A2(n14123), .ZN(n14124) );
  AOI22_X1 U15838 ( .A1(n15828), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U15839 ( .A1(n14136), .A2(n15024), .ZN(n14127) );
  OAI211_X1 U15840 ( .C1(n15830), .C2(n17963), .A(n14128), .B(n14127), .ZN(
        n15445) );
  NAND2_X1 U15841 ( .A1(n15446), .A2(n15445), .ZN(n14773) );
  NAND2_X1 U15842 ( .A1(n15805), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U15843 ( .A1(n15828), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14130) );
  NAND2_X1 U15844 ( .A1(n14136), .A2(n15201), .ZN(n14129) );
  NAND2_X1 U15845 ( .A1(n15805), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n14134) );
  AOI22_X1 U15846 ( .A1(n15828), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14133) );
  NAND2_X1 U15847 ( .A1(n14136), .A2(n15334), .ZN(n14132) );
  AOI22_X1 U15848 ( .A1(n15828), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14138) );
  NAND2_X1 U15849 ( .A1(n14136), .A2(n15365), .ZN(n14137) );
  OAI211_X1 U15850 ( .C1(n15830), .C2(n17965), .A(n14138), .B(n14137), .ZN(
        n15001) );
  AOI22_X1 U15851 ( .A1(n15828), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14139) );
  OAI21_X1 U15852 ( .B1(n15830), .B2(n17966), .A(n14139), .ZN(n16806) );
  NAND2_X1 U15853 ( .A1(n15805), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n14141) );
  AOI22_X1 U15854 ( .A1(n15828), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14140) );
  NAND2_X1 U15855 ( .A1(n15805), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n14143) );
  AOI22_X1 U15856 ( .A1(n15828), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14142) );
  NAND2_X1 U15857 ( .A1(n15805), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U15858 ( .A1(n15828), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U15859 ( .A1(n15828), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14146) );
  OAI21_X1 U15860 ( .B1(n15830), .B2(n17970), .A(n14146), .ZN(n16643) );
  NAND2_X1 U15861 ( .A1(n16644), .A2(n16643), .ZN(n16626) );
  NAND2_X1 U15862 ( .A1(n15805), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14148) );
  AOI22_X1 U15863 ( .A1(n15828), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14147) );
  AND2_X1 U15864 ( .A1(n14148), .A2(n14147), .ZN(n16627) );
  NAND2_X1 U15865 ( .A1(n15805), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U15866 ( .A1(n15828), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U15867 ( .A1(n15828), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14151) );
  OAI21_X1 U15868 ( .B1(n15830), .B2(n17971), .A(n14151), .ZN(n16779) );
  AOI22_X1 U15869 ( .A1(n15828), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14152) );
  OAI21_X1 U15870 ( .B1(n15830), .B2(n16862), .A(n14152), .ZN(n16769) );
  NAND2_X1 U15871 ( .A1(n15805), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n14154) );
  AOI22_X1 U15872 ( .A1(n15828), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14153) );
  AND2_X1 U15873 ( .A1(n14154), .A2(n14153), .ZN(n16763) );
  NAND2_X1 U15874 ( .A1(n15805), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U15875 ( .A1(n15828), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14155) );
  AND2_X1 U15876 ( .A1(n14156), .A2(n14155), .ZN(n16757) );
  AOI22_X1 U15877 ( .A1(n15828), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14157) );
  OAI21_X1 U15878 ( .B1(n15830), .B2(n19207), .A(n14157), .ZN(n16748) );
  AOI22_X1 U15879 ( .A1(n15828), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14158) );
  OAI21_X1 U15880 ( .B1(n15830), .B2(n14159), .A(n14158), .ZN(n14161) );
  NOR2_X1 U15881 ( .A1(n14160), .A2(n14161), .ZN(n14162) );
  OR2_X1 U15882 ( .A1(n15808), .A2(n14162), .ZN(n19225) );
  INV_X1 U15883 ( .A(n17098), .ZN(n14191) );
  INV_X1 U15884 ( .A(n14212), .ZN(n14163) );
  NAND2_X1 U15885 ( .A1(n14163), .A2(n19294), .ZN(n19275) );
  INV_X1 U15886 ( .A(n19275), .ZN(n17378) );
  NAND2_X1 U15887 ( .A1(n14212), .A2(n15101), .ZN(n17352) );
  OR2_X1 U15888 ( .A1(n14166), .A2(n12030), .ZN(n14181) );
  NAND3_X1 U15889 ( .A1(n14167), .A2(n12006), .A3(n14043), .ZN(n14168) );
  NAND2_X1 U15890 ( .A1(n14168), .A2(n19017), .ZN(n15068) );
  NAND2_X1 U15891 ( .A1(n15068), .A2(n14169), .ZN(n14179) );
  INV_X1 U15892 ( .A(n14171), .ZN(n14365) );
  NAND2_X1 U15893 ( .A1(n12030), .A2(n20125), .ZN(n14173) );
  NAND2_X1 U15894 ( .A1(n14175), .A2(n14174), .ZN(n14508) );
  NAND3_X1 U15895 ( .A1(n14170), .A2(n14176), .A3(n14508), .ZN(n14177) );
  AOI21_X1 U15896 ( .B1(n14179), .B2(n14178), .A(n14177), .ZN(n14180) );
  AND2_X1 U15897 ( .A1(n14181), .A2(n14180), .ZN(n15075) );
  NAND2_X1 U15898 ( .A1(n15075), .A2(n15061), .ZN(n14182) );
  NAND2_X1 U15899 ( .A1(n14212), .A2(n14182), .ZN(n17326) );
  NAND2_X1 U15900 ( .A1(n17352), .A2(n17326), .ZN(n19279) );
  INV_X1 U15901 ( .A(n17295), .ZN(n14190) );
  OR2_X1 U15902 ( .A1(n14183), .A2(n16881), .ZN(n17132) );
  NAND3_X1 U15903 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n17341) );
  NOR2_X1 U15904 ( .A1(n17342), .A2(n17341), .ZN(n17323) );
  INV_X1 U15905 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19290) );
  NOR2_X1 U15906 ( .A1(n19307), .A2(n19290), .ZN(n19289) );
  NAND2_X1 U15907 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17379) );
  INV_X1 U15908 ( .A(n17379), .ZN(n17358) );
  NOR2_X1 U15909 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17358), .ZN(
        n15266) );
  INV_X1 U15910 ( .A(n15266), .ZN(n17354) );
  AND3_X1 U15911 ( .A1(n17323), .A2(n19289), .A3(n17354), .ZN(n14192) );
  OAI21_X1 U15912 ( .B1(n17352), .B2(n14192), .A(n19275), .ZN(n17169) );
  INV_X1 U15913 ( .A(n17323), .ZN(n14184) );
  NAND2_X1 U15914 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n17358), .ZN(
        n17353) );
  NOR2_X1 U15915 ( .A1(n14184), .A2(n17353), .ZN(n17327) );
  NAND2_X1 U15916 ( .A1(n19289), .A2(n17327), .ZN(n17170) );
  INV_X1 U15917 ( .A(n17170), .ZN(n14193) );
  NOR2_X1 U15918 ( .A1(n17326), .A2(n14193), .ZN(n14185) );
  INV_X1 U15919 ( .A(n17247), .ZN(n14189) );
  NOR2_X1 U15920 ( .A1(n14187), .A2(n14186), .ZN(n14188) );
  NAND2_X1 U15921 ( .A1(n14189), .A2(n14188), .ZN(n17210) );
  NOR3_X1 U15922 ( .A1(n17317), .A2(n17157), .A3(n17210), .ZN(n17156) );
  AOI21_X1 U15923 ( .B1(n17156), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n17295), .ZN(n17150) );
  AOI211_X1 U15924 ( .C1(n19279), .C2(n17132), .A(n12345), .B(n17150), .ZN(
        n17125) );
  NOR2_X1 U15925 ( .A1(n17125), .A2(n17295), .ZN(n17115) );
  AOI21_X1 U15926 ( .B1(n14191), .B2(n14190), .A(n17115), .ZN(n17092) );
  INV_X1 U15927 ( .A(n17092), .ZN(n15870) );
  NAND2_X1 U15928 ( .A1(n15870), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14201) );
  NAND2_X1 U15929 ( .A1(n17328), .A2(n14192), .ZN(n14195) );
  NAND2_X1 U15930 ( .A1(n17361), .A2(n14193), .ZN(n14194) );
  NAND2_X1 U15931 ( .A1(n14195), .A2(n14194), .ZN(n17285) );
  INV_X1 U15932 ( .A(n17210), .ZN(n17167) );
  NOR2_X1 U15933 ( .A1(n17157), .A2(n17158), .ZN(n14196) );
  NAND2_X1 U15934 ( .A1(n17238), .A2(n14196), .ZN(n17148) );
  NOR2_X1 U15935 ( .A1(n17132), .A2(n17148), .ZN(n17124) );
  NAND2_X1 U15936 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17124), .ZN(
        n17099) );
  INV_X1 U15937 ( .A(n17099), .ZN(n17110) );
  NAND2_X1 U15938 ( .A1(n17098), .A2(n17110), .ZN(n17079) );
  INV_X1 U15939 ( .A(n17079), .ZN(n17088) );
  XNOR2_X1 U15940 ( .A(n14197), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14199) );
  AOI21_X1 U15941 ( .B1(n17088), .B2(n14199), .A(n14198), .ZN(n14200) );
  OAI211_X1 U15942 ( .C1(n17371), .C2(n19225), .A(n14201), .B(n14200), .ZN(
        n14209) );
  NAND2_X1 U15943 ( .A1(n15072), .A2(n15109), .ZN(n14204) );
  INV_X1 U15944 ( .A(n14202), .ZN(n14203) );
  NAND2_X1 U15945 ( .A1(n14204), .A2(n14203), .ZN(n14205) );
  NOR2_X1 U15946 ( .A1(n14209), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U15947 ( .A1(n14696), .A2(n14712), .ZN(n14218) );
  NAND2_X1 U15948 ( .A1(n15908), .A2(n14817), .ZN(n14214) );
  NOR2_X1 U15949 ( .A1(n14215), .A2(n14214), .ZN(n14217) );
  NAND2_X1 U15950 ( .A1(n14217), .A2(n14216), .ZN(n14623) );
  NAND2_X1 U15951 ( .A1(n14218), .A2(n14623), .ZN(n14220) );
  AND2_X1 U15952 ( .A1(n14222), .A2(n15163), .ZN(n14219) );
  NAND2_X2 U15953 ( .A1(n14809), .A2(n14886), .ZN(n14316) );
  NAND2_X2 U15954 ( .A1(n14316), .A2(n14226), .ZN(n15918) );
  INV_X1 U15955 ( .A(n14222), .ZN(n15917) );
  OAI22_X1 U15956 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n15917), .B2(P1_EBX_REG_30__SCAN_IN), .ZN(n15916) );
  OR2_X1 U15957 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14224) );
  MUX2_X1 U15958 ( .A(n14321), .B(n14226), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n14223) );
  INV_X1 U15959 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14225) );
  OR2_X1 U15960 ( .A1(n14316), .A2(n14225), .ZN(n14228) );
  NAND2_X1 U15961 ( .A1(n14327), .A2(n14225), .ZN(n14227) );
  NAND2_X1 U15962 ( .A1(n14228), .A2(n14227), .ZN(n14551) );
  XNOR2_X1 U15963 ( .A(n14229), .B(n14551), .ZN(n14573) );
  MUX2_X1 U15964 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n14231) );
  OR2_X1 U15965 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14230) );
  AND2_X1 U15966 ( .A1(n14231), .A2(n14230), .ZN(n14667) );
  NAND2_X1 U15967 ( .A1(n14668), .A2(n14667), .ZN(n14740) );
  OR2_X1 U15968 ( .A1(n14326), .A2(P1_EBX_REG_3__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U15969 ( .A1(n14316), .A2(n21992), .ZN(n14233) );
  INV_X1 U15970 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n17620) );
  NAND2_X1 U15971 ( .A1(n14222), .A2(n17620), .ZN(n14232) );
  NAND3_X1 U15972 ( .A1(n14233), .A2(n14313), .A3(n14232), .ZN(n14234) );
  AND2_X1 U15973 ( .A1(n14235), .A2(n14234), .ZN(n14741) );
  MUX2_X1 U15974 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n14236) );
  OAI21_X1 U15975 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15918), .A(
        n14236), .ZN(n20571) );
  OR2_X1 U15976 ( .A1(n14326), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n14242) );
  NAND2_X1 U15977 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14237) );
  NAND2_X1 U15978 ( .A1(n14316), .A2(n14237), .ZN(n14240) );
  INV_X1 U15979 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U15980 ( .A1(n14222), .A2(n14238), .ZN(n14239) );
  NAND2_X1 U15981 ( .A1(n14240), .A2(n14239), .ZN(n14241) );
  NAND2_X1 U15982 ( .A1(n14242), .A2(n14241), .ZN(n15161) );
  AND2_X2 U15983 ( .A1(n20569), .A2(n15161), .ZN(n15160) );
  MUX2_X1 U15984 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n14243) );
  OAI21_X1 U15985 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15918), .A(
        n14243), .ZN(n20552) );
  INV_X1 U15986 ( .A(n20552), .ZN(n14244) );
  OR2_X1 U15987 ( .A1(n14326), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n14250) );
  NAND2_X1 U15988 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14245) );
  NAND2_X1 U15989 ( .A1(n14316), .A2(n14245), .ZN(n14248) );
  INV_X1 U15990 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U15991 ( .A1(n14222), .A2(n14246), .ZN(n14247) );
  NAND2_X1 U15992 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  MUX2_X1 U15993 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n14251) );
  OAI21_X1 U15994 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15918), .A(
        n14251), .ZN(n15305) );
  OR2_X1 U15995 ( .A1(n14326), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n14256) );
  NAND2_X1 U15996 ( .A1(n14316), .A2(n22038), .ZN(n14254) );
  INV_X1 U15997 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14252) );
  NAND3_X1 U15998 ( .A1(n14254), .A2(n14313), .A3(n14253), .ZN(n14255) );
  NAND2_X1 U15999 ( .A1(n14256), .A2(n14255), .ZN(n15356) );
  MUX2_X1 U16000 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14257) );
  OAI21_X1 U16001 ( .B1(n15918), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n14257), .ZN(n14258) );
  INV_X1 U16002 ( .A(n14258), .ZN(n20559) );
  OR2_X1 U16003 ( .A1(n14326), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n14264) );
  NAND2_X1 U16004 ( .A1(n14316), .A2(n14259), .ZN(n14262) );
  INV_X1 U16005 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U16006 ( .A1(n14222), .A2(n14260), .ZN(n14261) );
  NAND3_X1 U16007 ( .A1(n14262), .A2(n14313), .A3(n14261), .ZN(n14263) );
  INV_X1 U16008 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n20558) );
  NAND2_X1 U16009 ( .A1(n14222), .A2(n20558), .ZN(n14266) );
  NAND2_X1 U16010 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14265) );
  NAND3_X1 U16011 ( .A1(n14266), .A2(n14316), .A3(n14265), .ZN(n14267) );
  OAI21_X1 U16012 ( .B1(n14321), .B2(P1_EBX_REG_12__SCAN_IN), .A(n14267), .ZN(
        n20556) );
  OR2_X1 U16013 ( .A1(n14326), .A2(P1_EBX_REG_13__SCAN_IN), .ZN(n14272) );
  NAND2_X1 U16014 ( .A1(n14316), .A2(n14268), .ZN(n14270) );
  INV_X1 U16015 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n17789) );
  NAND2_X1 U16016 ( .A1(n14222), .A2(n17789), .ZN(n14269) );
  NAND3_X1 U16017 ( .A1(n14270), .A2(n14226), .A3(n14269), .ZN(n14271) );
  NAND2_X1 U16018 ( .A1(n14272), .A2(n14271), .ZN(n16086) );
  NAND2_X1 U16019 ( .A1(n20554), .A2(n16086), .ZN(n16088) );
  INV_X1 U16020 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n17794) );
  NAND2_X1 U16021 ( .A1(n14222), .A2(n17794), .ZN(n14274) );
  NAND2_X1 U16022 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14273) );
  NAND3_X1 U16023 ( .A1(n14274), .A2(n14316), .A3(n14273), .ZN(n14275) );
  OAI21_X1 U16024 ( .B1(n14321), .B2(P1_EBX_REG_14__SCAN_IN), .A(n14275), .ZN(
        n15620) );
  OR2_X1 U16025 ( .A1(n14326), .A2(P1_EBX_REG_15__SCAN_IN), .ZN(n14279) );
  INV_X1 U16026 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16347) );
  NAND2_X1 U16027 ( .A1(n14316), .A2(n16347), .ZN(n14277) );
  INV_X1 U16028 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n17481) );
  NAND3_X1 U16029 ( .A1(n14277), .A2(n14226), .A3(n14276), .ZN(n14278) );
  MUX2_X1 U16030 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n14280) );
  OAI21_X1 U16031 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15918), .A(
        n14280), .ZN(n16133) );
  OR2_X1 U16032 ( .A1(n14326), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U16033 ( .A1(n14316), .A2(n14281), .ZN(n14283) );
  INV_X1 U16034 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n22248) );
  NAND2_X1 U16035 ( .A1(n14222), .A2(n22248), .ZN(n14282) );
  NAND3_X1 U16036 ( .A1(n14283), .A2(n14313), .A3(n14282), .ZN(n14284) );
  MUX2_X1 U16037 ( .A(n14321), .B(n14226), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14287) );
  OR2_X1 U16038 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14286) );
  NAND2_X1 U16039 ( .A1(n14287), .A2(n14286), .ZN(n16072) );
  NOR2_X1 U16040 ( .A1(n20566), .A2(n16072), .ZN(n14288) );
  OR2_X1 U16041 ( .A1(n14326), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14292) );
  NAND2_X1 U16042 ( .A1(n14316), .A2(n16529), .ZN(n14290) );
  INV_X1 U16043 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n17782) );
  NAND2_X1 U16044 ( .A1(n14222), .A2(n17782), .ZN(n14289) );
  NAND3_X1 U16045 ( .A1(n14290), .A2(n14226), .A3(n14289), .ZN(n14291) );
  NAND2_X1 U16046 ( .A1(n14292), .A2(n14291), .ZN(n16125) );
  MUX2_X1 U16047 ( .A(n14321), .B(n14226), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14293) );
  OAI21_X1 U16048 ( .B1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15918), .A(
        n14293), .ZN(n16060) );
  OR2_X2 U16049 ( .A1(n11185), .A2(n16060), .ZN(n16062) );
  OR2_X1 U16050 ( .A1(n14326), .A2(P1_EBX_REG_21__SCAN_IN), .ZN(n14297) );
  NAND2_X1 U16051 ( .A1(n14316), .A2(n16510), .ZN(n14295) );
  INV_X1 U16052 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n17638) );
  NAND2_X1 U16053 ( .A1(n14222), .A2(n17638), .ZN(n14294) );
  NAND3_X1 U16054 ( .A1(n14295), .A2(n14226), .A3(n14294), .ZN(n14296) );
  MUX2_X1 U16055 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14299) );
  OR2_X1 U16056 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14298) );
  AND2_X1 U16057 ( .A1(n14299), .A2(n14298), .ZN(n16037) );
  OR2_X1 U16058 ( .A1(n14326), .A2(P1_EBX_REG_23__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U16059 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14300) );
  NAND2_X1 U16060 ( .A1(n14316), .A2(n14300), .ZN(n14302) );
  INV_X1 U16061 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n17598) );
  NAND2_X1 U16062 ( .A1(n14222), .A2(n17598), .ZN(n14301) );
  NAND2_X1 U16063 ( .A1(n14302), .A2(n14301), .ZN(n14303) );
  AND2_X1 U16064 ( .A1(n14304), .A2(n14303), .ZN(n16005) );
  MUX2_X1 U16065 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14306) );
  OR2_X1 U16066 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14305) );
  NAND2_X1 U16067 ( .A1(n14306), .A2(n14305), .ZN(n16006) );
  NOR2_X1 U16068 ( .A1(n16005), .A2(n16006), .ZN(n14307) );
  OR2_X1 U16069 ( .A1(n14326), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n14312) );
  NAND2_X1 U16070 ( .A1(n14316), .A2(n16471), .ZN(n14310) );
  INV_X1 U16071 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14308) );
  NAND2_X1 U16072 ( .A1(n14222), .A2(n14308), .ZN(n14309) );
  NAND3_X1 U16073 ( .A1(n14310), .A2(n14313), .A3(n14309), .ZN(n14311) );
  AND2_X1 U16074 ( .A1(n14312), .A2(n14311), .ZN(n16002) );
  MUX2_X1 U16075 ( .A(n14321), .B(n14226), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14314) );
  OAI21_X1 U16076 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15918), .A(
        n14314), .ZN(n15981) );
  OR2_X2 U16077 ( .A1(n11189), .A2(n15981), .ZN(n15982) );
  OR2_X1 U16078 ( .A1(n14326), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U16079 ( .A1(n14226), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14315) );
  NAND2_X1 U16080 ( .A1(n14316), .A2(n14315), .ZN(n14318) );
  INV_X1 U16081 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n17596) );
  NAND2_X1 U16082 ( .A1(n14222), .A2(n17596), .ZN(n14317) );
  NAND2_X1 U16083 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  MUX2_X1 U16084 ( .A(n14321), .B(n14313), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14323) );
  OR2_X1 U16085 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14322) );
  AND2_X1 U16086 ( .A1(n14323), .A2(n14322), .ZN(n15956) );
  OR2_X1 U16087 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14325) );
  INV_X1 U16088 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n16112) );
  NAND2_X1 U16089 ( .A1(n14222), .A2(n16112), .ZN(n14324) );
  NAND2_X1 U16090 ( .A1(n14325), .A2(n14324), .ZN(n14328) );
  OAI22_X1 U16091 ( .A1(n14328), .A2(n14327), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14326), .ZN(n15944) );
  NAND2_X1 U16092 ( .A1(n11220), .A2(n14327), .ZN(n14329) );
  INV_X1 U16093 ( .A(n15945), .ZN(n15955) );
  AOI22_X1 U16094 ( .A1(n14329), .A2(n14328), .B1(n15955), .B2(n14313), .ZN(
        n14330) );
  XOR2_X1 U16095 ( .A(n15916), .B(n14330), .Z(n15933) );
  INV_X1 U16096 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n17640) );
  OR2_X1 U16097 ( .A1(n20574), .A2(n17640), .ZN(n14331) );
  OAI21_X1 U16098 ( .B1(n15933), .B2(n16143), .A(n14331), .ZN(n14332) );
  INV_X1 U16099 ( .A(n14332), .ZN(n14333) );
  NOR2_X1 U16100 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14336) );
  NOR4_X1 U16101 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14335) );
  NAND4_X1 U16102 ( .A1(n14336), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14335), .ZN(n14358) );
  NOR4_X1 U16103 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n14340) );
  NOR4_X1 U16104 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n14339) );
  NOR4_X1 U16105 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n14338) );
  NOR4_X1 U16106 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n14337) );
  AND4_X1 U16107 ( .A1(n14340), .A2(n14339), .A3(n14338), .A4(n14337), .ZN(
        n14345) );
  NOR4_X1 U16108 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n14343) );
  NOR4_X1 U16109 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n14342) );
  NOR4_X1 U16110 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n14341) );
  INV_X1 U16111 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20482) );
  AND4_X1 U16112 ( .A1(n14343), .A2(n14342), .A3(n14341), .A4(n20482), .ZN(
        n14344) );
  NAND2_X1 U16113 ( .A1(n14345), .A2(n14344), .ZN(n14346) );
  INV_X1 U16114 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n22851) );
  NOR3_X1 U16115 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n22851), .ZN(n14348) );
  NOR4_X1 U16116 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14347) );
  NAND4_X1 U16117 ( .A1(n15823), .A2(P1_W_R_N_REG_SCAN_IN), .A3(n14348), .A4(
        n14347), .ZN(U214) );
  NOR4_X1 U16118 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14352) );
  NOR4_X1 U16119 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14351) );
  NOR4_X1 U16120 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14350) );
  NOR4_X1 U16121 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14349) );
  NAND4_X1 U16122 ( .A1(n14352), .A2(n14351), .A3(n14350), .A4(n14349), .ZN(
        n14357) );
  NOR4_X1 U16123 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14355) );
  NOR4_X1 U16124 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14354) );
  NOR4_X1 U16125 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14353) );
  INV_X1 U16126 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17953) );
  NAND4_X1 U16127 ( .A1(n14355), .A2(n14354), .A3(n14353), .A4(n17953), .ZN(
        n14356) );
  OAI21_X1 U16128 ( .B1(n14357), .B2(n14356), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14371) );
  NOR2_X1 U16129 ( .A1(n15601), .A2(n14358), .ZN(n20639) );
  NAND2_X1 U16130 ( .A1(n20639), .A2(U214), .ZN(U212) );
  NAND2_X1 U16131 ( .A1(n14042), .A2(n19014), .ZN(n14359) );
  INV_X1 U16132 ( .A(n15591), .ZN(n19030) );
  INV_X1 U16133 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14363) );
  INV_X1 U16134 ( .A(n17840), .ZN(n14362) );
  NAND2_X1 U16135 ( .A1(n17416), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n14360) );
  OR2_X1 U16136 ( .A1(n14361), .A2(n14360), .ZN(n14368) );
  OAI211_X1 U16137 ( .C1(n19030), .C2(n14363), .A(n14362), .B(n15399), .ZN(
        P2_U2814) );
  OAI21_X1 U16138 ( .B1(n17840), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19012), 
        .ZN(n14364) );
  OAI21_X1 U16139 ( .B1(n14365), .B2(n19012), .A(n14364), .ZN(P2_U3612) );
  INV_X1 U16140 ( .A(n15399), .ZN(n14366) );
  INV_X1 U16141 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14373) );
  INV_X1 U16142 ( .A(n14367), .ZN(n14370) );
  NOR2_X1 U16143 ( .A1(n14368), .A2(n15109), .ZN(n14369) );
  NAND2_X1 U16144 ( .A1(n14370), .A2(n14369), .ZN(n14458) );
  AOI22_X1 U16145 ( .A1(n15596), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15601), .ZN(n15047) );
  NOR2_X1 U16146 ( .A1(n14458), .A2(n15047), .ZN(n14439) );
  AOI21_X1 U16147 ( .B1(n14463), .B2(P2_EAX_REG_1__SCAN_IN), .A(n14439), .ZN(
        n14372) );
  OAI21_X1 U16148 ( .B1(n14388), .B2(n14373), .A(n14372), .ZN(P2_U2968) );
  INV_X1 U16149 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14375) );
  OAI22_X1 U16150 ( .A1(n15601), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15596), .ZN(n20024) );
  NOR2_X1 U16151 ( .A1(n14458), .A2(n20024), .ZN(n14428) );
  AOI21_X1 U16152 ( .B1(n14463), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14428), .ZN(
        n14374) );
  OAI21_X1 U16153 ( .B1(n14388), .B2(n14375), .A(n14374), .ZN(P2_U2973) );
  INV_X1 U16154 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14377) );
  AOI22_X1 U16155 ( .A1(n15596), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15601), .ZN(n16771) );
  NOR2_X1 U16156 ( .A1(n14458), .A2(n16771), .ZN(n14446) );
  AOI21_X1 U16157 ( .B1(n14463), .B2(P2_EAX_REG_8__SCAN_IN), .A(n14446), .ZN(
        n14376) );
  OAI21_X1 U16158 ( .B1(n14388), .B2(n14377), .A(n14376), .ZN(P2_U2975) );
  INV_X1 U16159 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14379) );
  AOI22_X1 U16160 ( .A1(n15596), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15601), .ZN(n20072) );
  NOR2_X1 U16161 ( .A1(n14458), .A2(n20072), .ZN(n14455) );
  AOI21_X1 U16162 ( .B1(n14463), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14455), .ZN(
        n14378) );
  OAI21_X1 U16163 ( .B1(n14388), .B2(n14379), .A(n14378), .ZN(P2_U2972) );
  INV_X1 U16164 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14381) );
  AOI22_X1 U16165 ( .A1(n15596), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15601), .ZN(n20292) );
  NOR2_X1 U16166 ( .A1(n14458), .A2(n20292), .ZN(n14431) );
  AOI21_X1 U16167 ( .B1(n14463), .B2(P2_EAX_REG_0__SCAN_IN), .A(n14431), .ZN(
        n14380) );
  OAI21_X1 U16168 ( .B1(n14388), .B2(n14381), .A(n14380), .ZN(P2_U2967) );
  INV_X1 U16169 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14383) );
  AOI22_X1 U16170 ( .A1(n15596), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15601), .ZN(n20165) );
  NOR2_X1 U16171 ( .A1(n14458), .A2(n20165), .ZN(n14449) );
  AOI21_X1 U16172 ( .B1(n14463), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14449), .ZN(
        n14382) );
  OAI21_X1 U16173 ( .B1(n14388), .B2(n14383), .A(n14382), .ZN(P2_U2970) );
  INV_X1 U16174 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14385) );
  OAI22_X1 U16175 ( .A1(n15601), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n15596), .ZN(n20124) );
  NOR2_X1 U16176 ( .A1(n14458), .A2(n20124), .ZN(n14443) );
  AOI21_X1 U16177 ( .B1(n14463), .B2(P2_EAX_REG_4__SCAN_IN), .A(n14443), .ZN(
        n14384) );
  OAI21_X1 U16178 ( .B1(n14388), .B2(n14385), .A(n14384), .ZN(P2_U2971) );
  INV_X1 U16179 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14387) );
  AOI22_X1 U16180 ( .A1(n15596), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15601), .ZN(n20205) );
  NOR2_X1 U16181 ( .A1(n14458), .A2(n20205), .ZN(n14434) );
  AOI21_X1 U16182 ( .B1(n14463), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14434), .ZN(
        n14386) );
  OAI21_X1 U16183 ( .B1(n14388), .B2(n14387), .A(n14386), .ZN(P2_U2954) );
  INV_X1 U16184 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U16185 ( .A1(n14442), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14391) );
  INV_X1 U16186 ( .A(n14458), .ZN(n14407) );
  INV_X1 U16187 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20659) );
  OR2_X1 U16188 ( .A1(n15601), .A2(n20659), .ZN(n14390) );
  NAND2_X1 U16189 ( .A1(n15601), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14389) );
  NAND2_X1 U16190 ( .A1(n14390), .A2(n14389), .ZN(n19809) );
  NAND2_X1 U16191 ( .A1(n14407), .A2(n19809), .ZN(n14392) );
  OAI211_X1 U16192 ( .C1(n14599), .C2(n14477), .A(n14391), .B(n14392), .ZN(
        P2_U2964) );
  INV_X1 U16193 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n17942) );
  NAND2_X1 U16194 ( .A1(n14442), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14393) );
  OAI211_X1 U16195 ( .C1(n17942), .C2(n14477), .A(n14393), .B(n14392), .ZN(
        P2_U2979) );
  INV_X1 U16196 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14595) );
  NAND2_X1 U16197 ( .A1(n14442), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14396) );
  INV_X1 U16198 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20655) );
  OR2_X1 U16199 ( .A1(n15601), .A2(n20655), .ZN(n14395) );
  NAND2_X1 U16200 ( .A1(n15601), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14394) );
  NAND2_X1 U16201 ( .A1(n14395), .A2(n14394), .ZN(n19812) );
  NAND2_X1 U16202 ( .A1(n14407), .A2(n19812), .ZN(n14401) );
  OAI211_X1 U16203 ( .C1(n14595), .C2(n14477), .A(n14396), .B(n14401), .ZN(
        P2_U2962) );
  INV_X1 U16204 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14597) );
  NAND2_X1 U16205 ( .A1(n14442), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14397) );
  AOI22_X1 U16206 ( .A1(n15596), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15601), .ZN(n14748) );
  INV_X1 U16207 ( .A(n14748), .ZN(n16750) );
  NAND2_X1 U16208 ( .A1(n14407), .A2(n16750), .ZN(n14461) );
  OAI211_X1 U16209 ( .C1(n14477), .C2(n14597), .A(n14397), .B(n14461), .ZN(
        P2_U2963) );
  INV_X1 U16210 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14607) );
  NAND2_X1 U16211 ( .A1(n14442), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14398) );
  MUX2_X1 U16212 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n15601), .Z(n19806) );
  NAND2_X1 U16213 ( .A1(n14407), .A2(n19806), .ZN(n14399) );
  OAI211_X1 U16214 ( .C1(n14607), .C2(n14477), .A(n14398), .B(n14399), .ZN(
        P2_U2966) );
  INV_X1 U16215 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n17946) );
  NAND2_X1 U16216 ( .A1(n14442), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14400) );
  OAI211_X1 U16217 ( .C1(n17946), .C2(n14477), .A(n14400), .B(n14399), .ZN(
        P2_U2981) );
  INV_X1 U16218 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17938) );
  NAND2_X1 U16219 ( .A1(n14442), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14402) );
  OAI211_X1 U16220 ( .C1(n17938), .C2(n14477), .A(n14402), .B(n14401), .ZN(
        P2_U2977) );
  INV_X1 U16221 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14593) );
  NAND2_X1 U16222 ( .A1(n14442), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14403) );
  MUX2_X1 U16223 ( .A(BUF1_REG_9__SCAN_IN), .B(BUF2_REG_9__SCAN_IN), .S(n15601), .Z(n19815) );
  NAND2_X1 U16224 ( .A1(n14407), .A2(n19815), .ZN(n14404) );
  OAI211_X1 U16225 ( .C1(n14477), .C2(n14593), .A(n14403), .B(n14404), .ZN(
        P2_U2961) );
  INV_X1 U16226 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n17934) );
  NAND2_X1 U16227 ( .A1(n14442), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14405) );
  OAI211_X1 U16228 ( .C1(n17934), .C2(n14477), .A(n14405), .B(n14404), .ZN(
        P2_U2976) );
  INV_X1 U16229 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14601) );
  NAND2_X1 U16230 ( .A1(n14442), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14408) );
  AOI22_X1 U16231 ( .A1(n15596), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15601), .ZN(n16738) );
  INV_X1 U16232 ( .A(n16738), .ZN(n14406) );
  NAND2_X1 U16233 ( .A1(n14407), .A2(n14406), .ZN(n14465) );
  OAI211_X1 U16234 ( .C1(n14477), .C2(n14601), .A(n14408), .B(n14465), .ZN(
        P2_U2965) );
  INV_X1 U16235 ( .A(n14409), .ZN(n14521) );
  NAND2_X1 U16236 ( .A1(n14411), .A2(n14410), .ZN(n14412) );
  OR2_X1 U16237 ( .A1(n14413), .A2(n14412), .ZN(n14415) );
  AND2_X1 U16238 ( .A1(n14415), .A2(n14414), .ZN(n14620) );
  INV_X1 U16239 ( .A(n14620), .ZN(n15907) );
  NOR2_X1 U16240 ( .A1(n14521), .A2(n15907), .ZN(n15913) );
  AND2_X1 U16241 ( .A1(n15913), .A2(n15163), .ZN(n14416) );
  INV_X1 U16242 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n22852) );
  INV_X1 U16243 ( .A(n14549), .ZN(n15912) );
  NAND2_X1 U16244 ( .A1(n22559), .A2(n15308), .ZN(n15898) );
  OAI211_X1 U16245 ( .C1(n14416), .C2(n22852), .A(n15165), .B(n15898), .ZN(
        P1_U2801) );
  INV_X1 U16246 ( .A(n14417), .ZN(n14419) );
  NOR2_X1 U16247 ( .A1(n15582), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14418) );
  NOR2_X1 U16248 ( .A1(n14419), .A2(n14418), .ZN(n19277) );
  OR2_X1 U16249 ( .A1(n14420), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14421) );
  NAND2_X1 U16250 ( .A1(n14422), .A2(n14421), .ZN(n19287) );
  OR2_X1 U16251 ( .A1(n19294), .A2(n14423), .ZN(n19285) );
  OAI21_X1 U16252 ( .B1(n17873), .B2(n19287), .A(n19285), .ZN(n14424) );
  AOI21_X1 U16253 ( .B1(n17871), .B2(n19277), .A(n14424), .ZN(n14427) );
  OAI21_X1 U16254 ( .B1(n17057), .B2(n14425), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14426) );
  OAI211_X1 U16255 ( .C1(n17852), .C2(n15076), .A(n14427), .B(n14426), .ZN(
        P2_U3014) );
  INV_X1 U16256 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14430) );
  AOI21_X1 U16257 ( .B1(n14463), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14428), .ZN(
        n14429) );
  OAI21_X1 U16258 ( .B1(n14388), .B2(n14430), .A(n14429), .ZN(P2_U2958) );
  INV_X1 U16259 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14433) );
  AOI21_X1 U16260 ( .B1(n14463), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14431), .ZN(
        n14432) );
  OAI21_X1 U16261 ( .B1(n14467), .B2(n14433), .A(n14432), .ZN(P2_U2952) );
  INV_X1 U16262 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14436) );
  AOI21_X1 U16263 ( .B1(n14463), .B2(P2_EAX_REG_2__SCAN_IN), .A(n14434), .ZN(
        n14435) );
  OAI21_X1 U16264 ( .B1(n14467), .B2(n14436), .A(n14435), .ZN(P2_U2969) );
  INV_X1 U16265 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14438) );
  AOI22_X1 U16266 ( .A1(n15596), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15601), .ZN(n19818) );
  NOR2_X1 U16267 ( .A1(n14458), .A2(n19818), .ZN(n14452) );
  AOI21_X1 U16268 ( .B1(n14463), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14452), .ZN(
        n14437) );
  OAI21_X1 U16269 ( .B1(n14467), .B2(n14438), .A(n14437), .ZN(P2_U2974) );
  INV_X1 U16270 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n14441) );
  AOI21_X1 U16271 ( .B1(n14463), .B2(P2_EAX_REG_17__SCAN_IN), .A(n14439), .ZN(
        n14440) );
  OAI21_X1 U16272 ( .B1(n14467), .B2(n14441), .A(n14440), .ZN(P2_U2953) );
  INV_X1 U16273 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14445) );
  AOI21_X1 U16274 ( .B1(n14463), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14443), .ZN(
        n14444) );
  OAI21_X1 U16275 ( .B1(n14467), .B2(n14445), .A(n14444), .ZN(P2_U2956) );
  INV_X1 U16276 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14448) );
  AOI21_X1 U16277 ( .B1(n14463), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14446), .ZN(
        n14447) );
  OAI21_X1 U16278 ( .B1(n14467), .B2(n14448), .A(n14447), .ZN(P2_U2960) );
  INV_X1 U16279 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14451) );
  AOI21_X1 U16280 ( .B1(n14463), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14449), .ZN(
        n14450) );
  OAI21_X1 U16281 ( .B1(n14467), .B2(n14451), .A(n14450), .ZN(P2_U2955) );
  INV_X1 U16282 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14454) );
  AOI21_X1 U16283 ( .B1(n14463), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14452), .ZN(
        n14453) );
  OAI21_X1 U16284 ( .B1(n14467), .B2(n14454), .A(n14453), .ZN(P2_U2959) );
  INV_X1 U16285 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14457) );
  AOI21_X1 U16286 ( .B1(n14463), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14455), .ZN(
        n14456) );
  OAI21_X1 U16287 ( .B1(n14467), .B2(n14457), .A(n14456), .ZN(P2_U2957) );
  INV_X1 U16288 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14459) );
  AOI22_X1 U16289 ( .A1(n15596), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15601), .ZN(n15003) );
  INV_X1 U16290 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n17950) );
  OAI222_X1 U16291 ( .A1(n14388), .A2(n14459), .B1(n14458), .B2(n15003), .C1(
        n14477), .C2(n17950), .ZN(P2_U2982) );
  INV_X1 U16292 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U16293 ( .A1(n14463), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14460) );
  OAI211_X1 U16294 ( .C1(n14467), .C2(n14462), .A(n14461), .B(n14460), .ZN(
        P2_U2978) );
  INV_X1 U16295 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14466) );
  NAND2_X1 U16296 ( .A1(n14463), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14464) );
  OAI211_X1 U16297 ( .C1(n14467), .C2(n14466), .A(n14465), .B(n14464), .ZN(
        P2_U2980) );
  NOR2_X1 U16298 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14469) );
  OAI21_X1 U16299 ( .B1(n14470), .B2(n14469), .A(n14468), .ZN(n14471) );
  INV_X1 U16300 ( .A(n14471), .ZN(n14472) );
  MUX2_X1 U16301 ( .A(n14474), .B(n15076), .S(n16700), .Z(n14475) );
  OAI21_X1 U16302 ( .B1(n19825), .B2(n16732), .A(n14475), .ZN(P2_U2887) );
  INV_X1 U16303 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14481) );
  AND2_X1 U16304 ( .A1(n14042), .A2(n19017), .ZN(n14476) );
  NAND2_X1 U16305 ( .A1(n15038), .A2(n14476), .ZN(n15053) );
  OAI21_X1 U16306 ( .B1(n15053), .B2(n19332), .A(n14477), .ZN(n14478) );
  NAND2_X1 U16307 ( .A1(n17915), .A2(n14479), .ZN(n14609) );
  NOR2_X1 U16308 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15127), .ZN(n17936) );
  NOR2_X4 U16309 ( .A1(n17915), .A2(n17947), .ZN(n17935) );
  AOI22_X1 U16310 ( .A1(n17936), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14480) );
  OAI21_X1 U16311 ( .B1(n14481), .B2(n14609), .A(n14480), .ZN(P2_U2934) );
  INV_X1 U16312 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n15600) );
  AOI22_X1 U16313 ( .A1(n17936), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14482) );
  OAI21_X1 U16314 ( .B1(n15600), .B2(n14609), .A(n14482), .ZN(P2_U2933) );
  INV_X1 U16315 ( .A(n19842), .ZN(n17892) );
  MUX2_X1 U16316 ( .A(n14486), .B(n17372), .S(n16700), .Z(n14487) );
  OAI21_X1 U16317 ( .B1(n17892), .B2(n16732), .A(n14487), .ZN(P2_U2886) );
  MUX2_X1 U16318 ( .A(n15410), .B(n12110), .S(n16700), .Z(n14491) );
  OAI21_X1 U16319 ( .B1(n19940), .B2(n16732), .A(n14491), .ZN(P2_U2885) );
  OR2_X2 U16320 ( .A1(n15165), .A2(n15178), .ZN(n22484) );
  INV_X1 U16321 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14497) );
  INV_X1 U16322 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n14496) );
  NAND2_X1 U16323 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n22325) );
  INV_X1 U16324 ( .A(n15165), .ZN(n14492) );
  OAI21_X2 U16325 ( .B1(n17464), .B2(n22325), .A(n14492), .ZN(n22456) );
  NAND2_X1 U16326 ( .A1(n15178), .A2(n22325), .ZN(n14493) );
  INV_X1 U16327 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14494) );
  NOR2_X1 U16328 ( .A1(n16158), .A2(n14494), .ZN(n14495) );
  AOI21_X1 U16329 ( .B1(DATAI_15_), .B2(n16158), .A(n14495), .ZN(n16232) );
  OAI222_X1 U16330 ( .A1(n22484), .A2(n14497), .B1(n14496), .B2(n22414), .C1(
        n22478), .C2(n16232), .ZN(P1_U2967) );
  XNOR2_X1 U16331 ( .A(n14499), .B(n14498), .ZN(n15586) );
  NOR2_X1 U16332 ( .A1(n19825), .A2(n15586), .ZN(n14505) );
  OR2_X1 U16333 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  NAND2_X1 U16334 ( .A1(n14503), .A2(n14502), .ZN(n14758) );
  XNOR2_X1 U16335 ( .A(n19842), .B(n14758), .ZN(n14504) );
  NOR2_X1 U16336 ( .A1(n14504), .A2(n14505), .ZN(n14759) );
  AOI21_X1 U16337 ( .B1(n14505), .B2(n14504), .A(n14759), .ZN(n14513) );
  AND2_X1 U16338 ( .A1(n14171), .A2(n22349), .ZN(n15113) );
  NAND2_X1 U16339 ( .A1(n15112), .A2(n15113), .ZN(n14506) );
  NOR2_X1 U16340 ( .A1(n15115), .A2(n14506), .ZN(n14507) );
  AOI21_X1 U16341 ( .B1(n15038), .B2(n15101), .A(n14507), .ZN(n15056) );
  NAND2_X1 U16342 ( .A1(n15056), .A2(n14508), .ZN(n14509) );
  AOI22_X1 U16343 ( .A1(n20117), .A2(n14758), .B1(n20111), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14512) );
  AND2_X1 U16344 ( .A1(n14071), .A2(n12006), .ZN(n14510) );
  INV_X1 U16345 ( .A(n15047), .ZN(n16795) );
  NAND2_X1 U16346 ( .A1(n20064), .A2(n16795), .ZN(n14511) );
  OAI211_X1 U16347 ( .C1(n14513), .C2(n20065), .A(n14512), .B(n14511), .ZN(
        P2_U2918) );
  INV_X1 U16348 ( .A(n14514), .ZN(n14518) );
  INV_X1 U16349 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14517) );
  INV_X1 U16350 ( .A(n14515), .ZN(n14516) );
  AOI21_X1 U16351 ( .B1(n14518), .B2(n14517), .A(n14516), .ZN(n14582) );
  NAND2_X1 U16352 ( .A1(n14533), .A2(n14519), .ZN(n14520) );
  NAND2_X1 U16353 ( .A1(n14521), .A2(n14520), .ZN(n14718) );
  INV_X1 U16354 ( .A(n14522), .ZN(n14523) );
  NAND2_X1 U16355 ( .A1(n14523), .A2(n22343), .ZN(n22338) );
  NAND2_X1 U16356 ( .A1(n15178), .A2(n22338), .ZN(n14524) );
  NAND4_X1 U16357 ( .A1(n14620), .A2(n13156), .A3(n22325), .A4(n14524), .ZN(
        n14526) );
  NAND3_X1 U16358 ( .A1(n17436), .A2(n15178), .A3(n14712), .ZN(n14525) );
  NAND3_X1 U16359 ( .A1(n14718), .A2(n14526), .A3(n14525), .ZN(n14527) );
  NAND2_X1 U16360 ( .A1(n14527), .A2(n15163), .ZN(n14531) );
  NAND2_X1 U16361 ( .A1(n14797), .A2(n22338), .ZN(n15181) );
  NAND2_X1 U16362 ( .A1(n15181), .A2(n22325), .ZN(n14528) );
  OAI211_X1 U16363 ( .C1(n14686), .C2(n14528), .A(n14886), .B(n14629), .ZN(
        n14529) );
  NAND3_X1 U16364 ( .A1(n14883), .A2(n14529), .A3(n14839), .ZN(n14530) );
  INV_X1 U16365 ( .A(n14532), .ZN(n14535) );
  NAND2_X1 U16366 ( .A1(n14533), .A2(n14537), .ZN(n14534) );
  NAND2_X1 U16367 ( .A1(n14696), .A2(n15911), .ZN(n14714) );
  AND2_X1 U16368 ( .A1(n14534), .A2(n14714), .ZN(n15903) );
  OAI211_X1 U16369 ( .C1(n14817), .C2(n14547), .A(n14535), .B(n15903), .ZN(
        n14536) );
  NAND2_X1 U16370 ( .A1(n14537), .A2(n14725), .ZN(n14538) );
  NAND2_X1 U16371 ( .A1(n14538), .A2(n15177), .ZN(n14539) );
  AND2_X1 U16372 ( .A1(n14540), .A2(n14539), .ZN(n14543) );
  OAI211_X1 U16373 ( .C1(n14797), .C2(n14543), .A(n14542), .B(n14541), .ZN(
        n14690) );
  NOR2_X1 U16374 ( .A1(n14544), .A2(n14886), .ZN(n14545) );
  OR2_X1 U16375 ( .A1(n14690), .A2(n14545), .ZN(n14546) );
  INV_X1 U16376 ( .A(n16550), .ZN(n16397) );
  AND2_X1 U16377 ( .A1(n14696), .A2(n14222), .ZN(n15904) );
  AND2_X1 U16378 ( .A1(n16397), .A2(n22049), .ZN(n14612) );
  OAI22_X1 U16379 ( .A1(n14549), .A2(n15178), .B1(n14548), .B2(n14547), .ZN(
        n14550) );
  INV_X1 U16380 ( .A(n14551), .ZN(n14553) );
  OR2_X1 U16381 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14552) );
  NAND2_X1 U16382 ( .A1(n14553), .A2(n14552), .ZN(n15322) );
  INV_X1 U16383 ( .A(n15322), .ZN(n14554) );
  AND2_X1 U16384 ( .A1(n22108), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14581) );
  AOI21_X1 U16385 ( .B1(n22098), .B2(n14554), .A(n14581), .ZN(n14559) );
  NOR2_X1 U16386 ( .A1(n13115), .A2(n15195), .ZN(n14555) );
  NOR2_X1 U16387 ( .A1(n14557), .A2(n22108), .ZN(n14611) );
  OAI21_X1 U16388 ( .B1(n16548), .B2(n14611), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14558) );
  OAI211_X1 U16389 ( .C1(n14612), .C2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n14559), .B(n14558), .ZN(n14560) );
  AOI21_X1 U16390 ( .B1(n14582), .B2(n22099), .A(n14560), .ZN(n14561) );
  INV_X1 U16391 ( .A(n14561), .ZN(P1_U3031) );
  XNOR2_X1 U16392 ( .A(n19836), .B(n15586), .ZN(n14562) );
  NAND2_X1 U16393 ( .A1(n14562), .A2(n20119), .ZN(n14564) );
  INV_X1 U16394 ( .A(n15586), .ZN(n19280) );
  AOI22_X1 U16395 ( .A1(n20117), .A2(n19280), .B1(n20111), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14563) );
  OAI211_X1 U16396 ( .C1(n20292), .C2(n15004), .A(n14564), .B(n14563), .ZN(
        P2_U2919) );
  NOR2_X1 U16397 ( .A1(n16700), .A2(n12071), .ZN(n14569) );
  AOI21_X1 U16398 ( .B1(n12116), .B2(n16700), .A(n14569), .ZN(n14570) );
  OAI21_X1 U16399 ( .B1(n19941), .B2(n16732), .A(n14570), .ZN(P2_U2884) );
  OAI21_X1 U16400 ( .B1(n14572), .B2(n14571), .A(n14661), .ZN(n16097) );
  INV_X1 U16401 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n17805) );
  XNOR2_X1 U16402 ( .A(n14573), .B(n15917), .ZN(n16104) );
  OAI222_X1 U16403 ( .A1(n16097), .A2(n16146), .B1(n20574), .B2(n17805), .C1(
        n16104), .C2(n16143), .ZN(P1_U2871) );
  INV_X1 U16404 ( .A(n20614), .ZN(n20630) );
  INV_X1 U16405 ( .A(n14574), .ZN(n14577) );
  OAI21_X1 U16406 ( .B1(n14577), .B2(n14576), .A(n14575), .ZN(n15326) );
  INV_X1 U16407 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14578) );
  AOI21_X1 U16408 ( .B1(n16384), .B2(n14579), .A(n14578), .ZN(n14580) );
  AOI211_X1 U16409 ( .C1(n14582), .C2(n20595), .A(n14581), .B(n14580), .ZN(
        n14583) );
  OAI21_X1 U16410 ( .B1(n20630), .B2(n15326), .A(n14583), .ZN(P1_U2999) );
  INV_X1 U16411 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16412 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n17947), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17935), .ZN(n14584) );
  OAI21_X1 U16413 ( .B1(n14585), .B2(n14609), .A(n14584), .ZN(P2_U2935) );
  INV_X1 U16414 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U16415 ( .A1(n17947), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14586) );
  OAI21_X1 U16416 ( .B1(n14587), .B2(n14609), .A(n14586), .ZN(P2_U2929) );
  INV_X1 U16417 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14589) );
  AOI22_X1 U16418 ( .A1(n17947), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14588) );
  OAI21_X1 U16419 ( .B1(n14589), .B2(n14609), .A(n14588), .ZN(P2_U2928) );
  INV_X1 U16420 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U16421 ( .A1(n17947), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14590) );
  OAI21_X1 U16422 ( .B1(n14591), .B2(n14609), .A(n14590), .ZN(P2_U2931) );
  AOI22_X1 U16423 ( .A1(n17947), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14592) );
  OAI21_X1 U16424 ( .B1(n14593), .B2(n14609), .A(n14592), .ZN(P2_U2926) );
  AOI22_X1 U16425 ( .A1(n17947), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14594) );
  OAI21_X1 U16426 ( .B1(n14595), .B2(n14609), .A(n14594), .ZN(P2_U2925) );
  AOI22_X1 U16427 ( .A1(n17947), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14596) );
  OAI21_X1 U16428 ( .B1(n14597), .B2(n14609), .A(n14596), .ZN(P2_U2924) );
  AOI22_X1 U16429 ( .A1(n17947), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14598) );
  OAI21_X1 U16430 ( .B1(n14599), .B2(n14609), .A(n14598), .ZN(P2_U2923) );
  AOI22_X1 U16431 ( .A1(n17947), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14600) );
  OAI21_X1 U16432 ( .B1(n14601), .B2(n14609), .A(n14600), .ZN(P2_U2922) );
  INV_X1 U16433 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14603) );
  AOI22_X1 U16434 ( .A1(n17947), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U16435 ( .B1(n14603), .B2(n14609), .A(n14602), .ZN(P2_U2930) );
  INV_X1 U16436 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14605) );
  AOI22_X1 U16437 ( .A1(n17947), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14604) );
  OAI21_X1 U16438 ( .B1(n14605), .B2(n14609), .A(n14604), .ZN(P2_U2927) );
  AOI22_X1 U16439 ( .A1(n17936), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14606) );
  OAI21_X1 U16440 ( .B1(n14607), .B2(n14609), .A(n14606), .ZN(P2_U2921) );
  INV_X1 U16441 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15641) );
  AOI22_X1 U16442 ( .A1(n17936), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14608) );
  OAI21_X1 U16443 ( .B1(n15641), .B2(n14609), .A(n14608), .ZN(P2_U2932) );
  NOR2_X1 U16444 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16548), .ZN(
        n16407) );
  NOR3_X1 U16445 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n16407), .A3(
        n22071), .ZN(n14615) );
  NOR2_X1 U16446 ( .A1(n22067), .A2(n16104), .ZN(n14614) );
  INV_X1 U16447 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n14610) );
  NOR2_X1 U16448 ( .A1(n22044), .A2(n14610), .ZN(n15029) );
  INV_X1 U16449 ( .A(n14611), .ZN(n16552) );
  INV_X1 U16450 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21969) );
  AOI221_X1 U16451 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n16552), .C1(
        n14612), .C2(n16552), .A(n21969), .ZN(n14613) );
  NOR4_X1 U16452 ( .A1(n14615), .A2(n14614), .A3(n15029), .A4(n14613), .ZN(
        n14618) );
  OR2_X1 U16453 ( .A1(n14616), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15031) );
  NAND3_X1 U16454 ( .A1(n15031), .A2(n15030), .A3(n22099), .ZN(n14617) );
  NAND2_X1 U16455 ( .A1(n14618), .A2(n14617), .ZN(P1_U3030) );
  INV_X1 U16456 ( .A(n14688), .ZN(n17454) );
  NAND2_X1 U16457 ( .A1(n17454), .A2(n14620), .ZN(n14709) );
  NOR2_X1 U16458 ( .A1(n14686), .A2(n14712), .ZN(n17465) );
  NAND2_X1 U16459 ( .A1(n17465), .A2(n14222), .ZN(n14621) );
  NAND2_X1 U16460 ( .A1(n14709), .A2(n14621), .ZN(n14622) );
  NAND2_X1 U16461 ( .A1(n14622), .A2(n22325), .ZN(n14710) );
  OR2_X1 U16462 ( .A1(n14623), .A2(n15175), .ZN(n14624) );
  AOI21_X1 U16463 ( .B1(n14710), .B2(n14624), .A(n22303), .ZN(n14627) );
  NOR2_X1 U16464 ( .A1(n14714), .A2(n14625), .ZN(n14626) );
  AND2_X1 U16465 ( .A1(n14825), .A2(n14628), .ZN(n14634) );
  INV_X1 U16466 ( .A(n14634), .ZN(n14630) );
  AND2_X1 U16467 ( .A1(n14630), .A2(n14629), .ZN(n14631) );
  NAND2_X2 U16468 ( .A1(n16231), .A2(n14631), .ZN(n16243) );
  OR2_X1 U16469 ( .A1(n16158), .A2(n20641), .ZN(n14633) );
  NAND2_X1 U16470 ( .A1(n16158), .A2(DATAI_0_), .ZN(n14632) );
  AND2_X1 U16471 ( .A1(n14633), .A2(n14632), .ZN(n22386) );
  INV_X1 U16472 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n22391) );
  OAI222_X1 U16473 ( .A1(n15326), .A2(n16243), .B1(n22386), .B2(n16233), .C1(
        n16231), .C2(n22391), .ZN(P1_U2904) );
  OAI222_X1 U16474 ( .A1(n15322), .A2(n16143), .B1(n14225), .B2(n20574), .C1(
        n15326), .C2(n16146), .ZN(P1_U2872) );
  NAND2_X1 U16475 ( .A1(n13173), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16565) );
  NAND2_X1 U16476 ( .A1(n14638), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22560) );
  INV_X1 U16477 ( .A(n22560), .ZN(n22513) );
  AOI211_X1 U16478 ( .C1(n14778), .C2(n22590), .A(n22607), .B(n22513), .ZN(
        n14639) );
  AOI21_X1 U16479 ( .B1(n16565), .B2(n22593), .A(n14639), .ZN(n14645) );
  NOR2_X1 U16480 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22297) );
  INV_X1 U16481 ( .A(n22297), .ZN(n14640) );
  NAND2_X1 U16482 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16559) );
  INV_X1 U16483 ( .A(n13032), .ZN(n16579) );
  NAND2_X1 U16484 ( .A1(n16579), .A2(n14641), .ZN(n14642) );
  AOI21_X1 U16485 ( .B1(n14642), .B2(n13350), .A(P1_FLUSH_REG_SCAN_IN), .ZN(
        n16560) );
  NOR2_X1 U16486 ( .A1(n17473), .A2(n16559), .ZN(n14720) );
  OAI21_X1 U16487 ( .B1(n16560), .B2(P1_FLUSH_REG_SCAN_IN), .A(n14720), .ZN(
        n14643) );
  NAND2_X1 U16488 ( .A1(n16592), .A2(n14643), .ZN(n17476) );
  INV_X1 U16489 ( .A(n17476), .ZN(n14676) );
  NAND2_X1 U16490 ( .A1(n14676), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14644) );
  OAI21_X1 U16491 ( .B1(n14645), .B2(n14676), .A(n14644), .ZN(P1_U3477) );
  OR2_X1 U16492 ( .A1(n14648), .A2(n14647), .ZN(n14649) );
  NAND2_X1 U16493 ( .A1(n14646), .A2(n14649), .ZN(n20066) );
  INV_X1 U16494 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14653) );
  OAI21_X1 U16495 ( .B1(n14652), .B2(n14651), .A(n14650), .ZN(n15382) );
  MUX2_X1 U16496 ( .A(n14653), .B(n15382), .S(n16700), .Z(n14654) );
  OAI21_X1 U16497 ( .B1(n20066), .B2(n16732), .A(n14654), .ZN(P2_U2883) );
  XOR2_X1 U16498 ( .A(n14646), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14659)
         );
  AOI21_X1 U16499 ( .B1(n14656), .B2(n14650), .A(n14655), .ZN(n19040) );
  NOR2_X1 U16500 ( .A1(n16700), .A2(n12445), .ZN(n14657) );
  AOI21_X1 U16501 ( .B1(n19040), .B2(n16700), .A(n14657), .ZN(n14658) );
  OAI21_X1 U16502 ( .B1(n14659), .B2(n16732), .A(n14658), .ZN(P2_U2882) );
  NAND2_X1 U16503 ( .A1(n14660), .A2(n14661), .ZN(n14662) );
  AND2_X1 U16504 ( .A1(n14663), .A2(n14662), .ZN(n22119) );
  INV_X1 U16505 ( .A(n22119), .ZN(n14670) );
  INV_X1 U16506 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n14664) );
  OR2_X1 U16507 ( .A1(n16158), .A2(n14664), .ZN(n14666) );
  NAND2_X1 U16508 ( .A1(n16158), .A2(DATAI_2_), .ZN(n14665) );
  AND2_X1 U16509 ( .A1(n14666), .A2(n14665), .ZN(n22398) );
  INV_X1 U16510 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n22403) );
  OAI222_X1 U16511 ( .A1(n14670), .A2(n16243), .B1(n22398), .B2(n16233), .C1(
        n16231), .C2(n22403), .ZN(P1_U2902) );
  OR2_X1 U16512 ( .A1(n14668), .A2(n14667), .ZN(n14669) );
  NAND2_X1 U16513 ( .A1(n14740), .A2(n14669), .ZN(n22111) );
  INV_X1 U16514 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n14671) );
  OAI222_X1 U16515 ( .A1(n22111), .A2(n16143), .B1(n14671), .B2(n20574), .C1(
        n14670), .C2(n16146), .ZN(P1_U2870) );
  INV_X1 U16516 ( .A(n14673), .ZN(n15208) );
  AOI21_X1 U16517 ( .B1(n13936), .B2(n22513), .A(n22607), .ZN(n22611) );
  INV_X1 U16518 ( .A(n22611), .ZN(n16567) );
  AOI21_X1 U16519 ( .B1(n11647), .B2(n22560), .A(n16567), .ZN(n14674) );
  AOI21_X1 U16520 ( .B1(n16565), .B2(n15208), .A(n14674), .ZN(n14677) );
  NAND2_X1 U16521 ( .A1(n14676), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14675) );
  OAI21_X1 U16522 ( .B1(n14677), .B2(n14676), .A(n14675), .ZN(P1_U3476) );
  NOR2_X1 U16523 ( .A1(n14646), .A2(n12788), .ZN(n14678) );
  OAI211_X1 U16524 ( .C1(n14678), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16724), .B(n14765), .ZN(n14682) );
  OAI21_X1 U16525 ( .B1(n14680), .B2(n14655), .A(n14679), .ZN(n17851) );
  INV_X1 U16526 ( .A(n17851), .ZN(n19052) );
  NAND2_X1 U16527 ( .A1(n16700), .A2(n19052), .ZN(n14681) );
  OAI211_X1 U16528 ( .C1(n16700), .C2(n19044), .A(n14682), .B(n14681), .ZN(
        P2_U2881) );
  INV_X1 U16529 ( .A(n16564), .ZN(n14705) );
  INV_X1 U16530 ( .A(n14683), .ZN(n14685) );
  AND3_X1 U16531 ( .A1(n14686), .A2(n14685), .A3(n14684), .ZN(n14687) );
  NAND2_X1 U16532 ( .A1(n14688), .A2(n14687), .ZN(n14689) );
  NOR2_X1 U16533 ( .A1(n14690), .A2(n14689), .ZN(n16570) );
  INV_X1 U16534 ( .A(n14694), .ZN(n14691) );
  OAI21_X1 U16535 ( .B1(n16572), .B2(n13305), .A(n14691), .ZN(n14693) );
  NOR2_X1 U16536 ( .A1(n14693), .A2(n14692), .ZN(n14706) );
  NOR2_X1 U16537 ( .A1(n14725), .A2(n14706), .ZN(n14695) );
  INV_X1 U16538 ( .A(n16572), .ZN(n16578) );
  AOI21_X1 U16539 ( .B1(n16570), .B2(n14695), .A(n11716), .ZN(n14704) );
  NAND2_X1 U16540 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14700) );
  INV_X1 U16541 ( .A(n14700), .ZN(n14699) );
  AND2_X1 U16542 ( .A1(n15195), .A2(n21947), .ZN(n15914) );
  NAND2_X1 U16543 ( .A1(n16578), .A2(n14697), .ZN(n14698) );
  AOI22_X1 U16544 ( .A1(n17439), .A2(n14699), .B1(n11731), .B2(n14698), .ZN(
        n14702) );
  NAND2_X1 U16545 ( .A1(n17439), .A2(n14700), .ZN(n14701) );
  MUX2_X1 U16546 ( .A(n14702), .B(n14701), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14703) );
  OAI211_X1 U16547 ( .C1(n14705), .C2(n16570), .A(n14704), .B(n14703), .ZN(
        n17435) );
  INV_X1 U16548 ( .A(n22289), .ZN(n17401) );
  INV_X1 U16549 ( .A(n14706), .ZN(n14707) );
  AOI22_X1 U16550 ( .A1(n17435), .A2(n17401), .B1(n22298), .B2(n14707), .ZN(
        n14724) );
  NAND2_X1 U16551 ( .A1(n17439), .A2(n15910), .ZN(n14708) );
  NAND2_X1 U16552 ( .A1(n14709), .A2(n14708), .ZN(n15164) );
  INV_X1 U16553 ( .A(n22325), .ZN(n22327) );
  OAI21_X1 U16554 ( .B1(n22327), .B2(n22338), .A(n14710), .ZN(n14711) );
  OAI21_X1 U16555 ( .B1(n17465), .B2(n15164), .A(n14711), .ZN(n14719) );
  INV_X1 U16556 ( .A(n15904), .ZN(n14713) );
  MUX2_X1 U16557 ( .A(n14714), .B(n14713), .S(n14712), .Z(n14717) );
  INV_X1 U16558 ( .A(n15195), .ZN(n14715) );
  NAND2_X1 U16559 ( .A1(n14715), .A2(n14839), .ZN(n14716) );
  NAND4_X1 U16560 ( .A1(n14719), .A2(n14718), .A3(n14717), .A4(n14716), .ZN(
        n17457) );
  INV_X1 U16561 ( .A(n17457), .ZN(n14722) );
  INV_X1 U16562 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n14721) );
  INV_X1 U16563 ( .A(n14720), .ZN(n22294) );
  OAI22_X1 U16564 ( .A1(n14722), .A2(n22303), .B1(n14721), .B2(n22294), .ZN(
        n17400) );
  NAND2_X1 U16565 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n22286), .ZN(
        n14723) );
  OAI21_X1 U16566 ( .B1(n14724), .B2(n22286), .A(n14723), .ZN(P1_U3469) );
  XNOR2_X1 U16567 ( .A(n16572), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14731) );
  NOR2_X1 U16568 ( .A1(n14725), .A2(n14731), .ZN(n14726) );
  AOI22_X1 U16569 ( .A1(n16570), .A2(n14726), .B1(n11731), .B2(n14731), .ZN(
        n14730) );
  NAND2_X1 U16570 ( .A1(n17439), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14728) );
  NAND2_X1 U16571 ( .A1(n17439), .A2(n14727), .ZN(n16571) );
  MUX2_X1 U16572 ( .A(n14728), .B(n16571), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n14729) );
  OAI211_X1 U16573 ( .C1(n14673), .C2(n16570), .A(n14730), .B(n14729), .ZN(
        n17434) );
  INV_X1 U16574 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16415) );
  OAI22_X1 U16575 ( .A1(n16415), .A2(n21969), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16576) );
  INV_X1 U16576 ( .A(n16576), .ZN(n14733) );
  NOR2_X1 U16577 ( .A1(n15308), .A2(n14517), .ZN(n16577) );
  INV_X1 U16578 ( .A(n14731), .ZN(n14732) );
  AOI222_X1 U16579 ( .A1(n17434), .A2(n17401), .B1(n14733), .B2(n16577), .C1(
        n22298), .C2(n14732), .ZN(n14735) );
  NAND2_X1 U16580 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n22286), .ZN(
        n14734) );
  OAI21_X1 U16581 ( .B1(n14735), .B2(n22286), .A(n14734), .ZN(P1_U3472) );
  OAI21_X1 U16582 ( .B1(n14738), .B2(n14737), .A(n14950), .ZN(n15199) );
  INV_X1 U16583 ( .A(n20570), .ZN(n14739) );
  AOI21_X1 U16584 ( .B1(n14741), .B2(n14740), .A(n14739), .ZN(n21989) );
  INV_X1 U16585 ( .A(n20574), .ZN(n16119) );
  AOI22_X1 U16586 ( .A1(n21989), .A2(n20572), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n16119), .ZN(n14742) );
  OAI21_X1 U16587 ( .B1(n15199), .B2(n16146), .A(n14742), .ZN(P1_U2869) );
  INV_X1 U16588 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n14743) );
  OR2_X1 U16589 ( .A1(n16158), .A2(n14743), .ZN(n14745) );
  NAND2_X1 U16590 ( .A1(n16158), .A2(DATAI_1_), .ZN(n14744) );
  AND2_X1 U16591 ( .A1(n14745), .A2(n14744), .ZN(n22392) );
  INV_X1 U16592 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n22397) );
  OAI222_X1 U16593 ( .A1(n16097), .A2(n16243), .B1(n22392), .B2(n16233), .C1(
        n16231), .C2(n22397), .ZN(P1_U2903) );
  AND2_X1 U16594 ( .A1(n17299), .A2(n14746), .ZN(n14747) );
  OR2_X1 U16595 ( .A1(n14747), .A2(n15446), .ZN(n19070) );
  INV_X1 U16596 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n17940) );
  OAI222_X1 U16597 ( .A1(n15004), .A2(n14748), .B1(n19070), .B2(n20071), .C1(
        n17940), .C2(n15640), .ZN(P2_U2908) );
  XNOR2_X1 U16598 ( .A(n14749), .B(n14750), .ZN(n19056) );
  INV_X1 U16599 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n17928) );
  OAI222_X1 U16600 ( .A1(n15004), .A2(n20024), .B1(n19056), .B2(n20071), .C1(
        n17928), .C2(n15640), .ZN(P2_U2913) );
  INV_X1 U16601 ( .A(n14752), .ZN(n14753) );
  XNOR2_X1 U16602 ( .A(n14751), .B(n14753), .ZN(n15490) );
  INV_X1 U16603 ( .A(n15490), .ZN(n17330) );
  INV_X1 U16604 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n17930) );
  OAI222_X1 U16605 ( .A1(n15004), .A2(n19818), .B1(n17330), .B2(n20071), .C1(
        n17930), .C2(n15640), .ZN(P2_U2912) );
  NOR2_X1 U16606 ( .A1(n14756), .A2(n14755), .ZN(n14757) );
  OR2_X1 U16607 ( .A1(n14754), .A2(n14757), .ZN(n15480) );
  INV_X1 U16608 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17932) );
  OAI222_X1 U16609 ( .A1(n15004), .A2(n16771), .B1(n15480), .B2(n20071), .C1(
        n17932), .C2(n15640), .ZN(P2_U2911) );
  INV_X1 U16610 ( .A(n14758), .ZN(n19026) );
  AOI21_X1 U16611 ( .B1(n19026), .B2(n17892), .A(n14759), .ZN(n14893) );
  XNOR2_X1 U16612 ( .A(n14761), .B(n14760), .ZN(n17360) );
  INV_X1 U16613 ( .A(n17360), .ZN(n17886) );
  XNOR2_X1 U16614 ( .A(n14893), .B(n17886), .ZN(n14892) );
  XNOR2_X1 U16615 ( .A(n14892), .B(n19940), .ZN(n14762) );
  NAND2_X1 U16616 ( .A1(n14762), .A2(n20119), .ZN(n14764) );
  AOI22_X1 U16617 ( .A1(n20117), .A2(n17360), .B1(n20111), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n14763) );
  OAI211_X1 U16618 ( .C1(n20205), .C2(n15004), .A(n14764), .B(n14763), .ZN(
        P2_U2917) );
  XOR2_X1 U16619 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n14765), .Z(n14770)
         );
  OR2_X1 U16620 ( .A1(n14767), .A2(n14766), .ZN(n14768) );
  NAND2_X1 U16621 ( .A1(n14903), .A2(n14768), .ZN(n17331) );
  MUX2_X1 U16622 ( .A(n12451), .B(n17331), .S(n16700), .Z(n14769) );
  OAI21_X1 U16623 ( .B1(n14770), .B2(n16732), .A(n14769), .ZN(P2_U2880) );
  INV_X1 U16624 ( .A(n14771), .ZN(n15551) );
  NAND2_X1 U16625 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  NAND2_X1 U16626 ( .A1(n15551), .A2(n14774), .ZN(n19089) );
  INV_X1 U16627 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n17944) );
  OAI222_X1 U16628 ( .A1(n15004), .A2(n16738), .B1(n19089), .B2(n20071), .C1(
        n17944), .C2(n15640), .ZN(P2_U2906) );
  INV_X1 U16629 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n14775) );
  OR2_X1 U16630 ( .A1(n16158), .A2(n14775), .ZN(n14777) );
  NAND2_X1 U16631 ( .A1(n16158), .A2(DATAI_3_), .ZN(n14776) );
  AND2_X1 U16632 ( .A1(n14777), .A2(n14776), .ZN(n22404) );
  INV_X1 U16633 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n22409) );
  OAI222_X1 U16634 ( .A1(n15199), .A2(n16243), .B1(n22404), .B2(n16233), .C1(
        n16231), .C2(n22409), .ZN(P1_U2901) );
  NOR3_X1 U16635 ( .A1(n22585), .A2(n22586), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n22570) );
  NAND2_X1 U16636 ( .A1(n13936), .A2(n14778), .ZN(n14848) );
  INV_X1 U16637 ( .A(n22582), .ZN(n22486) );
  INV_X1 U16638 ( .A(n22607), .ZN(n22563) );
  INV_X1 U16639 ( .A(n14849), .ZN(n17397) );
  INV_X1 U16640 ( .A(n15210), .ZN(n14953) );
  NAND2_X1 U16641 ( .A1(n22604), .A2(n14953), .ZN(n14781) );
  INV_X1 U16642 ( .A(n22570), .ZN(n14779) );
  NOR2_X1 U16643 ( .A1(n22571), .A2(n14779), .ZN(n14841) );
  INV_X1 U16644 ( .A(n14841), .ZN(n14780) );
  NAND2_X1 U16645 ( .A1(n14781), .A2(n14780), .ZN(n14789) );
  INV_X1 U16646 ( .A(n14789), .ZN(n14782) );
  OAI211_X1 U16647 ( .C1(n14785), .C2(n22590), .A(n22563), .B(n14782), .ZN(
        n14783) );
  OAI211_X1 U16648 ( .C1(n22559), .C2(n22570), .A(n14783), .B(n22613), .ZN(
        n14784) );
  INV_X1 U16649 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14796) );
  NAND2_X1 U16650 ( .A1(n20614), .A2(n15823), .ZN(n14838) );
  NAND2_X1 U16651 ( .A1(n16158), .A2(n20614), .ZN(n14837) );
  INV_X1 U16652 ( .A(n14837), .ZN(n14836) );
  AOI22_X1 U16653 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n14835), .B1(DATAI_31_), 
        .B2(n14836), .ZN(n22849) );
  INV_X1 U16654 ( .A(n22849), .ZN(n22833) );
  AOI22_X1 U16655 ( .A1(DATAI_23_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n22838) );
  INV_X1 U16656 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n14786) );
  OR2_X1 U16657 ( .A1(n16158), .A2(n14786), .ZN(n14788) );
  NAND2_X1 U16658 ( .A1(n16158), .A2(DATAI_7_), .ZN(n14787) );
  NAND2_X1 U16659 ( .A1(n14788), .A2(n14787), .ZN(n16181) );
  NAND2_X1 U16660 ( .A1(n14789), .A2(n22563), .ZN(n14791) );
  NAND2_X1 U16661 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22570), .ZN(n14790) );
  NAND2_X1 U16662 ( .A1(n14791), .A2(n14790), .ZN(n14842) );
  AOI22_X1 U16663 ( .A1(n22841), .A2(n14842), .B1(n22839), .B2(n14841), .ZN(
        n14793) );
  OAI21_X1 U16664 ( .B1(n22591), .B2(n22838), .A(n14793), .ZN(n14794) );
  AOI21_X1 U16665 ( .B1(n14828), .B2(n22833), .A(n14794), .ZN(n14795) );
  OAI21_X1 U16666 ( .B1(n14847), .B2(n14796), .A(n14795), .ZN(P1_U3144) );
  INV_X1 U16667 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U16668 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14835), .B1(DATAI_25_), 
        .B2(n14836), .ZN(n22646) );
  AOI22_X1 U16669 ( .A1(DATAI_17_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n22640) );
  NOR2_X1 U16670 ( .A1(n14840), .A2(n14797), .ZN(n22641) );
  AOI22_X1 U16671 ( .A1(n22642), .A2(n14842), .B1(n22641), .B2(n14841), .ZN(
        n14798) );
  OAI21_X1 U16672 ( .B1(n22591), .B2(n22640), .A(n14798), .ZN(n14799) );
  AOI21_X1 U16673 ( .B1(n14828), .B2(n22637), .A(n14799), .ZN(n14800) );
  OAI21_X1 U16674 ( .B1(n14847), .B2(n14801), .A(n14800), .ZN(P1_U3138) );
  INV_X1 U16675 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14808) );
  AOI22_X1 U16676 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14835), .B1(DATAI_30_), 
        .B2(n14836), .ZN(n22781) );
  AOI22_X1 U16677 ( .A1(DATAI_22_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n22775) );
  OR2_X1 U16678 ( .A1(n16158), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14803) );
  INV_X1 U16679 ( .A(DATAI_6_), .ZN(n17690) );
  NAND2_X1 U16680 ( .A1(n16158), .A2(n17690), .ZN(n14802) );
  AND2_X1 U16681 ( .A1(n14803), .A2(n14802), .ZN(n16187) );
  NAND2_X1 U16682 ( .A1(n14816), .A2(n16187), .ZN(n22771) );
  INV_X1 U16683 ( .A(n22771), .ZN(n22777) );
  AOI22_X1 U16684 ( .A1(n22777), .A2(n14842), .B1(n22776), .B2(n14841), .ZN(
        n14805) );
  OAI21_X1 U16685 ( .B1(n22591), .B2(n22775), .A(n14805), .ZN(n14806) );
  AOI21_X1 U16686 ( .B1(n14828), .B2(n22772), .A(n14806), .ZN(n14807) );
  OAI21_X1 U16687 ( .B1(n14847), .B2(n14808), .A(n14807), .ZN(P1_U3143) );
  INV_X1 U16688 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14813) );
  AOI22_X1 U16689 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14835), .B1(DATAI_27_), 
        .B2(n14836), .ZN(n22700) );
  INV_X1 U16690 ( .A(n22700), .ZN(n22691) );
  AOI22_X1 U16691 ( .A1(DATAI_19_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n22694) );
  AOI22_X1 U16692 ( .A1(n22696), .A2(n14842), .B1(n22695), .B2(n14841), .ZN(
        n14810) );
  OAI21_X1 U16693 ( .B1(n22591), .B2(n22694), .A(n14810), .ZN(n14811) );
  AOI21_X1 U16694 ( .B1(n14828), .B2(n22691), .A(n14811), .ZN(n14812) );
  OAI21_X1 U16695 ( .B1(n14847), .B2(n14813), .A(n14812), .ZN(P1_U3140) );
  INV_X1 U16696 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14821) );
  AOI22_X1 U16697 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14835), .B1(DATAI_28_), 
        .B2(n14836), .ZN(n22727) );
  INV_X1 U16698 ( .A(n22727), .ZN(n22718) );
  AOI22_X1 U16699 ( .A1(DATAI_20_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n22721) );
  OR2_X1 U16700 ( .A1(n16158), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14815) );
  INV_X1 U16701 ( .A(DATAI_4_), .ZN(n17527) );
  NAND2_X1 U16702 ( .A1(n16158), .A2(n17527), .ZN(n14814) );
  AND2_X1 U16703 ( .A1(n14815), .A2(n14814), .ZN(n22410) );
  NAND2_X1 U16704 ( .A1(n14816), .A2(n22410), .ZN(n22717) );
  INV_X1 U16705 ( .A(n22717), .ZN(n22723) );
  AOI22_X1 U16706 ( .A1(n22723), .A2(n14842), .B1(n22722), .B2(n14841), .ZN(
        n14818) );
  OAI21_X1 U16707 ( .B1(n22591), .B2(n22721), .A(n14818), .ZN(n14819) );
  AOI21_X1 U16708 ( .B1(n14828), .B2(n22718), .A(n14819), .ZN(n14820) );
  OAI21_X1 U16709 ( .B1(n14847), .B2(n14821), .A(n14820), .ZN(P1_U3141) );
  INV_X1 U16710 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16711 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14835), .B1(DATAI_29_), 
        .B2(n14836), .ZN(n22754) );
  INV_X1 U16712 ( .A(n22754), .ZN(n22745) );
  AOI22_X1 U16713 ( .A1(DATAI_21_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n22748) );
  INV_X1 U16714 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n14822) );
  OR2_X1 U16715 ( .A1(n16158), .A2(n14822), .ZN(n14824) );
  NAND2_X1 U16716 ( .A1(n16158), .A2(DATAI_5_), .ZN(n14823) );
  AND2_X1 U16717 ( .A1(n14824), .A2(n14823), .ZN(n22418) );
  AOI22_X1 U16718 ( .A1(n22750), .A2(n14842), .B1(n22749), .B2(n14841), .ZN(
        n14826) );
  OAI21_X1 U16719 ( .B1(n22591), .B2(n22748), .A(n14826), .ZN(n14827) );
  AOI21_X1 U16720 ( .B1(n14828), .B2(n22745), .A(n14827), .ZN(n14829) );
  OAI21_X1 U16721 ( .B1(n14847), .B2(n14830), .A(n14829), .ZN(P1_U3142) );
  INV_X1 U16722 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14834) );
  AOI22_X1 U16723 ( .A1(DATAI_16_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n22601) );
  INV_X1 U16724 ( .A(n22601), .ZN(n22616) );
  AOI22_X1 U16725 ( .A1(DATAI_24_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n22619) );
  AOI22_X1 U16726 ( .A1(n22609), .A2(n14842), .B1(n22608), .B2(n14841), .ZN(
        n14831) );
  OAI21_X1 U16727 ( .B1(n22823), .B2(n22619), .A(n14831), .ZN(n14832) );
  AOI21_X1 U16728 ( .B1(n22834), .B2(n22616), .A(n14832), .ZN(n14833) );
  OAI21_X1 U16729 ( .B1(n14847), .B2(n14834), .A(n14833), .ZN(P1_U3137) );
  INV_X1 U16730 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U16731 ( .A1(DATAI_18_), .A2(n14836), .B1(n14835), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n22667) );
  INV_X1 U16732 ( .A(n22667), .ZN(n22670) );
  INV_X1 U16733 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20688) );
  INV_X1 U16734 ( .A(DATAI_26_), .ZN(n17652) );
  OAI22_X1 U16735 ( .A1(n20688), .A2(n14838), .B1(n17652), .B2(n14837), .ZN(
        n22664) );
  INV_X1 U16736 ( .A(n22664), .ZN(n22673) );
  AOI22_X1 U16737 ( .A1(n22669), .A2(n14842), .B1(n22668), .B2(n14841), .ZN(
        n14843) );
  OAI21_X1 U16738 ( .B1(n22823), .B2(n22673), .A(n14843), .ZN(n14844) );
  AOI21_X1 U16739 ( .B1(n22834), .B2(n22670), .A(n14844), .ZN(n14845) );
  OAI21_X1 U16740 ( .B1(n14847), .B2(n14846), .A(n14845), .ZN(P1_U3139) );
  NOR3_X1 U16741 ( .A1(n22585), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14854) );
  OR2_X1 U16742 ( .A1(n14673), .A2(n14849), .ZN(n22528) );
  INV_X1 U16743 ( .A(n14854), .ZN(n16583) );
  NOR2_X1 U16744 ( .A1(n22571), .A2(n16583), .ZN(n14852) );
  AOI21_X1 U16745 ( .B1(n16590), .B2(n14953), .A(n14852), .ZN(n14853) );
  OAI211_X1 U16746 ( .C1(n14851), .C2(n22590), .A(n22563), .B(n14853), .ZN(
        n14850) );
  NAND2_X1 U16747 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n14858) );
  INV_X1 U16748 ( .A(n22775), .ZN(n22778) );
  INV_X1 U16749 ( .A(n22776), .ZN(n22767) );
  INV_X1 U16750 ( .A(n14852), .ZN(n14879) );
  INV_X1 U16751 ( .A(n14853), .ZN(n14855) );
  AOI22_X1 U16752 ( .A1(n14855), .A2(n22563), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14854), .ZN(n14878) );
  OAI22_X1 U16753 ( .A1(n22767), .A2(n14879), .B1(n14878), .B2(n22771), .ZN(
        n14856) );
  AOI21_X1 U16754 ( .B1(n22802), .B2(n22778), .A(n14856), .ZN(n14857) );
  OAI211_X1 U16755 ( .C1(n22781), .C2(n16588), .A(n14858), .B(n14857), .ZN(
        P1_U3079) );
  NAND2_X1 U16756 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n14861) );
  INV_X1 U16757 ( .A(n22640), .ZN(n22643) );
  INV_X1 U16758 ( .A(n22641), .ZN(n22632) );
  OAI22_X1 U16759 ( .A1(n22632), .A2(n14879), .B1(n14878), .B2(n22636), .ZN(
        n14859) );
  AOI21_X1 U16760 ( .B1(n22802), .B2(n22643), .A(n14859), .ZN(n14860) );
  OAI211_X1 U16761 ( .C1(n22646), .C2(n16588), .A(n14861), .B(n14860), .ZN(
        P1_U3074) );
  NAND2_X1 U16762 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n14864) );
  INV_X1 U16763 ( .A(n22838), .ZN(n22843) );
  INV_X1 U16764 ( .A(n22839), .ZN(n22821) );
  INV_X1 U16765 ( .A(n22841), .ZN(n22829) );
  OAI22_X1 U16766 ( .A1(n22821), .A2(n14879), .B1(n14878), .B2(n22829), .ZN(
        n14862) );
  AOI21_X1 U16767 ( .B1(n22802), .B2(n22843), .A(n14862), .ZN(n14863) );
  OAI211_X1 U16768 ( .C1(n22849), .C2(n16588), .A(n14864), .B(n14863), .ZN(
        P1_U3080) );
  NAND2_X1 U16769 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n14867) );
  INV_X1 U16770 ( .A(n22668), .ZN(n22659) );
  OAI22_X1 U16771 ( .A1(n22659), .A2(n14879), .B1(n14878), .B2(n22663), .ZN(
        n14865) );
  AOI21_X1 U16772 ( .B1(n16621), .B2(n22664), .A(n14865), .ZN(n14866) );
  OAI211_X1 U16773 ( .C1(n22667), .C2(n22526), .A(n14867), .B(n14866), .ZN(
        P1_U3075) );
  NAND2_X1 U16774 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n14870) );
  INV_X1 U16775 ( .A(n22748), .ZN(n22751) );
  INV_X1 U16776 ( .A(n22749), .ZN(n22740) );
  OAI22_X1 U16777 ( .A1(n22740), .A2(n14879), .B1(n14878), .B2(n22744), .ZN(
        n14868) );
  AOI21_X1 U16778 ( .B1(n22802), .B2(n22751), .A(n14868), .ZN(n14869) );
  OAI211_X1 U16779 ( .C1(n22754), .C2(n16588), .A(n14870), .B(n14869), .ZN(
        P1_U3078) );
  NAND2_X1 U16780 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n14873) );
  INV_X1 U16781 ( .A(n22694), .ZN(n22697) );
  INV_X1 U16782 ( .A(n22695), .ZN(n22686) );
  OAI22_X1 U16783 ( .A1(n22686), .A2(n14879), .B1(n14878), .B2(n22690), .ZN(
        n14871) );
  AOI21_X1 U16784 ( .B1(n22802), .B2(n22697), .A(n14871), .ZN(n14872) );
  OAI211_X1 U16785 ( .C1(n22700), .C2(n16588), .A(n14873), .B(n14872), .ZN(
        P1_U3076) );
  NAND2_X1 U16786 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n14876) );
  INV_X1 U16787 ( .A(n22619), .ZN(n22598) );
  INV_X1 U16788 ( .A(n22608), .ZN(n22572) );
  OAI22_X1 U16789 ( .A1(n22572), .A2(n14879), .B1(n14878), .B2(n22581), .ZN(
        n14874) );
  AOI21_X1 U16790 ( .B1(n16621), .B2(n22598), .A(n14874), .ZN(n14875) );
  OAI211_X1 U16791 ( .C1(n22601), .C2(n22526), .A(n14876), .B(n14875), .ZN(
        P1_U3073) );
  NAND2_X1 U16792 ( .A1(n14877), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n14882) );
  INV_X1 U16793 ( .A(n22721), .ZN(n22724) );
  INV_X1 U16794 ( .A(n22722), .ZN(n22713) );
  OAI22_X1 U16795 ( .A1(n22713), .A2(n14879), .B1(n14878), .B2(n22717), .ZN(
        n14880) );
  AOI21_X1 U16796 ( .B1(n22802), .B2(n22724), .A(n14880), .ZN(n14881) );
  OAI211_X1 U16797 ( .C1(n22727), .C2(n16588), .A(n14882), .B(n14881), .ZN(
        P1_U3077) );
  INV_X1 U16798 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n22400) );
  NAND2_X1 U16799 ( .A1(n17439), .A2(n14883), .ZN(n14884) );
  INV_X1 U16800 ( .A(n22338), .ZN(n17463) );
  NAND2_X1 U16801 ( .A1(n20463), .A2(n14886), .ZN(n15318) );
  NOR2_X1 U16802 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16559), .ZN(n15290) );
  NOR2_X4 U16803 ( .A1(n21945), .A2(n20463), .ZN(n20474) );
  AOI22_X1 U16804 ( .A1(n15290), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14887) );
  OAI21_X1 U16805 ( .B1(n22400), .B2(n15318), .A(n14887), .ZN(P1_U2918) );
  INV_X1 U16806 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n22394) );
  AOI22_X1 U16807 ( .A1(n15290), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14888) );
  OAI21_X1 U16808 ( .B1(n22394), .B2(n15318), .A(n14888), .ZN(P1_U2919) );
  OR2_X1 U16809 ( .A1(n11572), .A2(n14889), .ZN(n14891) );
  NAND2_X1 U16810 ( .A1(n14891), .A2(n14890), .ZN(n17896) );
  NAND2_X1 U16811 ( .A1(n14892), .A2(n17897), .ZN(n14896) );
  XNOR2_X1 U16812 ( .A(n19960), .B(n17896), .ZN(n14894) );
  NAND2_X1 U16813 ( .A1(n14893), .A2(n17360), .ZN(n14895) );
  NAND3_X1 U16814 ( .A1(n14896), .A2(n14894), .A3(n14895), .ZN(n14976) );
  INV_X1 U16815 ( .A(n14976), .ZN(n14898) );
  AOI21_X1 U16816 ( .B1(n14896), .B2(n14895), .A(n14894), .ZN(n14897) );
  OAI21_X1 U16817 ( .B1(n14898), .B2(n14897), .A(n20119), .ZN(n14901) );
  INV_X1 U16818 ( .A(n20165), .ZN(n14899) );
  AOI22_X1 U16819 ( .A1(n20064), .A2(n14899), .B1(n20111), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n14900) );
  OAI211_X1 U16820 ( .C1(n17896), .C2(n16790), .A(n14901), .B(n14900), .ZN(
        P2_U2916) );
  NAND2_X1 U16821 ( .A1(n14903), .A2(n14902), .ZN(n14904) );
  AND2_X1 U16822 ( .A1(n14911), .A2(n14904), .ZN(n19297) );
  INV_X1 U16823 ( .A(n19297), .ZN(n15487) );
  OAI211_X1 U16824 ( .C1(n14907), .C2(n14906), .A(n14905), .B(n16724), .ZN(
        n14909) );
  NAND2_X1 U16825 ( .A1(n15538), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U16826 ( .C1(n15487), .C2(n15538), .A(n14909), .B(n14908), .ZN(
        P2_U2879) );
  XNOR2_X1 U16827 ( .A(n14905), .B(n14982), .ZN(n14915) );
  AND2_X1 U16828 ( .A1(n14911), .A2(n14910), .ZN(n14912) );
  NOR2_X1 U16829 ( .A1(n14981), .A2(n14912), .ZN(n17311) );
  NOR2_X1 U16830 ( .A1(n16700), .A2(n12462), .ZN(n14913) );
  AOI21_X1 U16831 ( .B1(n17311), .B2(n16700), .A(n14913), .ZN(n14914) );
  OAI21_X1 U16832 ( .B1(n14915), .B2(n16732), .A(n14914), .ZN(P2_U2878) );
  INV_X1 U16833 ( .A(n22487), .ZN(n22554) );
  INV_X1 U16834 ( .A(n14917), .ZN(n14916) );
  NOR3_X1 U16835 ( .A1(n22585), .A2(n22584), .A3(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n22530) );
  NAND2_X1 U16836 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14924) );
  NAND2_X1 U16837 ( .A1(n14638), .A2(n11155), .ZN(n22501) );
  NAND2_X1 U16838 ( .A1(n14918), .A2(n22586), .ZN(n14945) );
  AND2_X1 U16839 ( .A1(n11610), .A2(n17438), .ZN(n22603) );
  INV_X1 U16840 ( .A(n22603), .ZN(n14920) );
  OAI21_X1 U16841 ( .B1(n22528), .B2(n14920), .A(n14945), .ZN(n14921) );
  AOI22_X1 U16842 ( .A1(n14921), .A2(n22563), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n22530), .ZN(n14944) );
  OAI22_X1 U16843 ( .A1(n22821), .A2(n14945), .B1(n14944), .B2(n22829), .ZN(
        n14922) );
  AOI21_X1 U16844 ( .B1(n22803), .B2(n22833), .A(n14922), .ZN(n14923) );
  OAI211_X1 U16845 ( .C1(n22838), .C2(n17833), .A(n14924), .B(n14923), .ZN(
        P1_U3096) );
  NAND2_X1 U16846 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14927) );
  OAI22_X1 U16847 ( .A1(n22767), .A2(n14945), .B1(n22771), .B2(n14944), .ZN(
        n14925) );
  AOI21_X1 U16848 ( .B1(n22803), .B2(n22772), .A(n14925), .ZN(n14926) );
  OAI211_X1 U16849 ( .C1(n22775), .C2(n17833), .A(n14927), .B(n14926), .ZN(
        P1_U3095) );
  NAND2_X1 U16850 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14930) );
  OAI22_X1 U16851 ( .A1(n22713), .A2(n14945), .B1(n22717), .B2(n14944), .ZN(
        n14928) );
  AOI21_X1 U16852 ( .B1(n22803), .B2(n22718), .A(n14928), .ZN(n14929) );
  OAI211_X1 U16853 ( .C1(n22721), .C2(n17833), .A(n14930), .B(n14929), .ZN(
        P1_U3093) );
  NAND2_X1 U16854 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14933) );
  OAI22_X1 U16855 ( .A1(n22740), .A2(n14945), .B1(n14944), .B2(n22744), .ZN(
        n14931) );
  AOI21_X1 U16856 ( .B1(n22803), .B2(n22745), .A(n14931), .ZN(n14932) );
  OAI211_X1 U16857 ( .C1(n22748), .C2(n17833), .A(n14933), .B(n14932), .ZN(
        P1_U3094) );
  NAND2_X1 U16858 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14936) );
  OAI22_X1 U16859 ( .A1(n22686), .A2(n14945), .B1(n14944), .B2(n22690), .ZN(
        n14934) );
  AOI21_X1 U16860 ( .B1(n22803), .B2(n22691), .A(n14934), .ZN(n14935) );
  OAI211_X1 U16861 ( .C1(n22694), .C2(n17833), .A(n14936), .B(n14935), .ZN(
        P1_U3092) );
  NAND2_X1 U16862 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14939) );
  OAI22_X1 U16863 ( .A1(n22632), .A2(n14945), .B1(n14944), .B2(n22636), .ZN(
        n14937) );
  AOI21_X1 U16864 ( .B1(n22803), .B2(n22637), .A(n14937), .ZN(n14938) );
  OAI211_X1 U16865 ( .C1(n22640), .C2(n17833), .A(n14939), .B(n14938), .ZN(
        P1_U3090) );
  NAND2_X1 U16866 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14942) );
  OAI22_X1 U16867 ( .A1(n22659), .A2(n14945), .B1(n14944), .B2(n22663), .ZN(
        n14940) );
  AOI21_X1 U16868 ( .B1(n22803), .B2(n22664), .A(n14940), .ZN(n14941) );
  OAI211_X1 U16869 ( .C1(n22667), .C2(n17833), .A(n14942), .B(n14941), .ZN(
        P1_U3091) );
  NAND2_X1 U16870 ( .A1(n14943), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14948) );
  OAI22_X1 U16871 ( .A1(n22572), .A2(n14945), .B1(n14944), .B2(n22581), .ZN(
        n14946) );
  AOI21_X1 U16872 ( .B1(n22803), .B2(n22598), .A(n14946), .ZN(n14947) );
  OAI211_X1 U16873 ( .C1(n22601), .C2(n17833), .A(n14948), .B(n14947), .ZN(
        P1_U3089) );
  XOR2_X1 U16874 ( .A(n14950), .B(n14949), .Z(n22136) );
  INV_X1 U16875 ( .A(n22136), .ZN(n14952) );
  AOI22_X1 U16876 ( .A1(n16241), .A2(n22410), .B1(P1_EAX_REG_4__SCAN_IN), .B2(
        n16240), .ZN(n14951) );
  OAI21_X1 U16877 ( .B1(n14952), .B2(n16243), .A(n14951), .ZN(P1_U2900) );
  NOR3_X1 U16878 ( .A1(n22586), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14956) );
  NAND2_X1 U16879 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n22555), .ZN(n14954) );
  AND2_X1 U16880 ( .A1(n16564), .A2(n14673), .ZN(n22556) );
  INV_X1 U16881 ( .A(n14956), .ZN(n15129) );
  NOR2_X1 U16882 ( .A1(n22571), .A2(n15129), .ZN(n15008) );
  AOI21_X1 U16883 ( .B1(n22556), .B2(n14953), .A(n15008), .ZN(n14958) );
  NAND3_X1 U16884 ( .A1(n14954), .A2(n14958), .A3(n22563), .ZN(n14955) );
  OAI211_X1 U16885 ( .C1(n22563), .C2(n14956), .A(n14955), .B(n22613), .ZN(
        n15007) );
  AOI22_X1 U16886 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22637), .ZN(n14960) );
  OAI22_X1 U16887 ( .A1(n14958), .A2(n22607), .B1(n15129), .B2(n22605), .ZN(
        n15009) );
  AOI22_X1 U16888 ( .A1(n15009), .A2(n22642), .B1(n11263), .B2(n15008), .ZN(
        n14959) );
  OAI211_X1 U16889 ( .C1(n22640), .C2(n22540), .A(n14960), .B(n14959), .ZN(
        P1_U3106) );
  AOI22_X1 U16890 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22772), .ZN(n14962) );
  AOI22_X1 U16891 ( .A1(n15009), .A2(n22777), .B1(n11123), .B2(n15008), .ZN(
        n14961) );
  OAI211_X1 U16892 ( .C1(n22775), .C2(n22540), .A(n14962), .B(n14961), .ZN(
        P1_U3111) );
  AOI22_X1 U16893 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22718), .ZN(n14964) );
  AOI22_X1 U16894 ( .A1(n15009), .A2(n22723), .B1(n22722), .B2(n15008), .ZN(
        n14963) );
  OAI211_X1 U16895 ( .C1(n22721), .C2(n22540), .A(n14964), .B(n14963), .ZN(
        P1_U3109) );
  AOI22_X1 U16896 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22745), .ZN(n14966) );
  AOI22_X1 U16897 ( .A1(n15009), .A2(n22750), .B1(n11122), .B2(n15008), .ZN(
        n14965) );
  OAI211_X1 U16898 ( .C1(n22748), .C2(n22540), .A(n14966), .B(n14965), .ZN(
        P1_U3110) );
  AOI22_X1 U16899 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22691), .ZN(n14968) );
  AOI22_X1 U16900 ( .A1(n15009), .A2(n22696), .B1(n22695), .B2(n15008), .ZN(
        n14967) );
  OAI211_X1 U16901 ( .C1(n22694), .C2(n22540), .A(n14968), .B(n14967), .ZN(
        P1_U3108) );
  AOI22_X1 U16902 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n15007), .B1(
        n15130), .B2(n22833), .ZN(n14970) );
  AOI22_X1 U16903 ( .A1(n15009), .A2(n22841), .B1(n22839), .B2(n15008), .ZN(
        n14969) );
  OAI211_X1 U16904 ( .C1(n22838), .C2(n22540), .A(n14970), .B(n14969), .ZN(
        P1_U3112) );
  NAND2_X1 U16905 ( .A1(n19941), .A2(n17896), .ZN(n14975) );
  INV_X1 U16906 ( .A(n14890), .ZN(n14971) );
  OR2_X1 U16907 ( .A1(n14972), .A2(n14971), .ZN(n14974) );
  INV_X1 U16908 ( .A(n15516), .ZN(n14973) );
  NAND2_X1 U16909 ( .A1(n14974), .A2(n14973), .ZN(n15346) );
  INV_X1 U16910 ( .A(n15346), .ZN(n15402) );
  AOI21_X1 U16911 ( .B1(n14976), .B2(n14975), .A(n15402), .ZN(n20067) );
  XNOR2_X1 U16912 ( .A(n20067), .B(n20066), .ZN(n14979) );
  INV_X1 U16913 ( .A(n20124), .ZN(n20112) );
  AOI22_X1 U16914 ( .A1(n20064), .A2(n20112), .B1(n20111), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n14978) );
  NAND2_X1 U16915 ( .A1(n20117), .A2(n15402), .ZN(n14977) );
  OAI211_X1 U16916 ( .C1(n14979), .C2(n20065), .A(n14978), .B(n14977), .ZN(
        P2_U2915) );
  OAI21_X1 U16917 ( .B1(n14981), .B2(n14980), .A(n15015), .ZN(n19064) );
  NOR2_X1 U16918 ( .A1(n14905), .A2(n14982), .ZN(n14985) );
  OR2_X1 U16919 ( .A1(n14905), .A2(n14983), .ZN(n15013) );
  OAI211_X1 U16920 ( .C1(n14985), .C2(n14984), .A(n16724), .B(n15013), .ZN(
        n14987) );
  NAND2_X1 U16921 ( .A1(n15538), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n14986) );
  OAI211_X1 U16922 ( .C1(n19064), .C2(n15538), .A(n14987), .B(n14986), .ZN(
        P2_U2877) );
  OAI21_X1 U16923 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n21987) );
  INV_X1 U16924 ( .A(n15199), .ZN(n14993) );
  AOI22_X1 U16925 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n14991) );
  OAI21_X1 U16926 ( .B1(n20634), .B2(n15186), .A(n14991), .ZN(n14992) );
  AOI21_X1 U16927 ( .B1(n14993), .B2(n20614), .A(n14992), .ZN(n14994) );
  OAI21_X1 U16928 ( .B1(n22280), .B2(n21987), .A(n14994), .ZN(P1_U2996) );
  OAI21_X1 U16929 ( .B1(n14997), .B2(n14996), .A(n14995), .ZN(n21968) );
  AOI22_X1 U16930 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14998) );
  OAI21_X1 U16931 ( .B1(n20634), .B2(n22113), .A(n14998), .ZN(n14999) );
  AOI21_X1 U16932 ( .B1(n22119), .B2(n20614), .A(n14999), .ZN(n15000) );
  OAI21_X1 U16933 ( .B1(n22280), .B2(n21968), .A(n15000), .ZN(P1_U2997) );
  NOR2_X1 U16934 ( .A1(n11713), .A2(n15001), .ZN(n15002) );
  OR2_X1 U16935 ( .A1(n16807), .A2(n15002), .ZN(n17236) );
  OAI222_X1 U16936 ( .A1(n15004), .A2(n15003), .B1(n17236), .B2(n20071), .C1(
        n17950), .C2(n15640), .ZN(P2_U2904) );
  AOI22_X1 U16937 ( .A1(n22809), .A2(n22616), .B1(n15007), .B2(
        P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15006) );
  AOI22_X1 U16938 ( .A1(n15009), .A2(n22609), .B1(n22608), .B2(n15008), .ZN(
        n15005) );
  OAI211_X1 U16939 ( .C1(n22619), .C2(n17834), .A(n15006), .B(n15005), .ZN(
        P1_U3105) );
  AOI22_X1 U16940 ( .A1(n22809), .A2(n22670), .B1(n15007), .B2(
        P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U16941 ( .A1(n15009), .A2(n22669), .B1(n22668), .B2(n15008), .ZN(
        n15010) );
  OAI211_X1 U16942 ( .C1(n22673), .C2(n17834), .A(n15011), .B(n15010), .ZN(
        P1_U3107) );
  XNOR2_X1 U16943 ( .A(n15013), .B(n15012), .ZN(n15019) );
  NAND2_X1 U16944 ( .A1(n15538), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n15018) );
  INV_X1 U16945 ( .A(n15014), .ZN(n15021) );
  AOI21_X1 U16946 ( .B1(n15016), .B2(n15015), .A(n15014), .ZN(n19069) );
  NAND2_X1 U16947 ( .A1(n19069), .A2(n16700), .ZN(n15017) );
  OAI211_X1 U16948 ( .C1(n15019), .C2(n16732), .A(n15018), .B(n15017), .ZN(
        P2_U2876) );
  AND2_X1 U16949 ( .A1(n15021), .A2(n15020), .ZN(n15022) );
  NOR2_X1 U16950 ( .A1(n15204), .A2(n15022), .ZN(n17001) );
  INV_X1 U16951 ( .A(n17001), .ZN(n17275) );
  OAI211_X1 U16952 ( .C1(n15025), .C2(n15024), .A(n15023), .B(n16724), .ZN(
        n15027) );
  NAND2_X1 U16953 ( .A1(n15538), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15026) );
  OAI211_X1 U16954 ( .C1(n17275), .C2(n15538), .A(n15027), .B(n15026), .ZN(
        P2_U2875) );
  NOR2_X1 U16955 ( .A1(n20634), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15028) );
  AOI211_X1 U16956 ( .C1(n20628), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15029), .B(n15028), .ZN(n15033) );
  NAND3_X1 U16957 ( .A1(n15031), .A2(n15030), .A3(n20595), .ZN(n15032) );
  OAI211_X1 U16958 ( .C1(n16097), .C2(n20630), .A(n15033), .B(n15032), .ZN(
        P1_U2998) );
  OR2_X1 U16959 ( .A1(n15035), .A2(n15036), .ZN(n15296) );
  INV_X1 U16960 ( .A(n15296), .ZN(n15034) );
  AOI21_X1 U16961 ( .B1(n15036), .B2(n15035), .A(n15034), .ZN(n22148) );
  INV_X1 U16962 ( .A(n22148), .ZN(n15162) );
  OAI222_X1 U16963 ( .A1(n15162), .A2(n16243), .B1(n22418), .B2(n16233), .C1(
        n16231), .C2(n13399), .ZN(P1_U2899) );
  AND2_X1 U16964 ( .A1(n19842), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n17884) );
  INV_X1 U16965 ( .A(n17884), .ZN(n17885) );
  NAND3_X1 U16966 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19826) );
  OAI21_X1 U16967 ( .B1(n19843), .B2(n17885), .A(n19826), .ZN(n15044) );
  OAI21_X1 U16968 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n19322), .ZN(n19319) );
  INV_X1 U16969 ( .A(n19319), .ZN(n19016) );
  NAND2_X1 U16970 ( .A1(n19975), .A2(n15039), .ZN(n19962) );
  INV_X1 U16971 ( .A(n15037), .ZN(n19992) );
  INV_X1 U16972 ( .A(n20008), .ZN(n20295) );
  OAI21_X1 U16973 ( .B1(n19992), .B2(n20295), .A(n20009), .ZN(n15042) );
  OAI21_X1 U16974 ( .B1(n12178), .B2(n19962), .A(n15042), .ZN(n15043) );
  NAND2_X1 U16975 ( .A1(n15044), .A2(n15043), .ZN(n20300) );
  INV_X1 U16976 ( .A(n12178), .ZN(n15045) );
  OAI21_X1 U16977 ( .B1(n15045), .B2(n20295), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15046) );
  OAI21_X1 U16978 ( .B1(n19826), .B2(n15037), .A(n15046), .ZN(n20296) );
  NOR2_X2 U16979 ( .A1(n15047), .A2(n20291), .ZN(n20286) );
  NOR2_X2 U16980 ( .A1(n15109), .A2(n20293), .ZN(n20283) );
  INV_X1 U16981 ( .A(n20283), .ZN(n15049) );
  AOI22_X1 U16982 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20297), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n20298), .ZN(n20280) );
  AOI22_X1 U16983 ( .A1(n20285), .A2(n20277), .B1(n20299), .B2(n20284), .ZN(
        n15048) );
  OAI21_X1 U16984 ( .B1(n15049), .B2(n20008), .A(n15048), .ZN(n15050) );
  AOI21_X1 U16985 ( .B1(n20296), .B2(n20286), .A(n15050), .ZN(n15051) );
  OAI21_X1 U16986 ( .B1(n20210), .B2(n15052), .A(n15051), .ZN(P2_U3169) );
  INV_X1 U16987 ( .A(n15053), .ZN(n15054) );
  NAND2_X1 U16988 ( .A1(n15054), .A2(n15395), .ZN(n15058) );
  AND4_X1 U16989 ( .A1(n15058), .A2(n15057), .A3(n15056), .A4(n15055), .ZN(
        n15530) );
  INV_X1 U16990 ( .A(n15075), .ZN(n15094) );
  NOR2_X1 U16991 ( .A1(n15101), .A2(n15059), .ZN(n15090) );
  NOR2_X1 U16992 ( .A1(n15089), .A2(n15085), .ZN(n15063) );
  NOR2_X1 U16993 ( .A1(n15090), .A2(n15063), .ZN(n15067) );
  INV_X1 U16994 ( .A(n15060), .ZN(n15087) );
  NAND2_X1 U16995 ( .A1(n15072), .A2(n15087), .ZN(n15084) );
  NOR2_X1 U16996 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15065) );
  INV_X1 U16997 ( .A(n15061), .ZN(n15062) );
  NOR2_X1 U16998 ( .A1(n14202), .A2(n15062), .ZN(n15086) );
  INV_X1 U16999 ( .A(n15063), .ZN(n15064) );
  OAI22_X1 U17000 ( .A1(n15084), .A2(n15065), .B1(n15086), .B2(n15064), .ZN(
        n15066) );
  AOI211_X1 U17001 ( .C1(n12098), .C2(n15094), .A(n15067), .B(n15066), .ZN(
        n17384) );
  NOR2_X1 U17002 ( .A1(n17384), .A2(n15530), .ZN(n15082) );
  NAND2_X1 U17003 ( .A1(n15068), .A2(n13022), .ZN(n15071) );
  AOI22_X1 U17004 ( .A1(n15072), .A2(n11741), .B1(n15069), .B2(n15071), .ZN(
        n15070) );
  OAI21_X1 U17005 ( .B1(n17372), .B2(n15075), .A(n15070), .ZN(n15578) );
  NAND2_X1 U17006 ( .A1(n15578), .A2(n19985), .ZN(n15078) );
  INV_X1 U17007 ( .A(n15071), .ZN(n15073) );
  INV_X1 U17008 ( .A(n15072), .ZN(n15088) );
  MUX2_X1 U17009 ( .A(n15073), .B(n15088), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15074) );
  OAI21_X1 U17010 ( .B1(n15076), .B2(n15075), .A(n15074), .ZN(n15529) );
  OAI22_X1 U17011 ( .A1(n15578), .A2(n19985), .B1(n19987), .B2(n15529), .ZN(
        n15077) );
  NAND2_X1 U17012 ( .A1(n15078), .A2(n15077), .ZN(n15081) );
  INV_X1 U17013 ( .A(n15081), .ZN(n15079) );
  AOI21_X1 U17014 ( .B1(n15530), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n15082), .ZN(n15119) );
  OAI21_X1 U17015 ( .B1(n15530), .B2(n15079), .A(n15119), .ZN(n15080) );
  OAI221_X1 U17016 ( .B1(n19871), .B2(n15082), .C1(n19871), .C2(n15081), .A(
        n15080), .ZN(n15095) );
  INV_X1 U17017 ( .A(n15089), .ZN(n15083) );
  OAI211_X1 U17018 ( .C1(n15086), .C2(n15085), .A(n15084), .B(n15083), .ZN(
        n15092) );
  OAI22_X1 U17019 ( .A1(n15090), .A2(n15089), .B1(n15088), .B2(n15087), .ZN(
        n15091) );
  MUX2_X1 U17020 ( .A(n15092), .B(n15091), .S(n11777), .Z(n15093) );
  AOI211_X1 U17021 ( .C1(n12116), .C2(n15094), .A(n12143), .B(n15093), .ZN(
        n17388) );
  MUX2_X1 U17022 ( .A(n17388), .B(n11777), .S(n15530), .Z(n15118) );
  OR2_X1 U17023 ( .A1(n15095), .A2(n15118), .ZN(n15096) );
  AOI221_X1 U17024 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15096), 
        .C1(n15095), .C2(n15118), .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n15121) );
  INV_X1 U17025 ( .A(n15097), .ZN(n15106) );
  NOR2_X1 U17026 ( .A1(n15100), .A2(n15098), .ZN(n15099) );
  AOI21_X1 U17027 ( .B1(n15101), .B2(n15100), .A(n15099), .ZN(n15105) );
  AOI22_X1 U17028 ( .A1(n15115), .A2(n15112), .B1(n15103), .B2(n15102), .ZN(
        n15104) );
  OAI211_X1 U17029 ( .C1(n19318), .C2(n15106), .A(n15105), .B(n15104), .ZN(
        n19334) );
  INV_X1 U17030 ( .A(n15107), .ZN(n15108) );
  AND2_X1 U17031 ( .A1(n15109), .A2(n15108), .ZN(n15110) );
  AND2_X1 U17032 ( .A1(n14042), .A2(n15110), .ZN(n19270) );
  NOR3_X1 U17033 ( .A1(n19334), .A2(n19270), .A3(n15111), .ZN(n15117) );
  INV_X1 U17034 ( .A(n15112), .ZN(n15114) );
  NOR4_X1 U17035 ( .A1(n15115), .A2(n15114), .A3(n15395), .A4(n15113), .ZN(
        n19333) );
  OAI21_X1 U17036 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n19333), .ZN(n15116) );
  OAI211_X1 U17037 ( .C1(n15119), .C2(n15118), .A(n15117), .B(n15116), .ZN(
        n15120) );
  AOI211_X1 U17038 ( .C1(n15530), .C2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n15121), .B(n15120), .ZN(n19324) );
  AND3_X1 U17039 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19324), .A3(n17416), 
        .ZN(n15125) );
  AND2_X1 U17040 ( .A1(n15395), .A2(n19841), .ZN(n15389) );
  NAND3_X1 U17041 ( .A1(n15122), .A2(n15109), .A3(n15389), .ZN(n15123) );
  OAI21_X1 U17042 ( .B1(n15125), .B2(n15124), .A(n15123), .ZN(n15126) );
  INV_X1 U17043 ( .A(n15126), .ZN(n19321) );
  OAI21_X1 U17044 ( .B1(n19321), .B2(n19322), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n15128) );
  NOR2_X1 U17045 ( .A1(n19322), .A2(n15127), .ZN(n17415) );
  INV_X1 U17046 ( .A(n17415), .ZN(n19330) );
  NAND2_X1 U17047 ( .A1(n15128), .A2(n19330), .ZN(P2_U3593) );
  NOR2_X1 U17048 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n15129), .ZN(
        n15137) );
  OAI21_X1 U17049 ( .B1(n15130), .B2(n15157), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n15131) );
  AOI21_X1 U17050 ( .B1(n22556), .B2(n14636), .A(n15137), .ZN(n15133) );
  NAND2_X1 U17051 ( .A1(n15131), .A2(n15133), .ZN(n15132) );
  AND2_X1 U17052 ( .A1(n15135), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n22569) );
  NAND2_X1 U17053 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n15140) );
  INV_X1 U17054 ( .A(n15133), .ZN(n15136) );
  INV_X1 U17055 ( .A(n16585), .ZN(n15134) );
  INV_X1 U17056 ( .A(n22542), .ZN(n16584) );
  NOR2_X1 U17057 ( .A1(n15134), .A2(n16584), .ZN(n22578) );
  NOR2_X1 U17058 ( .A1(n15135), .A2(n22605), .ZN(n22544) );
  AOI22_X1 U17059 ( .A1(n15136), .A2(n22563), .B1(n22578), .B2(n22544), .ZN(
        n17832) );
  INV_X1 U17060 ( .A(n15137), .ZN(n17831) );
  OAI22_X1 U17061 ( .A1(n17832), .A2(n22690), .B1(n17831), .B2(n22686), .ZN(
        n15138) );
  AOI21_X1 U17062 ( .B1(n15157), .B2(n22691), .A(n15138), .ZN(n15139) );
  OAI211_X1 U17063 ( .C1(n22694), .C2(n17834), .A(n15140), .B(n15139), .ZN(
        P1_U3100) );
  NAND2_X1 U17064 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n15143) );
  OAI22_X1 U17065 ( .A1(n17832), .A2(n22717), .B1(n17831), .B2(n22713), .ZN(
        n15141) );
  AOI21_X1 U17066 ( .B1(n15157), .B2(n22718), .A(n15141), .ZN(n15142) );
  OAI211_X1 U17067 ( .C1(n22721), .C2(n17834), .A(n15143), .B(n15142), .ZN(
        P1_U3101) );
  NAND2_X1 U17068 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n15146) );
  OAI22_X1 U17069 ( .A1(n17832), .A2(n22636), .B1(n17831), .B2(n22632), .ZN(
        n15144) );
  AOI21_X1 U17070 ( .B1(n15157), .B2(n22637), .A(n15144), .ZN(n15145) );
  OAI211_X1 U17071 ( .C1(n22640), .C2(n17834), .A(n15146), .B(n15145), .ZN(
        P1_U3098) );
  NAND2_X1 U17072 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n15149) );
  OAI22_X1 U17073 ( .A1(n17832), .A2(n22744), .B1(n17831), .B2(n22740), .ZN(
        n15147) );
  AOI21_X1 U17074 ( .B1(n15157), .B2(n22745), .A(n15147), .ZN(n15148) );
  OAI211_X1 U17075 ( .C1(n22748), .C2(n17834), .A(n15149), .B(n15148), .ZN(
        P1_U3102) );
  NAND2_X1 U17076 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n15152) );
  OAI22_X1 U17077 ( .A1(n17832), .A2(n22771), .B1(n17831), .B2(n22767), .ZN(
        n15150) );
  AOI21_X1 U17078 ( .B1(n15157), .B2(n22772), .A(n15150), .ZN(n15151) );
  OAI211_X1 U17079 ( .C1(n22775), .C2(n17834), .A(n15152), .B(n15151), .ZN(
        P1_U3103) );
  NAND2_X1 U17080 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n15155) );
  OAI22_X1 U17081 ( .A1(n17832), .A2(n22829), .B1(n17831), .B2(n22821), .ZN(
        n15153) );
  AOI21_X1 U17082 ( .B1(n15157), .B2(n22833), .A(n15153), .ZN(n15154) );
  OAI211_X1 U17083 ( .C1(n22838), .C2(n17834), .A(n15155), .B(n15154), .ZN(
        P1_U3104) );
  NAND2_X1 U17084 ( .A1(n17837), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n15159) );
  OAI22_X1 U17085 ( .A1(n17832), .A2(n22581), .B1(n17831), .B2(n22572), .ZN(
        n15156) );
  AOI21_X1 U17086 ( .B1(n15157), .B2(n22598), .A(n15156), .ZN(n15158) );
  OAI211_X1 U17087 ( .C1(n22601), .C2(n17834), .A(n15159), .B(n15158), .ZN(
        P1_U3097) );
  INV_X1 U17088 ( .A(n15160), .ZN(n20551) );
  OAI21_X1 U17089 ( .B1(n20569), .B2(n15161), .A(n20551), .ZN(n22145) );
  OAI222_X1 U17090 ( .A1(n22145), .A2(n16143), .B1(n20574), .B2(n14238), .C1(
        n15162), .C2(n16146), .ZN(P1_U2867) );
  NAND2_X1 U17091 ( .A1(n15164), .A2(n15163), .ZN(n15166) );
  NAND2_X1 U17092 ( .A1(n15167), .A2(n17473), .ZN(n17470) );
  NAND2_X1 U17093 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n22297), .ZN(n17469) );
  OAI22_X1 U17094 ( .A1(n15308), .A2(n17470), .B1(n17473), .B2(n17469), .ZN(
        n15168) );
  INV_X1 U17095 ( .A(n15170), .ZN(n15171) );
  NAND2_X1 U17096 ( .A1(n15171), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15173) );
  INV_X1 U17097 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15172) );
  XNOR2_X1 U17098 ( .A(n15173), .B(n15172), .ZN(n15846) );
  NOR2_X1 U17099 ( .A1(n15846), .A2(n15308), .ZN(n15174) );
  NOR2_X1 U17100 ( .A1(n15196), .A2(n15175), .ZN(n15176) );
  INV_X1 U17101 ( .A(n22147), .ZN(n15325) );
  OR2_X1 U17102 ( .A1(n15196), .A2(n15177), .ZN(n15188) );
  AND2_X1 U17103 ( .A1(n15178), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n15182) );
  NAND2_X1 U17104 ( .A1(n22325), .A2(n22590), .ZN(n15180) );
  NAND2_X1 U17105 ( .A1(n15182), .A2(n15180), .ZN(n15179) );
  INV_X1 U17106 ( .A(n15180), .ZN(n17462) );
  NAND2_X1 U17107 ( .A1(n15181), .A2(n17462), .ZN(n15187) );
  INV_X1 U17108 ( .A(n15182), .ZN(n15183) );
  NAND2_X1 U17109 ( .A1(n15187), .A2(n15183), .ZN(n15184) );
  NOR2_X2 U17110 ( .A1(n15188), .A2(n15184), .ZN(n22272) );
  AND2_X1 U17111 ( .A1(n15846), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15185) );
  INV_X1 U17112 ( .A(n15186), .ZN(n15190) );
  OAI221_X1 U17113 ( .B1(n22200), .B2(P1_REIP_REG_1__SCAN_IN), .C1(n22200), 
        .C2(P1_REIP_REG_2__SCAN_IN), .A(n16102), .ZN(n15189) );
  AOI22_X1 U17114 ( .A1(n22253), .A2(n15190), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n15189), .ZN(n15192) );
  NAND2_X1 U17115 ( .A1(n22263), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15191) );
  OAI211_X1 U17116 ( .C1(n22249), .C2(n17620), .A(n15192), .B(n15191), .ZN(
        n15194) );
  INV_X1 U17117 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n22124) );
  NOR4_X1 U17118 ( .A1(n22200), .A2(n14610), .A3(P1_REIP_REG_3__SCAN_IN), .A4(
        n22124), .ZN(n15193) );
  AOI211_X1 U17119 ( .C1(n21989), .C2(n22255), .A(n15194), .B(n15193), .ZN(
        n15198) );
  NOR2_X1 U17120 ( .A1(n15196), .A2(n15195), .ZN(n22131) );
  NAND2_X1 U17121 ( .A1(n16564), .A2(n22131), .ZN(n15197) );
  OAI211_X1 U17122 ( .C1(n15199), .C2(n15325), .A(n15198), .B(n15197), .ZN(
        P1_U2837) );
  INV_X1 U17123 ( .A(n15023), .ZN(n15202) );
  OAI211_X1 U17124 ( .C1(n15202), .C2(n15201), .A(n16724), .B(n15331), .ZN(
        n15207) );
  NOR2_X1 U17125 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  OR2_X1 U17126 ( .A1(n15329), .A2(n15205), .ZN(n19090) );
  INV_X1 U17127 ( .A(n19090), .ZN(n17261) );
  NAND2_X1 U17128 ( .A1(n17261), .A2(n16700), .ZN(n15206) );
  OAI211_X1 U17129 ( .C1(n16700), .C2(n11908), .A(n15207), .B(n15206), .ZN(
        P2_U2874) );
  NOR3_X1 U17130 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15216) );
  INV_X1 U17131 ( .A(n15216), .ZN(n22492) );
  INV_X1 U17132 ( .A(n22613), .ZN(n15212) );
  OR2_X1 U17133 ( .A1(n16564), .A2(n15208), .ZN(n22515) );
  NOR2_X1 U17134 ( .A1(n22571), .A2(n22492), .ZN(n15247) );
  INV_X1 U17135 ( .A(n15247), .ZN(n15209) );
  OAI21_X1 U17136 ( .B1(n22515), .B2(n15210), .A(n15209), .ZN(n15215) );
  AOI211_X1 U17137 ( .C1(n15214), .C2(P1_STATEBS16_REG_SCAN_IN), .A(n22607), 
        .B(n15215), .ZN(n15211) );
  INV_X1 U17138 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15222) );
  NAND2_X1 U17139 ( .A1(n15214), .A2(n11155), .ZN(n22490) );
  NAND2_X1 U17140 ( .A1(n15215), .A2(n22563), .ZN(n15218) );
  NAND2_X1 U17141 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15216), .ZN(n15217) );
  NAND2_X1 U17142 ( .A1(n15218), .A2(n15217), .ZN(n15248) );
  AOI22_X1 U17143 ( .A1(n15248), .A2(n22696), .B1(n22695), .B2(n15247), .ZN(
        n15219) );
  OAI21_X1 U17144 ( .B1(n22502), .B2(n22694), .A(n15219), .ZN(n15220) );
  AOI21_X1 U17145 ( .B1(n22783), .B2(n22691), .A(n15220), .ZN(n15221) );
  OAI21_X1 U17146 ( .B1(n15253), .B2(n15222), .A(n15221), .ZN(P1_U3044) );
  INV_X1 U17147 ( .A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15226) );
  AOI22_X1 U17148 ( .A1(n15248), .A2(n22777), .B1(n22776), .B2(n15247), .ZN(
        n15223) );
  OAI21_X1 U17149 ( .B1(n22502), .B2(n22775), .A(n15223), .ZN(n15224) );
  AOI21_X1 U17150 ( .B1(n22783), .B2(n22772), .A(n15224), .ZN(n15225) );
  OAI21_X1 U17151 ( .B1(n15253), .B2(n15226), .A(n15225), .ZN(P1_U3047) );
  INV_X1 U17152 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15230) );
  AOI22_X1 U17153 ( .A1(n15248), .A2(n22609), .B1(n22608), .B2(n15247), .ZN(
        n15227) );
  OAI21_X1 U17154 ( .B1(n22490), .B2(n22619), .A(n15227), .ZN(n15228) );
  AOI21_X1 U17155 ( .B1(n22789), .B2(n22616), .A(n15228), .ZN(n15229) );
  OAI21_X1 U17156 ( .B1(n15253), .B2(n15230), .A(n15229), .ZN(P1_U3041) );
  INV_X1 U17157 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15234) );
  AOI22_X1 U17158 ( .A1(n15248), .A2(n22750), .B1(n22749), .B2(n15247), .ZN(
        n15231) );
  OAI21_X1 U17159 ( .B1(n22502), .B2(n22748), .A(n15231), .ZN(n15232) );
  AOI21_X1 U17160 ( .B1(n22783), .B2(n22745), .A(n15232), .ZN(n15233) );
  OAI21_X1 U17161 ( .B1(n15253), .B2(n15234), .A(n15233), .ZN(P1_U3046) );
  INV_X1 U17162 ( .A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15238) );
  AOI22_X1 U17163 ( .A1(n15248), .A2(n22723), .B1(n22722), .B2(n15247), .ZN(
        n15235) );
  OAI21_X1 U17164 ( .B1(n22502), .B2(n22721), .A(n15235), .ZN(n15236) );
  AOI21_X1 U17165 ( .B1(n22783), .B2(n22718), .A(n15236), .ZN(n15237) );
  OAI21_X1 U17166 ( .B1(n15253), .B2(n15238), .A(n15237), .ZN(P1_U3045) );
  INV_X1 U17167 ( .A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15242) );
  AOI22_X1 U17168 ( .A1(n15248), .A2(n22841), .B1(n22839), .B2(n15247), .ZN(
        n15239) );
  OAI21_X1 U17169 ( .B1(n22502), .B2(n22838), .A(n15239), .ZN(n15240) );
  AOI21_X1 U17170 ( .B1(n22783), .B2(n22833), .A(n15240), .ZN(n15241) );
  OAI21_X1 U17171 ( .B1(n15253), .B2(n15242), .A(n15241), .ZN(P1_U3048) );
  INV_X1 U17172 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15246) );
  AOI22_X1 U17173 ( .A1(n15248), .A2(n22642), .B1(n22641), .B2(n15247), .ZN(
        n15243) );
  OAI21_X1 U17174 ( .B1(n22502), .B2(n22640), .A(n15243), .ZN(n15244) );
  AOI21_X1 U17175 ( .B1(n22783), .B2(n22637), .A(n15244), .ZN(n15245) );
  OAI21_X1 U17176 ( .B1(n15253), .B2(n15246), .A(n15245), .ZN(P1_U3042) );
  INV_X1 U17177 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n15252) );
  AOI22_X1 U17178 ( .A1(n15248), .A2(n22669), .B1(n22668), .B2(n15247), .ZN(
        n15249) );
  OAI21_X1 U17179 ( .B1(n22490), .B2(n22673), .A(n15249), .ZN(n15250) );
  AOI21_X1 U17180 ( .B1(n22789), .B2(n22670), .A(n15250), .ZN(n15251) );
  OAI21_X1 U17181 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(P1_U3043) );
  OR2_X1 U17182 ( .A1(n15256), .A2(n15255), .ZN(n15257) );
  AND2_X1 U17183 ( .A1(n15254), .A2(n15257), .ZN(n22171) );
  INV_X1 U17184 ( .A(n22171), .ZN(n15260) );
  NAND2_X1 U17185 ( .A1(n20549), .A2(n15258), .ZN(n15259) );
  AND2_X1 U17186 ( .A1(n15306), .A2(n15259), .ZN(n22017) );
  INV_X1 U17187 ( .A(n22017), .ZN(n22169) );
  OAI222_X1 U17188 ( .A1(n15260), .A2(n16146), .B1(n20574), .B2(n14246), .C1(
        n22169), .C2(n16143), .ZN(P1_U2865) );
  INV_X1 U17189 ( .A(n16181), .ZN(n22428) );
  OAI222_X1 U17190 ( .A1(n15260), .A2(n16243), .B1(n22428), .B2(n16233), .C1(
        n16231), .C2(n13411), .ZN(P1_U2897) );
  XNOR2_X1 U17191 ( .A(n15337), .B(n12070), .ZN(n15339) );
  XNOR2_X1 U17192 ( .A(n15339), .B(n15338), .ZN(n15282) );
  NOR2_X1 U17193 ( .A1(n15262), .A2(n15261), .ZN(n15278) );
  NOR2_X1 U17194 ( .A1(n15278), .A2(n19302), .ZN(n15272) );
  INV_X1 U17195 ( .A(n17353), .ZN(n15264) );
  NAND2_X1 U17196 ( .A1(n17361), .A2(n15264), .ZN(n15265) );
  OAI21_X1 U17197 ( .B1(n15266), .B2(n17352), .A(n15265), .ZN(n17344) );
  AOI21_X1 U17198 ( .B1(n17328), .B2(n15266), .A(n17378), .ZN(n17324) );
  OAI21_X1 U17199 ( .B1(n17379), .B2(n17362), .A(n17361), .ZN(n15267) );
  NAND3_X1 U17200 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17324), .A3(
        n15267), .ZN(n15343) );
  OAI21_X1 U17201 ( .B1(n17344), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n15343), .ZN(n15270) );
  NOR2_X1 U17202 ( .A1(n19294), .A2(n15268), .ZN(n15277) );
  AOI21_X1 U17203 ( .B1(n19298), .B2(n12116), .A(n15277), .ZN(n15269) );
  OAI211_X1 U17204 ( .C1(n17896), .C2(n17371), .A(n15270), .B(n15269), .ZN(
        n15271) );
  AOI21_X1 U17205 ( .B1(n15272), .B2(n15263), .A(n15271), .ZN(n15273) );
  OAI21_X1 U17206 ( .B1(n15282), .B2(n17351), .A(n15273), .ZN(P2_U3043) );
  INV_X1 U17207 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15422) );
  OAI21_X1 U17208 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n15274), .A(
        n15275), .ZN(n15419) );
  OAI22_X1 U17209 ( .A1(n15422), .A2(n17877), .B1(n17042), .B2(n15419), .ZN(
        n15276) );
  AOI211_X1 U17210 ( .C1(n17870), .C2(n12116), .A(n15277), .B(n15276), .ZN(
        n15281) );
  INV_X1 U17211 ( .A(n15278), .ZN(n15279) );
  NAND3_X1 U17212 ( .A1(n15279), .A2(n17843), .A3(n15263), .ZN(n15280) );
  OAI211_X1 U17213 ( .C1(n15282), .C2(n17853), .A(n15281), .B(n15280), .ZN(
        P2_U3011) );
  INV_X1 U17214 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n22436) );
  AOI22_X1 U17215 ( .A1(n15290), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n15283) );
  OAI21_X1 U17216 ( .B1(n22436), .B2(n15318), .A(n15283), .ZN(P1_U2912) );
  INV_X1 U17217 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n22420) );
  AOI22_X1 U17218 ( .A1(n15290), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15284) );
  OAI21_X1 U17219 ( .B1(n22420), .B2(n15318), .A(n15284), .ZN(P1_U2915) );
  INV_X1 U17220 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n22443) );
  AOI22_X1 U17221 ( .A1(n15290), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n15285) );
  OAI21_X1 U17222 ( .B1(n22443), .B2(n15318), .A(n15285), .ZN(P1_U2911) );
  INV_X1 U17223 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n22450) );
  AOI22_X1 U17224 ( .A1(n15290), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n15286) );
  OAI21_X1 U17225 ( .B1(n22450), .B2(n15318), .A(n15286), .ZN(P1_U2910) );
  INV_X1 U17226 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n22413) );
  AOI22_X1 U17227 ( .A1(n15290), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15287) );
  OAI21_X1 U17228 ( .B1(n22413), .B2(n15318), .A(n15287), .ZN(P1_U2916) );
  INV_X1 U17229 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n22458) );
  AOI22_X1 U17230 ( .A1(n15290), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15288) );
  OAI21_X1 U17231 ( .B1(n22458), .B2(n15318), .A(n15288), .ZN(P1_U2909) );
  INV_X1 U17232 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n22406) );
  AOI22_X1 U17233 ( .A1(n15290), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15289) );
  OAI21_X1 U17234 ( .B1(n22406), .B2(n15318), .A(n15289), .ZN(P1_U2917) );
  INV_X1 U17235 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n22425) );
  AOI22_X1 U17236 ( .A1(n15290), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U17237 ( .B1(n22425), .B2(n15318), .A(n15291), .ZN(P1_U2914) );
  INV_X1 U17238 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n22481) );
  AOI22_X1 U17239 ( .A1(n21945), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15292) );
  OAI21_X1 U17240 ( .B1(n22481), .B2(n15318), .A(n15292), .ZN(P1_U2906) );
  INV_X1 U17241 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n22472) );
  AOI22_X1 U17242 ( .A1(n21945), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15293) );
  OAI21_X1 U17243 ( .B1(n22472), .B2(n15318), .A(n15293), .ZN(P1_U2907) );
  INV_X1 U17244 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n22430) );
  AOI22_X1 U17245 ( .A1(n21945), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n15294) );
  OAI21_X1 U17246 ( .B1(n22430), .B2(n15318), .A(n15294), .ZN(P1_U2913) );
  INV_X1 U17247 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n22465) );
  AOI22_X1 U17248 ( .A1(n21945), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15295) );
  OAI21_X1 U17249 ( .B1(n22465), .B2(n15318), .A(n15295), .ZN(P1_U2908) );
  INV_X1 U17250 ( .A(n16187), .ZN(n22423) );
  XOR2_X1 U17251 ( .A(n15297), .B(n15296), .Z(n22159) );
  INV_X1 U17252 ( .A(n22159), .ZN(n15298) );
  OAI222_X1 U17253 ( .A1(n16231), .A2(n15299), .B1(n22423), .B2(n16233), .C1(
        n16243), .C2(n15298), .ZN(P1_U2898) );
  XOR2_X1 U17254 ( .A(n15300), .B(n15254), .Z(n15503) );
  INV_X1 U17255 ( .A(n15503), .ZN(n15351) );
  INV_X1 U17256 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n15301) );
  OR2_X1 U17257 ( .A1(n16158), .A2(n15301), .ZN(n15303) );
  NAND2_X1 U17258 ( .A1(n16158), .A2(DATAI_8_), .ZN(n15302) );
  NAND2_X1 U17259 ( .A1(n15303), .A2(n15302), .ZN(n22433) );
  AOI22_X1 U17260 ( .A1(n16241), .A2(n22433), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16240), .ZN(n15304) );
  OAI21_X1 U17261 ( .B1(n15351), .B2(n16243), .A(n15304), .ZN(P1_U2896) );
  NAND4_X1 U17262 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_4__SCAN_IN), .ZN(n22139)
         );
  INV_X1 U17263 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n22150) );
  NOR2_X1 U17264 ( .A1(n22139), .A2(n22150), .ZN(n22152) );
  NAND2_X1 U17265 ( .A1(n22152), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n22163) );
  INV_X1 U17266 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n22173) );
  NOR2_X1 U17267 ( .A1(n22163), .A2(n22173), .ZN(n15311) );
  NAND2_X1 U17268 ( .A1(n15311), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n22175) );
  AOI21_X1 U17269 ( .B1(n22214), .B2(n22175), .A(n22190), .ZN(n22186) );
  INV_X1 U17270 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n17753) );
  AND2_X1 U17271 ( .A1(n15306), .A2(n15305), .ZN(n15307) );
  NOR2_X1 U17272 ( .A1(n15357), .A2(n15307), .ZN(n22021) );
  AOI22_X1 U17273 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n22263), .B1(
        n22255), .B2(n22021), .ZN(n15310) );
  AND2_X1 U17274 ( .A1(n22559), .A2(n15308), .ZN(n15309) );
  NAND2_X1 U17275 ( .A1(n16102), .A2(n15309), .ZN(n22264) );
  OAI211_X1 U17276 ( .C1(n22186), .C2(n17753), .A(n15310), .B(n22264), .ZN(
        n15315) );
  AND3_X1 U17277 ( .A1(n22214), .A2(n22175), .A3(n15311), .ZN(n15314) );
  INV_X1 U17278 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15312) );
  OAI22_X1 U17279 ( .A1(n22249), .A2(n15312), .B1(n15501), .B2(n22267), .ZN(
        n15313) );
  NOR3_X1 U17280 ( .A1(n15315), .A2(n15314), .A3(n15313), .ZN(n15316) );
  OAI21_X1 U17281 ( .B1(n15351), .B2(n22268), .A(n15316), .ZN(P1_U2832) );
  INV_X1 U17282 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n22388) );
  AOI22_X1 U17283 ( .A1(n21945), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20474), .ZN(n15317) );
  OAI21_X1 U17284 ( .B1(n22388), .B2(n15318), .A(n15317), .ZN(P1_U2920) );
  NAND2_X1 U17285 ( .A1(n22273), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n15321) );
  NAND2_X1 U17286 ( .A1(n22246), .A2(n22267), .ZN(n15319) );
  AOI22_X1 U17287 ( .A1(n22272), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n15319), .B2(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15320) );
  OAI211_X1 U17288 ( .C1(n22278), .C2(n15322), .A(n15321), .B(n15320), .ZN(
        n15323) );
  AOI21_X1 U17289 ( .B1(n17438), .B2(n22131), .A(n15323), .ZN(n15324) );
  OAI21_X1 U17290 ( .B1(n15326), .B2(n15325), .A(n15324), .ZN(P1_U2840) );
  OR2_X1 U17291 ( .A1(n15329), .A2(n15328), .ZN(n15330) );
  NAND2_X1 U17292 ( .A1(n15327), .A2(n15330), .ZN(n16980) );
  INV_X1 U17293 ( .A(n15332), .ZN(n15333) );
  OAI211_X1 U17294 ( .C1(n15200), .C2(n15334), .A(n15333), .B(n16724), .ZN(
        n15336) );
  NAND2_X1 U17295 ( .A1(n15538), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15335) );
  OAI211_X1 U17296 ( .C1(n16980), .C2(n15538), .A(n15336), .B(n15335), .ZN(
        P2_U2873) );
  AOI22_X1 U17297 ( .A1(n15339), .A2(n15338), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15337), .ZN(n15341) );
  XNOR2_X1 U17298 ( .A(n15404), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n15340) );
  XNOR2_X1 U17299 ( .A(n15341), .B(n15340), .ZN(n17846) );
  INV_X1 U17300 ( .A(n17846), .ZN(n15350) );
  XNOR2_X1 U17301 ( .A(n15342), .B(n15521), .ZN(n17844) );
  NAND2_X1 U17302 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17344), .ZN(
        n15520) );
  INV_X1 U17303 ( .A(n17324), .ZN(n15344) );
  OAI21_X1 U17304 ( .B1(n19279), .B2(n15344), .A(n15343), .ZN(n15515) );
  NAND2_X1 U17305 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19124), .ZN(n15345) );
  OAI221_X1 U17306 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15520), .C1(
        n15521), .C2(n15515), .A(n15345), .ZN(n15348) );
  OAI22_X1 U17307 ( .A1(n15382), .A2(n14207), .B1(n17371), .B2(n15346), .ZN(
        n15347) );
  AOI211_X1 U17308 ( .C1(n17844), .C2(n17377), .A(n15348), .B(n15347), .ZN(
        n15349) );
  OAI21_X1 U17309 ( .B1(n15350), .B2(n17351), .A(n15349), .ZN(P2_U3042) );
  INV_X1 U17310 ( .A(n22021), .ZN(n15352) );
  OAI222_X1 U17311 ( .A1(n15352), .A2(n16143), .B1(n20574), .B2(n15312), .C1(
        n16146), .C2(n15351), .ZN(P1_U2864) );
  AND2_X1 U17312 ( .A1(n15354), .A2(n15353), .ZN(n15355) );
  OR2_X1 U17313 ( .A1(n15355), .A2(n11160), .ZN(n22181) );
  INV_X1 U17314 ( .A(n15356), .ZN(n15359) );
  INV_X1 U17315 ( .A(n15357), .ZN(n15358) );
  AOI21_X1 U17316 ( .B1(n15359), .B2(n15358), .A(n20560), .ZN(n22179) );
  AOI22_X1 U17317 ( .A1(n22179), .A2(n20572), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n16119), .ZN(n15360) );
  OAI21_X1 U17318 ( .B1(n22181), .B2(n16146), .A(n15360), .ZN(P1_U2863) );
  INV_X1 U17319 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20653) );
  OR2_X1 U17320 ( .A1(n16158), .A2(n20653), .ZN(n15362) );
  NAND2_X1 U17321 ( .A1(n16158), .A2(DATAI_9_), .ZN(n15361) );
  NAND2_X1 U17322 ( .A1(n15362), .A2(n15361), .ZN(n22440) );
  AOI22_X1 U17323 ( .A1(n16241), .A2(n22440), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16240), .ZN(n15363) );
  OAI21_X1 U17324 ( .B1(n22181), .B2(n16243), .A(n15363), .ZN(P1_U2895) );
  OAI211_X1 U17325 ( .C1(n15332), .C2(n15365), .A(n15364), .B(n16724), .ZN(
        n15369) );
  INV_X1 U17326 ( .A(n15327), .ZN(n15367) );
  OAI21_X1 U17327 ( .B1(n15367), .B2(n11529), .A(n15539), .ZN(n16970) );
  INV_X1 U17328 ( .A(n16970), .ZN(n17234) );
  NAND2_X1 U17329 ( .A1(n17234), .A2(n16700), .ZN(n15368) );
  OAI211_X1 U17330 ( .C1(n16700), .C2(n12483), .A(n15369), .B(n15368), .ZN(
        P2_U2872) );
  NOR2_X1 U17331 ( .A1(n11160), .A2(n15372), .ZN(n15373) );
  OR2_X1 U17332 ( .A1(n15371), .A2(n15373), .ZN(n22195) );
  MUX2_X1 U17333 ( .A(BUF1_REG_10__SCAN_IN), .B(DATAI_10_), .S(n16158), .Z(
        n22447) );
  AOI22_X1 U17334 ( .A1(n16241), .A2(n22447), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16240), .ZN(n15374) );
  OAI21_X1 U17335 ( .B1(n22195), .B2(n16243), .A(n15374), .ZN(P1_U2894) );
  AOI21_X1 U17336 ( .B1(n17849), .B2(n15275), .A(n15375), .ZN(n17842) );
  INV_X1 U17337 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15871) );
  XNOR2_X1 U17338 ( .A(n15377), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15880) );
  AOI21_X1 U17339 ( .B1(n15895), .B2(n17049), .A(n15274), .ZN(n15892) );
  AOI22_X1 U17340 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19322), .ZN(n15378) );
  INV_X1 U17341 ( .A(n15378), .ZN(n15583) );
  OAI22_X1 U17342 ( .A1(n19322), .A2(n17052), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15577) );
  OR2_X1 U17343 ( .A1(n15583), .A2(n15577), .ZN(n15408) );
  NOR2_X1 U17344 ( .A1(n15892), .A2(n15408), .ZN(n15418) );
  NAND2_X1 U17345 ( .A1(n15418), .A2(n15419), .ZN(n15438) );
  AND2_X1 U17346 ( .A1(n15795), .A2(n15438), .ZN(n15381) );
  NOR4_X1 U17347 ( .A1(n17416), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n15379)
         );
  INV_X1 U17348 ( .A(n19244), .ZN(n19316) );
  AOI21_X1 U17349 ( .B1(n17842), .B2(n15381), .A(n19316), .ZN(n15380) );
  OAI21_X1 U17350 ( .B1(n17842), .B2(n15381), .A(n15380), .ZN(n15407) );
  INV_X1 U17351 ( .A(n15382), .ZN(n17845) );
  NOR2_X1 U17352 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n22359), .ZN(n15394) );
  NAND2_X1 U17353 ( .A1(n15383), .A2(n15394), .ZN(n15384) );
  INV_X1 U17354 ( .A(n19012), .ZN(n15388) );
  INV_X1 U17355 ( .A(n15394), .ZN(n15385) );
  NAND2_X1 U17356 ( .A1(n15385), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n15386) );
  NOR2_X1 U17357 ( .A1(n12031), .A2(n15386), .ZN(n15387) );
  NAND2_X1 U17358 ( .A1(n15390), .A2(n15389), .ZN(n15391) );
  NOR2_X2 U17359 ( .A1(n19012), .A2(n15391), .ZN(n19241) );
  NAND2_X1 U17360 ( .A1(n19903), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19313) );
  OR3_X1 U17361 ( .A1(n19975), .A2(n19313), .A3(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n19328) );
  INV_X1 U17362 ( .A(n19328), .ZN(n15392) );
  NOR3_X1 U17363 ( .A1(n15392), .A2(n19124), .A3(n19244), .ZN(n15393) );
  NOR2_X1 U17364 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n15394), .ZN(n15397) );
  NAND2_X1 U17365 ( .A1(n15395), .A2(n19841), .ZN(n15396) );
  OAI21_X1 U17366 ( .B1(n15109), .B2(n15397), .A(n15396), .ZN(n15398) );
  AOI22_X1 U17367 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19237), .ZN(n15400) );
  OAI211_X1 U17368 ( .C1(n17849), .C2(n19208), .A(n19294), .B(n15400), .ZN(
        n15401) );
  AOI21_X1 U17369 ( .B1(n19241), .B2(n15402), .A(n15401), .ZN(n15403) );
  OAI21_X1 U17370 ( .B1(n15404), .B2(n19215), .A(n15403), .ZN(n15405) );
  AOI21_X1 U17371 ( .B1(n17845), .B2(n19227), .A(n15405), .ZN(n15406) );
  OAI211_X1 U17372 ( .C1(n15591), .C2(n20066), .A(n15407), .B(n15406), .ZN(
        P2_U2851) );
  NAND2_X1 U17373 ( .A1(n15795), .A2(n15408), .ZN(n15576) );
  XNOR2_X1 U17374 ( .A(n15892), .B(n15576), .ZN(n15409) );
  NAND2_X1 U17375 ( .A1(n15409), .A2(n19244), .ZN(n15417) );
  OAI22_X1 U17376 ( .A1(n15410), .A2(n19210), .B1(n12060), .B2(n19256), .ZN(
        n15412) );
  NOR2_X1 U17377 ( .A1(n19208), .A2(n15895), .ZN(n15411) );
  AOI211_X1 U17378 ( .C1(n19261), .C2(n15413), .A(n15412), .B(n15411), .ZN(
        n15414) );
  OAI21_X1 U17379 ( .B1(n17886), .B2(n19268), .A(n15414), .ZN(n15415) );
  AOI21_X1 U17380 ( .B1(n12095), .B2(n19251), .A(n15415), .ZN(n15416) );
  OAI211_X1 U17381 ( .C1(n19940), .C2(n15591), .A(n15417), .B(n15416), .ZN(
        P2_U2853) );
  NOR2_X1 U17382 ( .A1(n15794), .A2(n15418), .ZN(n15420) );
  XNOR2_X1 U17383 ( .A(n15420), .B(n15419), .ZN(n15421) );
  NAND2_X1 U17384 ( .A1(n15421), .A2(n19244), .ZN(n15429) );
  OAI22_X1 U17385 ( .A1(n12071), .A2(n19210), .B1(n15268), .B2(n19256), .ZN(
        n15423) );
  AOI21_X1 U17386 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n19239), .A(
        n15423), .ZN(n15424) );
  OAI21_X1 U17387 ( .B1(n19215), .B2(n15425), .A(n15424), .ZN(n15427) );
  NOR2_X1 U17388 ( .A1(n17896), .A2(n19268), .ZN(n15426) );
  AOI211_X1 U17389 ( .C1(n19227), .C2(n12116), .A(n15427), .B(n15426), .ZN(
        n15428) );
  OAI211_X1 U17390 ( .C1(n19941), .C2(n15591), .A(n15429), .B(n15428), .ZN(
        P2_U2852) );
  AND2_X1 U17391 ( .A1(n15442), .A2(n16999), .ZN(n15430) );
  NOR2_X1 U17392 ( .A1(n15468), .A2(n15430), .ZN(n15467) );
  INV_X1 U17393 ( .A(n15467), .ZN(n17003) );
  OR2_X1 U17394 ( .A1(n15431), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15433) );
  NAND2_X1 U17395 ( .A1(n15433), .A2(n15432), .ZN(n19058) );
  INV_X1 U17396 ( .A(n19058), .ZN(n15440) );
  AOI21_X1 U17397 ( .B1(n17878), .B2(n15434), .A(n15435), .ZN(n17861) );
  AOI21_X1 U17398 ( .B1(n17860), .B2(n15436), .A(n15437), .ZN(n19051) );
  NOR2_X1 U17399 ( .A1(n17842), .A2(n15438), .ZN(n19037) );
  OAI21_X1 U17400 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n15375), .A(
        n15436), .ZN(n19038) );
  NAND2_X1 U17401 ( .A1(n19037), .A2(n19038), .ZN(n19049) );
  NOR2_X1 U17402 ( .A1(n19051), .A2(n19049), .ZN(n15488) );
  OAI21_X1 U17403 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n15437), .A(
        n15434), .ZN(n17041) );
  NAND2_X1 U17404 ( .A1(n15488), .A2(n17041), .ZN(n15478) );
  NOR2_X1 U17405 ( .A1(n17861), .A2(n15478), .ZN(n15453) );
  NOR2_X1 U17406 ( .A1(n15435), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15439) );
  OR2_X1 U17407 ( .A1(n15431), .A2(n15439), .ZN(n17032) );
  NAND2_X1 U17408 ( .A1(n15453), .A2(n17032), .ZN(n19057) );
  NOR2_X1 U17409 ( .A1(n15440), .A2(n19057), .ZN(n19080) );
  NAND2_X1 U17410 ( .A1(n15432), .A2(n19072), .ZN(n15441) );
  NAND2_X1 U17411 ( .A1(n15442), .A2(n15441), .ZN(n19083) );
  NAND2_X1 U17412 ( .A1(n19080), .A2(n19083), .ZN(n19079) );
  NAND2_X1 U17413 ( .A1(n15795), .A2(n19079), .ZN(n15443) );
  XOR2_X1 U17414 ( .A(n17003), .B(n15443), .Z(n15444) );
  NAND2_X1 U17415 ( .A1(n15444), .A2(n19244), .ZN(n15451) );
  XNOR2_X1 U17416 ( .A(n15446), .B(n15445), .ZN(n19811) );
  OAI22_X1 U17417 ( .A1(n16999), .A2(n19208), .B1(n17963), .B2(n19256), .ZN(
        n15447) );
  AOI211_X1 U17418 ( .C1(n11121), .C2(P2_EBX_REG_12__SCAN_IN), .A(n19124), .B(
        n15447), .ZN(n15448) );
  OAI21_X1 U17419 ( .B1(n19268), .B2(n19811), .A(n15448), .ZN(n15449) );
  AOI21_X1 U17420 ( .B1(n17001), .B2(n19227), .A(n15449), .ZN(n15450) );
  OAI211_X1 U17421 ( .C1(n19215), .C2(n15452), .A(n15451), .B(n15450), .ZN(
        P2_U2843) );
  NOR2_X1 U17422 ( .A1(n15794), .A2(n15453), .ZN(n15454) );
  XNOR2_X1 U17423 ( .A(n17032), .B(n15454), .ZN(n15455) );
  NAND2_X1 U17424 ( .A1(n15455), .A2(n19244), .ZN(n15462) );
  OAI21_X1 U17425 ( .B1(n14754), .B2(n15457), .A(n15456), .ZN(n19817) );
  INV_X1 U17426 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17031) );
  OAI22_X1 U17427 ( .A1(n17031), .A2(n19208), .B1(n17961), .B2(n19256), .ZN(
        n15458) );
  AOI211_X1 U17428 ( .C1(n11121), .C2(P2_EBX_REG_9__SCAN_IN), .A(n19124), .B(
        n15458), .ZN(n15459) );
  OAI21_X1 U17429 ( .B1(n19268), .B2(n19817), .A(n15459), .ZN(n15460) );
  AOI21_X1 U17430 ( .B1(n19251), .B2(n17311), .A(n15460), .ZN(n15461) );
  OAI211_X1 U17431 ( .C1(n19215), .C2(n15463), .A(n15462), .B(n15461), .ZN(
        P2_U2846) );
  AOI21_X1 U17432 ( .B1(n16966), .B2(n11225), .A(n15464), .ZN(n16968) );
  OR2_X1 U17433 ( .A1(n15465), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15466) );
  NAND2_X1 U17434 ( .A1(n15466), .A2(n11225), .ZN(n15545) );
  INV_X1 U17435 ( .A(n15545), .ZN(n16977) );
  NOR2_X1 U17436 ( .A1(n15467), .A2(n19079), .ZN(n19094) );
  NOR2_X1 U17437 ( .A1(n15468), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15469) );
  OR2_X1 U17438 ( .A1(n15465), .A2(n15469), .ZN(n19093) );
  NAND2_X1 U17439 ( .A1(n19094), .A2(n19093), .ZN(n15546) );
  NOR2_X1 U17440 ( .A1(n16977), .A2(n15546), .ZN(n15790) );
  NOR2_X1 U17441 ( .A1(n15794), .A2(n15790), .ZN(n15470) );
  XOR2_X1 U17442 ( .A(n16968), .B(n15470), .Z(n15471) );
  NAND2_X1 U17443 ( .A1(n15471), .A2(n19244), .ZN(n15476) );
  OAI22_X1 U17444 ( .A1(n16966), .A2(n19208), .B1(n17965), .B2(n19256), .ZN(
        n15472) );
  AOI211_X1 U17445 ( .C1(n11121), .C2(P2_EBX_REG_15__SCAN_IN), .A(n19124), .B(
        n15472), .ZN(n15473) );
  OAI21_X1 U17446 ( .B1(n17236), .B2(n19268), .A(n15473), .ZN(n15474) );
  AOI21_X1 U17447 ( .B1(n17234), .B2(n19227), .A(n15474), .ZN(n15475) );
  OAI211_X1 U17448 ( .C1(n19215), .C2(n15477), .A(n15476), .B(n15475), .ZN(
        P2_U2840) );
  INV_X1 U17449 ( .A(n19227), .ZN(n19166) );
  NAND2_X1 U17450 ( .A1(n15795), .A2(n15478), .ZN(n15479) );
  XNOR2_X1 U17451 ( .A(n17861), .B(n15479), .ZN(n15481) );
  INV_X1 U17452 ( .A(n15480), .ZN(n19291) );
  AOI22_X1 U17453 ( .A1(n19244), .A2(n15481), .B1(n19241), .B2(n19291), .ZN(
        n15486) );
  AOI22_X1 U17454 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n19261), .B2(n15482), .ZN(n15483) );
  OAI21_X1 U17455 ( .B1(n14116), .B2(n19256), .A(n15483), .ZN(n15484) );
  AOI211_X1 U17456 ( .C1(n11121), .C2(P2_EBX_REG_8__SCAN_IN), .A(n19124), .B(
        n15484), .ZN(n15485) );
  OAI211_X1 U17457 ( .C1(n19166), .C2(n15487), .A(n15486), .B(n15485), .ZN(
        P2_U2847) );
  NOR2_X1 U17458 ( .A1(n15794), .A2(n15488), .ZN(n15489) );
  XNOR2_X1 U17459 ( .A(n15489), .B(n17041), .ZN(n15491) );
  AOI22_X1 U17460 ( .A1(n19244), .A2(n15491), .B1(n19241), .B2(n15490), .ZN(
        n15496) );
  AOI22_X1 U17461 ( .A1(n15492), .A2(n19261), .B1(n19239), .B2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n15493) );
  OAI211_X1 U17462 ( .C1(n12451), .C2(n19210), .A(n15493), .B(n19294), .ZN(
        n15494) );
  AOI21_X1 U17463 ( .B1(P2_REIP_REG_7__SCAN_IN), .B2(n19237), .A(n15494), .ZN(
        n15495) );
  OAI211_X1 U17464 ( .C1(n19166), .C2(n17331), .A(n15496), .B(n15495), .ZN(
        P2_U2848) );
  OAI21_X1 U17465 ( .B1(n15499), .B2(n15498), .A(n15497), .ZN(n22022) );
  NAND2_X1 U17466 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15500) );
  NAND2_X1 U17467 ( .A1(n22108), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n22019) );
  OAI211_X1 U17468 ( .C1(n20634), .C2(n15501), .A(n15500), .B(n22019), .ZN(
        n15502) );
  AOI21_X1 U17469 ( .B1(n15503), .B2(n20614), .A(n15502), .ZN(n15504) );
  OAI21_X1 U17470 ( .B1(n22022), .B2(n22280), .A(n15504), .ZN(P1_U2991) );
  XNOR2_X1 U17471 ( .A(n15505), .B(n15506), .ZN(n15528) );
  NAND2_X1 U17472 ( .A1(n15508), .A2(n15522), .ZN(n15513) );
  NAND3_X1 U17473 ( .A1(n15514), .A2(n17843), .A3(n15513), .ZN(n15512) );
  NAND2_X1 U17474 ( .A1(n19124), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n15518) );
  INV_X1 U17475 ( .A(n15518), .ZN(n15510) );
  OAI22_X1 U17476 ( .A1(n11561), .A2(n17877), .B1(n17042), .B2(n19038), .ZN(
        n15509) );
  AOI211_X1 U17477 ( .C1(n17870), .C2(n19040), .A(n15510), .B(n15509), .ZN(
        n15511) );
  OAI211_X1 U17478 ( .C1(n15528), .C2(n17853), .A(n15512), .B(n15511), .ZN(
        P2_U3009) );
  NAND3_X1 U17479 ( .A1(n15514), .A2(n17377), .A3(n15513), .ZN(n15527) );
  INV_X1 U17480 ( .A(n15515), .ZN(n15525) );
  XNOR2_X1 U17481 ( .A(n15517), .B(n15516), .ZN(n20070) );
  NAND2_X1 U17482 ( .A1(n19298), .A2(n19040), .ZN(n15519) );
  OAI211_X1 U17483 ( .C1(n17371), .C2(n20070), .A(n15519), .B(n15518), .ZN(
        n15524) );
  AOI221_X1 U17484 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n15522), .C2(n15521), .A(
        n15520), .ZN(n15523) );
  AOI211_X1 U17485 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15525), .A(
        n15524), .B(n15523), .ZN(n15526) );
  OAI211_X1 U17486 ( .C1(n15528), .C2(n17351), .A(n15527), .B(n15526), .ZN(
        P2_U3041) );
  INV_X1 U17487 ( .A(n19311), .ZN(n19271) );
  AOI22_X1 U17488 ( .A1(n15794), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n15583), .B2(n15795), .ZN(n15575) );
  AOI222_X1 U17489 ( .A1(n15529), .A2(n19271), .B1(n19836), .B2(n19320), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15575), .ZN(n15535) );
  OR2_X1 U17490 ( .A1(n15530), .A2(n19332), .ZN(n15533) );
  OAI22_X1 U17491 ( .A1(n19330), .A2(n12377), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19975), .ZN(n15531) );
  INV_X1 U17492 ( .A(n15531), .ZN(n15532) );
  NAND2_X1 U17493 ( .A1(n15533), .A2(n15532), .ZN(n19274) );
  INV_X1 U17494 ( .A(n19274), .ZN(n15580) );
  NAND2_X1 U17495 ( .A1(n15580), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15534) );
  OAI21_X1 U17496 ( .B1(n15535), .B2(n15580), .A(n15534), .ZN(P2_U3601) );
  INV_X1 U17497 ( .A(n15364), .ZN(n15537) );
  OAI21_X1 U17498 ( .B1(n15537), .B2(n15536), .A(n15571), .ZN(n16804) );
  INV_X1 U17499 ( .A(n15539), .ZN(n15542) );
  INV_X1 U17500 ( .A(n15540), .ZN(n15541) );
  OAI21_X1 U17501 ( .B1(n15542), .B2(n15541), .A(n15568), .ZN(n19106) );
  NOR2_X1 U17502 ( .A1(n19106), .A2(n15538), .ZN(n15543) );
  AOI21_X1 U17503 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n15538), .A(n15543), .ZN(
        n15544) );
  OAI21_X1 U17504 ( .B1(n16804), .B2(n16732), .A(n15544), .ZN(P2_U2871) );
  AND2_X1 U17505 ( .A1(n19265), .A2(n15546), .ZN(n19092) );
  AOI22_X1 U17506 ( .A1(n15545), .A2(n19092), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19239), .ZN(n15556) );
  INV_X1 U17507 ( .A(n16980), .ZN(n17250) );
  INV_X1 U17508 ( .A(n15546), .ZN(n15547) );
  OAI211_X1 U17509 ( .C1(n15547), .C2(n15794), .A(n16977), .B(n19244), .ZN(
        n15548) );
  OAI211_X1 U17510 ( .C1(n15549), .C2(n19210), .A(n15548), .B(n19294), .ZN(
        n15554) );
  AND2_X1 U17511 ( .A1(n15551), .A2(n15550), .ZN(n15552) );
  OR2_X1 U17512 ( .A1(n11713), .A2(n15552), .ZN(n19808) );
  OAI22_X1 U17513 ( .A1(n19808), .A2(n19268), .B1(n17964), .B2(n19256), .ZN(
        n15553) );
  AOI211_X1 U17514 ( .C1(n17250), .C2(n19251), .A(n15554), .B(n15553), .ZN(
        n15555) );
  OAI211_X1 U17515 ( .C1(n15557), .C2(n19215), .A(n15556), .B(n15555), .ZN(
        P2_U2841) );
  OAI21_X1 U17516 ( .B1(n15371), .B2(n15559), .A(n15558), .ZN(n16083) );
  INV_X1 U17517 ( .A(n15560), .ZN(n16082) );
  XNOR2_X1 U17518 ( .A(n16083), .B(n16082), .ZN(n22205) );
  INV_X1 U17519 ( .A(n20555), .ZN(n15561) );
  AOI21_X1 U17520 ( .B1(n15562), .B2(n20562), .A(n15561), .ZN(n22202) );
  AOI22_X1 U17521 ( .A1(n22202), .A2(n20572), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n16119), .ZN(n15563) );
  OAI21_X1 U17522 ( .B1(n22205), .B2(n16146), .A(n15563), .ZN(P1_U2861) );
  INV_X1 U17523 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20657) );
  OR2_X1 U17524 ( .A1(n16158), .A2(n20657), .ZN(n15565) );
  NAND2_X1 U17525 ( .A1(n16158), .A2(DATAI_11_), .ZN(n15564) );
  NAND2_X1 U17526 ( .A1(n15565), .A2(n15564), .ZN(n22454) );
  AOI22_X1 U17527 ( .A1(n16241), .A2(n22454), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16240), .ZN(n15566) );
  OAI21_X1 U17528 ( .B1(n22205), .B2(n16243), .A(n15566), .ZN(P1_U2893) );
  INV_X1 U17529 ( .A(n15611), .ZN(n15570) );
  NAND2_X1 U17530 ( .A1(n15568), .A2(n15567), .ZN(n15569) );
  NAND2_X1 U17531 ( .A1(n15570), .A2(n15569), .ZN(n19118) );
  AOI21_X1 U17532 ( .B1(n15572), .B2(n15571), .A(n15595), .ZN(n16794) );
  NAND2_X1 U17533 ( .A1(n16794), .A2(n16724), .ZN(n15574) );
  NAND2_X1 U17534 ( .A1(n15538), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15573) );
  OAI211_X1 U17535 ( .C1(n19118), .C2(n15538), .A(n15574), .B(n15573), .ZN(
        P2_U2870) );
  NOR2_X1 U17536 ( .A1(n15575), .A2(n17416), .ZN(n17383) );
  AOI21_X1 U17537 ( .B1(n15583), .B2(n15577), .A(n15576), .ZN(n19031) );
  AOI21_X1 U17538 ( .B1(n15794), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19031), .ZN(n17385) );
  AOI222_X1 U17539 ( .A1(n15578), .A2(n19271), .B1(n17383), .B2(n17385), .C1(
        n19842), .C2(n19320), .ZN(n15581) );
  NAND2_X1 U17540 ( .A1(n15580), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15579) );
  OAI21_X1 U17541 ( .B1(n15581), .B2(n15580), .A(n15579), .ZN(P2_U3600) );
  NOR2_X1 U17542 ( .A1(n19316), .A2(n15795), .ZN(n19086) );
  OAI21_X1 U17543 ( .B1(n19239), .B2(n19086), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15590) );
  INV_X1 U17544 ( .A(n15582), .ZN(n15585) );
  AOI22_X1 U17545 ( .A1(n11121), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n15583), .B2(
        n19265), .ZN(n15584) );
  OAI21_X1 U17546 ( .B1(n19215), .B2(n15585), .A(n15584), .ZN(n15588) );
  OAI22_X1 U17547 ( .A1(n19268), .A2(n15586), .B1(n19256), .B2(n14423), .ZN(
        n15587) );
  AOI211_X1 U17548 ( .C1(n19276), .C2(n19251), .A(n15588), .B(n15587), .ZN(
        n15589) );
  OAI211_X1 U17549 ( .C1(n15591), .C2(n19825), .A(n15590), .B(n15589), .ZN(
        P2_U2855) );
  INV_X1 U17550 ( .A(n15592), .ZN(n15593) );
  OAI21_X1 U17551 ( .B1(n15595), .B2(n15594), .A(n15593), .ZN(n15615) );
  AND2_X1 U17552 ( .A1(n15602), .A2(n15596), .ZN(n15597) );
  NAND2_X1 U17553 ( .A1(n16799), .A2(n15598), .ZN(n15599) );
  NAND2_X1 U17554 ( .A1(n15639), .A2(n15599), .ZN(n19136) );
  OAI22_X1 U17555 ( .A1(n16790), .A2(n19136), .B1(n15640), .B2(n15600), .ZN(
        n15608) );
  AND2_X1 U17556 ( .A1(n15602), .A2(n15601), .ZN(n15603) );
  INV_X1 U17557 ( .A(n20114), .ZN(n15606) );
  INV_X1 U17558 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15605) );
  INV_X1 U17559 ( .A(n20113), .ZN(n16737) );
  OAI22_X1 U17560 ( .A1(n15606), .A2(n15605), .B1(n16737), .B2(n20205), .ZN(
        n15607) );
  AOI211_X1 U17561 ( .C1(n20115), .C2(BUF1_REG_18__SCAN_IN), .A(n15608), .B(
        n15607), .ZN(n15609) );
  OAI21_X1 U17562 ( .B1(n15615), .B2(n20065), .A(n15609), .ZN(P2_U2901) );
  OR2_X1 U17563 ( .A1(n15611), .A2(n15610), .ZN(n15612) );
  NAND2_X1 U17564 ( .A1(n11228), .A2(n15612), .ZN(n19128) );
  NOR2_X1 U17565 ( .A1(n19128), .A2(n15538), .ZN(n15613) );
  AOI21_X1 U17566 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n15538), .A(n15613), .ZN(
        n15614) );
  OAI21_X1 U17567 ( .B1(n15615), .B2(n16732), .A(n15614), .ZN(P2_U2869) );
  NAND2_X1 U17568 ( .A1(n15617), .A2(n15616), .ZN(n16084) );
  AOI21_X1 U17569 ( .B1(n15619), .B2(n16084), .A(n11633), .ZN(n16373) );
  INV_X1 U17570 ( .A(n16373), .ZN(n15632) );
  NAND2_X1 U17571 ( .A1(n16088), .A2(n15620), .ZN(n15621) );
  AND2_X1 U17572 ( .A1(n16139), .A2(n15621), .ZN(n21952) );
  INV_X1 U17573 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n17751) );
  INV_X1 U17574 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n22185) );
  NOR2_X1 U17575 ( .A1(n22175), .A2(n22185), .ZN(n22188) );
  NAND2_X1 U17576 ( .A1(n22188), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n22201) );
  INV_X1 U17577 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n22211) );
  NOR2_X1 U17578 ( .A1(n22201), .A2(n22211), .ZN(n22215) );
  NAND2_X1 U17579 ( .A1(n22215), .A2(P1_REIP_REG_12__SCAN_IN), .ZN(n16090) );
  NOR3_X1 U17580 ( .A1(n22200), .A2(n17751), .A3(n16090), .ZN(n15622) );
  NAND2_X1 U17581 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15622), .ZN(n22225) );
  OAI211_X1 U17582 ( .C1(P1_REIP_REG_14__SCAN_IN), .C2(n15622), .A(n22273), 
        .B(n22225), .ZN(n15628) );
  INV_X1 U17583 ( .A(n16371), .ZN(n15623) );
  NAND2_X1 U17584 ( .A1(n22253), .A2(n15623), .ZN(n15625) );
  NAND2_X1 U17585 ( .A1(n22263), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15624) );
  NAND3_X1 U17586 ( .A1(n15625), .A2(n15624), .A3(n22264), .ZN(n15626) );
  AOI21_X1 U17587 ( .B1(n22272), .B2(P1_EBX_REG_14__SCAN_IN), .A(n15626), .ZN(
        n15627) );
  NAND2_X1 U17588 ( .A1(n15628), .A2(n15627), .ZN(n15629) );
  AOI21_X1 U17589 ( .B1(n21952), .B2(n22255), .A(n15629), .ZN(n15630) );
  OAI21_X1 U17590 ( .B1(n15632), .B2(n22268), .A(n15630), .ZN(P1_U2826) );
  MUX2_X1 U17591 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n16158), .Z(
        n22476) );
  AOI22_X1 U17592 ( .A1(n16241), .A2(n22476), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16240), .ZN(n15631) );
  OAI21_X1 U17593 ( .B1(n15632), .B2(n16243), .A(n15631), .ZN(P1_U2890) );
  NAND2_X1 U17594 ( .A1(n16373), .A2(n14221), .ZN(n15634) );
  NAND2_X1 U17595 ( .A1(n21952), .A2(n20572), .ZN(n15633) );
  OAI211_X1 U17596 ( .C1(n17794), .C2(n20574), .A(n15634), .B(n15633), .ZN(
        P1_U2858) );
  OAI21_X1 U17597 ( .B1(n15592), .B2(n15636), .A(n15635), .ZN(n16733) );
  AOI22_X1 U17598 ( .A1(n20114), .A2(BUF2_REG_19__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15644) );
  INV_X1 U17599 ( .A(n15637), .ZN(n15638) );
  XNOR2_X1 U17600 ( .A(n15639), .B(n15638), .ZN(n19138) );
  OAI22_X1 U17601 ( .A1(n16737), .A2(n20165), .B1(n15641), .B2(n15640), .ZN(
        n15642) );
  AOI21_X1 U17602 ( .B1(n20117), .B2(n19138), .A(n15642), .ZN(n15643) );
  OAI211_X1 U17603 ( .C1(n16733), .C2(n20065), .A(n15644), .B(n15643), .ZN(
        P2_U2900) );
  NOR3_X4 U17604 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n15645), .ZN(n18407) );
  BUF_X4 U17605 ( .A(n18407), .Z(n18434) );
  AOI22_X1 U17606 ( .A1(n18434), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15649) );
  NOR2_X2 U17607 ( .A1(n15651), .A2(n15650), .ZN(n15716) );
  AOI22_X1 U17608 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U17609 ( .A1(n11127), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15647) );
  NOR2_X2 U17610 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n21401), .ZN(
        n15725) );
  AOI22_X1 U17611 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n15646) );
  NAND4_X1 U17612 ( .A1(n15649), .A2(n15648), .A3(n15647), .A4(n15646), .ZN(
        n15658) );
  AOI22_X1 U17613 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15656) );
  AOI22_X1 U17614 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11131), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n15655) );
  AOI22_X1 U17615 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n15654) );
  NAND3_X1 U17616 ( .A1(n21888), .A2(n21891), .A3(n20764), .ZN(n15724) );
  OR2_X2 U17617 ( .A1(n15652), .A2(n21411), .ZN(n18202) );
  AOI22_X1 U17618 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n15653) );
  NAND4_X1 U17619 ( .A1(n15656), .A2(n15655), .A3(n15654), .A4(n15653), .ZN(
        n15657) );
  AOI22_X1 U17620 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15662) );
  AOI22_X1 U17621 ( .A1(n18434), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15661) );
  AOI22_X1 U17622 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15660) );
  AOI22_X1 U17623 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15659) );
  NAND4_X1 U17624 ( .A1(n15662), .A2(n15661), .A3(n15660), .A4(n15659), .ZN(
        n15668) );
  AOI22_X1 U17625 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15666) );
  AOI22_X1 U17626 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15665) );
  AOI22_X1 U17627 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15664) );
  AOI22_X1 U17628 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11132), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15663) );
  NAND4_X1 U17629 ( .A1(n15666), .A2(n15665), .A3(n15664), .A4(n15663), .ZN(
        n15667) );
  AOI22_X1 U17630 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15672) );
  INV_X2 U17631 ( .A(n20786), .ZN(n18423) );
  AOI22_X1 U17632 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15671) );
  AOI22_X1 U17633 ( .A1(n11126), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15670) );
  AOI22_X1 U17634 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15669) );
  NAND4_X1 U17635 ( .A1(n15672), .A2(n15671), .A3(n15670), .A4(n15669), .ZN(
        n15678) );
  AOI22_X1 U17636 ( .A1(n15715), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15676) );
  AOI22_X1 U17637 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n15675) );
  AOI22_X1 U17638 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15674) );
  AOI22_X1 U17639 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15673) );
  NAND4_X1 U17640 ( .A1(n15676), .A2(n15675), .A3(n15674), .A4(n15673), .ZN(
        n15677) );
  AOI22_X1 U17641 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18407), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15682) );
  INV_X2 U17642 ( .A(n18086), .ZN(n18453) );
  AOI22_X1 U17643 ( .A1(n11131), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15681) );
  AOI22_X1 U17644 ( .A1(n11126), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15680) );
  AOI22_X1 U17645 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n15679) );
  NAND4_X1 U17646 ( .A1(n15682), .A2(n15681), .A3(n15680), .A4(n15679), .ZN(
        n15688) );
  AOI22_X1 U17647 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15686) );
  AOI22_X1 U17648 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15685) );
  AOI22_X1 U17649 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15684) );
  AOI22_X1 U17650 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n15683) );
  NAND4_X1 U17651 ( .A1(n15686), .A2(n15685), .A3(n15684), .A4(n15683), .ZN(
        n15687) );
  AOI22_X1 U17652 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15692) );
  AOI22_X1 U17653 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15691) );
  AOI22_X1 U17654 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15690) );
  AOI22_X1 U17655 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15689) );
  NAND4_X1 U17656 ( .A1(n15692), .A2(n15691), .A3(n15690), .A4(n15689), .ZN(
        n15698) );
  AOI22_X1 U17657 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15696) );
  AOI22_X1 U17658 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15695) );
  AOI22_X1 U17659 ( .A1(n15715), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15694) );
  AOI22_X1 U17660 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15693) );
  NAND4_X1 U17661 ( .A1(n15696), .A2(n15695), .A3(n15694), .A4(n15693), .ZN(
        n15697) );
  AOI22_X1 U17662 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15708) );
  AOI22_X1 U17663 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15707) );
  AOI22_X1 U17664 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15699) );
  OAI21_X1 U17665 ( .B1(n15724), .B2(n19447), .A(n15699), .ZN(n15705) );
  AOI22_X1 U17666 ( .A1(n15715), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15703) );
  AOI22_X1 U17667 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15702) );
  AOI22_X1 U17668 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15701) );
  AOI22_X1 U17669 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15700) );
  NAND4_X1 U17670 ( .A1(n15703), .A2(n15702), .A3(n15701), .A4(n15700), .ZN(
        n15704) );
  NAND3_X2 U17671 ( .A1(n15708), .A2(n15707), .A3(n15706), .ZN(n21294) );
  NAND4_X1 U17672 ( .A1(n21439), .A2(n21442), .A3(n19572), .A4(n15743), .ZN(
        n21409) );
  AOI22_X1 U17673 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15712) );
  AOI22_X1 U17674 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15711) );
  AOI22_X1 U17675 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15710) );
  INV_X2 U17676 ( .A(n11184), .ZN(n20804) );
  AOI22_X1 U17677 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15709) );
  NAND4_X1 U17678 ( .A1(n15712), .A2(n15711), .A3(n15710), .A4(n15709), .ZN(
        n15722) );
  AOI22_X1 U17679 ( .A1(n15713), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15720) );
  AOI22_X1 U17680 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15719) );
  AOI22_X1 U17681 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15718) );
  AOI22_X1 U17682 ( .A1(n11132), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15717) );
  NAND4_X1 U17683 ( .A1(n15720), .A2(n15719), .A3(n15718), .A4(n15717), .ZN(
        n15721) );
  AOI22_X1 U17684 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U17685 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15733) );
  AOI22_X1 U17686 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18407), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n15723) );
  OAI21_X1 U17687 ( .B1(n15724), .B2(n19698), .A(n15723), .ZN(n15731) );
  AOI22_X1 U17688 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15729) );
  AOI22_X1 U17689 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15728) );
  AOI22_X1 U17690 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15727) );
  AOI22_X1 U17691 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15726) );
  NAND4_X1 U17692 ( .A1(n15729), .A2(n15728), .A3(n15727), .A4(n15726), .ZN(
        n15730) );
  INV_X1 U17693 ( .A(n19490), .ZN(n21254) );
  NOR3_X1 U17694 ( .A1(n21396), .A2(n15772), .A3(n15776), .ZN(n15736) );
  INV_X1 U17695 ( .A(n21442), .ZN(n17983) );
  NOR2_X1 U17696 ( .A1(n21440), .A2(n17983), .ZN(n15768) );
  AOI211_X1 U17697 ( .C1(n21433), .C2(n15768), .A(n19572), .B(n21438), .ZN(
        n15735) );
  NOR2_X1 U17698 ( .A1(n15736), .A2(n15735), .ZN(n15746) );
  NAND3_X1 U17699 ( .A1(n19490), .A2(n18488), .A3(n15746), .ZN(n15737) );
  NAND2_X1 U17700 ( .A1(n15747), .A2(n21440), .ZN(n15770) );
  NAND2_X1 U17701 ( .A1(n21435), .A2(n19708), .ZN(n17408) );
  NOR2_X1 U17702 ( .A1(n21435), .A2(n15737), .ZN(n21913) );
  INV_X1 U17703 ( .A(n21913), .ZN(n20710) );
  INV_X1 U17704 ( .A(n19572), .ZN(n15742) );
  NAND2_X1 U17705 ( .A1(n15772), .A2(n21395), .ZN(n17982) );
  INV_X1 U17706 ( .A(n17982), .ZN(n15739) );
  NAND2_X1 U17707 ( .A1(n19657), .A2(n19708), .ZN(n21192) );
  INV_X1 U17708 ( .A(n21192), .ZN(n15738) );
  NAND3_X1 U17709 ( .A1(n15739), .A2(n21294), .A3(n15738), .ZN(n15740) );
  AND2_X1 U17710 ( .A1(n17408), .A2(n21434), .ZN(n15769) );
  NAND2_X1 U17711 ( .A1(n11367), .A2(n19657), .ZN(n17409) );
  NOR2_X1 U17712 ( .A1(n21267), .A2(n21382), .ZN(n21197) );
  OAI21_X1 U17713 ( .B1(n21439), .B2(n21267), .A(n17983), .ZN(n15741) );
  OAI211_X1 U17714 ( .C1(n15743), .C2(n15742), .A(n15774), .B(n15741), .ZN(
        n15744) );
  INV_X1 U17715 ( .A(n15744), .ZN(n15745) );
  OAI211_X1 U17716 ( .C1(n21439), .C2(n15769), .A(n15746), .B(n15745), .ZN(
        n18489) );
  NAND2_X1 U17717 ( .A1(n15748), .A2(n17392), .ZN(n17391) );
  NAND2_X1 U17718 ( .A1(n18491), .A2(n17391), .ZN(n21910) );
  NOR2_X1 U17719 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21426) );
  INV_X1 U17720 ( .A(n21426), .ZN(n21402) );
  NOR2_X1 U17721 ( .A1(n21910), .A2(n21402), .ZN(n15778) );
  INV_X1 U17722 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n22369) );
  INV_X1 U17723 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n22320) );
  NAND2_X1 U17724 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n22320), .ZN(n22375) );
  INV_X2 U17725 ( .A(n19006), .ZN(n22323) );
  AOI21_X1 U17726 ( .B1(n19006), .B2(n22375), .A(n18997), .ZN(n21436) );
  NAND2_X1 U17727 ( .A1(n21436), .A2(n15749), .ZN(n17407) );
  OAI22_X1 U17728 ( .A1(n21392), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n21895), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U17729 ( .A1(n21892), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15762) );
  XNOR2_X1 U17730 ( .A(n15763), .B(n15762), .ZN(n15761) );
  NOR2_X1 U17731 ( .A1(n15762), .A2(n15763), .ZN(n15750) );
  INV_X1 U17732 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21900) );
  OAI22_X1 U17733 ( .A1(n21891), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n21900), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15755) );
  OAI21_X1 U17734 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21891), .A(
        n15751), .ZN(n15752) );
  OAI22_X1 U17735 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21904), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n15752), .ZN(n15758) );
  NOR2_X1 U17736 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21904), .ZN(
        n15753) );
  NAND2_X1 U17737 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n15752), .ZN(
        n15757) );
  AOI22_X1 U17738 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15758), .B1(
        n15753), .B2(n15757), .ZN(n15764) );
  NAND2_X1 U17739 ( .A1(n15756), .A2(n15755), .ZN(n15754) );
  AND2_X1 U17740 ( .A1(n15757), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15759) );
  OAI22_X1 U17741 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n17392), .B1(
        n15759), .B2(n15758), .ZN(n15760) );
  INV_X1 U17742 ( .A(n15760), .ZN(n15766) );
  AOI21_X1 U17743 ( .B1(n21194), .B2(n17407), .A(n21881), .ZN(n15777) );
  NAND2_X1 U17744 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n22370) );
  OAI21_X1 U17745 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21892), .A(
        n15762), .ZN(n18485) );
  INV_X1 U17746 ( .A(n15763), .ZN(n15765) );
  NAND2_X1 U17747 ( .A1(n15765), .A2(n15764), .ZN(n15767) );
  OAI211_X1 U17748 ( .C1(n18485), .C2(n15767), .A(n15766), .B(n18486), .ZN(
        n21877) );
  NAND3_X1 U17749 ( .A1(n18488), .A2(n21438), .A3(n21396), .ZN(n18487) );
  INV_X1 U17750 ( .A(n15768), .ZN(n15775) );
  OAI211_X1 U17751 ( .C1(n21442), .C2(n21382), .A(n18488), .B(n15769), .ZN(
        n15771) );
  OAI21_X1 U17752 ( .B1(n15772), .B2(n15771), .A(n15770), .ZN(n15773) );
  OAI211_X1 U17753 ( .C1(n15776), .C2(n15775), .A(n15774), .B(n15773), .ZN(
        n21444) );
  NAND2_X1 U17754 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n21936), .ZN(n19366) );
  NAND2_X1 U17755 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18359) );
  NOR2_X1 U17756 ( .A1(n21936), .A2(n18359), .ZN(n17405) );
  NAND2_X1 U17757 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n17405), .ZN(n17393) );
  OAI211_X1 U17758 ( .C1(n21909), .C2(n21937), .A(n19366), .B(n17393), .ZN(
        n21429) );
  INV_X1 U17759 ( .A(n21429), .ZN(n21431) );
  MUX2_X1 U17760 ( .A(n15778), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n21431), .Z(P3_U3284) );
  INV_X1 U17761 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n19209) );
  INV_X1 U17762 ( .A(n15799), .ZN(n15779) );
  AOI21_X1 U17763 ( .B1(n19209), .B2(n15779), .A(n14024), .ZN(n16829) );
  INV_X1 U17764 ( .A(n16829), .ZN(n19220) );
  OR2_X1 U17765 ( .A1(n11243), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15781) );
  NAND2_X1 U17766 ( .A1(n15780), .A2(n15781), .ZN(n19178) );
  INV_X1 U17767 ( .A(n19178), .ZN(n19180) );
  AOI21_X1 U17768 ( .B1(n16872), .B2(n15782), .A(n11243), .ZN(n19162) );
  NAND2_X1 U17769 ( .A1(n15785), .A2(n11556), .ZN(n15784) );
  NAND2_X1 U17770 ( .A1(n15782), .A2(n15784), .ZN(n16884) );
  INV_X1 U17771 ( .A(n16884), .ZN(n19154) );
  AOI21_X1 U17772 ( .B1(n16902), .B2(n11548), .A(n11143), .ZN(n16905) );
  OAI21_X1 U17773 ( .B1(n15786), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n11548), .ZN(n16911) );
  INV_X1 U17774 ( .A(n16911), .ZN(n16639) );
  AOI21_X1 U17775 ( .B1(n16919), .B2(n11235), .A(n15786), .ZN(n19142) );
  OAI21_X1 U17776 ( .B1(n15787), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11235), .ZN(n16931) );
  INV_X1 U17777 ( .A(n16931), .ZN(n19130) );
  OAI21_X1 U17778 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15464), .A(
        n15788), .ZN(n19100) );
  INV_X1 U17779 ( .A(n19100), .ZN(n15791) );
  INV_X1 U17780 ( .A(n16968), .ZN(n15789) );
  NAND2_X1 U17781 ( .A1(n15790), .A2(n15789), .ZN(n19099) );
  NOR2_X1 U17782 ( .A1(n15791), .A2(n19099), .ZN(n19112) );
  INV_X1 U17783 ( .A(n15787), .ZN(n15793) );
  NAND2_X1 U17784 ( .A1(n12538), .A2(n15788), .ZN(n15792) );
  NAND2_X1 U17785 ( .A1(n15793), .A2(n15792), .ZN(n19123) );
  NOR2_X1 U17786 ( .A1(n15794), .A2(n19129), .ZN(n19141) );
  NOR2_X1 U17787 ( .A1(n19142), .A2(n19141), .ZN(n19140) );
  NOR2_X1 U17788 ( .A1(n16639), .A2(n16638), .ZN(n16637) );
  NOR2_X1 U17789 ( .A1(n15794), .A2(n16637), .ZN(n16633) );
  NOR2_X1 U17790 ( .A1(n19162), .A2(n19161), .ZN(n19160) );
  AOI21_X1 U17791 ( .B1(n19180), .B2(n15795), .A(n19179), .ZN(n19192) );
  INV_X1 U17792 ( .A(n15798), .ZN(n15796) );
  AOI21_X1 U17793 ( .B1(n16852), .B2(n15780), .A(n15796), .ZN(n16854) );
  INV_X1 U17794 ( .A(n16854), .ZN(n19191) );
  NAND2_X1 U17795 ( .A1(n19190), .A2(n15795), .ZN(n19201) );
  AND2_X1 U17796 ( .A1(n15798), .A2(n15797), .ZN(n15800) );
  OR2_X1 U17797 ( .A1(n15800), .A2(n15799), .ZN(n19202) );
  NAND2_X1 U17798 ( .A1(n19201), .A2(n19202), .ZN(n19200) );
  NAND2_X1 U17799 ( .A1(n19200), .A2(n15795), .ZN(n19219) );
  NAND2_X1 U17800 ( .A1(n19220), .A2(n19219), .ZN(n19218) );
  NAND2_X1 U17801 ( .A1(n15795), .A2(n19218), .ZN(n19230) );
  NAND2_X1 U17802 ( .A1(n19230), .A2(n19231), .ZN(n19229) );
  NAND2_X1 U17803 ( .A1(n19229), .A2(n15795), .ZN(n19245) );
  NAND2_X1 U17804 ( .A1(n14023), .A2(n16818), .ZN(n15801) );
  AND2_X1 U17805 ( .A1(n15802), .A2(n15801), .ZN(n16820) );
  INV_X1 U17806 ( .A(n16820), .ZN(n19246) );
  NAND2_X1 U17807 ( .A1(n19245), .A2(n19246), .ZN(n19243) );
  NAND2_X1 U17808 ( .A1(n15795), .A2(n19243), .ZN(n19263) );
  AOI21_X1 U17809 ( .B1(n19264), .B2(n19263), .A(n19316), .ZN(n15804) );
  OR2_X1 U17810 ( .A1(n19263), .A2(n19264), .ZN(n15803) );
  AOI222_X1 U17811 ( .A1(n15805), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n15828), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n15806), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15809) );
  AOI22_X1 U17812 ( .A1(n15828), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15807) );
  OAI21_X1 U17813 ( .B1(n15830), .B2(n17974), .A(n15807), .ZN(n16734) );
  AOI21_X1 U17814 ( .B1(n15809), .B2(n11188), .A(n15832), .ZN(n17064) );
  NAND2_X1 U17815 ( .A1(n17064), .A2(n19241), .ZN(n15811) );
  AOI22_X1 U17816 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n11121), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19239), .ZN(n15810) );
  OAI211_X1 U17817 ( .C1(n17976), .C2(n19256), .A(n15811), .B(n15810), .ZN(
        n15812) );
  AOI21_X1 U17818 ( .B1(n17061), .B2(n19251), .A(n15812), .ZN(n15813) );
  OAI211_X1 U17819 ( .C1(n15815), .C2(n19215), .A(n15814), .B(n15813), .ZN(
        P2_U2825) );
  INV_X1 U17820 ( .A(n15824), .ZN(n15816) );
  INV_X1 U17821 ( .A(DATAI_31_), .ZN(n15827) );
  AOI22_X1 U17822 ( .A1(n13293), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n15818), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n15819) );
  INV_X1 U17823 ( .A(n15819), .ZN(n15820) );
  AND2_X1 U17824 ( .A1(n16231), .A2(n15908), .ZN(n15822) );
  AOI22_X1 U17825 ( .A1(n16229), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n16240), .ZN(n15825) );
  OAI211_X1 U17826 ( .C1(n16227), .C2(n15827), .A(n15826), .B(n15825), .ZN(
        P1_U2873) );
  INV_X1 U17827 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19255) );
  AOI22_X1 U17828 ( .A1(n15828), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n15806), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15829) );
  OAI21_X1 U17829 ( .B1(n15830), .B2(n19255), .A(n15829), .ZN(n15831) );
  XNOR2_X1 U17830 ( .A(n15832), .B(n15831), .ZN(n19269) );
  AOI22_X1 U17831 ( .A1(n20115), .A2(BUF1_REG_31__SCAN_IN), .B1(n20111), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n15834) );
  NAND2_X1 U17832 ( .A1(n20114), .A2(BUF2_REG_31__SCAN_IN), .ZN(n15833) );
  OAI211_X1 U17833 ( .C1(n19269), .C2(n16790), .A(n15834), .B(n15833), .ZN(
        P2_U2888) );
  INV_X1 U17834 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16414) );
  XNOR2_X1 U17835 ( .A(n20603), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15840) );
  INV_X1 U17836 ( .A(n15840), .ZN(n15836) );
  AOI21_X1 U17837 ( .B1(n16403), .B2(n16414), .A(n20603), .ZN(n15837) );
  INV_X1 U17838 ( .A(n15837), .ZN(n15835) );
  NAND2_X1 U17839 ( .A1(n15836), .A2(n15835), .ZN(n15843) );
  NAND2_X1 U17840 ( .A1(n20603), .A2(n16403), .ZN(n15839) );
  INV_X1 U17841 ( .A(n15839), .ZN(n15838) );
  OAI21_X1 U17842 ( .B1(n15838), .B2(n15837), .A(n16415), .ZN(n15842) );
  OAI211_X1 U17843 ( .C1(n15844), .C2(n15843), .A(n15842), .B(n15841), .ZN(
        n16421) );
  INV_X1 U17844 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20521) );
  NOR2_X1 U17845 ( .A1(n22044), .A2(n20521), .ZN(n16418) );
  AOI21_X1 U17846 ( .B1(n20628), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16418), .ZN(n15845) );
  OAI21_X1 U17847 ( .B1(n20634), .B2(n15846), .A(n15845), .ZN(n15847) );
  OAI21_X1 U17848 ( .B1(n22280), .B2(n16421), .A(n15848), .ZN(P1_U2968) );
  AOI22_X1 U17849 ( .A1(n20114), .A2(BUF2_REG_30__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15850) );
  AOI22_X1 U17850 ( .A1(n20113), .A2(n19806), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n20111), .ZN(n15849) );
  NAND2_X1 U17851 ( .A1(n15850), .A2(n15849), .ZN(n15851) );
  AOI21_X1 U17852 ( .B1(n17064), .B2(n20117), .A(n15851), .ZN(n15852) );
  OAI21_X1 U17853 ( .B1(n15853), .B2(n20065), .A(n15852), .ZN(P2_U2889) );
  NOR2_X1 U17854 ( .A1(n15856), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n15858) );
  MUX2_X1 U17855 ( .A(n12260), .B(n15858), .S(n15857), .Z(n19262) );
  NAND2_X1 U17856 ( .A1(n19262), .A2(n15859), .ZN(n15860) );
  XNOR2_X1 U17857 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n15861), .ZN(
        n15862) );
  INV_X1 U17858 ( .A(n15862), .ZN(n15882) );
  NAND2_X1 U17859 ( .A1(n15864), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15867) );
  AOI22_X1 U17860 ( .A1(n15865), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n15866) );
  OAI211_X1 U17861 ( .C1(n15868), .C2(n19255), .A(n15867), .B(n15866), .ZN(
        n15869) );
  NAND2_X1 U17862 ( .A1(n17092), .A2(n11602), .ZN(n17078) );
  OAI22_X1 U17863 ( .A1(n17078), .A2(n17065), .B1(n19279), .B2(n15870), .ZN(
        n17066) );
  INV_X1 U17864 ( .A(n15872), .ZN(n15875) );
  NOR2_X1 U17865 ( .A1(n19294), .A2(n19255), .ZN(n15878) );
  INV_X1 U17866 ( .A(n15878), .ZN(n15873) );
  OAI21_X1 U17867 ( .B1(n15886), .B2(n17351), .A(n15877), .ZN(P2_U3015) );
  AOI21_X1 U17868 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15878), .ZN(n15879) );
  OAI21_X1 U17869 ( .B1(n17042), .B2(n15880), .A(n15879), .ZN(n15881) );
  NAND2_X1 U17870 ( .A1(n15862), .A2(n17843), .ZN(n15883) );
  OAI21_X1 U17871 ( .B1(n15886), .B2(n17853), .A(n15885), .ZN(P2_U2983) );
  XOR2_X1 U17872 ( .A(n15888), .B(n15887), .Z(n17357) );
  AOI21_X1 U17873 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(n17356) );
  NOR2_X1 U17874 ( .A1(n19294), .A2(n12060), .ZN(n17364) );
  AOI21_X1 U17875 ( .B1(n17843), .B2(n17356), .A(n17364), .ZN(n15894) );
  NAND2_X1 U17876 ( .A1(n17862), .A2(n15892), .ZN(n15893) );
  OAI211_X1 U17877 ( .C1(n15895), .C2(n17877), .A(n15894), .B(n15893), .ZN(
        n15896) );
  AOI21_X1 U17878 ( .B1(n17357), .B2(n17871), .A(n15896), .ZN(n15897) );
  OAI21_X1 U17879 ( .B1(n12110), .B2(n17852), .A(n15897), .ZN(P2_U3012) );
  INV_X1 U17880 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20701) );
  NAND2_X1 U17881 ( .A1(n15898), .A2(n20701), .ZN(n15901) );
  INV_X1 U17882 ( .A(n15899), .ZN(n15900) );
  MUX2_X1 U17883 ( .A(n15901), .B(n15900), .S(n21943), .Z(P1_U3487) );
  NAND2_X1 U17884 ( .A1(n15903), .A2(n15902), .ZN(n15905) );
  MUX2_X1 U17885 ( .A(n15905), .B(n15904), .S(n15910), .Z(n15906) );
  AOI21_X1 U17886 ( .B1(n14409), .B2(n15907), .A(n15906), .ZN(n15909) );
  NOR2_X1 U17887 ( .A1(n15909), .A2(n15908), .ZN(n17450) );
  OAI22_X1 U17888 ( .A1(n15913), .A2(n15912), .B1(n15911), .B2(n15910), .ZN(
        n20635) );
  INV_X1 U17889 ( .A(n15914), .ZN(n15915) );
  AOI21_X1 U17890 ( .B1(n15915), .B2(n22338), .A(n22327), .ZN(n21946) );
  NOR2_X1 U17891 ( .A1(n20635), .A2(n21946), .ZN(n17453) );
  NOR2_X1 U17892 ( .A1(n17453), .A2(n22303), .ZN(n22281) );
  MUX2_X1 U17893 ( .A(P1_MORE_REG_SCAN_IN), .B(n17450), .S(n22281), .Z(
        P1_U3484) );
  OAI22_X1 U17894 ( .A1(n15918), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n15917), .B2(P1_EBX_REG_31__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U17895 ( .A1(n15921), .A2(n22256), .ZN(n15931) );
  NAND2_X1 U17896 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16031) );
  NAND2_X1 U17897 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n16032) );
  INV_X1 U17898 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n17744) );
  NOR4_X1 U17899 ( .A1(n16031), .A2(n16032), .A3(n17751), .A4(n17744), .ZN(
        n15922) );
  NAND3_X1 U17900 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(n15922), .ZN(n16050) );
  INV_X1 U17901 ( .A(n16050), .ZN(n15923) );
  NAND3_X1 U17902 ( .A1(n15923), .A2(P1_REIP_REG_21__SCAN_IN), .A3(
        P1_REIP_REG_22__SCAN_IN), .ZN(n15924) );
  NOR2_X1 U17903 ( .A1(n16090), .A2(n15924), .ZN(n15925) );
  AND2_X1 U17904 ( .A1(n22214), .A2(n15925), .ZN(n16021) );
  INV_X1 U17905 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n17643) );
  INV_X1 U17906 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n17734) );
  NOR2_X1 U17907 ( .A1(n17643), .A2(n17734), .ZN(n15985) );
  NAND3_X1 U17908 ( .A1(n16012), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n15985), 
        .ZN(n15984) );
  INV_X1 U17909 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20513) );
  NOR2_X1 U17910 ( .A1(n15984), .A2(n20513), .ZN(n15973) );
  NAND2_X1 U17911 ( .A1(n15973), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15957) );
  INV_X1 U17912 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20517) );
  NOR2_X1 U17913 ( .A1(n15957), .A2(n20517), .ZN(n15935) );
  AND2_X1 U17914 ( .A1(n15935), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n15926) );
  INV_X1 U17915 ( .A(n22273), .ZN(n15995) );
  NOR2_X1 U17916 ( .A1(n15926), .A2(n15995), .ZN(n15934) );
  INV_X1 U17917 ( .A(n15926), .ZN(n15928) );
  AOI22_X1 U17918 ( .A1(n22272), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n22263), .ZN(n15927) );
  OAI21_X1 U17919 ( .B1(n15928), .B2(P1_REIP_REG_31__SCAN_IN), .A(n15927), 
        .ZN(n15929) );
  AOI21_X1 U17920 ( .B1(n15934), .B2(P1_REIP_REG_31__SCAN_IN), .A(n15929), 
        .ZN(n15930) );
  OAI211_X1 U17921 ( .C1(n16396), .C2(n22278), .A(n15931), .B(n15930), .ZN(
        P1_U2809) );
  INV_X1 U17922 ( .A(n15933), .ZN(n16427) );
  OAI21_X1 U17923 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n15935), .A(n15934), 
        .ZN(n15938) );
  AOI22_X1 U17924 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n15936), .ZN(n15937) );
  OAI211_X1 U17925 ( .C1(n17640), .C2(n22249), .A(n15938), .B(n15937), .ZN(
        n15939) );
  AOI21_X1 U17926 ( .B1(n16427), .B2(n22255), .A(n15939), .ZN(n15940) );
  OAI21_X1 U17927 ( .B1(n16150), .B2(n22268), .A(n15940), .ZN(P1_U2810) );
  INV_X1 U17928 ( .A(n16250), .ZN(n16113) );
  XNOR2_X1 U17929 ( .A(n15945), .B(n15944), .ZN(n16111) );
  INV_X1 U17930 ( .A(n16111), .ZN(n16434) );
  NAND3_X1 U17931 ( .A1(n15957), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n22273), 
        .ZN(n15949) );
  OAI22_X1 U17932 ( .A1(n15946), .A2(n22246), .B1(n22267), .B2(n16248), .ZN(
        n15947) );
  AOI21_X1 U17933 ( .B1(n22272), .B2(P1_EBX_REG_29__SCAN_IN), .A(n15947), .ZN(
        n15948) );
  OAI211_X1 U17934 ( .C1(n15957), .C2(P1_REIP_REG_29__SCAN_IN), .A(n15949), 
        .B(n15948), .ZN(n15950) );
  AOI21_X1 U17935 ( .B1(n16434), .B2(n22255), .A(n15950), .ZN(n15951) );
  OAI21_X1 U17936 ( .B1(n16113), .B2(n22268), .A(n15951), .ZN(P1_U2811) );
  BUF_X1 U17937 ( .A(n15952), .Z(n15953) );
  OAI21_X1 U17938 ( .B1(n15956), .B2(n15965), .A(n15955), .ZN(n16447) );
  INV_X1 U17939 ( .A(n16447), .ZN(n15963) );
  AOI21_X1 U17940 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n22273), .A(n15973), 
        .ZN(n15961) );
  INV_X1 U17941 ( .A(n15957), .ZN(n15960) );
  AOI22_X1 U17942 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16254), .ZN(n15959) );
  NAND2_X1 U17943 ( .A1(n22272), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n15958) );
  OAI211_X1 U17944 ( .C1(n15961), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        n15962) );
  AOI21_X1 U17945 ( .B1(n15963), .B2(n22255), .A(n15962), .ZN(n15964) );
  OAI21_X1 U17946 ( .B1(n16265), .B2(n22268), .A(n15964), .ZN(P1_U2812) );
  INV_X1 U17947 ( .A(n15965), .ZN(n15968) );
  NAND2_X1 U17948 ( .A1(n15982), .A2(n15966), .ZN(n15967) );
  NAND2_X1 U17949 ( .A1(n15968), .A2(n15967), .ZN(n16448) );
  INV_X1 U17950 ( .A(n15969), .ZN(n15970) );
  AOI21_X2 U17951 ( .B1(n15971), .B2(n15970), .A(n15953), .ZN(n16272) );
  NAND2_X1 U17952 ( .A1(n16272), .A2(n22256), .ZN(n15978) );
  OAI22_X1 U17953 ( .A1(n15972), .A2(n22246), .B1(n22267), .B2(n16270), .ZN(
        n15976) );
  NAND2_X1 U17954 ( .A1(n22273), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15974) );
  AOI21_X1 U17955 ( .B1(n15984), .B2(n15974), .A(n15973), .ZN(n15975) );
  AOI211_X1 U17956 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n22272), .A(n15976), .B(
        n15975), .ZN(n15977) );
  OAI211_X1 U17957 ( .C1(n16448), .C2(n22278), .A(n15978), .B(n15977), .ZN(
        P1_U2813) );
  XNOR2_X1 U17958 ( .A(n15979), .B(n15980), .ZN(n16281) );
  INV_X1 U17959 ( .A(n11189), .ZN(n16001) );
  INV_X1 U17960 ( .A(n15981), .ZN(n15983) );
  OAI21_X1 U17961 ( .B1(n16001), .B2(n15983), .A(n15982), .ZN(n16115) );
  INV_X1 U17962 ( .A(n16115), .ZN(n16466) );
  INV_X1 U17963 ( .A(n15984), .ZN(n15989) );
  AOI22_X1 U17964 ( .A1(n16012), .A2(n15985), .B1(P1_REIP_REG_26__SCAN_IN), 
        .B2(n22273), .ZN(n15988) );
  AOI22_X1 U17965 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16276), .ZN(n15987) );
  NAND2_X1 U17966 ( .A1(n22272), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n15986) );
  OAI211_X1 U17967 ( .C1(n15989), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        n15990) );
  AOI21_X1 U17968 ( .B1(n16466), .B2(n22255), .A(n15990), .ZN(n15991) );
  OAI21_X1 U17969 ( .B1(n16281), .B2(n22268), .A(n15991), .ZN(P1_U2814) );
  OAI21_X1 U17970 ( .B1(n15993), .B2(n15994), .A(n15979), .ZN(n16286) );
  NOR2_X1 U17971 ( .A1(n16012), .A2(n15995), .ZN(n16020) );
  INV_X1 U17972 ( .A(n16012), .ZN(n15999) );
  XNOR2_X1 U17973 ( .A(P1_REIP_REG_24__SCAN_IN), .B(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15998) );
  AOI22_X1 U17974 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16289), .ZN(n15997) );
  NAND2_X1 U17975 ( .A1(n22272), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U17976 ( .C1(n15999), .C2(n15998), .A(n15997), .B(n15996), .ZN(
        n16000) );
  AOI21_X1 U17977 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(n16020), .A(n16000), 
        .ZN(n16004) );
  AOI21_X1 U17978 ( .B1(n16002), .B2(n11229), .A(n16001), .ZN(n16474) );
  NAND2_X1 U17979 ( .A1(n16474), .A2(n22255), .ZN(n16003) );
  OAI211_X1 U17980 ( .C1(n16286), .C2(n22268), .A(n16004), .B(n16003), .ZN(
        P1_U2815) );
  INV_X1 U17981 ( .A(n16005), .ZN(n16019) );
  NAND2_X1 U17982 ( .A1(n16035), .A2(n16019), .ZN(n16007) );
  NAND2_X1 U17983 ( .A1(n16007), .A2(n16006), .ZN(n16008) );
  NAND2_X1 U17984 ( .A1(n16008), .A2(n11229), .ZN(n16477) );
  INV_X1 U17985 ( .A(n15993), .ZN(n16010) );
  OAI21_X1 U17986 ( .B1(n16011), .B2(n16009), .A(n16010), .ZN(n16295) );
  INV_X1 U17987 ( .A(n16295), .ZN(n16176) );
  NAND2_X1 U17988 ( .A1(n16176), .A2(n22256), .ZN(n16017) );
  INV_X1 U17989 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n17775) );
  NAND2_X1 U17990 ( .A1(n16012), .A2(n17643), .ZN(n16014) );
  AOI22_X1 U17991 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16298), .ZN(n16013) );
  OAI211_X1 U17992 ( .C1(n17775), .C2(n22249), .A(n16014), .B(n16013), .ZN(
        n16015) );
  AOI21_X1 U17993 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n16020), .A(n16015), 
        .ZN(n16016) );
  OAI211_X1 U17994 ( .C1(n16477), .C2(n22278), .A(n16017), .B(n16016), .ZN(
        P1_U2816) );
  AOI21_X1 U17995 ( .B1(n16018), .B2(n11163), .A(n16009), .ZN(n16305) );
  INV_X1 U17996 ( .A(n16305), .ZN(n16185) );
  XNOR2_X1 U17997 ( .A(n16035), .B(n16019), .ZN(n16117) );
  INV_X1 U17998 ( .A(n16117), .ZN(n16495) );
  OAI21_X1 U17999 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(n16021), .A(n16020), 
        .ZN(n16024) );
  INV_X1 U18000 ( .A(n16303), .ZN(n16022) );
  AOI22_X1 U18001 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16022), .ZN(n16023) );
  OAI211_X1 U18002 ( .C1(n17598), .C2(n22249), .A(n16024), .B(n16023), .ZN(
        n16025) );
  AOI21_X1 U18003 ( .B1(n16495), .B2(n22255), .A(n16025), .ZN(n16026) );
  OAI21_X1 U18004 ( .B1(n16185), .B2(n22268), .A(n16026), .ZN(P1_U2817) );
  INV_X1 U18005 ( .A(n16027), .ZN(n16030) );
  INV_X1 U18006 ( .A(n16028), .ZN(n16029) );
  OAI21_X1 U18007 ( .B1(n16030), .B2(n16029), .A(n11163), .ZN(n16186) );
  NOR2_X1 U18008 ( .A1(n17744), .A2(n22225), .ZN(n22235) );
  NAND2_X1 U18009 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(n22235), .ZN(n16071) );
  NOR2_X1 U18010 ( .A1(n16031), .A2(n16071), .ZN(n22275) );
  INV_X1 U18011 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20504) );
  NOR3_X1 U18012 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n20504), .A3(n16032), 
        .ZN(n16042) );
  NAND2_X1 U18013 ( .A1(n22214), .A2(n20504), .ZN(n16051) );
  INV_X1 U18014 ( .A(n16090), .ZN(n16033) );
  NAND2_X1 U18015 ( .A1(n16102), .A2(n16033), .ZN(n16089) );
  OR2_X1 U18016 ( .A1(n16089), .A2(n16050), .ZN(n16034) );
  NAND2_X1 U18017 ( .A1(n22273), .A2(n16034), .ZN(n16064) );
  INV_X1 U18018 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n17737) );
  AOI21_X1 U18019 ( .B1(n16051), .B2(n16064), .A(n17737), .ZN(n16041) );
  INV_X1 U18020 ( .A(n16035), .ZN(n16036) );
  OAI21_X1 U18021 ( .B1(n16037), .B2(n16047), .A(n16036), .ZN(n22096) );
  AOI22_X1 U18022 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16311), .ZN(n16039) );
  NAND2_X1 U18023 ( .A1(n22272), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n16038) );
  OAI211_X1 U18024 ( .C1(n22096), .C2(n22278), .A(n16039), .B(n16038), .ZN(
        n16040) );
  AOI211_X1 U18025 ( .C1(n22275), .C2(n16042), .A(n16041), .B(n16040), .ZN(
        n16043) );
  OAI21_X1 U18026 ( .B1(n16186), .B2(n22268), .A(n16043), .ZN(P1_U2818) );
  OAI21_X1 U18027 ( .B1(n16045), .B2(n16046), .A(n16027), .ZN(n16322) );
  AOI21_X1 U18028 ( .B1(n16048), .B2(n16062), .A(n16047), .ZN(n16505) );
  INV_X1 U18029 ( .A(n16325), .ZN(n16049) );
  OAI22_X1 U18030 ( .A1(n16321), .A2(n22246), .B1(n22267), .B2(n16049), .ZN(
        n16053) );
  NOR3_X1 U18031 ( .A1(n16051), .A2(n16090), .A3(n16050), .ZN(n16052) );
  AOI211_X1 U18032 ( .C1(n22272), .C2(P1_EBX_REG_21__SCAN_IN), .A(n16053), .B(
        n16052), .ZN(n16054) );
  OAI21_X1 U18033 ( .B1(n20504), .B2(n16064), .A(n16054), .ZN(n16055) );
  AOI21_X1 U18034 ( .B1(n16505), .B2(n22255), .A(n16055), .ZN(n16056) );
  OAI21_X1 U18035 ( .B1(n16322), .B2(n22268), .A(n16056), .ZN(P1_U2819) );
  INV_X1 U18036 ( .A(n16045), .ZN(n16058) );
  OAI21_X1 U18037 ( .B1(n16059), .B2(n16057), .A(n16058), .ZN(n16331) );
  NAND2_X1 U18038 ( .A1(n11185), .A2(n16060), .ZN(n16061) );
  NAND2_X1 U18039 ( .A1(n16062), .A2(n16061), .ZN(n16121) );
  INV_X1 U18040 ( .A(n16121), .ZN(n16516) );
  AOI21_X1 U18041 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n22275), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n16063) );
  NOR2_X1 U18042 ( .A1(n16064), .A2(n16063), .ZN(n16067) );
  INV_X1 U18043 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n17605) );
  AOI22_X1 U18044 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16334), .ZN(n16065) );
  OAI21_X1 U18045 ( .B1(n22249), .B2(n17605), .A(n16065), .ZN(n16066) );
  AOI211_X1 U18046 ( .C1(n16516), .C2(n22255), .A(n16067), .B(n16066), .ZN(
        n16068) );
  OAI21_X1 U18047 ( .B1(n16331), .B2(n22268), .A(n16068), .ZN(P1_U2820) );
  OAI21_X1 U18048 ( .B1(n16069), .B2(n11726), .A(n16123), .ZN(n16208) );
  INV_X1 U18049 ( .A(n16071), .ZN(n22259) );
  NAND2_X1 U18050 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n22259), .ZN(n16078) );
  AND2_X1 U18051 ( .A1(n22273), .A2(n16078), .ZN(n22258) );
  INV_X1 U18052 ( .A(n20566), .ZN(n16074) );
  INV_X1 U18053 ( .A(n16072), .ZN(n16073) );
  AOI21_X1 U18054 ( .B1(n20567), .B2(n16074), .A(n16073), .ZN(n16075) );
  OR2_X1 U18055 ( .A1(n16126), .A2(n16075), .ZN(n22066) );
  AOI21_X1 U18056 ( .B1(n22263), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n22251), .ZN(n16076) );
  OAI21_X1 U18057 ( .B1(n22066), .B2(n22278), .A(n16076), .ZN(n16080) );
  AOI22_X1 U18058 ( .A1(n22272), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n16339), 
        .B2(n22253), .ZN(n16077) );
  OAI21_X1 U18059 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n16078), .A(n16077), 
        .ZN(n16079) );
  AOI211_X1 U18060 ( .C1(n22258), .C2(P1_REIP_REG_18__SCAN_IN), .A(n16080), 
        .B(n16079), .ZN(n16081) );
  OAI21_X1 U18061 ( .B1(n16208), .B2(n22268), .A(n16081), .ZN(P1_U2822) );
  OAI21_X1 U18062 ( .B1(n16083), .B2(n16082), .A(n15558), .ZN(n16235) );
  OR2_X1 U18063 ( .A1(n20554), .A2(n16086), .ZN(n16087) );
  NAND2_X1 U18064 ( .A1(n16088), .A2(n16087), .ZN(n16554) );
  NAND2_X1 U18065 ( .A1(n22273), .A2(n16089), .ZN(n22217) );
  OAI22_X1 U18066 ( .A1(n22278), .A2(n16554), .B1(n17751), .B2(n22217), .ZN(
        n16095) );
  NOR2_X1 U18067 ( .A1(n22200), .A2(n16090), .ZN(n16091) );
  AOI21_X1 U18068 ( .B1(n16091), .B2(n17751), .A(n22251), .ZN(n16093) );
  AOI22_X1 U18069 ( .A1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n16388), .ZN(n16092) );
  OAI211_X1 U18070 ( .C1(n22249), .C2(n17789), .A(n16093), .B(n16092), .ZN(
        n16094) );
  NOR2_X1 U18071 ( .A1(n16095), .A2(n16094), .ZN(n16096) );
  OAI21_X1 U18072 ( .B1(n16385), .B2(n22268), .A(n16096), .ZN(P1_U2827) );
  INV_X1 U18073 ( .A(n16097), .ZN(n16098) );
  NAND2_X1 U18074 ( .A1(n16098), .A2(n22147), .ZN(n16109) );
  NAND2_X1 U18075 ( .A1(n22263), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16101) );
  INV_X1 U18076 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16099) );
  NAND2_X1 U18077 ( .A1(n22253), .A2(n16099), .ZN(n16100) );
  OAI211_X1 U18078 ( .C1(n14610), .C2(n16102), .A(n16101), .B(n16100), .ZN(
        n16103) );
  AOI21_X1 U18079 ( .B1(n22272), .B2(P1_EBX_REG_1__SCAN_IN), .A(n16103), .ZN(
        n16108) );
  INV_X1 U18080 ( .A(n16104), .ZN(n16105) );
  AOI22_X1 U18081 ( .A1(n22255), .A2(n16105), .B1(n22214), .B2(n14610), .ZN(
        n16107) );
  INV_X1 U18082 ( .A(n22131), .ZN(n22117) );
  OR2_X1 U18083 ( .A1(n14636), .A2(n22117), .ZN(n16106) );
  NAND4_X1 U18084 ( .A1(n16109), .A2(n16108), .A3(n16107), .A4(n16106), .ZN(
        P1_U2839) );
  INV_X1 U18085 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n16110) );
  OAI22_X1 U18086 ( .A1(n16396), .A2(n16143), .B1(n20574), .B2(n16110), .ZN(
        P1_U2841) );
  OAI222_X1 U18087 ( .A1(n16113), .A2(n16146), .B1(n16112), .B2(n20574), .C1(
        n16143), .C2(n16111), .ZN(P1_U2843) );
  INV_X1 U18088 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n17594) );
  OAI222_X1 U18089 ( .A1(n16146), .A2(n16265), .B1(n17594), .B2(n20574), .C1(
        n16447), .C2(n16143), .ZN(P1_U2844) );
  INV_X1 U18090 ( .A(n16272), .ZN(n16114) );
  OAI222_X1 U18091 ( .A1(n16114), .A2(n16146), .B1(n17596), .B2(n20574), .C1(
        n16448), .C2(n16143), .ZN(P1_U2845) );
  INV_X1 U18092 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n17772) );
  OAI222_X1 U18093 ( .A1(n16115), .A2(n16143), .B1(n17772), .B2(n20574), .C1(
        n16281), .C2(n16146), .ZN(P1_U2846) );
  AOI22_X1 U18094 ( .A1(n16474), .A2(n20572), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n16119), .ZN(n16116) );
  OAI21_X1 U18095 ( .B1(n16286), .B2(n16146), .A(n16116), .ZN(P1_U2847) );
  OAI222_X1 U18096 ( .A1(n16295), .A2(n16146), .B1(n17775), .B2(n20574), .C1(
        n16477), .C2(n16143), .ZN(P1_U2848) );
  OAI222_X1 U18097 ( .A1(n16185), .A2(n16146), .B1(n17598), .B2(n20574), .C1(
        n16143), .C2(n16117), .ZN(P1_U2849) );
  INV_X1 U18098 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n16118) );
  OAI222_X1 U18099 ( .A1(n16186), .A2(n16146), .B1(n16118), .B2(n20574), .C1(
        n22096), .C2(n16143), .ZN(P1_U2850) );
  AOI22_X1 U18100 ( .A1(n16505), .A2(n20572), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n16119), .ZN(n16120) );
  OAI21_X1 U18101 ( .B1(n16322), .B2(n16146), .A(n16120), .ZN(P1_U2851) );
  OAI222_X1 U18102 ( .A1(n16331), .A2(n16146), .B1(n20574), .B2(n17605), .C1(
        n16121), .C2(n16143), .ZN(P1_U2852) );
  AND2_X1 U18103 ( .A1(n16123), .A2(n16122), .ZN(n16124) );
  OR2_X1 U18104 ( .A1(n16124), .A2(n16057), .ZN(n22269) );
  OR2_X1 U18105 ( .A1(n16126), .A2(n16125), .ZN(n16127) );
  NAND2_X1 U18106 ( .A1(n11185), .A2(n16127), .ZN(n22279) );
  OAI22_X1 U18107 ( .A1(n22279), .A2(n16143), .B1(n17782), .B2(n20574), .ZN(
        n16128) );
  INV_X1 U18108 ( .A(n16128), .ZN(n16129) );
  OAI21_X1 U18109 ( .B1(n22269), .B2(n16146), .A(n16129), .ZN(P1_U2853) );
  INV_X1 U18110 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n16130) );
  OAI222_X1 U18111 ( .A1(n16208), .A2(n16146), .B1(n16130), .B2(n20574), .C1(
        n22066), .C2(n16143), .ZN(P1_U2854) );
  AND2_X1 U18112 ( .A1(n16135), .A2(n16131), .ZN(n16132) );
  OR2_X1 U18113 ( .A1(n16132), .A2(n16217), .ZN(n22241) );
  INV_X1 U18114 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n22237) );
  AND2_X1 U18115 ( .A1(n11234), .A2(n16133), .ZN(n16134) );
  NOR2_X1 U18116 ( .A1(n20567), .A2(n16134), .ZN(n22086) );
  INV_X1 U18117 ( .A(n22086), .ZN(n22240) );
  OAI222_X1 U18118 ( .A1(n22241), .A2(n16146), .B1(n22237), .B2(n20574), .C1(
        n22240), .C2(n16143), .ZN(P1_U2856) );
  INV_X1 U18119 ( .A(n16135), .ZN(n16136) );
  AOI21_X1 U18120 ( .B1(n16137), .B2(n15618), .A(n16136), .ZN(n16361) );
  NAND2_X1 U18121 ( .A1(n16139), .A2(n16138), .ZN(n16140) );
  NAND2_X1 U18122 ( .A1(n11234), .A2(n16140), .ZN(n22228) );
  OAI22_X1 U18123 ( .A1(n22228), .A2(n16143), .B1(n17481), .B2(n20574), .ZN(
        n16141) );
  AOI21_X1 U18124 ( .B1(n16361), .B2(n14221), .A(n16141), .ZN(n16142) );
  INV_X1 U18125 ( .A(n16142), .ZN(P1_U2857) );
  OAI22_X1 U18126 ( .A1(n16554), .A2(n16143), .B1(n17789), .B2(n20574), .ZN(
        n16144) );
  INV_X1 U18127 ( .A(n16144), .ZN(n16145) );
  OAI21_X1 U18128 ( .B1(n16385), .B2(n16146), .A(n16145), .ZN(P1_U2859) );
  AOI22_X1 U18129 ( .A1(n16225), .A2(n22476), .B1(n16240), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n16147) );
  OAI21_X1 U18130 ( .B1(n16227), .B2(n17654), .A(n16147), .ZN(n16148) );
  AOI21_X1 U18131 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n16229), .A(n16148), .ZN(
        n16149) );
  OAI21_X1 U18132 ( .B1(n16150), .B2(n16243), .A(n16149), .ZN(P1_U2874) );
  NAND2_X1 U18133 ( .A1(n16250), .A2(n16209), .ZN(n16156) );
  INV_X1 U18134 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20661) );
  OR2_X1 U18135 ( .A1(n16158), .A2(n20661), .ZN(n16152) );
  NAND2_X1 U18136 ( .A1(n16158), .A2(DATAI_13_), .ZN(n16151) );
  NAND2_X1 U18137 ( .A1(n16152), .A2(n16151), .ZN(n22469) );
  AOI22_X1 U18138 ( .A1(n16225), .A2(n22469), .B1(n16240), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n16155) );
  NAND2_X1 U18139 ( .A1(n16229), .A2(BUF1_REG_29__SCAN_IN), .ZN(n16154) );
  NAND2_X1 U18140 ( .A1(n16211), .A2(DATAI_29_), .ZN(n16153) );
  NAND4_X1 U18141 ( .A1(n16156), .A2(n16155), .A3(n16154), .A4(n16153), .ZN(
        P1_U2875) );
  INV_X1 U18142 ( .A(n16265), .ZN(n16157) );
  NAND2_X1 U18143 ( .A1(n16157), .A2(n16209), .ZN(n16164) );
  OR2_X1 U18144 ( .A1(n16158), .A2(n20659), .ZN(n16160) );
  NAND2_X1 U18145 ( .A1(n16158), .A2(DATAI_12_), .ZN(n16159) );
  NAND2_X1 U18146 ( .A1(n16160), .A2(n16159), .ZN(n22462) );
  AOI22_X1 U18147 ( .A1(n16225), .A2(n22462), .B1(n16240), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n16163) );
  NAND2_X1 U18148 ( .A1(n16229), .A2(BUF1_REG_28__SCAN_IN), .ZN(n16162) );
  NAND2_X1 U18149 ( .A1(n16211), .A2(DATAI_28_), .ZN(n16161) );
  NAND4_X1 U18150 ( .A1(n16164), .A2(n16163), .A3(n16162), .A4(n16161), .ZN(
        P1_U2876) );
  NAND2_X1 U18151 ( .A1(n16272), .A2(n16209), .ZN(n16168) );
  AOI22_X1 U18152 ( .A1(n16225), .A2(n22454), .B1(n16240), .B2(
        P1_EAX_REG_27__SCAN_IN), .ZN(n16167) );
  NAND2_X1 U18153 ( .A1(n16229), .A2(BUF1_REG_27__SCAN_IN), .ZN(n16166) );
  NAND2_X1 U18154 ( .A1(n16211), .A2(DATAI_27_), .ZN(n16165) );
  NAND4_X1 U18155 ( .A1(n16168), .A2(n16167), .A3(n16166), .A4(n16165), .ZN(
        P1_U2877) );
  AOI22_X1 U18156 ( .A1(n16225), .A2(n22447), .B1(n16240), .B2(
        P1_EAX_REG_26__SCAN_IN), .ZN(n16169) );
  OAI21_X1 U18157 ( .B1(n16227), .B2(n17652), .A(n16169), .ZN(n16170) );
  AOI21_X1 U18158 ( .B1(n16229), .B2(BUF1_REG_26__SCAN_IN), .A(n16170), .ZN(
        n16171) );
  OAI21_X1 U18159 ( .B1(n16281), .B2(n16243), .A(n16171), .ZN(P1_U2878) );
  INV_X1 U18160 ( .A(DATAI_25_), .ZN(n17651) );
  AOI22_X1 U18161 ( .A1(n16225), .A2(n22440), .B1(n16240), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n16172) );
  OAI21_X1 U18162 ( .B1(n16227), .B2(n17651), .A(n16172), .ZN(n16174) );
  NOR2_X1 U18163 ( .A1(n16286), .A2(n16243), .ZN(n16173) );
  AOI211_X1 U18164 ( .C1(n16229), .C2(BUF1_REG_25__SCAN_IN), .A(n16174), .B(
        n16173), .ZN(n16175) );
  INV_X1 U18165 ( .A(n16175), .ZN(P1_U2879) );
  NAND2_X1 U18166 ( .A1(n16176), .A2(n16209), .ZN(n16180) );
  AOI22_X1 U18167 ( .A1(n16225), .A2(n22433), .B1(n16240), .B2(
        P1_EAX_REG_24__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U18168 ( .A1(n16229), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16178) );
  NAND2_X1 U18169 ( .A1(n16211), .A2(DATAI_24_), .ZN(n16177) );
  NAND4_X1 U18170 ( .A1(n16180), .A2(n16179), .A3(n16178), .A4(n16177), .ZN(
        P1_U2880) );
  INV_X1 U18171 ( .A(DATAI_23_), .ZN(n17663) );
  AOI22_X1 U18172 ( .A1(n16225), .A2(n16181), .B1(n16240), .B2(
        P1_EAX_REG_23__SCAN_IN), .ZN(n16182) );
  OAI21_X1 U18173 ( .B1(n16227), .B2(n17663), .A(n16182), .ZN(n16183) );
  AOI21_X1 U18174 ( .B1(n16229), .B2(BUF1_REG_23__SCAN_IN), .A(n16183), .ZN(
        n16184) );
  OAI21_X1 U18175 ( .B1(n16185), .B2(n16243), .A(n16184), .ZN(P1_U2881) );
  INV_X1 U18176 ( .A(n16186), .ZN(n16315) );
  NAND2_X1 U18177 ( .A1(n16315), .A2(n16209), .ZN(n16191) );
  AOI22_X1 U18178 ( .A1(n16225), .A2(n16187), .B1(n16240), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n16190) );
  NAND2_X1 U18179 ( .A1(n16229), .A2(BUF1_REG_22__SCAN_IN), .ZN(n16189) );
  NAND2_X1 U18180 ( .A1(n16211), .A2(DATAI_22_), .ZN(n16188) );
  NAND4_X1 U18181 ( .A1(n16191), .A2(n16190), .A3(n16189), .A4(n16188), .ZN(
        P1_U2882) );
  INV_X1 U18182 ( .A(DATAI_21_), .ZN(n16194) );
  INV_X1 U18183 ( .A(n22418), .ZN(n16192) );
  AOI22_X1 U18184 ( .A1(n16225), .A2(n16192), .B1(n16240), .B2(
        P1_EAX_REG_21__SCAN_IN), .ZN(n16193) );
  OAI21_X1 U18185 ( .B1(n16227), .B2(n16194), .A(n16193), .ZN(n16196) );
  NOR2_X1 U18186 ( .A1(n16322), .A2(n16243), .ZN(n16195) );
  AOI211_X1 U18187 ( .C1(n16229), .C2(BUF1_REG_21__SCAN_IN), .A(n16196), .B(
        n16195), .ZN(n16197) );
  INV_X1 U18188 ( .A(n16197), .ZN(P1_U2883) );
  INV_X1 U18189 ( .A(DATAI_20_), .ZN(n16199) );
  AOI22_X1 U18190 ( .A1(n16225), .A2(n22410), .B1(n16240), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n16198) );
  OAI21_X1 U18191 ( .B1(n16227), .B2(n16199), .A(n16198), .ZN(n16201) );
  NOR2_X1 U18192 ( .A1(n16331), .A2(n16243), .ZN(n16200) );
  AOI211_X1 U18193 ( .C1(n16229), .C2(BUF1_REG_20__SCAN_IN), .A(n16201), .B(
        n16200), .ZN(n16202) );
  INV_X1 U18194 ( .A(n16202), .ZN(P1_U2884) );
  INV_X1 U18195 ( .A(DATAI_19_), .ZN(n17665) );
  INV_X1 U18196 ( .A(n22404), .ZN(n16203) );
  AOI22_X1 U18197 ( .A1(n16225), .A2(n16203), .B1(n16240), .B2(
        P1_EAX_REG_19__SCAN_IN), .ZN(n16204) );
  OAI21_X1 U18198 ( .B1(n17665), .B2(n16227), .A(n16204), .ZN(n16206) );
  NOR2_X1 U18199 ( .A1(n22269), .A2(n16243), .ZN(n16205) );
  AOI211_X1 U18200 ( .C1(n16229), .C2(BUF1_REG_19__SCAN_IN), .A(n16206), .B(
        n16205), .ZN(n16207) );
  INV_X1 U18201 ( .A(n16207), .ZN(P1_U2885) );
  INV_X1 U18202 ( .A(n16208), .ZN(n16343) );
  NAND2_X1 U18203 ( .A1(n16343), .A2(n16209), .ZN(n16215) );
  INV_X1 U18204 ( .A(n22398), .ZN(n16210) );
  AOI22_X1 U18205 ( .A1(n16225), .A2(n16210), .B1(n16240), .B2(
        P1_EAX_REG_18__SCAN_IN), .ZN(n16214) );
  NAND2_X1 U18206 ( .A1(n16229), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16213) );
  NAND2_X1 U18207 ( .A1(n16211), .A2(DATAI_18_), .ZN(n16212) );
  NAND4_X1 U18208 ( .A1(n16215), .A2(n16214), .A3(n16213), .A4(n16212), .ZN(
        P1_U2886) );
  INV_X1 U18209 ( .A(n16217), .ZN(n16218) );
  INV_X1 U18210 ( .A(n22257), .ZN(n16223) );
  INV_X1 U18211 ( .A(DATAI_17_), .ZN(n17667) );
  INV_X1 U18212 ( .A(n22392), .ZN(n16219) );
  AOI22_X1 U18213 ( .A1(n16225), .A2(n16219), .B1(n16240), .B2(
        P1_EAX_REG_17__SCAN_IN), .ZN(n16220) );
  OAI21_X1 U18214 ( .B1(n17667), .B2(n16227), .A(n16220), .ZN(n16221) );
  AOI21_X1 U18215 ( .B1(n16229), .B2(BUF1_REG_17__SCAN_IN), .A(n16221), .ZN(
        n16222) );
  OAI21_X1 U18216 ( .B1(n16223), .B2(n16243), .A(n16222), .ZN(P1_U2887) );
  INV_X1 U18217 ( .A(DATAI_16_), .ZN(n17673) );
  INV_X1 U18218 ( .A(n22386), .ZN(n16224) );
  AOI22_X1 U18219 ( .A1(n16225), .A2(n16224), .B1(n16240), .B2(
        P1_EAX_REG_16__SCAN_IN), .ZN(n16226) );
  OAI21_X1 U18220 ( .B1(n17673), .B2(n16227), .A(n16226), .ZN(n16228) );
  AOI21_X1 U18221 ( .B1(n16229), .B2(BUF1_REG_16__SCAN_IN), .A(n16228), .ZN(
        n16230) );
  OAI21_X1 U18222 ( .B1(n22241), .B2(n16243), .A(n16230), .ZN(P1_U2888) );
  INV_X1 U18223 ( .A(n16361), .ZN(n22229) );
  OAI222_X1 U18224 ( .A1(n22229), .A2(n16243), .B1(n16233), .B2(n16232), .C1(
        n16231), .C2(n14497), .ZN(P1_U2889) );
  AOI22_X1 U18225 ( .A1(n16241), .A2(n22469), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n16240), .ZN(n16234) );
  OAI21_X1 U18226 ( .B1(n16385), .B2(n16243), .A(n16234), .ZN(P1_U2891) );
  INV_X1 U18227 ( .A(n16235), .ZN(n16239) );
  INV_X1 U18228 ( .A(n16236), .ZN(n16238) );
  INV_X1 U18229 ( .A(n22220), .ZN(n16244) );
  AOI22_X1 U18230 ( .A1(n16241), .A2(n22462), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n16240), .ZN(n16242) );
  OAI21_X1 U18231 ( .B1(n16244), .B2(n16243), .A(n16242), .ZN(P1_U2892) );
  XOR2_X1 U18232 ( .A(n16246), .B(n16245), .Z(n16437) );
  NOR2_X1 U18233 ( .A1(n22044), .A2(n20517), .ZN(n16432) );
  AOI21_X1 U18234 ( .B1(n20628), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16432), .ZN(n16247) );
  OAI21_X1 U18235 ( .B1(n20634), .B2(n16248), .A(n16247), .ZN(n16249) );
  AOI21_X1 U18236 ( .B1(n16250), .B2(n20614), .A(n16249), .ZN(n16251) );
  OAI21_X1 U18237 ( .B1(n22280), .B2(n16437), .A(n16251), .ZN(P1_U2970) );
  NAND2_X1 U18238 ( .A1(n22108), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n16439) );
  OAI21_X1 U18239 ( .B1(n16384), .B2(n16252), .A(n16439), .ZN(n16253) );
  AOI21_X1 U18240 ( .B1(n16254), .B2(n20625), .A(n16253), .ZN(n16264) );
  NAND2_X1 U18241 ( .A1(n16255), .A2(n16256), .ZN(n16257) );
  INV_X1 U18242 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16453) );
  MUX2_X1 U18243 ( .A(n20603), .B(n16257), .S(n16453), .Z(n16261) );
  OAI21_X1 U18244 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16258), .A(
        n16257), .ZN(n16260) );
  INV_X1 U18245 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16460) );
  NAND2_X1 U18246 ( .A1(n20603), .A2(n16460), .ZN(n16259) );
  NAND3_X1 U18247 ( .A1(n16261), .A2(n16260), .A3(n16259), .ZN(n16262) );
  XNOR2_X1 U18248 ( .A(n16262), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16438) );
  NAND2_X1 U18249 ( .A1(n16438), .A2(n20595), .ZN(n16263) );
  OAI211_X1 U18250 ( .C1(n16265), .C2(n20630), .A(n16264), .B(n16263), .ZN(
        P1_U2971) );
  NAND2_X1 U18251 ( .A1(n16274), .A2(n16266), .ZN(n16268) );
  XNOR2_X1 U18252 ( .A(n20603), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16267) );
  XNOR2_X1 U18253 ( .A(n16268), .B(n16267), .ZN(n16458) );
  NOR2_X1 U18254 ( .A1(n22044), .A2(n20513), .ZN(n16450) );
  AOI21_X1 U18255 ( .B1(n20628), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16450), .ZN(n16269) );
  OAI21_X1 U18256 ( .B1(n20634), .B2(n16270), .A(n16269), .ZN(n16271) );
  AOI21_X1 U18257 ( .B1(n16272), .B2(n20614), .A(n16271), .ZN(n16273) );
  OAI21_X1 U18258 ( .B1(n16458), .B2(n22280), .A(n16273), .ZN(P1_U2972) );
  OAI21_X1 U18259 ( .B1(n16275), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16274), .ZN(n16468) );
  AND2_X1 U18260 ( .A1(n22108), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n16461) );
  AOI21_X1 U18261 ( .B1(n20628), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16461), .ZN(n16278) );
  NAND2_X1 U18262 ( .A1(n20625), .A2(n16276), .ZN(n16277) );
  OAI211_X1 U18263 ( .C1(n16468), .C2(n22280), .A(n16278), .B(n16277), .ZN(
        n16279) );
  INV_X1 U18264 ( .A(n16279), .ZN(n16280) );
  OAI21_X1 U18265 ( .B1(n16281), .B2(n20630), .A(n16280), .ZN(P1_U2973) );
  NOR2_X1 U18266 ( .A1(n16255), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16283) );
  NAND2_X1 U18267 ( .A1(n20617), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16300) );
  OAI211_X1 U18268 ( .C1(n16283), .C2(n16459), .A(n16282), .B(n16300), .ZN(
        n16284) );
  XNOR2_X1 U18269 ( .A(n16284), .B(n16471), .ZN(n16476) );
  NAND2_X1 U18270 ( .A1(n22108), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n16470) );
  OAI21_X1 U18271 ( .B1(n16384), .B2(n16285), .A(n16470), .ZN(n16288) );
  NOR2_X1 U18272 ( .A1(n16286), .A2(n20630), .ZN(n16287) );
  AOI211_X1 U18273 ( .C1(n20625), .C2(n16289), .A(n16288), .B(n16287), .ZN(
        n16290) );
  OAI21_X1 U18274 ( .B1(n22280), .B2(n16476), .A(n16290), .ZN(P1_U2974) );
  AND2_X1 U18275 ( .A1(n16255), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16292) );
  NOR2_X1 U18276 ( .A1(n16255), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16291) );
  MUX2_X1 U18277 ( .A(n16292), .B(n16291), .S(n20617), .Z(n16293) );
  XNOR2_X1 U18278 ( .A(n16293), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16488) );
  INV_X1 U18279 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16294) );
  NAND2_X1 U18280 ( .A1(n22108), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16482) );
  OAI21_X1 U18281 ( .B1(n16384), .B2(n16294), .A(n16482), .ZN(n16297) );
  NOR2_X1 U18282 ( .A1(n16295), .A2(n20630), .ZN(n16296) );
  AOI211_X1 U18283 ( .C1(n20625), .C2(n16298), .A(n16297), .B(n16296), .ZN(
        n16299) );
  OAI21_X1 U18284 ( .B1(n22280), .B2(n16488), .A(n16299), .ZN(P1_U2975) );
  OAI21_X1 U18285 ( .B1(n20617), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16300), .ZN(n16301) );
  XOR2_X1 U18286 ( .A(n16301), .B(n16255), .Z(n16497) );
  NAND2_X1 U18287 ( .A1(n22108), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n16491) );
  NAND2_X1 U18288 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16302) );
  OAI211_X1 U18289 ( .C1(n20634), .C2(n16303), .A(n16491), .B(n16302), .ZN(
        n16304) );
  AOI21_X1 U18290 ( .B1(n16305), .B2(n20614), .A(n16304), .ZN(n16306) );
  OAI21_X1 U18291 ( .B1(n16497), .B2(n22280), .A(n16306), .ZN(P1_U2976) );
  INV_X1 U18292 ( .A(n16255), .ZN(n16310) );
  INV_X1 U18293 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n22101) );
  AOI21_X1 U18294 ( .B1(n16307), .B2(n16309), .A(n22101), .ZN(n16308) );
  AOI21_X1 U18295 ( .B1(n16310), .B2(n16309), .A(n16308), .ZN(n22095) );
  INV_X1 U18296 ( .A(n16311), .ZN(n16313) );
  AOI22_X1 U18297 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n16312) );
  OAI21_X1 U18298 ( .B1(n20634), .B2(n16313), .A(n16312), .ZN(n16314) );
  AOI21_X1 U18299 ( .B1(n16315), .B2(n20614), .A(n16314), .ZN(n16316) );
  OAI21_X1 U18300 ( .B1(n22095), .B2(n22280), .A(n16316), .ZN(P1_U2977) );
  XNOR2_X1 U18301 ( .A(n20603), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16337) );
  NAND2_X1 U18302 ( .A1(n16338), .A2(n16337), .ZN(n16336) );
  NAND2_X1 U18303 ( .A1(n20617), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16317) );
  NAND2_X1 U18304 ( .A1(n16336), .A2(n16317), .ZN(n16524) );
  MUX2_X1 U18305 ( .A(n16524), .B(n16529), .S(n20603), .Z(n16318) );
  MUX2_X1 U18306 ( .A(n16529), .B(n16524), .S(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(n16319) );
  NAND2_X1 U18307 ( .A1(n16327), .A2(n16319), .ZN(n16320) );
  XNOR2_X1 U18308 ( .A(n16320), .B(n16510), .ZN(n16512) );
  NAND2_X1 U18309 ( .A1(n22108), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16503) );
  OAI21_X1 U18310 ( .B1(n16384), .B2(n16321), .A(n16503), .ZN(n16324) );
  NOR2_X1 U18311 ( .A1(n16322), .A2(n20630), .ZN(n16323) );
  AOI211_X1 U18312 ( .C1(n20625), .C2(n16325), .A(n16324), .B(n16323), .ZN(
        n16326) );
  OAI21_X1 U18313 ( .B1(n22280), .B2(n16512), .A(n16326), .ZN(P1_U2978) );
  OAI21_X1 U18314 ( .B1(n16529), .B2(n16524), .A(n16327), .ZN(n16329) );
  XNOR2_X1 U18315 ( .A(n16329), .B(n16328), .ZN(n16522) );
  INV_X1 U18316 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16330) );
  NAND2_X1 U18317 ( .A1(n22108), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16513) );
  OAI21_X1 U18318 ( .B1(n16384), .B2(n16330), .A(n16513), .ZN(n16333) );
  NOR2_X1 U18319 ( .A1(n16331), .A2(n20630), .ZN(n16332) );
  AOI211_X1 U18320 ( .C1(n20625), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16335) );
  OAI21_X1 U18321 ( .B1(n22280), .B2(n16522), .A(n16335), .ZN(P1_U2979) );
  OAI21_X1 U18322 ( .B1(n16338), .B2(n16337), .A(n16336), .ZN(n22068) );
  INV_X1 U18323 ( .A(n16339), .ZN(n16341) );
  AOI22_X1 U18324 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n16340) );
  OAI21_X1 U18325 ( .B1(n16341), .B2(n20634), .A(n16340), .ZN(n16342) );
  AOI21_X1 U18326 ( .B1(n16343), .B2(n20614), .A(n16342), .ZN(n16344) );
  OAI21_X1 U18327 ( .B1(n22280), .B2(n22068), .A(n16344), .ZN(P1_U2981) );
  OAI21_X1 U18328 ( .B1(n16363), .B2(n16346), .A(n16345), .ZN(n16356) );
  MUX2_X1 U18329 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n16347), .S(
        n20603), .Z(n16357) );
  NOR2_X1 U18330 ( .A1(n16356), .A2(n16357), .ZN(n16355) );
  AOI21_X1 U18331 ( .B1(n20603), .B2(n16347), .A(n16355), .ZN(n16350) );
  INV_X1 U18332 ( .A(n16348), .ZN(n20622) );
  AOI21_X1 U18333 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n20603), .A(
        n20622), .ZN(n16349) );
  XNOR2_X1 U18334 ( .A(n16350), .B(n16349), .ZN(n22087) );
  AOI22_X1 U18335 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16352) );
  NAND2_X1 U18336 ( .A1(n22239), .A2(n20625), .ZN(n16351) );
  OAI211_X1 U18337 ( .C1(n22241), .C2(n20630), .A(n16352), .B(n16351), .ZN(
        n16353) );
  AOI21_X1 U18338 ( .B1(n22087), .B2(n20595), .A(n16353), .ZN(n16354) );
  INV_X1 U18339 ( .A(n16354), .ZN(P1_U2983) );
  AOI21_X1 U18340 ( .B1(n16357), .B2(n16356), .A(n16355), .ZN(n16542) );
  NAND2_X1 U18341 ( .A1(n22108), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16539) );
  NAND2_X1 U18342 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16358) );
  OAI211_X1 U18343 ( .C1(n16359), .C2(n20634), .A(n16539), .B(n16358), .ZN(
        n16360) );
  AOI21_X1 U18344 ( .B1(n16361), .B2(n20614), .A(n16360), .ZN(n16362) );
  OAI21_X1 U18345 ( .B1(n16542), .B2(n22280), .A(n16362), .ZN(P1_U2984) );
  OAI21_X1 U18346 ( .B1(n20620), .B2(n16365), .A(n16364), .ZN(n16367) );
  NAND2_X1 U18347 ( .A1(n16367), .A2(n16366), .ZN(n16369) );
  XNOR2_X1 U18348 ( .A(n20603), .B(n21957), .ZN(n16368) );
  XNOR2_X1 U18349 ( .A(n16369), .B(n16368), .ZN(n21953) );
  INV_X1 U18350 ( .A(n21953), .ZN(n16375) );
  AOI22_X1 U18351 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16370) );
  OAI21_X1 U18352 ( .B1(n20634), .B2(n16371), .A(n16370), .ZN(n16372) );
  AOI21_X1 U18353 ( .B1(n16373), .B2(n20614), .A(n16372), .ZN(n16374) );
  OAI21_X1 U18354 ( .B1(n16375), .B2(n22280), .A(n16374), .ZN(P1_U2985) );
  INV_X1 U18355 ( .A(n16376), .ZN(n16377) );
  AOI21_X1 U18356 ( .B1(n20620), .B2(n16378), .A(n16377), .ZN(n20612) );
  AND2_X1 U18357 ( .A1(n16379), .A2(n16380), .ZN(n20611) );
  NAND2_X1 U18358 ( .A1(n20612), .A2(n20611), .ZN(n20610) );
  NAND2_X1 U18359 ( .A1(n20610), .A2(n16380), .ZN(n16382) );
  XNOR2_X1 U18360 ( .A(n16382), .B(n16381), .ZN(n16558) );
  INV_X1 U18361 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16383) );
  OAI22_X1 U18362 ( .A1(n16384), .A2(n16383), .B1(n22044), .B2(n17751), .ZN(
        n16387) );
  NOR2_X1 U18363 ( .A1(n16385), .A2(n20630), .ZN(n16386) );
  AOI211_X1 U18364 ( .C1(n20625), .C2(n16388), .A(n16387), .B(n16386), .ZN(
        n16389) );
  OAI21_X1 U18365 ( .B1(n22280), .B2(n16558), .A(n16389), .ZN(P1_U2986) );
  OAI21_X1 U18366 ( .B1(n16391), .B2(n16390), .A(n20604), .ZN(n22034) );
  NAND2_X1 U18367 ( .A1(n22034), .A2(n20595), .ZN(n16395) );
  NAND2_X1 U18368 ( .A1(n20628), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16392) );
  NAND2_X1 U18369 ( .A1(n22108), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n22031) );
  NAND2_X1 U18370 ( .A1(n16392), .A2(n22031), .ZN(n16393) );
  AOI21_X1 U18371 ( .B1(n20625), .B2(n22183), .A(n16393), .ZN(n16394) );
  OAI211_X1 U18372 ( .C1(n20630), .C2(n22181), .A(n16395), .B(n16394), .ZN(
        P1_U2990) );
  NOR2_X1 U18373 ( .A1(n16396), .A2(n22067), .ZN(n16419) );
  INV_X1 U18374 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n22024) );
  NOR3_X1 U18375 ( .A1(n22030), .A2(n22024), .A3(n21999), .ZN(n22033) );
  NAND3_X1 U18376 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n22033), .ZN(n22046) );
  NOR2_X1 U18377 ( .A1(n14259), .A2(n22046), .ZN(n22051) );
  NAND2_X1 U18378 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n22051), .ZN(
        n16506) );
  INV_X1 U18379 ( .A(n16506), .ZN(n21958) );
  NOR2_X1 U18380 ( .A1(n21986), .A2(n21992), .ZN(n21981) );
  OAI21_X1 U18381 ( .B1(n14517), .B2(n21969), .A(n21974), .ZN(n21978) );
  NAND2_X1 U18382 ( .A1(n21981), .A2(n21978), .ZN(n22002) );
  NOR2_X1 U18383 ( .A1(n21954), .A2(n22002), .ZN(n22012) );
  NAND2_X1 U18384 ( .A1(n21958), .A2(n22012), .ZN(n16531) );
  NOR2_X1 U18385 ( .A1(n14281), .A2(n22078), .ZN(n22073) );
  NAND4_X1 U18386 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(n22073), .ZN(n16508) );
  NOR2_X1 U18387 ( .A1(n16531), .A2(n16508), .ZN(n16499) );
  NAND2_X1 U18388 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21977) );
  INV_X1 U18389 ( .A(n21977), .ZN(n21980) );
  NAND2_X1 U18390 ( .A1(n21980), .A2(n21981), .ZN(n21995) );
  NOR3_X1 U18391 ( .A1(n21954), .A2(n16506), .A3(n21995), .ZN(n16546) );
  NAND2_X1 U18392 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16546), .ZN(
        n16547) );
  NOR2_X1 U18393 ( .A1(n21957), .A2(n16547), .ZN(n16537) );
  NAND3_X1 U18394 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16537), .A3(
        n22073), .ZN(n16406) );
  OAI21_X1 U18395 ( .B1(n16397), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n16552), .ZN(n22015) );
  AOI21_X1 U18396 ( .B1(n16406), .B2(n22045), .A(n22015), .ZN(n16398) );
  OAI21_X1 U18397 ( .B1(n16499), .B2(n22049), .A(n16398), .ZN(n16525) );
  NOR2_X1 U18398 ( .A1(n22104), .A2(n22101), .ZN(n16409) );
  OAI22_X1 U18399 ( .A1(n22071), .A2(n16409), .B1(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n22049), .ZN(n16399) );
  OR2_X1 U18400 ( .A1(n16525), .A2(n16399), .ZN(n16490) );
  OAI22_X1 U18401 ( .A1(n16532), .A2(n16459), .B1(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n22049), .ZN(n16400) );
  NOR2_X1 U18402 ( .A1(n16490), .A2(n16400), .ZN(n16472) );
  NAND2_X1 U18403 ( .A1(n16472), .A2(n22071), .ZN(n16404) );
  INV_X1 U18404 ( .A(n16404), .ZN(n16405) );
  INV_X1 U18405 ( .A(n16430), .ZN(n16440) );
  INV_X1 U18406 ( .A(n16472), .ZN(n16402) );
  NAND2_X1 U18407 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16401) );
  OAI21_X1 U18408 ( .B1(n16402), .B2(n16401), .A(n16404), .ZN(n16454) );
  OAI21_X1 U18409 ( .B1(n16405), .B2(n16440), .A(n16454), .ZN(n16433) );
  AOI211_X1 U18410 ( .C1(n16414), .C2(n16404), .A(n16403), .B(n16433), .ZN(
        n16425) );
  NOR3_X1 U18411 ( .A1(n16425), .A2(n16405), .A3(n16415), .ZN(n16417) );
  INV_X1 U18412 ( .A(n16406), .ZN(n16498) );
  NAND2_X1 U18413 ( .A1(n16498), .A2(n21979), .ZN(n16509) );
  INV_X1 U18414 ( .A(n16509), .ZN(n16408) );
  NAND2_X1 U18415 ( .A1(n16408), .A2(n16409), .ZN(n16478) );
  NAND2_X1 U18416 ( .A1(n16499), .A2(n16409), .ZN(n16410) );
  OR2_X1 U18417 ( .A1(n22049), .A2(n16410), .ZN(n16411) );
  NAND2_X1 U18418 ( .A1(n16478), .A2(n16411), .ZN(n16489) );
  INV_X1 U18419 ( .A(n16412), .ZN(n16413) );
  NAND2_X1 U18420 ( .A1(n16489), .A2(n16413), .ZN(n16463) );
  NOR3_X1 U18421 ( .A1(n16449), .A2(n16414), .A3(n16430), .ZN(n16422) );
  AND3_X1 U18422 ( .A1(n16422), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16415), .ZN(n16416) );
  NOR4_X1 U18423 ( .A1(n16419), .A2(n16418), .A3(n16417), .A4(n16416), .ZN(
        n16420) );
  OAI21_X1 U18424 ( .B1(n16421), .B2(n22084), .A(n16420), .ZN(P1_U3000) );
  NOR2_X1 U18425 ( .A1(n16422), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16424) );
  OAI21_X1 U18426 ( .B1(n16425), .B2(n16424), .A(n16423), .ZN(n16426) );
  AOI21_X1 U18427 ( .B1(n16427), .B2(n22098), .A(n16426), .ZN(n16428) );
  OAI21_X1 U18428 ( .B1(n16429), .B2(n22084), .A(n16428), .ZN(P1_U3001) );
  NOR3_X1 U18429 ( .A1(n16449), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n16430), .ZN(n16431) );
  AOI211_X1 U18430 ( .C1(n16433), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16432), .B(n16431), .ZN(n16436) );
  NAND2_X1 U18431 ( .A1(n16434), .A2(n22098), .ZN(n16435) );
  OAI211_X1 U18432 ( .C1(n16437), .C2(n22084), .A(n16436), .B(n16435), .ZN(
        P1_U3002) );
  NAND2_X1 U18433 ( .A1(n16438), .A2(n22099), .ZN(n16446) );
  INV_X1 U18434 ( .A(n16454), .ZN(n16444) );
  INV_X1 U18435 ( .A(n16439), .ZN(n16443) );
  NOR3_X1 U18436 ( .A1(n16449), .A2(n16441), .A3(n16440), .ZN(n16442) );
  AOI211_X1 U18437 ( .C1(n16444), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16443), .B(n16442), .ZN(n16445) );
  OAI211_X1 U18438 ( .C1(n22067), .C2(n16447), .A(n16446), .B(n16445), .ZN(
        P1_U3003) );
  INV_X1 U18439 ( .A(n16448), .ZN(n16456) );
  INV_X1 U18440 ( .A(n16449), .ZN(n16451) );
  AOI21_X1 U18441 ( .B1(n16451), .B2(n16453), .A(n16450), .ZN(n16452) );
  OAI21_X1 U18442 ( .B1(n16454), .B2(n16453), .A(n16452), .ZN(n16455) );
  AOI21_X1 U18443 ( .B1(n16456), .B2(n22098), .A(n16455), .ZN(n16457) );
  OAI21_X1 U18444 ( .B1(n16458), .B2(n22084), .A(n16457), .ZN(P1_U3004) );
  NAND3_X1 U18445 ( .A1(n16489), .A2(n16459), .A3(n16471), .ZN(n16469) );
  AOI21_X1 U18446 ( .B1(n16469), .B2(n16472), .A(n16460), .ZN(n16465) );
  INV_X1 U18447 ( .A(n16461), .ZN(n16462) );
  OAI21_X1 U18448 ( .B1(n16463), .B2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16462), .ZN(n16464) );
  AOI211_X1 U18449 ( .C1(n16466), .C2(n22098), .A(n16465), .B(n16464), .ZN(
        n16467) );
  OAI21_X1 U18450 ( .B1(n16468), .B2(n22084), .A(n16467), .ZN(P1_U3005) );
  OAI211_X1 U18451 ( .C1(n16472), .C2(n16471), .A(n16470), .B(n16469), .ZN(
        n16473) );
  AOI21_X1 U18452 ( .B1(n16474), .B2(n22098), .A(n16473), .ZN(n16475) );
  OAI21_X1 U18453 ( .B1(n16476), .B2(n22084), .A(n16475), .ZN(P1_U3006) );
  INV_X1 U18454 ( .A(n16477), .ZN(n16486) );
  INV_X1 U18455 ( .A(n16478), .ZN(n16480) );
  AOI21_X1 U18456 ( .B1(n16480), .B2(n16479), .A(n16490), .ZN(n16484) );
  NAND3_X1 U18457 ( .A1(n16489), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16483), .ZN(n16481) );
  OAI211_X1 U18458 ( .C1(n16484), .C2(n16483), .A(n16482), .B(n16481), .ZN(
        n16485) );
  AOI21_X1 U18459 ( .B1(n16486), .B2(n22098), .A(n16485), .ZN(n16487) );
  OAI21_X1 U18460 ( .B1(n16488), .B2(n22084), .A(n16487), .ZN(P1_U3007) );
  INV_X1 U18461 ( .A(n16489), .ZN(n16493) );
  NAND2_X1 U18462 ( .A1(n16490), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16492) );
  OAI211_X1 U18463 ( .C1(n16493), .C2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16492), .B(n16491), .ZN(n16494) );
  AOI21_X1 U18464 ( .B1(n16495), .B2(n22098), .A(n16494), .ZN(n16496) );
  OAI21_X1 U18465 ( .B1(n16497), .B2(n22084), .A(n16496), .ZN(P1_U3008) );
  AOI21_X1 U18466 ( .B1(n16532), .B2(n16499), .A(n16498), .ZN(n16501) );
  NAND2_X1 U18467 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16500) );
  OR2_X1 U18468 ( .A1(n16501), .A2(n16500), .ZN(n16502) );
  INV_X1 U18469 ( .A(n22071), .ZN(n22014) );
  AOI21_X1 U18470 ( .B1(n16502), .B2(n22014), .A(n22015), .ZN(n22102) );
  OAI21_X1 U18471 ( .B1(n22102), .B2(n16510), .A(n16503), .ZN(n16504) );
  AOI21_X1 U18472 ( .B1(n16505), .B2(n22098), .A(n16504), .ZN(n16511) );
  NAND2_X1 U18473 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16546), .ZN(
        n16549) );
  INV_X1 U18474 ( .A(n16549), .ZN(n16507) );
  INV_X1 U18475 ( .A(n22012), .ZN(n22004) );
  NOR3_X1 U18476 ( .A1(n16506), .A2(n22049), .A3(n22004), .ZN(n16535) );
  AOI21_X1 U18477 ( .B1(n16507), .B2(n16550), .A(n16535), .ZN(n16543) );
  OR2_X1 U18478 ( .A1(n16508), .A2(n16543), .ZN(n16518) );
  NAND2_X1 U18479 ( .A1(n16518), .A2(n16509), .ZN(n16528) );
  NAND4_X1 U18480 ( .A1(n16528), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n16510), .ZN(n22103) );
  OAI211_X1 U18481 ( .C1(n16512), .C2(n22084), .A(n16511), .B(n22103), .ZN(
        P1_U3010) );
  INV_X1 U18482 ( .A(n16513), .ZN(n16515) );
  INV_X1 U18483 ( .A(n16528), .ZN(n22105) );
  NOR3_X1 U18484 ( .A1(n22105), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16529), .ZN(n16514) );
  AOI211_X1 U18485 ( .C1(n22098), .C2(n16516), .A(n16515), .B(n16514), .ZN(
        n16521) );
  INV_X1 U18486 ( .A(n16548), .ZN(n16517) );
  AOI21_X1 U18487 ( .B1(n16518), .B2(n16517), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16519) );
  OAI21_X1 U18488 ( .B1(n16519), .B2(n16525), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16520) );
  OAI211_X1 U18489 ( .C1(n16522), .C2(n22084), .A(n16521), .B(n16520), .ZN(
        P1_U3011) );
  XNOR2_X1 U18490 ( .A(n20603), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n16523) );
  XNOR2_X1 U18491 ( .A(n16524), .B(n16523), .ZN(n20629) );
  AOI22_X1 U18492 ( .A1(n16525), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n22108), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n16526) );
  OAI21_X1 U18493 ( .B1(n22279), .B2(n22067), .A(n16526), .ZN(n16527) );
  AOI21_X1 U18494 ( .B1(n16529), .B2(n16528), .A(n16527), .ZN(n16530) );
  OAI21_X1 U18495 ( .B1(n20629), .B2(n22084), .A(n16530), .ZN(P1_U3012) );
  NAND2_X1 U18496 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16534) );
  NAND2_X1 U18497 ( .A1(n22005), .A2(n16531), .ZN(n16551) );
  OAI21_X1 U18498 ( .B1(n16537), .B2(n16532), .A(n16551), .ZN(n16533) );
  AOI211_X1 U18499 ( .C1(n22005), .C2(n16534), .A(n22015), .B(n16533), .ZN(
        n22070) );
  INV_X1 U18500 ( .A(n22070), .ZN(n22088) );
  INV_X1 U18501 ( .A(n16534), .ZN(n16536) );
  AOI22_X1 U18502 ( .A1(n16537), .A2(n21979), .B1(n16536), .B2(n16535), .ZN(
        n22079) );
  NOR2_X1 U18503 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n22079), .ZN(
        n22089) );
  INV_X1 U18504 ( .A(n22089), .ZN(n16538) );
  OAI211_X1 U18505 ( .C1(n22228), .C2(n22067), .A(n16539), .B(n16538), .ZN(
        n16540) );
  AOI21_X1 U18506 ( .B1(n22088), .B2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n16540), .ZN(n16541) );
  OAI21_X1 U18507 ( .B1(n16542), .B2(n22084), .A(n16541), .ZN(P1_U3016) );
  AND2_X1 U18508 ( .A1(n16548), .A2(n16547), .ZN(n16545) );
  NOR2_X1 U18509 ( .A1(n22044), .A2(n17751), .ZN(n16544) );
  NOR2_X1 U18510 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16543), .ZN(
        n21960) );
  AOI211_X1 U18511 ( .C1(n16546), .C2(n16545), .A(n16544), .B(n21960), .ZN(
        n16557) );
  AOI22_X1 U18512 ( .A1(n16550), .A2(n16549), .B1(n16548), .B2(n16547), .ZN(
        n16553) );
  NAND3_X1 U18513 ( .A1(n16553), .A2(n16552), .A3(n16551), .ZN(n21959) );
  INV_X1 U18514 ( .A(n16554), .ZN(n16555) );
  AOI22_X1 U18515 ( .A1(n21959), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16555), .B2(n22098), .ZN(n16556) );
  OAI211_X1 U18516 ( .C1(n16558), .C2(n22084), .A(n16557), .B(n16556), .ZN(
        P1_U3018) );
  NOR2_X1 U18517 ( .A1(n16560), .A2(n16559), .ZN(n22301) );
  AOI21_X1 U18518 ( .B1(n17438), .B2(n16565), .A(n22301), .ZN(n16561) );
  OAI21_X1 U18519 ( .B1(n11155), .B2(n22607), .A(n16561), .ZN(n16563) );
  MUX2_X1 U18520 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16563), .S(
        n17476), .Z(P1_U3478) );
  AOI21_X1 U18521 ( .B1(n16565), .B2(n16564), .A(n22612), .ZN(n16566) );
  OAI21_X1 U18522 ( .B1(n16568), .B2(n16567), .A(n16566), .ZN(n16569) );
  MUX2_X1 U18523 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16569), .S(
        n17476), .Z(P1_U3475) );
  INV_X1 U18524 ( .A(n16570), .ZN(n17437) );
  INV_X1 U18525 ( .A(n16571), .ZN(n16575) );
  NOR3_X1 U18526 ( .A1(n16573), .A2(n16572), .A3(n13032), .ZN(n16574) );
  AOI211_X1 U18527 ( .C1(n22593), .C2(n17437), .A(n16575), .B(n16574), .ZN(
        n17440) );
  NAND2_X1 U18528 ( .A1(n16577), .A2(n16576), .ZN(n16581) );
  NAND3_X1 U18529 ( .A1(n16579), .A2(n22298), .A3(n16578), .ZN(n16580) );
  OAI211_X1 U18530 ( .C1(n17440), .C2(n22289), .A(n16581), .B(n16580), .ZN(
        n16582) );
  MUX2_X1 U18531 ( .A(n16582), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n22286), .Z(P1_U3473) );
  NOR2_X1 U18532 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16583), .ZN(
        n16594) );
  INV_X1 U18533 ( .A(n16594), .ZN(n16619) );
  INV_X1 U18534 ( .A(n22569), .ZN(n22589) );
  NOR2_X1 U18535 ( .A1(n16585), .A2(n16584), .ZN(n22493) );
  INV_X1 U18536 ( .A(n22493), .ZN(n16587) );
  NAND3_X1 U18537 ( .A1(n16590), .A2(n22563), .A3(n14636), .ZN(n16586) );
  OAI21_X1 U18538 ( .B1(n22589), .B2(n16587), .A(n16586), .ZN(n16617) );
  AOI21_X1 U18539 ( .B1(n16623), .B2(n16588), .A(n22590), .ZN(n16589) );
  AOI21_X1 U18540 ( .B1(n16590), .B2(n14636), .A(n16589), .ZN(n16591) );
  NOR2_X1 U18541 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n16591), .ZN(n16593) );
  AOI22_X1 U18542 ( .A1(n16617), .A2(n22609), .B1(
        P1_INSTQUEUE_REG_4__0__SCAN_IN), .B2(n16616), .ZN(n16595) );
  OAI21_X1 U18543 ( .B1(n22572), .B2(n16619), .A(n16595), .ZN(n16596) );
  AOI21_X1 U18544 ( .B1(n16621), .B2(n22616), .A(n16596), .ZN(n16597) );
  OAI21_X1 U18545 ( .B1(n16623), .B2(n22619), .A(n16597), .ZN(P1_U3065) );
  AOI22_X1 U18546 ( .A1(n16617), .A2(n22642), .B1(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n16616), .ZN(n16598) );
  OAI21_X1 U18547 ( .B1(n22632), .B2(n16619), .A(n16598), .ZN(n16599) );
  AOI21_X1 U18548 ( .B1(n16621), .B2(n22643), .A(n16599), .ZN(n16600) );
  OAI21_X1 U18549 ( .B1(n16623), .B2(n22646), .A(n16600), .ZN(P1_U3066) );
  AOI22_X1 U18550 ( .A1(n16617), .A2(n22669), .B1(
        P1_INSTQUEUE_REG_4__2__SCAN_IN), .B2(n16616), .ZN(n16601) );
  OAI21_X1 U18551 ( .B1(n22659), .B2(n16619), .A(n16601), .ZN(n16602) );
  AOI21_X1 U18552 ( .B1(n16621), .B2(n22670), .A(n16602), .ZN(n16603) );
  OAI21_X1 U18553 ( .B1(n16623), .B2(n22673), .A(n16603), .ZN(P1_U3067) );
  AOI22_X1 U18554 ( .A1(n16617), .A2(n22696), .B1(
        P1_INSTQUEUE_REG_4__3__SCAN_IN), .B2(n16616), .ZN(n16604) );
  OAI21_X1 U18555 ( .B1(n22686), .B2(n16619), .A(n16604), .ZN(n16605) );
  AOI21_X1 U18556 ( .B1(n16621), .B2(n22697), .A(n16605), .ZN(n16606) );
  OAI21_X1 U18557 ( .B1(n16623), .B2(n22700), .A(n16606), .ZN(P1_U3068) );
  AOI22_X1 U18558 ( .A1(n16617), .A2(n22723), .B1(
        P1_INSTQUEUE_REG_4__4__SCAN_IN), .B2(n16616), .ZN(n16607) );
  OAI21_X1 U18559 ( .B1(n22713), .B2(n16619), .A(n16607), .ZN(n16608) );
  AOI21_X1 U18560 ( .B1(n16621), .B2(n22724), .A(n16608), .ZN(n16609) );
  OAI21_X1 U18561 ( .B1(n16623), .B2(n22727), .A(n16609), .ZN(P1_U3069) );
  AOI22_X1 U18562 ( .A1(n16617), .A2(n22750), .B1(
        P1_INSTQUEUE_REG_4__5__SCAN_IN), .B2(n16616), .ZN(n16610) );
  OAI21_X1 U18563 ( .B1(n22740), .B2(n16619), .A(n16610), .ZN(n16611) );
  AOI21_X1 U18564 ( .B1(n16621), .B2(n22751), .A(n16611), .ZN(n16612) );
  OAI21_X1 U18565 ( .B1(n16623), .B2(n22754), .A(n16612), .ZN(P1_U3070) );
  AOI22_X1 U18566 ( .A1(n16617), .A2(n22777), .B1(
        P1_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n16616), .ZN(n16613) );
  OAI21_X1 U18567 ( .B1(n22767), .B2(n16619), .A(n16613), .ZN(n16614) );
  AOI21_X1 U18568 ( .B1(n16621), .B2(n22778), .A(n16614), .ZN(n16615) );
  OAI21_X1 U18569 ( .B1(n16623), .B2(n22781), .A(n16615), .ZN(P1_U3071) );
  AOI22_X1 U18570 ( .A1(n16617), .A2(n22841), .B1(
        P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n16616), .ZN(n16618) );
  OAI21_X1 U18571 ( .B1(n22821), .B2(n16619), .A(n16618), .ZN(n16620) );
  AOI21_X1 U18572 ( .B1(n16621), .B2(n22843), .A(n16620), .ZN(n16622) );
  OAI21_X1 U18573 ( .B1(n16623), .B2(n22849), .A(n16622), .ZN(P1_U3072) );
  OAI21_X1 U18574 ( .B1(n16624), .B2(n16625), .A(n16710), .ZN(n17155) );
  NAND2_X1 U18575 ( .A1(n16626), .A2(n16627), .ZN(n16628) );
  NAND2_X1 U18576 ( .A1(n11161), .A2(n16628), .ZN(n17161) );
  AOI22_X1 U18577 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19237), .ZN(n16631) );
  AOI22_X1 U18578 ( .A1(n16629), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16630) );
  OAI211_X1 U18579 ( .C1(n17161), .C2(n19268), .A(n16631), .B(n16630), .ZN(
        n16635) );
  AOI211_X1 U18580 ( .C1(n16905), .C2(n16633), .A(n16632), .B(n19316), .ZN(
        n16634) );
  NOR2_X1 U18581 ( .A1(n16635), .A2(n16634), .ZN(n16636) );
  OAI21_X1 U18582 ( .B1(n17155), .B2(n19166), .A(n16636), .ZN(P2_U2834) );
  AOI211_X1 U18583 ( .C1(n16639), .C2(n16638), .A(n16637), .B(n19316), .ZN(
        n16640) );
  INV_X1 U18584 ( .A(n16640), .ZN(n16651) );
  AND2_X1 U18585 ( .A1(n11182), .A2(n16641), .ZN(n16642) );
  NOR2_X1 U18586 ( .A1(n16624), .A2(n16642), .ZN(n17178) );
  OAI21_X1 U18587 ( .B1(n16644), .B2(n16643), .A(n16626), .ZN(n20116) );
  NAND2_X1 U18588 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19239), .ZN(
        n16645) );
  OAI21_X1 U18589 ( .B1(n19210), .B2(n16646), .A(n16645), .ZN(n16647) );
  AOI21_X1 U18590 ( .B1(P2_REIP_REG_20__SCAN_IN), .B2(n19237), .A(n16647), 
        .ZN(n16648) );
  OAI21_X1 U18591 ( .B1(n20116), .B2(n19268), .A(n16648), .ZN(n16649) );
  AOI21_X1 U18592 ( .B1(n17178), .B2(n19251), .A(n16649), .ZN(n16650) );
  OAI211_X1 U18593 ( .C1(n19215), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        P2_U2835) );
  MUX2_X1 U18594 ( .A(n19252), .B(P2_EBX_REG_31__SCAN_IN), .S(n15538), .Z(
        P2_U2856) );
  XOR2_X1 U18595 ( .A(n16654), .B(n16653), .Z(n16655) );
  XNOR2_X1 U18596 ( .A(n16656), .B(n16655), .ZN(n16741) );
  OAI21_X1 U18597 ( .B1(n16659), .B2(n16658), .A(n16657), .ZN(n17072) );
  NOR2_X1 U18598 ( .A1(n17072), .A2(n15538), .ZN(n16660) );
  AOI21_X1 U18599 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n15538), .A(n16660), .ZN(
        n16661) );
  OAI21_X1 U18600 ( .B1(n16741), .B2(n16732), .A(n16661), .ZN(P2_U2858) );
  NOR2_X1 U18601 ( .A1(n11186), .A2(n16662), .ZN(n16664) );
  XNOR2_X1 U18602 ( .A(n16664), .B(n16663), .ZN(n16746) );
  NAND2_X1 U18603 ( .A1(n15538), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16666) );
  NAND2_X1 U18604 ( .A1(n19228), .A2(n16700), .ZN(n16665) );
  OAI211_X1 U18605 ( .C1(n16746), .C2(n16732), .A(n16666), .B(n16665), .ZN(
        P2_U2859) );
  XOR2_X1 U18606 ( .A(n16670), .B(n16669), .Z(n16755) );
  NAND2_X1 U18607 ( .A1(n15538), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16675) );
  INV_X1 U18608 ( .A(n16671), .ZN(n16672) );
  AOI21_X1 U18609 ( .B1(n16673), .B2(n16680), .A(n16672), .ZN(n19213) );
  NAND2_X1 U18610 ( .A1(n19213), .A2(n16700), .ZN(n16674) );
  OAI211_X1 U18611 ( .C1(n16755), .C2(n16732), .A(n16675), .B(n16674), .ZN(
        P2_U2860) );
  OAI21_X1 U18612 ( .B1(n16678), .B2(n16677), .A(n16676), .ZN(n16756) );
  INV_X1 U18613 ( .A(n16680), .ZN(n16681) );
  AOI21_X1 U18614 ( .B1(n16682), .B2(n16679), .A(n16681), .ZN(n19199) );
  INV_X1 U18615 ( .A(n19199), .ZN(n17105) );
  NOR2_X1 U18616 ( .A1(n17105), .A2(n15538), .ZN(n16683) );
  AOI21_X1 U18617 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n15538), .A(n16683), .ZN(
        n16684) );
  OAI21_X1 U18618 ( .B1(n16756), .B2(n16732), .A(n16684), .ZN(P2_U2861) );
  OAI21_X1 U18619 ( .B1(n16687), .B2(n16686), .A(n16685), .ZN(n16768) );
  OR2_X1 U18620 ( .A1(n16697), .A2(n16688), .ZN(n16689) );
  NAND2_X1 U18621 ( .A1(n16679), .A2(n16689), .ZN(n19186) );
  NOR2_X1 U18622 ( .A1(n19186), .A2(n15538), .ZN(n16690) );
  AOI21_X1 U18623 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n15538), .A(n16690), .ZN(
        n16691) );
  OAI21_X1 U18624 ( .B1(n16768), .B2(n16732), .A(n16691), .ZN(P2_U2862) );
  OAI21_X1 U18625 ( .B1(n16694), .B2(n16693), .A(n16692), .ZN(n16777) );
  NAND2_X1 U18626 ( .A1(n15538), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16702) );
  INV_X1 U18627 ( .A(n16695), .ZN(n16699) );
  INV_X1 U18628 ( .A(n16696), .ZN(n16698) );
  AOI21_X1 U18629 ( .B1(n16699), .B2(n16698), .A(n16697), .ZN(n19176) );
  NAND2_X1 U18630 ( .A1(n19176), .A2(n16700), .ZN(n16701) );
  OAI211_X1 U18631 ( .C1(n16777), .C2(n16732), .A(n16702), .B(n16701), .ZN(
        P2_U2863) );
  XNOR2_X1 U18632 ( .A(n16703), .B(n16704), .ZN(n16787) );
  AND2_X1 U18633 ( .A1(n11183), .A2(n16705), .ZN(n16706) );
  OR2_X1 U18634 ( .A1(n16706), .A2(n16696), .ZN(n19167) );
  NOR2_X1 U18635 ( .A1(n19167), .A2(n15538), .ZN(n16707) );
  AOI21_X1 U18636 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15538), .A(n16707), .ZN(
        n16708) );
  OAI21_X1 U18637 ( .B1(n16787), .B2(n16732), .A(n16708), .ZN(P2_U2864) );
  NAND2_X1 U18638 ( .A1(n16710), .A2(n16709), .ZN(n16711) );
  AND2_X1 U18639 ( .A1(n11183), .A2(n16711), .ZN(n19152) );
  INV_X1 U18640 ( .A(n19152), .ZN(n16716) );
  OR2_X1 U18641 ( .A1(n16717), .A2(n16712), .ZN(n16713) );
  AND2_X1 U18642 ( .A1(n16703), .A2(n16713), .ZN(n20020) );
  NAND2_X1 U18643 ( .A1(n20020), .A2(n16724), .ZN(n16715) );
  NAND2_X1 U18644 ( .A1(n15538), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16714) );
  OAI211_X1 U18645 ( .C1(n16716), .C2(n15538), .A(n16715), .B(n16714), .ZN(
        P2_U2865) );
  AOI21_X1 U18646 ( .B1(n16718), .B2(n16721), .A(n16717), .ZN(n16792) );
  NAND2_X1 U18647 ( .A1(n16792), .A2(n16724), .ZN(n16720) );
  NAND2_X1 U18648 ( .A1(n15538), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n16719) );
  OAI211_X1 U18649 ( .C1(n15538), .C2(n17155), .A(n16720), .B(n16719), .ZN(
        P2_U2866) );
  INV_X1 U18650 ( .A(n17178), .ZN(n16727) );
  INV_X1 U18651 ( .A(n16721), .ZN(n16722) );
  AOI21_X1 U18652 ( .B1(n16723), .B2(n15635), .A(n16722), .ZN(n20120) );
  NAND2_X1 U18653 ( .A1(n20120), .A2(n16724), .ZN(n16726) );
  NAND2_X1 U18654 ( .A1(n15538), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n16725) );
  OAI211_X1 U18655 ( .C1(n15538), .C2(n16727), .A(n16726), .B(n16725), .ZN(
        P2_U2867) );
  NAND2_X1 U18656 ( .A1(n11228), .A2(n16728), .ZN(n16729) );
  NAND2_X1 U18657 ( .A1(n11182), .A2(n16729), .ZN(n19137) );
  NOR2_X1 U18658 ( .A1(n19137), .A2(n15538), .ZN(n16730) );
  AOI21_X1 U18659 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15538), .A(n16730), .ZN(
        n16731) );
  OAI21_X1 U18660 ( .B1(n16733), .B2(n16732), .A(n16731), .ZN(P2_U2868) );
  XOR2_X1 U18661 ( .A(n16734), .B(n15808), .Z(n19240) );
  AOI22_X1 U18662 ( .A1(n20114), .A2(BUF2_REG_29__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U18663 ( .A1(n20111), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n16735) );
  OAI211_X1 U18664 ( .C1(n16738), .C2(n16737), .A(n16736), .B(n16735), .ZN(
        n16739) );
  AOI21_X1 U18665 ( .B1(n19240), .B2(n20117), .A(n16739), .ZN(n16740) );
  OAI21_X1 U18666 ( .B1(n16741), .B2(n20065), .A(n16740), .ZN(P2_U2890) );
  AOI22_X1 U18667 ( .A1(n20113), .A2(n19809), .B1(n20111), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16743) );
  AOI22_X1 U18668 ( .A1(n20114), .A2(BUF2_REG_28__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n16742) );
  OAI211_X1 U18669 ( .C1(n19225), .C2(n16790), .A(n16743), .B(n16742), .ZN(
        n16744) );
  INV_X1 U18670 ( .A(n16744), .ZN(n16745) );
  OAI21_X1 U18671 ( .B1(n16746), .B2(n20065), .A(n16745), .ZN(P2_U2891) );
  NOR2_X1 U18672 ( .A1(n16747), .A2(n16748), .ZN(n16749) );
  OR2_X1 U18673 ( .A1(n14160), .A2(n16749), .ZN(n19223) );
  AOI22_X1 U18674 ( .A1(n20113), .A2(n16750), .B1(n20111), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16752) );
  AOI22_X1 U18675 ( .A1(n20114), .A2(BUF2_REG_27__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n16751) );
  OAI211_X1 U18676 ( .C1(n19223), .C2(n16790), .A(n16752), .B(n16751), .ZN(
        n16753) );
  INV_X1 U18677 ( .A(n16753), .ZN(n16754) );
  OAI21_X1 U18678 ( .B1(n16755), .B2(n20065), .A(n16754), .ZN(P2_U2892) );
  OR2_X1 U18679 ( .A1(n16756), .A2(n20065), .ZN(n16762) );
  AOI22_X1 U18680 ( .A1(n20113), .A2(n19812), .B1(n20111), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16761) );
  AOI22_X1 U18681 ( .A1(n20114), .A2(BUF2_REG_26__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n16760) );
  AND2_X1 U18682 ( .A1(n11162), .A2(n16757), .ZN(n16758) );
  NOR2_X1 U18683 ( .A1(n16747), .A2(n16758), .ZN(n19198) );
  NAND2_X1 U18684 ( .A1(n19198), .A2(n20117), .ZN(n16759) );
  NAND4_X1 U18685 ( .A1(n16762), .A2(n16761), .A3(n16760), .A4(n16759), .ZN(
        P2_U2893) );
  XNOR2_X1 U18686 ( .A(n11208), .B(n16763), .ZN(n19187) );
  AOI22_X1 U18687 ( .A1(n20113), .A2(n19815), .B1(n20111), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16765) );
  AOI22_X1 U18688 ( .A1(n20114), .A2(BUF2_REG_25__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n16764) );
  OAI211_X1 U18689 ( .C1(n19187), .C2(n16790), .A(n16765), .B(n16764), .ZN(
        n16766) );
  INV_X1 U18690 ( .A(n16766), .ZN(n16767) );
  OAI21_X1 U18691 ( .B1(n16768), .B2(n20065), .A(n16767), .ZN(P2_U2894) );
  OR2_X1 U18692 ( .A1(n16781), .A2(n16769), .ZN(n16770) );
  NAND2_X1 U18693 ( .A1(n11208), .A2(n16770), .ZN(n19174) );
  INV_X1 U18694 ( .A(n16771), .ZN(n16772) );
  AOI22_X1 U18695 ( .A1(n20113), .A2(n16772), .B1(n20111), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16774) );
  AOI22_X1 U18696 ( .A1(n20114), .A2(BUF2_REG_24__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16773) );
  OAI211_X1 U18697 ( .C1(n19174), .C2(n16790), .A(n16774), .B(n16773), .ZN(
        n16775) );
  INV_X1 U18698 ( .A(n16775), .ZN(n16776) );
  OAI21_X1 U18699 ( .B1(n16777), .B2(n20065), .A(n16776), .ZN(P2_U2895) );
  NOR2_X1 U18700 ( .A1(n16778), .A2(n16779), .ZN(n16780) );
  OR2_X1 U18701 ( .A1(n16781), .A2(n16780), .ZN(n19165) );
  INV_X1 U18702 ( .A(n19818), .ZN(n16782) );
  AOI22_X1 U18703 ( .A1(n20113), .A2(n16782), .B1(n20111), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16784) );
  AOI22_X1 U18704 ( .A1(n20114), .A2(BUF2_REG_23__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n16783) );
  OAI211_X1 U18705 ( .C1(n19165), .C2(n16790), .A(n16784), .B(n16783), .ZN(
        n16785) );
  INV_X1 U18706 ( .A(n16785), .ZN(n16786) );
  OAI21_X1 U18707 ( .B1(n16787), .B2(n20065), .A(n16786), .ZN(P2_U2896) );
  AOI22_X1 U18708 ( .A1(n20114), .A2(BUF2_REG_21__SCAN_IN), .B1(n20115), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16789) );
  INV_X1 U18709 ( .A(n20072), .ZN(n20063) );
  AOI22_X1 U18710 ( .A1(n20113), .A2(n20063), .B1(n20111), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16788) );
  OAI211_X1 U18711 ( .C1(n17161), .C2(n16790), .A(n16789), .B(n16788), .ZN(
        n16791) );
  AOI21_X1 U18712 ( .B1(n16792), .B2(n20119), .A(n16791), .ZN(n16793) );
  INV_X1 U18713 ( .A(n16793), .ZN(P2_U2898) );
  NAND2_X1 U18714 ( .A1(n16794), .A2(n20119), .ZN(n16803) );
  AOI22_X1 U18715 ( .A1(n20114), .A2(BUF2_REG_17__SCAN_IN), .B1(n20113), .B2(
        n16795), .ZN(n16802) );
  NAND2_X1 U18716 ( .A1(n16796), .A2(n16797), .ZN(n16798) );
  AND2_X1 U18717 ( .A1(n16799), .A2(n16798), .ZN(n19116) );
  AOI22_X1 U18718 ( .A1(n19116), .A2(n20117), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n20111), .ZN(n16801) );
  NAND2_X1 U18719 ( .A1(n20115), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16800) );
  NAND4_X1 U18720 ( .A1(n16803), .A2(n16802), .A3(n16801), .A4(n16800), .ZN(
        P2_U2902) );
  OR2_X1 U18721 ( .A1(n16804), .A2(n20065), .ZN(n16812) );
  INV_X1 U18722 ( .A(n20292), .ZN(n16805) );
  AOI22_X1 U18723 ( .A1(n20114), .A2(BUF2_REG_16__SCAN_IN), .B1(n20113), .B2(
        n16805), .ZN(n16811) );
  OR2_X1 U18724 ( .A1(n16807), .A2(n16806), .ZN(n16808) );
  AND2_X1 U18725 ( .A1(n16796), .A2(n16808), .ZN(n19104) );
  AOI22_X1 U18726 ( .A1(n20117), .A2(n19104), .B1(n20111), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n16810) );
  NAND2_X1 U18727 ( .A1(n20115), .A2(BUF1_REG_16__SCAN_IN), .ZN(n16809) );
  NAND4_X1 U18728 ( .A1(n16812), .A2(n16811), .A3(n16810), .A4(n16809), .ZN(
        P2_U2903) );
  NOR2_X1 U18729 ( .A1(n16814), .A2(n16813), .ZN(n16816) );
  XOR2_X1 U18730 ( .A(n16816), .B(n16815), .Z(n17086) );
  AOI21_X1 U18731 ( .B1(n16828), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16817) );
  NOR2_X1 U18732 ( .A1(n16817), .A2(n11200), .ZN(n17083) );
  NAND2_X1 U18733 ( .A1(n19124), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n17074) );
  OAI21_X1 U18734 ( .B1(n17877), .B2(n16818), .A(n17074), .ZN(n16819) );
  AOI21_X1 U18735 ( .B1(n17862), .B2(n16820), .A(n16819), .ZN(n16821) );
  OAI21_X1 U18736 ( .B1(n17072), .B2(n17852), .A(n16821), .ZN(n16822) );
  AOI21_X1 U18737 ( .B1(n17083), .B2(n17843), .A(n16822), .ZN(n16823) );
  OAI21_X1 U18738 ( .B1(n17086), .B2(n17853), .A(n16823), .ZN(P2_U2985) );
  INV_X1 U18739 ( .A(n16824), .ZN(n16825) );
  NOR2_X1 U18740 ( .A1(n16826), .A2(n16825), .ZN(n16827) );
  XNOR2_X1 U18741 ( .A(n16827), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17097) );
  AOI21_X1 U18742 ( .B1(n17091), .B2(n16840), .A(n16828), .ZN(n17087) );
  NAND2_X1 U18743 ( .A1(n17087), .A2(n17843), .ZN(n16833) );
  NAND2_X1 U18744 ( .A1(n17862), .A2(n16829), .ZN(n16830) );
  NAND2_X1 U18745 ( .A1(n19124), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n17090) );
  OAI211_X1 U18746 ( .C1(n17877), .C2(n19209), .A(n16830), .B(n17090), .ZN(
        n16831) );
  AOI21_X1 U18747 ( .B1(n19213), .B2(n17870), .A(n16831), .ZN(n16832) );
  OAI211_X1 U18748 ( .C1(n17097), .C2(n17853), .A(n16833), .B(n16832), .ZN(
        P2_U2987) );
  AOI21_X1 U18749 ( .B1(n16851), .B2(n16847), .A(n16848), .ZN(n16836) );
  MUX2_X1 U18750 ( .A(n16847), .B(n16836), .S(n16835), .Z(n16839) );
  INV_X1 U18751 ( .A(n16837), .ZN(n16838) );
  NAND2_X1 U18752 ( .A1(n16839), .A2(n16838), .ZN(n17109) );
  INV_X1 U18753 ( .A(n16840), .ZN(n16842) );
  AOI21_X1 U18754 ( .B1(n11197), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16841) );
  NOR2_X1 U18755 ( .A1(n16842), .A2(n16841), .ZN(n17107) );
  NAND2_X1 U18756 ( .A1(n19199), .A2(n17870), .ZN(n16844) );
  NOR2_X1 U18757 ( .A1(n19294), .A2(n17973), .ZN(n17102) );
  AOI21_X1 U18758 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17102), .ZN(n16843) );
  OAI211_X1 U18759 ( .C1(n17042), .C2(n19202), .A(n16844), .B(n16843), .ZN(
        n16845) );
  AOI21_X1 U18760 ( .B1(n17107), .B2(n17843), .A(n16845), .ZN(n16846) );
  OAI21_X1 U18761 ( .B1(n17853), .B2(n17109), .A(n16846), .ZN(P2_U2988) );
  XNOR2_X1 U18762 ( .A(n11197), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17120) );
  INV_X1 U18763 ( .A(n16847), .ZN(n16849) );
  NOR2_X1 U18764 ( .A1(n16849), .A2(n16848), .ZN(n16850) );
  XNOR2_X1 U18765 ( .A(n16851), .B(n16850), .ZN(n17118) );
  NAND2_X1 U18766 ( .A1(n19124), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n17113) );
  OAI21_X1 U18767 ( .B1(n17877), .B2(n16852), .A(n17113), .ZN(n16853) );
  AOI21_X1 U18768 ( .B1(n17862), .B2(n16854), .A(n16853), .ZN(n16855) );
  OAI21_X1 U18769 ( .B1(n19186), .B2(n17852), .A(n16855), .ZN(n16856) );
  AOI21_X1 U18770 ( .B1(n17118), .B2(n17871), .A(n16856), .ZN(n16857) );
  OAI21_X1 U18771 ( .B1(n17120), .B2(n17873), .A(n16857), .ZN(P2_U2989) );
  XNOR2_X1 U18772 ( .A(n16858), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16859) );
  XNOR2_X1 U18773 ( .A(n16860), .B(n16859), .ZN(n17131) );
  AOI21_X1 U18774 ( .B1(n12345), .B2(n16861), .A(n11197), .ZN(n17121) );
  NAND2_X1 U18775 ( .A1(n17121), .A2(n17843), .ZN(n16866) );
  NOR2_X1 U18776 ( .A1(n19294), .A2(n16862), .ZN(n17122) );
  AOI21_X1 U18777 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n17122), .ZN(n16863) );
  OAI21_X1 U18778 ( .B1(n17042), .B2(n19178), .A(n16863), .ZN(n16864) );
  AOI21_X1 U18779 ( .B1(n19176), .B2(n17870), .A(n16864), .ZN(n16865) );
  OAI211_X1 U18780 ( .C1(n17131), .C2(n17853), .A(n16866), .B(n16865), .ZN(
        P2_U2990) );
  OAI21_X1 U18781 ( .B1(n11215), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16861), .ZN(n17141) );
  INV_X1 U18782 ( .A(n16867), .ZN(n16868) );
  NOR2_X1 U18783 ( .A1(n16869), .A2(n16868), .ZN(n16870) );
  XNOR2_X1 U18784 ( .A(n16871), .B(n16870), .ZN(n17139) );
  NAND2_X1 U18785 ( .A1(n19124), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n17134) );
  OAI21_X1 U18786 ( .B1(n17877), .B2(n16872), .A(n17134), .ZN(n16873) );
  AOI21_X1 U18787 ( .B1(n17862), .B2(n19162), .A(n16873), .ZN(n16874) );
  OAI21_X1 U18788 ( .B1(n19167), .B2(n17852), .A(n16874), .ZN(n16875) );
  AOI21_X1 U18789 ( .B1(n17139), .B2(n17871), .A(n16875), .ZN(n16876) );
  OAI21_X1 U18790 ( .B1(n17141), .B2(n17873), .A(n16876), .ZN(P2_U2991) );
  XNOR2_X1 U18791 ( .A(n16877), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16878) );
  XNOR2_X1 U18792 ( .A(n16879), .B(n16878), .ZN(n17153) );
  AOI21_X1 U18793 ( .B1(n16881), .B2(n16880), .A(n11215), .ZN(n17142) );
  NAND2_X1 U18794 ( .A1(n17142), .A2(n17843), .ZN(n16887) );
  NOR2_X1 U18795 ( .A1(n19294), .A2(n16882), .ZN(n17145) );
  AOI21_X1 U18796 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n17145), .ZN(n16883) );
  OAI21_X1 U18797 ( .B1(n17042), .B2(n16884), .A(n16883), .ZN(n16885) );
  AOI21_X1 U18798 ( .B1(n19152), .B2(n17870), .A(n16885), .ZN(n16886) );
  OAI211_X1 U18799 ( .C1(n17153), .C2(n17853), .A(n16887), .B(n16886), .ZN(
        P2_U2992) );
  OAI21_X1 U18800 ( .B1(n16888), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16880), .ZN(n17166) );
  NAND2_X1 U18801 ( .A1(n16890), .A2(n16889), .ZN(n16900) );
  INV_X1 U18802 ( .A(n17007), .ZN(n16892) );
  AND4_X1 U18803 ( .A1(n16962), .A2(n16956), .A3(n16957), .A4(n16960), .ZN(
        n16893) );
  OAI21_X1 U18804 ( .B1(n16994), .B2(n16894), .A(n16893), .ZN(n16948) );
  NAND2_X1 U18805 ( .A1(n17154), .A2(n17871), .ZN(n16907) );
  OR2_X1 U18806 ( .A1(n19294), .A2(n16901), .ZN(n17159) );
  OAI21_X1 U18807 ( .B1(n17877), .B2(n16902), .A(n17159), .ZN(n16904) );
  NOR2_X1 U18808 ( .A1(n17155), .A2(n17852), .ZN(n16903) );
  AOI211_X1 U18809 ( .C1(n17862), .C2(n16905), .A(n16904), .B(n16903), .ZN(
        n16906) );
  OAI211_X1 U18810 ( .C1(n17873), .C2(n17166), .A(n16907), .B(n16906), .ZN(
        P2_U2993) );
  XNOR2_X1 U18811 ( .A(n16908), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17185) );
  NAND2_X1 U18812 ( .A1(n17178), .A2(n17870), .ZN(n16910) );
  NOR2_X1 U18813 ( .A1(n19294), .A2(n17970), .ZN(n17177) );
  AOI21_X1 U18814 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17177), .ZN(n16909) );
  OAI211_X1 U18815 ( .C1(n17042), .C2(n16911), .A(n16910), .B(n16909), .ZN(
        n16912) );
  XNOR2_X1 U18816 ( .A(n16924), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n17197) );
  INV_X1 U18817 ( .A(n16928), .ZN(n16913) );
  NOR2_X1 U18818 ( .A1(n16914), .A2(n16913), .ZN(n16918) );
  NAND2_X1 U18819 ( .A1(n16916), .A2(n16915), .ZN(n16917) );
  XNOR2_X1 U18820 ( .A(n16918), .B(n16917), .ZN(n17195) );
  NOR2_X1 U18821 ( .A1(n19294), .A2(n17969), .ZN(n17187) );
  NOR2_X1 U18822 ( .A1(n17877), .A2(n16919), .ZN(n16920) );
  AOI211_X1 U18823 ( .C1(n19142), .C2(n17862), .A(n17187), .B(n16920), .ZN(
        n16921) );
  OAI21_X1 U18824 ( .B1(n19137), .B2(n17852), .A(n16921), .ZN(n16922) );
  AOI21_X1 U18825 ( .B1(n17195), .B2(n17871), .A(n16922), .ZN(n16923) );
  OAI21_X1 U18826 ( .B1(n17197), .B2(n17873), .A(n16923), .ZN(P2_U2995) );
  INV_X1 U18827 ( .A(n16924), .ZN(n16926) );
  OAI21_X1 U18828 ( .B1(n17209), .B2(n17222), .A(n17203), .ZN(n16925) );
  NAND2_X1 U18829 ( .A1(n16926), .A2(n16925), .ZN(n17208) );
  NAND2_X1 U18830 ( .A1(n16928), .A2(n16927), .ZN(n16930) );
  XOR2_X1 U18831 ( .A(n16930), .B(n16929), .Z(n17206) );
  NOR2_X1 U18832 ( .A1(n19294), .A2(n17968), .ZN(n17199) );
  NOR2_X1 U18833 ( .A1(n17042), .A2(n16931), .ZN(n16932) );
  AOI211_X1 U18834 ( .C1(n17057), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17199), .B(n16932), .ZN(n16933) );
  OAI21_X1 U18835 ( .B1(n19128), .B2(n17852), .A(n16933), .ZN(n16934) );
  AOI21_X1 U18836 ( .B1(n17206), .B2(n17871), .A(n16934), .ZN(n16935) );
  OAI21_X1 U18837 ( .B1(n17208), .B2(n17873), .A(n16935), .ZN(P2_U2996) );
  XNOR2_X1 U18838 ( .A(n17209), .B(n17222), .ZN(n16945) );
  INV_X1 U18839 ( .A(n16936), .ZN(n16938) );
  NAND2_X1 U18840 ( .A1(n16938), .A2(n16937), .ZN(n16939) );
  XNOR2_X1 U18841 ( .A(n16940), .B(n16939), .ZN(n17220) );
  NOR2_X1 U18842 ( .A1(n19294), .A2(n17967), .ZN(n17214) );
  NOR2_X1 U18843 ( .A1(n17042), .A2(n19123), .ZN(n16941) );
  AOI211_X1 U18844 ( .C1(n17057), .C2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17214), .B(n16941), .ZN(n16942) );
  OAI21_X1 U18845 ( .B1(n19118), .B2(n17852), .A(n16942), .ZN(n16943) );
  AOI21_X1 U18846 ( .B1(n17220), .B2(n17871), .A(n16943), .ZN(n16944) );
  OAI21_X1 U18847 ( .B1(n16945), .B2(n17873), .A(n16944), .ZN(P2_U2997) );
  XNOR2_X1 U18848 ( .A(n17216), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16954) );
  INV_X1 U18849 ( .A(n19106), .ZN(n16952) );
  NAND2_X1 U18850 ( .A1(n19124), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n17224) );
  NAND2_X1 U18851 ( .A1(n17057), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16946) );
  OAI211_X1 U18852 ( .C1(n17042), .C2(n19100), .A(n17224), .B(n16946), .ZN(
        n16951) );
  NOR2_X1 U18853 ( .A1(n16948), .A2(n16947), .ZN(n17226) );
  INV_X1 U18854 ( .A(n16949), .ZN(n17225) );
  NOR3_X1 U18855 ( .A1(n17226), .A2(n17225), .A3(n17853), .ZN(n16950) );
  AOI211_X1 U18856 ( .C1(n17870), .C2(n16952), .A(n16951), .B(n16950), .ZN(
        n16953) );
  OAI21_X1 U18857 ( .B1(n17873), .B2(n16954), .A(n16953), .ZN(P2_U2998) );
  INV_X1 U18858 ( .A(n16996), .ZN(n16955) );
  AOI21_X1 U18859 ( .B1(n16994), .B2(n16956), .A(n16955), .ZN(n16985) );
  NAND2_X1 U18860 ( .A1(n16958), .A2(n16957), .ZN(n16984) );
  NOR2_X1 U18861 ( .A1(n16985), .A2(n16984), .ZN(n16983) );
  INV_X1 U18862 ( .A(n16983), .ZN(n16959) );
  NAND2_X1 U18863 ( .A1(n16959), .A2(n16958), .ZN(n16976) );
  AND2_X1 U18864 ( .A1(n16961), .A2(n16960), .ZN(n16975) );
  NAND2_X1 U18865 ( .A1(n16976), .A2(n16975), .ZN(n16974) );
  NAND2_X1 U18866 ( .A1(n16974), .A2(n16961), .ZN(n16965) );
  NAND2_X1 U18867 ( .A1(n16963), .A2(n16962), .ZN(n16964) );
  XNOR2_X1 U18868 ( .A(n16965), .B(n16964), .ZN(n17245) );
  AOI21_X1 U18869 ( .B1(n17240), .B2(n16973), .A(n17216), .ZN(n17243) );
  NOR2_X1 U18870 ( .A1(n19294), .A2(n17965), .ZN(n17233) );
  NOR2_X1 U18871 ( .A1(n17877), .A2(n16966), .ZN(n16967) );
  AOI211_X1 U18872 ( .C1(n16968), .C2(n17862), .A(n17233), .B(n16967), .ZN(
        n16969) );
  OAI21_X1 U18873 ( .B1(n16970), .B2(n17852), .A(n16969), .ZN(n16971) );
  AOI21_X1 U18874 ( .B1(n17243), .B2(n17843), .A(n16971), .ZN(n16972) );
  OAI21_X1 U18875 ( .B1(n17853), .B2(n17245), .A(n16972), .ZN(P2_U2999) );
  OAI21_X1 U18876 ( .B1(n16987), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16973), .ZN(n17256) );
  OAI21_X1 U18877 ( .B1(n16976), .B2(n16975), .A(n16974), .ZN(n17246) );
  NOR2_X1 U18878 ( .A1(n19294), .A2(n17964), .ZN(n17249) );
  AOI21_X1 U18879 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17249), .ZN(n16979) );
  NAND2_X1 U18880 ( .A1(n17862), .A2(n16977), .ZN(n16978) );
  OAI211_X1 U18881 ( .C1(n16980), .C2(n17852), .A(n16979), .B(n16978), .ZN(
        n16981) );
  AOI21_X1 U18882 ( .B1(n17246), .B2(n17871), .A(n16981), .ZN(n16982) );
  OAI21_X1 U18883 ( .B1(n17873), .B2(n17256), .A(n16982), .ZN(P2_U3000) );
  AOI21_X1 U18884 ( .B1(n16985), .B2(n16984), .A(n16983), .ZN(n17268) );
  NAND2_X1 U18885 ( .A1(n17030), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17017) );
  NOR2_X2 U18886 ( .A1(n17017), .A2(n17283), .ZN(n17012) );
  AOI21_X1 U18887 ( .B1(n17012), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16988) );
  NOR2_X1 U18888 ( .A1(n16988), .A2(n16987), .ZN(n17257) );
  NAND2_X1 U18889 ( .A1(n17257), .A2(n17843), .ZN(n16992) );
  INV_X1 U18890 ( .A(n19093), .ZN(n19087) );
  NOR2_X1 U18891 ( .A1(n19294), .A2(n19084), .ZN(n17260) );
  AOI21_X1 U18892 ( .B1(n17057), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17260), .ZN(n16989) );
  OAI21_X1 U18893 ( .B1(n19090), .B2(n17852), .A(n16989), .ZN(n16990) );
  AOI21_X1 U18894 ( .B1(n17862), .B2(n19087), .A(n16990), .ZN(n16991) );
  OAI211_X1 U18895 ( .C1(n17268), .C2(n17853), .A(n16992), .B(n16991), .ZN(
        P2_U3001) );
  XNOR2_X1 U18896 ( .A(n17012), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17280) );
  NAND2_X1 U18897 ( .A1(n16994), .A2(n16993), .ZN(n16998) );
  NAND2_X1 U18898 ( .A1(n16996), .A2(n16995), .ZN(n16997) );
  XNOR2_X1 U18899 ( .A(n16998), .B(n16997), .ZN(n17278) );
  NOR2_X1 U18900 ( .A1(n19294), .A2(n17963), .ZN(n17271) );
  NOR2_X1 U18901 ( .A1(n17877), .A2(n16999), .ZN(n17000) );
  AOI211_X1 U18902 ( .C1(n17001), .C2(n17870), .A(n17271), .B(n17000), .ZN(
        n17002) );
  OAI21_X1 U18903 ( .B1(n17042), .B2(n17003), .A(n17002), .ZN(n17004) );
  AOI21_X1 U18904 ( .B1(n17278), .B2(n17871), .A(n17004), .ZN(n17005) );
  OAI21_X1 U18905 ( .B1(n17280), .B2(n17873), .A(n17005), .ZN(P2_U3002) );
  NAND2_X1 U18906 ( .A1(n17007), .A2(n17006), .ZN(n17011) );
  NAND2_X1 U18907 ( .A1(n17009), .A2(n17008), .ZN(n17010) );
  XOR2_X1 U18908 ( .A(n17011), .B(n17010), .Z(n17293) );
  AOI21_X1 U18909 ( .B1(n17283), .B2(n17017), .A(n17012), .ZN(n17281) );
  NAND2_X1 U18910 ( .A1(n17281), .A2(n17843), .ZN(n17016) );
  NAND2_X1 U18911 ( .A1(n19124), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n17287) );
  OAI21_X1 U18912 ( .B1(n17877), .B2(n19072), .A(n17287), .ZN(n17014) );
  NOR2_X1 U18913 ( .A1(n17042), .A2(n19083), .ZN(n17013) );
  AOI211_X1 U18914 ( .C1(n17870), .C2(n19069), .A(n17014), .B(n17013), .ZN(
        n17015) );
  OAI211_X1 U18915 ( .C1(n17293), .C2(n17853), .A(n17016), .B(n17015), .ZN(
        P2_U3003) );
  OAI21_X1 U18916 ( .B1(n17030), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17017), .ZN(n17308) );
  NAND2_X1 U18917 ( .A1(n17019), .A2(n17018), .ZN(n17020) );
  XNOR2_X1 U18918 ( .A(n17021), .B(n17020), .ZN(n17306) );
  NOR2_X1 U18919 ( .A1(n19294), .A2(n17962), .ZN(n17300) );
  NOR2_X1 U18920 ( .A1(n17852), .A2(n19064), .ZN(n17022) );
  AOI211_X1 U18921 ( .C1(n17057), .C2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17300), .B(n17022), .ZN(n17023) );
  OAI21_X1 U18922 ( .B1(n17042), .B2(n19058), .A(n17023), .ZN(n17024) );
  AOI21_X1 U18923 ( .B1(n17306), .B2(n17871), .A(n17024), .ZN(n17025) );
  OAI21_X1 U18924 ( .B1(n17308), .B2(n17873), .A(n17025), .ZN(P2_U3004) );
  NAND2_X1 U18925 ( .A1(n17027), .A2(n17026), .ZN(n17029) );
  XOR2_X1 U18926 ( .A(n17029), .B(n17028), .Z(n17320) );
  INV_X1 U18927 ( .A(n17030), .ZN(n17310) );
  NAND2_X1 U18928 ( .A1(n11147), .A2(n17282), .ZN(n17309) );
  NAND3_X1 U18929 ( .A1(n17310), .A2(n17843), .A3(n17309), .ZN(n17036) );
  NAND2_X1 U18930 ( .A1(n19124), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n17313) );
  OAI21_X1 U18931 ( .B1(n17877), .B2(n17031), .A(n17313), .ZN(n17034) );
  NOR2_X1 U18932 ( .A1(n17042), .A2(n17032), .ZN(n17033) );
  AOI211_X1 U18933 ( .C1(n17870), .C2(n17311), .A(n17034), .B(n17033), .ZN(
        n17035) );
  OAI211_X1 U18934 ( .C1(n17320), .C2(n17853), .A(n17036), .B(n17035), .ZN(
        P2_U3005) );
  OR2_X1 U18935 ( .A1(n17038), .A2(n17037), .ZN(n17322) );
  NAND3_X1 U18936 ( .A1(n17322), .A2(n17843), .A3(n17321), .ZN(n17048) );
  XOR2_X1 U18937 ( .A(n17039), .B(n17040), .Z(n17334) );
  INV_X1 U18938 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17043) );
  OAI22_X1 U18939 ( .A1(n17043), .A2(n17877), .B1(n17042), .B2(n17041), .ZN(
        n17046) );
  OAI22_X1 U18940 ( .A1(n17852), .A2(n17331), .B1(n17044), .B2(n19294), .ZN(
        n17045) );
  AOI211_X1 U18941 ( .C1(n17334), .C2(n17871), .A(n17046), .B(n17045), .ZN(
        n17047) );
  NAND2_X1 U18942 ( .A1(n17048), .A2(n17047), .ZN(P2_U3007) );
  AOI22_X1 U18943 ( .A1(n17049), .A2(n17862), .B1(n17870), .B2(n19029), .ZN(
        n17060) );
  AOI21_X1 U18944 ( .B1(n17052), .B2(n17051), .A(n17050), .ZN(n17376) );
  NOR2_X1 U18945 ( .A1(n19294), .A2(n17053), .ZN(n17374) );
  AOI21_X1 U18946 ( .B1(n17843), .B2(n17376), .A(n17374), .ZN(n17059) );
  NOR2_X1 U18947 ( .A1(n17055), .A2(n17054), .ZN(n17056) );
  XOR2_X1 U18948 ( .A(n17056), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17375) );
  AOI22_X1 U18949 ( .A1(n17375), .A2(n17871), .B1(n17057), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17058) );
  NAND3_X1 U18950 ( .A1(n17060), .A2(n17059), .A3(n17058), .ZN(P2_U3013) );
  INV_X1 U18951 ( .A(n17061), .ZN(n17068) );
  NOR3_X1 U18952 ( .A1(n17079), .A2(n17076), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17062) );
  INV_X1 U18953 ( .A(n17069), .ZN(n17070) );
  OAI21_X1 U18954 ( .B1(n17071), .B2(n17351), .A(n17070), .ZN(P2_U3016) );
  INV_X1 U18955 ( .A(n17072), .ZN(n19242) );
  NAND2_X1 U18956 ( .A1(n19240), .A2(n19292), .ZN(n17073) );
  OAI211_X1 U18957 ( .C1(n17092), .C2(n17075), .A(n17074), .B(n17073), .ZN(
        n17082) );
  AOI22_X1 U18958 ( .A1(n17078), .A2(n17077), .B1(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17076), .ZN(n17080) );
  NOR2_X1 U18959 ( .A1(n17080), .A2(n17079), .ZN(n17081) );
  AOI211_X1 U18960 ( .C1(n19242), .C2(n19298), .A(n17082), .B(n17081), .ZN(
        n17085) );
  NAND2_X1 U18961 ( .A1(n17083), .A2(n17377), .ZN(n17084) );
  OAI211_X1 U18962 ( .C1(n17086), .C2(n17351), .A(n17085), .B(n17084), .ZN(
        P2_U3017) );
  NAND2_X1 U18963 ( .A1(n17087), .A2(n17377), .ZN(n17096) );
  NAND2_X1 U18964 ( .A1(n17088), .A2(n17091), .ZN(n17089) );
  OAI211_X1 U18965 ( .C1(n19223), .C2(n17371), .A(n17090), .B(n17089), .ZN(
        n17094) );
  NOR2_X1 U18966 ( .A1(n17092), .A2(n17091), .ZN(n17093) );
  AOI211_X1 U18967 ( .C1(n19213), .C2(n19298), .A(n17094), .B(n17093), .ZN(
        n17095) );
  OAI211_X1 U18968 ( .C1(n17097), .C2(n17351), .A(n17096), .B(n17095), .ZN(
        P2_U3019) );
  AOI211_X1 U18969 ( .C1(n17111), .C2(n17100), .A(n17099), .B(n17098), .ZN(
        n17101) );
  AOI211_X1 U18970 ( .C1(n19198), .C2(n19292), .A(n17102), .B(n17101), .ZN(
        n17104) );
  NAND2_X1 U18971 ( .A1(n17115), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17103) );
  OAI211_X1 U18972 ( .C1(n17105), .C2(n14207), .A(n17104), .B(n17103), .ZN(
        n17106) );
  AOI21_X1 U18973 ( .B1(n17107), .B2(n17377), .A(n17106), .ZN(n17108) );
  OAI21_X1 U18974 ( .B1(n17351), .B2(n17109), .A(n17108), .ZN(P2_U3020) );
  NAND2_X1 U18975 ( .A1(n17111), .A2(n17110), .ZN(n17112) );
  OAI211_X1 U18976 ( .C1(n19187), .C2(n17371), .A(n17113), .B(n17112), .ZN(
        n17114) );
  AOI21_X1 U18977 ( .B1(n17115), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17114), .ZN(n17116) );
  OAI21_X1 U18978 ( .B1(n19186), .B2(n14207), .A(n17116), .ZN(n17117) );
  AOI21_X1 U18979 ( .B1(n17118), .B2(n19299), .A(n17117), .ZN(n17119) );
  OAI21_X1 U18980 ( .B1(n17120), .B2(n19302), .A(n17119), .ZN(P2_U3021) );
  NAND2_X1 U18981 ( .A1(n17121), .A2(n17377), .ZN(n17130) );
  INV_X1 U18982 ( .A(n17122), .ZN(n17123) );
  OAI21_X1 U18983 ( .B1(n19174), .B2(n17371), .A(n17123), .ZN(n17128) );
  INV_X1 U18984 ( .A(n17124), .ZN(n17126) );
  AOI21_X1 U18985 ( .B1(n17126), .B2(n12345), .A(n17125), .ZN(n17127) );
  AOI211_X1 U18986 ( .C1(n19298), .C2(n19176), .A(n17128), .B(n17127), .ZN(
        n17129) );
  OAI211_X1 U18987 ( .C1(n17131), .C2(n17351), .A(n17130), .B(n17129), .ZN(
        P2_U3022) );
  INV_X1 U18988 ( .A(n17148), .ZN(n17133) );
  OAI211_X1 U18989 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n17133), .B(n17132), .ZN(
        n17135) );
  OAI211_X1 U18990 ( .C1(n19165), .C2(n17371), .A(n17135), .B(n17134), .ZN(
        n17136) );
  AOI21_X1 U18991 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17150), .A(
        n17136), .ZN(n17137) );
  OAI21_X1 U18992 ( .B1(n19167), .B2(n14207), .A(n17137), .ZN(n17138) );
  AOI21_X1 U18993 ( .B1(n17139), .B2(n19299), .A(n17138), .ZN(n17140) );
  OAI21_X1 U18994 ( .B1(n17141), .B2(n19302), .A(n17140), .ZN(P2_U3023) );
  NAND2_X1 U18995 ( .A1(n17142), .A2(n17377), .ZN(n17152) );
  NAND2_X1 U18996 ( .A1(n19152), .A2(n19298), .ZN(n17147) );
  AND2_X1 U18997 ( .A1(n11161), .A2(n17143), .ZN(n17144) );
  NOR2_X1 U18998 ( .A1(n16778), .A2(n17144), .ZN(n20019) );
  AOI21_X1 U18999 ( .B1(n20019), .B2(n19292), .A(n17145), .ZN(n17146) );
  OAI211_X1 U19000 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17148), .A(
        n17147), .B(n17146), .ZN(n17149) );
  AOI21_X1 U19001 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17150), .A(
        n17149), .ZN(n17151) );
  OAI211_X1 U19002 ( .C1(n17153), .C2(n17351), .A(n17152), .B(n17151), .ZN(
        P2_U3024) );
  INV_X1 U19003 ( .A(n17155), .ZN(n17164) );
  NOR3_X1 U19004 ( .A1(n17156), .A2(n17295), .A3(n17158), .ZN(n17163) );
  NAND3_X1 U19005 ( .A1(n17238), .A2(n11605), .A3(n17158), .ZN(n17160) );
  OAI211_X1 U19006 ( .C1(n17371), .C2(n17161), .A(n17160), .B(n17159), .ZN(
        n17162) );
  AOI211_X1 U19007 ( .C1(n17164), .C2(n19298), .A(n17163), .B(n17162), .ZN(
        n17165) );
  NAND2_X1 U19008 ( .A1(n17238), .A2(n17171), .ZN(n17190) );
  OR2_X1 U19009 ( .A1(n17190), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17201) );
  NOR2_X1 U19010 ( .A1(n17352), .A2(n17167), .ZN(n17168) );
  NOR2_X1 U19011 ( .A1(n17169), .A2(n17168), .ZN(n17175) );
  NOR2_X1 U19012 ( .A1(n17170), .A2(n17210), .ZN(n17172) );
  OAI21_X1 U19013 ( .B1(n17326), .B2(n17172), .A(n17171), .ZN(n17173) );
  NAND2_X1 U19014 ( .A1(n17173), .A2(n19279), .ZN(n17174) );
  AND2_X1 U19015 ( .A1(n17175), .A2(n17174), .ZN(n17204) );
  AND2_X1 U19016 ( .A1(n17201), .A2(n17204), .ZN(n17186) );
  NOR2_X1 U19017 ( .A1(n20116), .A2(n17371), .ZN(n17176) );
  AOI211_X1 U19018 ( .C1(n17178), .C2(n19298), .A(n17177), .B(n17176), .ZN(
        n17182) );
  INV_X1 U19019 ( .A(n17190), .ZN(n17180) );
  OAI21_X1 U19020 ( .B1(n17203), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17179) );
  OAI211_X1 U19021 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n17180), .B(n17179), .ZN(
        n17181) );
  OAI211_X1 U19022 ( .C1(n17186), .C2(n17183), .A(n17182), .B(n17181), .ZN(
        n17184) );
  NOR2_X1 U19023 ( .A1(n17186), .A2(n17188), .ZN(n17194) );
  AOI21_X1 U19024 ( .B1(n19138), .B2(n19292), .A(n17187), .ZN(n17192) );
  NAND2_X1 U19025 ( .A1(n17188), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17189) );
  OR2_X1 U19026 ( .A1(n17190), .A2(n17189), .ZN(n17191) );
  OAI211_X1 U19027 ( .C1(n19137), .C2(n14207), .A(n17192), .B(n17191), .ZN(
        n17193) );
  AOI211_X1 U19028 ( .C1(n17195), .C2(n19299), .A(n17194), .B(n17193), .ZN(
        n17196) );
  OAI21_X1 U19029 ( .B1(n17197), .B2(n19302), .A(n17196), .ZN(P2_U3027) );
  INV_X1 U19030 ( .A(n19136), .ZN(n17200) );
  NOR2_X1 U19031 ( .A1(n19128), .A2(n14207), .ZN(n17198) );
  AOI211_X1 U19032 ( .C1(n19292), .C2(n17200), .A(n17199), .B(n17198), .ZN(
        n17202) );
  OAI211_X1 U19033 ( .C1(n17204), .C2(n17203), .A(n17202), .B(n17201), .ZN(
        n17205) );
  AOI21_X1 U19034 ( .B1(n17206), .B2(n19299), .A(n17205), .ZN(n17207) );
  OAI21_X1 U19035 ( .B1(n17208), .B2(n19302), .A(n17207), .ZN(P2_U3028) );
  OAI21_X1 U19036 ( .B1(n17377), .B2(n17328), .A(n17209), .ZN(n17213) );
  NAND2_X1 U19037 ( .A1(n19279), .A2(n17210), .ZN(n17211) );
  OAI21_X1 U19038 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17326), .A(
        n17211), .ZN(n17212) );
  NOR2_X1 U19039 ( .A1(n17317), .A2(n17212), .ZN(n17241) );
  NAND2_X1 U19040 ( .A1(n17213), .A2(n17241), .ZN(n17229) );
  AOI21_X1 U19041 ( .B1(n17217), .B2(n19279), .A(n17229), .ZN(n17223) );
  AOI21_X1 U19042 ( .B1(n19292), .B2(n19116), .A(n17214), .ZN(n17215) );
  OAI21_X1 U19043 ( .B1(n19118), .B2(n14207), .A(n17215), .ZN(n17219) );
  AOI22_X1 U19044 ( .A1(n17216), .A2(n17377), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17238), .ZN(n17232) );
  NOR3_X1 U19045 ( .A1(n17232), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n17217), .ZN(n17218) );
  AOI211_X1 U19046 ( .C1(n19299), .C2(n17220), .A(n17219), .B(n17218), .ZN(
        n17221) );
  OAI21_X1 U19047 ( .B1(n17223), .B2(n17222), .A(n17221), .ZN(P2_U3029) );
  OAI21_X1 U19048 ( .B1(n19106), .B2(n14207), .A(n17224), .ZN(n17228) );
  NOR3_X1 U19049 ( .A1(n17226), .A2(n17225), .A3(n17351), .ZN(n17227) );
  AOI211_X1 U19050 ( .C1(n19292), .C2(n19104), .A(n17228), .B(n17227), .ZN(
        n17231) );
  NAND2_X1 U19051 ( .A1(n17229), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n17230) );
  OAI211_X1 U19052 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17232), .A(
        n17231), .B(n17230), .ZN(P2_U3030) );
  AOI21_X1 U19053 ( .B1(n17234), .B2(n19298), .A(n17233), .ZN(n17235) );
  OAI21_X1 U19054 ( .B1(n17371), .B2(n17236), .A(n17235), .ZN(n17237) );
  AOI21_X1 U19055 ( .B1(n17238), .B2(n17240), .A(n17237), .ZN(n17239) );
  OAI21_X1 U19056 ( .B1(n17241), .B2(n17240), .A(n17239), .ZN(n17242) );
  AOI21_X1 U19057 ( .B1(n17243), .B2(n17377), .A(n17242), .ZN(n17244) );
  OAI21_X1 U19058 ( .B1(n17351), .B2(n17245), .A(n17244), .ZN(P2_U3031) );
  NAND2_X1 U19059 ( .A1(n17246), .A2(n19299), .ZN(n17255) );
  NOR2_X1 U19060 ( .A1(n17317), .A2(n17247), .ZN(n17270) );
  INV_X1 U19061 ( .A(n17285), .ZN(n17314) );
  NOR2_X1 U19062 ( .A1(n17314), .A2(n17247), .ZN(n17259) );
  NAND2_X1 U19063 ( .A1(n17259), .A2(n17269), .ZN(n17274) );
  OAI21_X1 U19064 ( .B1(n17295), .B2(n17270), .A(n17274), .ZN(n17265) );
  OAI21_X1 U19065 ( .B1(n17269), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17248) );
  OAI211_X1 U19066 ( .C1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n17259), .B(n17248), .ZN(
        n17252) );
  AOI21_X1 U19067 ( .B1(n17250), .B2(n19298), .A(n17249), .ZN(n17251) );
  OAI211_X1 U19068 ( .C1(n17371), .C2(n19808), .A(n17252), .B(n17251), .ZN(
        n17253) );
  AOI21_X1 U19069 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17265), .A(
        n17253), .ZN(n17254) );
  OAI211_X1 U19070 ( .C1(n17256), .C2(n19302), .A(n17255), .B(n17254), .ZN(
        P2_U3032) );
  NAND2_X1 U19071 ( .A1(n17257), .A2(n17377), .ZN(n17267) );
  NAND3_X1 U19072 ( .A1(n17259), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        n17258), .ZN(n17263) );
  AOI21_X1 U19073 ( .B1(n17261), .B2(n19298), .A(n17260), .ZN(n17262) );
  OAI211_X1 U19074 ( .C1(n17371), .C2(n19089), .A(n17263), .B(n17262), .ZN(
        n17264) );
  AOI21_X1 U19075 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17265), .A(
        n17264), .ZN(n17266) );
  OAI211_X1 U19076 ( .C1(n17268), .C2(n17351), .A(n17267), .B(n17266), .ZN(
        P2_U3033) );
  NOR3_X1 U19077 ( .A1(n17270), .A2(n17295), .A3(n17269), .ZN(n17277) );
  INV_X1 U19078 ( .A(n19811), .ZN(n17272) );
  AOI21_X1 U19079 ( .B1(n19292), .B2(n17272), .A(n17271), .ZN(n17273) );
  OAI211_X1 U19080 ( .C1(n17275), .C2(n14207), .A(n17274), .B(n17273), .ZN(
        n17276) );
  AOI211_X1 U19081 ( .C1(n17278), .C2(n19299), .A(n17277), .B(n17276), .ZN(
        n17279) );
  OAI21_X1 U19082 ( .B1(n17280), .B2(n19302), .A(n17279), .ZN(P2_U3034) );
  NAND2_X1 U19083 ( .A1(n17281), .A2(n17377), .ZN(n17292) );
  NOR2_X1 U19084 ( .A1(n17317), .A2(n17282), .ZN(n17296) );
  NAND3_X1 U19085 ( .A1(n17285), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n17294), .ZN(n17303) );
  OAI21_X1 U19086 ( .B1(n17296), .B2(n17295), .A(n17303), .ZN(n17290) );
  AND3_X1 U19087 ( .A1(n17285), .A2(n17284), .A3(n17283), .ZN(n17289) );
  NAND2_X1 U19088 ( .A1(n19298), .A2(n19069), .ZN(n17286) );
  OAI211_X1 U19089 ( .C1(n17371), .C2(n19070), .A(n17287), .B(n17286), .ZN(
        n17288) );
  AOI211_X1 U19090 ( .C1(n17290), .C2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17289), .B(n17288), .ZN(n17291) );
  OAI211_X1 U19091 ( .C1(n17293), .C2(n17351), .A(n17292), .B(n17291), .ZN(
        P2_U3035) );
  NOR3_X1 U19092 ( .A1(n17296), .A2(n17295), .A3(n17294), .ZN(n17305) );
  NAND2_X1 U19093 ( .A1(n15456), .A2(n17297), .ZN(n17298) );
  NAND2_X1 U19094 ( .A1(n17299), .A2(n17298), .ZN(n19814) );
  INV_X1 U19095 ( .A(n19064), .ZN(n17301) );
  AOI21_X1 U19096 ( .B1(n19298), .B2(n17301), .A(n17300), .ZN(n17302) );
  OAI211_X1 U19097 ( .C1(n17371), .C2(n19814), .A(n17303), .B(n17302), .ZN(
        n17304) );
  AOI211_X1 U19098 ( .C1(n17306), .C2(n19299), .A(n17305), .B(n17304), .ZN(
        n17307) );
  OAI21_X1 U19099 ( .B1(n17308), .B2(n19302), .A(n17307), .ZN(P2_U3036) );
  NAND3_X1 U19100 ( .A1(n17310), .A2(n17377), .A3(n17309), .ZN(n17319) );
  NAND2_X1 U19101 ( .A1(n19298), .A2(n17311), .ZN(n17312) );
  OAI211_X1 U19102 ( .C1(n17371), .C2(n19817), .A(n17313), .B(n17312), .ZN(
        n17316) );
  NOR2_X1 U19103 ( .A1(n17314), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17315) );
  AOI211_X1 U19104 ( .C1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n17317), .A(
        n17316), .B(n17315), .ZN(n17318) );
  OAI211_X1 U19105 ( .C1(n17320), .C2(n17351), .A(n17319), .B(n17318), .ZN(
        P2_U3037) );
  NAND3_X1 U19106 ( .A1(n17322), .A2(n17377), .A3(n17321), .ZN(n17336) );
  NAND2_X1 U19107 ( .A1(n17323), .A2(n17344), .ZN(n19288) );
  NAND2_X1 U19108 ( .A1(n17328), .A2(n17341), .ZN(n17325) );
  OAI211_X1 U19109 ( .C1(n17327), .C2(n17326), .A(n17325), .B(n17324), .ZN(
        n17348) );
  AOI21_X1 U19110 ( .B1(n17328), .B2(n17342), .A(n17348), .ZN(n19308) );
  NAND2_X1 U19111 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19124), .ZN(n17329) );
  OAI221_X1 U19112 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n19288), .C1(
        n19290), .C2(n19308), .A(n17329), .ZN(n17333) );
  OAI22_X1 U19113 ( .A1(n14207), .A2(n17331), .B1(n17371), .B2(n17330), .ZN(
        n17332) );
  AOI211_X1 U19114 ( .C1(n17334), .C2(n19299), .A(n17333), .B(n17332), .ZN(
        n17335) );
  NAND2_X1 U19115 ( .A1(n17336), .A2(n17335), .ZN(P2_U3039) );
  XNOR2_X1 U19116 ( .A(n17338), .B(n17337), .ZN(n17854) );
  NOR2_X1 U19117 ( .A1(n17339), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17850) );
  INV_X1 U19118 ( .A(n17850), .ZN(n17340) );
  NAND3_X1 U19119 ( .A1(n17340), .A2(n17377), .A3(n17856), .ZN(n17350) );
  INV_X1 U19120 ( .A(n17341), .ZN(n17343) );
  NAND3_X1 U19121 ( .A1(n17344), .A2(n17343), .A3(n17342), .ZN(n17346) );
  AOI22_X1 U19122 ( .A1(n19298), .A2(n19052), .B1(n19124), .B2(
        P2_REIP_REG_6__SCAN_IN), .ZN(n17345) );
  OAI211_X1 U19123 ( .C1(n17371), .C2(n19056), .A(n17346), .B(n17345), .ZN(
        n17347) );
  AOI21_X1 U19124 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17348), .A(
        n17347), .ZN(n17349) );
  OAI211_X1 U19125 ( .C1(n17854), .C2(n17351), .A(n17350), .B(n17349), .ZN(
        P2_U3040) );
  AOI21_X1 U19126 ( .B1(n17354), .B2(n17353), .A(n17352), .ZN(n17355) );
  INV_X1 U19127 ( .A(n17355), .ZN(n17370) );
  AOI22_X1 U19128 ( .A1(n19299), .A2(n17357), .B1(n17377), .B2(n17356), .ZN(
        n17369) );
  NAND3_X1 U19129 ( .A1(n17361), .A2(n17358), .A3(n17362), .ZN(n17359) );
  OAI21_X1 U19130 ( .B1(n14207), .B2(n12110), .A(n17359), .ZN(n17367) );
  AND2_X1 U19131 ( .A1(n19292), .A2(n17360), .ZN(n17366) );
  NAND2_X1 U19132 ( .A1(n17361), .A2(n17379), .ZN(n17363) );
  AOI21_X1 U19133 ( .B1(n19275), .B2(n17363), .A(n17362), .ZN(n17365) );
  NOR4_X1 U19134 ( .A1(n17367), .A2(n17366), .A3(n17365), .A4(n17364), .ZN(
        n17368) );
  NAND3_X1 U19135 ( .A1(n17370), .A2(n17369), .A3(n17368), .ZN(P2_U3044) );
  OAI22_X1 U19136 ( .A1(n17372), .A2(n14207), .B1(n17371), .B2(n19026), .ZN(
        n17373) );
  AOI211_X1 U19137 ( .C1(n19299), .C2(n17375), .A(n17374), .B(n17373), .ZN(
        n17382) );
  AOI22_X1 U19138 ( .A1(n17378), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n17377), .B2(n17376), .ZN(n17381) );
  OAI211_X1 U19139 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n19279), .B(n17379), .ZN(n17380) );
  NAND3_X1 U19140 ( .A1(n17382), .A2(n17381), .A3(n17380), .ZN(P2_U3045) );
  INV_X1 U19141 ( .A(n17383), .ZN(n17386) );
  OAI222_X1 U19142 ( .A1(n17389), .A2(n19940), .B1(n17386), .B2(n17385), .C1(
        n19311), .C2(n17384), .ZN(n17387) );
  MUX2_X1 U19143 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17387), .S(
        n19274), .Z(P2_U3599) );
  OAI22_X1 U19144 ( .A1(n19941), .A2(n17389), .B1(n17388), .B2(n19311), .ZN(
        n17390) );
  MUX2_X1 U19145 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17390), .S(
        n19274), .Z(P2_U3596) );
  NAND2_X1 U19146 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19363) );
  INV_X1 U19147 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n22314) );
  NOR2_X1 U19148 ( .A1(n21389), .A2(n22314), .ZN(n18568) );
  INV_X1 U19149 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21923) );
  NAND2_X1 U19150 ( .A1(n21923), .A2(n18359), .ZN(n20707) );
  NOR2_X1 U19151 ( .A1(n18568), .A2(n20707), .ZN(n17394) );
  NAND2_X1 U19152 ( .A1(n21892), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19364) );
  NOR2_X1 U19153 ( .A1(n18390), .A2(n17391), .ZN(n18361) );
  INV_X1 U19154 ( .A(n17405), .ZN(n21922) );
  INV_X1 U19155 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21915) );
  NAND2_X1 U19156 ( .A1(n21389), .A2(n21915), .ZN(n21927) );
  NAND2_X1 U19157 ( .A1(n17392), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n21926) );
  OAI211_X1 U19158 ( .C1(n18361), .C2(n21922), .A(n19571), .B(n17393), .ZN(
        n18358) );
  NAND2_X1 U19159 ( .A1(n19364), .A2(n18358), .ZN(n18921) );
  AOI221_X1 U19160 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19363), .C1(n17394), 
        .C2(n19363), .A(n18921), .ZN(n18920) );
  NOR2_X1 U19161 ( .A1(n21923), .A2(n21892), .ZN(n17395) );
  OAI21_X1 U19162 ( .B1(n17395), .B2(n17394), .A(n18358), .ZN(n18923) );
  INV_X1 U19163 ( .A(n18923), .ZN(n18918) );
  NAND3_X1 U19164 ( .A1(n21915), .A2(n21923), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n19389) );
  NAND2_X1 U19165 ( .A1(n21895), .A2(n19389), .ZN(n19421) );
  OAI21_X1 U19166 ( .B1(n18918), .B2(n18917), .A(n19421), .ZN(n17396) );
  AOI22_X1 U19167 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18920), .B1(
        n17396), .B2(n21900), .ZN(P3_U2865) );
  INV_X1 U19168 ( .A(n22286), .ZN(n22284) );
  NOR2_X1 U19169 ( .A1(n17398), .A2(n17397), .ZN(n17399) );
  XNOR2_X1 U19170 ( .A(n17399), .B(n13350), .ZN(n22132) );
  NAND4_X1 U19171 ( .A1(n22132), .A2(n17401), .A3(n17454), .A4(n17400), .ZN(
        n17402) );
  OAI21_X1 U19172 ( .B1(n22284), .B2(n13350), .A(n17402), .ZN(P1_U3468) );
  INV_X1 U19173 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17403) );
  AOI221_X1 U19174 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(n22369), .C1(
        P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n22323), 
        .ZN(n22317) );
  INV_X1 U19175 ( .A(BS16), .ZN(n17533) );
  INV_X1 U19176 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n22377) );
  NAND2_X1 U19177 ( .A1(n22377), .A2(n22369), .ZN(n22319) );
  AOI21_X1 U19178 ( .B1(n17533), .B2(n22319), .A(n17404), .ZN(n22313) );
  AOI21_X1 U19179 ( .B1(n17403), .B2(n17404), .A(n22313), .ZN(P3_U3280) );
  AND2_X1 U19180 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n17404), .ZN(P3_U3028) );
  AND2_X1 U19181 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n17404), .ZN(P3_U3027) );
  AND2_X1 U19182 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n17404), .ZN(P3_U3026) );
  AND2_X1 U19183 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n17404), .ZN(P3_U3025) );
  AND2_X1 U19184 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n17404), .ZN(P3_U3024) );
  AND2_X1 U19185 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n17404), .ZN(P3_U3023) );
  AND2_X1 U19186 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n17404), .ZN(P3_U3022) );
  AND2_X1 U19187 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n17404), .ZN(P3_U3021) );
  AND2_X1 U19188 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n17404), .ZN(
        P3_U3020) );
  AND2_X1 U19189 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n17404), .ZN(
        P3_U3019) );
  AND2_X1 U19190 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n17404), .ZN(
        P3_U3018) );
  AND2_X1 U19191 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n17404), .ZN(
        P3_U3017) );
  AND2_X1 U19192 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n17404), .ZN(
        P3_U3016) );
  AND2_X1 U19193 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n17404), .ZN(
        P3_U3015) );
  AND2_X1 U19194 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n17404), .ZN(
        P3_U3014) );
  AND2_X1 U19195 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n17404), .ZN(
        P3_U3013) );
  AND2_X1 U19196 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n17404), .ZN(
        P3_U3012) );
  AND2_X1 U19197 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n17404), .ZN(
        P3_U3011) );
  AND2_X1 U19198 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n17404), .ZN(
        P3_U3010) );
  AND2_X1 U19199 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n17404), .ZN(
        P3_U3009) );
  AND2_X1 U19200 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n17404), .ZN(
        P3_U3008) );
  AND2_X1 U19201 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n17404), .ZN(
        P3_U3007) );
  AND2_X1 U19202 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n17404), .ZN(
        P3_U3006) );
  AND2_X1 U19203 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n17404), .ZN(
        P3_U3005) );
  AND2_X1 U19204 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n17404), .ZN(
        P3_U3004) );
  AND2_X1 U19205 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n17404), .ZN(
        P3_U3003) );
  AND2_X1 U19206 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n17404), .ZN(
        P3_U3002) );
  AND2_X1 U19207 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n17404), .ZN(
        P3_U3001) );
  AND2_X1 U19208 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n17404), .ZN(
        P3_U3000) );
  AND2_X1 U19209 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n17404), .ZN(
        P3_U2999) );
  INV_X1 U19210 ( .A(n18568), .ZN(n18873) );
  AOI21_X1 U19211 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n17406)
         );
  NOR4_X1 U19212 ( .A1(n21389), .A2(n21936), .A3(n22370), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21872) );
  AOI211_X1 U19213 ( .C1(n18873), .C2(n17406), .A(n17405), .B(n21872), .ZN(
        P3_U2998) );
  NOR2_X1 U19214 ( .A1(n21904), .A2(n18358), .ZN(P3_U2867) );
  NAND2_X1 U19215 ( .A1(n21936), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18910) );
  AND2_X1 U19216 ( .A1(n18979), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NOR2_X1 U19217 ( .A1(n21927), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18522) );
  NOR2_X1 U19218 ( .A1(n18522), .A2(n20767), .ZN(n17410) );
  INV_X1 U19219 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18948) );
  NAND2_X1 U19220 ( .A1(n17409), .A2(n17408), .ZN(n20704) );
  AOI22_X1 U19221 ( .A1(n17410), .A2(n18948), .B1(n20767), .B2(n20704), .ZN(
        P3_U3298) );
  INV_X1 U19222 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18947) );
  NAND2_X1 U19223 ( .A1(n19708), .A2(n20767), .ZN(n21190) );
  INV_X1 U19224 ( .A(n21190), .ZN(n20803) );
  AOI21_X1 U19225 ( .B1(n17410), .B2(n18947), .A(n20803), .ZN(P3_U3299) );
  NOR2_X1 U19226 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n22348), .ZN(n22358) );
  INV_X1 U19227 ( .A(n22350), .ZN(n17411) );
  AOI21_X1 U19228 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22358), .A(n17411), 
        .ZN(n17412) );
  INV_X1 U19229 ( .A(n17412), .ZN(n22312) );
  INV_X1 U19230 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n17429) );
  NAND2_X1 U19231 ( .A1(n22354), .A2(n22348), .ZN(n22346) );
  AOI21_X1 U19232 ( .B1(n17533), .B2(n22346), .A(n17413), .ZN(n22309) );
  AOI21_X1 U19233 ( .B1(n17413), .B2(n17429), .A(n22309), .ZN(P2_U3591) );
  AND2_X1 U19234 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n17413), .ZN(P2_U3208) );
  AND2_X1 U19235 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n17413), .ZN(P2_U3207) );
  AND2_X1 U19236 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n17413), .ZN(P2_U3206) );
  AND2_X1 U19237 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n17413), .ZN(P2_U3205) );
  AND2_X1 U19238 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n17413), .ZN(P2_U3204) );
  AND2_X1 U19239 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n17413), .ZN(P2_U3203) );
  AND2_X1 U19240 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n17413), .ZN(P2_U3202) );
  AND2_X1 U19241 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n17413), .ZN(P2_U3201) );
  AND2_X1 U19242 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n17413), .ZN(
        P2_U3200) );
  AND2_X1 U19243 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n17413), .ZN(
        P2_U3199) );
  AND2_X1 U19244 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n17413), .ZN(
        P2_U3198) );
  AND2_X1 U19245 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n17413), .ZN(
        P2_U3197) );
  AND2_X1 U19246 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n17413), .ZN(
        P2_U3196) );
  AND2_X1 U19247 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n17413), .ZN(
        P2_U3195) );
  AND2_X1 U19248 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n17412), .ZN(
        P2_U3194) );
  AND2_X1 U19249 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n17412), .ZN(
        P2_U3193) );
  AND2_X1 U19250 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n17412), .ZN(
        P2_U3192) );
  AND2_X1 U19251 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n17412), .ZN(
        P2_U3191) );
  AND2_X1 U19252 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n17412), .ZN(
        P2_U3190) );
  AND2_X1 U19253 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n17412), .ZN(
        P2_U3189) );
  AND2_X1 U19254 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n17412), .ZN(
        P2_U3188) );
  AND2_X1 U19255 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n17412), .ZN(
        P2_U3187) );
  AND2_X1 U19256 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n17412), .ZN(
        P2_U3186) );
  AND2_X1 U19257 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n17412), .ZN(
        P2_U3185) );
  AND2_X1 U19258 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n17412), .ZN(
        P2_U3184) );
  AND2_X1 U19259 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n17412), .ZN(
        P2_U3183) );
  AND2_X1 U19260 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n17413), .ZN(
        P2_U3182) );
  AND2_X1 U19261 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n17413), .ZN(
        P2_U3181) );
  AND2_X1 U19262 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n17413), .ZN(
        P2_U3180) );
  AND2_X1 U19263 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n17413), .ZN(
        P2_U3179) );
  NAND2_X1 U19264 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n22349), .ZN(n19310) );
  AOI21_X1 U19265 ( .B1(n17414), .B2(n19322), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n17417) );
  AOI221_X1 U19266 ( .B1(n19310), .B2(n17417), .C1(n17416), .C2(n17417), .A(
        n17415), .ZN(P2_U3178) );
  OAI221_X1 U19267 ( .B1(n12377), .B2(n19330), .C1(n19318), .C2(n19330), .A(
        n20291), .ZN(n17901) );
  NOR2_X1 U19268 ( .A1(n17418), .A2(n17901), .ZN(P2_U3047) );
  AND2_X1 U19269 ( .A1(n17935), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U19270 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n17422) );
  NOR4_X1 U19271 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n17421) );
  NOR4_X1 U19272 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n17420) );
  NOR4_X1 U19273 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n17419) );
  NAND4_X1 U19274 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17428) );
  NOR4_X1 U19275 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n17426) );
  AOI211_X1 U19276 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17425) );
  NOR4_X1 U19277 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17424) );
  NOR4_X1 U19278 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17423) );
  NAND4_X1 U19279 ( .A1(n17426), .A2(n17425), .A3(n17424), .A4(n17423), .ZN(
        n17427) );
  NOR2_X1 U19280 ( .A1(n17428), .A2(n17427), .ZN(n17911) );
  INV_X1 U19281 ( .A(n17911), .ZN(n17909) );
  NOR2_X1 U19282 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17909), .ZN(n17904) );
  INV_X1 U19283 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22311) );
  NAND3_X1 U19284 ( .A1(n14423), .A2(n22311), .A3(n17429), .ZN(n17908) );
  INV_X1 U19285 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U19286 ( .A1(n17904), .A2(n17908), .B1(n17909), .B2(n17430), .ZN(
        P2_U2821) );
  INV_X1 U19287 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U19288 ( .A1(n17904), .A2(n14423), .B1(n17909), .B2(n17431), .ZN(
        P2_U2820) );
  INV_X1 U19289 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20536) );
  INV_X1 U19290 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n22334) );
  NOR2_X1 U19291 ( .A1(n22334), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n22324) );
  INV_X2 U19292 ( .A(n22853), .ZN(n22850) );
  OAI21_X1 U19293 ( .B1(n22324), .B2(n22343), .A(n22850), .ZN(n17433) );
  INV_X1 U19294 ( .A(n17433), .ZN(n22308) );
  AOI221_X1 U19295 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n17533), .C1(
        P1_STATE_REG_2__SCAN_IN), .C2(n17533), .A(n17432), .ZN(n22305) );
  AOI21_X1 U19296 ( .B1(n20536), .B2(n17432), .A(n22305), .ZN(P1_U3464) );
  AND2_X1 U19297 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n17432), .ZN(P1_U3193) );
  AND2_X1 U19298 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n17432), .ZN(P1_U3192) );
  AND2_X1 U19299 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n17432), .ZN(P1_U3191) );
  AND2_X1 U19300 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n17432), .ZN(P1_U3190) );
  AND2_X1 U19301 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n17432), .ZN(P1_U3189) );
  AND2_X1 U19302 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n17432), .ZN(P1_U3188) );
  AND2_X1 U19303 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n17432), .ZN(P1_U3187) );
  AND2_X1 U19304 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n17432), .ZN(P1_U3186) );
  AND2_X1 U19305 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n17432), .ZN(
        P1_U3185) );
  AND2_X1 U19306 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n17432), .ZN(
        P1_U3184) );
  AND2_X1 U19307 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n17432), .ZN(
        P1_U3183) );
  AND2_X1 U19308 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n17432), .ZN(
        P1_U3182) );
  AND2_X1 U19309 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n17432), .ZN(
        P1_U3181) );
  AND2_X1 U19310 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n17433), .ZN(
        P1_U3180) );
  AND2_X1 U19311 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n17433), .ZN(
        P1_U3179) );
  AND2_X1 U19312 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n17433), .ZN(
        P1_U3178) );
  AND2_X1 U19313 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n17433), .ZN(
        P1_U3177) );
  AND2_X1 U19314 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n17433), .ZN(
        P1_U3176) );
  AND2_X1 U19315 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n17433), .ZN(
        P1_U3175) );
  AND2_X1 U19316 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n17433), .ZN(
        P1_U3174) );
  AND2_X1 U19317 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n17433), .ZN(
        P1_U3173) );
  AND2_X1 U19318 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n17433), .ZN(
        P1_U3172) );
  AND2_X1 U19319 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n17433), .ZN(
        P1_U3171) );
  AND2_X1 U19320 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n17433), .ZN(
        P1_U3170) );
  AND2_X1 U19321 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n17433), .ZN(
        P1_U3169) );
  AND2_X1 U19322 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n17433), .ZN(
        P1_U3168) );
  AND2_X1 U19323 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n17432), .ZN(
        P1_U3167) );
  AND2_X1 U19324 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n17432), .ZN(
        P1_U3166) );
  AND2_X1 U19325 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n17432), .ZN(
        P1_U3165) );
  AND2_X1 U19326 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n17433), .ZN(
        P1_U3164) );
  MUX2_X1 U19327 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n17434), .S(
        n17457), .Z(n17461) );
  MUX2_X1 U19328 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n17435), .S(
        n17457), .Z(n17460) );
  INV_X1 U19329 ( .A(n17460), .ZN(n17448) );
  AOI22_X1 U19330 ( .A1(n17438), .A2(n17437), .B1(n17436), .B2(n13179), .ZN(
        n22283) );
  NAND2_X1 U19331 ( .A1(n17439), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n22288) );
  NAND3_X1 U19332 ( .A1(n22283), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(
        n22288), .ZN(n17442) );
  INV_X1 U19333 ( .A(n17440), .ZN(n17441) );
  OAI211_X1 U19334 ( .C1(n22584), .C2(n17442), .A(n17441), .B(n17457), .ZN(
        n17444) );
  NAND2_X1 U19335 ( .A1(n22584), .A2(n17442), .ZN(n17443) );
  NAND2_X1 U19336 ( .A1(n17444), .A2(n17443), .ZN(n17445) );
  AOI222_X1 U19337 ( .A1(n17461), .A2(n22585), .B1(n17461), .B2(n17445), .C1(
        n22585), .C2(n17445), .ZN(n17446) );
  OR2_X1 U19338 ( .A1(n17446), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n17447) );
  AOI221_X1 U19339 ( .B1(n17448), .B2(n17447), .C1(n17446), .C2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17459) );
  INV_X1 U19340 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17717) );
  NAND2_X1 U19341 ( .A1(n17717), .A2(n14721), .ZN(n17452) );
  INV_X1 U19342 ( .A(n17449), .ZN(n17451) );
  AOI211_X1 U19343 ( .C1(n17453), .C2(n17452), .A(n17451), .B(n17450), .ZN(
        n17456) );
  NAND2_X1 U19344 ( .A1(n17454), .A2(n22132), .ZN(n17455) );
  OAI211_X1 U19345 ( .C1(n13350), .C2(n17457), .A(n17456), .B(n17455), .ZN(
        n17458) );
  AOI211_X1 U19346 ( .C1(n17461), .C2(n17460), .A(n17459), .B(n17458), .ZN(
        n22304) );
  INV_X1 U19347 ( .A(n22304), .ZN(n17468) );
  NAND4_X1 U19348 ( .A1(n17465), .A2(n17464), .A3(n17463), .A4(n17462), .ZN(
        n17467) );
  OAI21_X1 U19349 ( .B1(n15308), .B2(n17473), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n22291) );
  INV_X1 U19350 ( .A(n22291), .ZN(n17466) );
  NAND2_X1 U19351 ( .A1(n22325), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n22293) );
  NAND3_X1 U19352 ( .A1(n17467), .A2(n17466), .A3(n22293), .ZN(n17471) );
  AOI221_X1 U19353 ( .B1(n17473), .B2(n15308), .C1(n17468), .C2(n15308), .A(
        n17471), .ZN(n22296) );
  NOR2_X1 U19354 ( .A1(n22296), .A2(n17473), .ZN(n22295) );
  OAI211_X1 U19355 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n22325), .A(n22295), 
        .B(n17469), .ZN(n22300) );
  NAND2_X1 U19356 ( .A1(n22327), .A2(n22605), .ZN(n17472) );
  OAI211_X1 U19357 ( .C1(n17473), .C2(n17472), .A(n17471), .B(n17470), .ZN(
        n17474) );
  NAND2_X1 U19358 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n17474), .ZN(n17475) );
  OAI21_X1 U19359 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n22300), .A(n17475), 
        .ZN(P1_U3162) );
  NOR2_X1 U19360 ( .A1(n17477), .A2(n17476), .ZN(P1_U3032) );
  AND2_X1 U19361 ( .A1(n20474), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19362 ( .A1(n22324), .A2(n22343), .ZN(n17478) );
  INV_X1 U19363 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17544) );
  AOI21_X1 U19364 ( .B1(n17478), .B2(n17544), .A(n22853), .ZN(P1_U2802) );
  XOR2_X1 U19365 ( .A(n22420), .B(keyinput_254), .Z(n17830) );
  OAI22_X1 U19366 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_237), .B1(
        P1_EBX_REG_5__SCAN_IN), .B2(keyinput_238), .ZN(n17479) );
  AOI221_X1 U19367 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_237), .C1(
        keyinput_238), .C2(P1_EBX_REG_5__SCAN_IN), .A(n17479), .ZN(n17627) );
  INV_X1 U19368 ( .A(keyinput_236), .ZN(n17616) );
  INV_X1 U19369 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n22191) );
  XNOR2_X1 U19370 ( .A(n22191), .B(keyinput_233), .ZN(n17487) );
  AOI22_X1 U19371 ( .A1(n17481), .A2(keyinput_228), .B1(keyinput_229), .B2(
        n17794), .ZN(n17480) );
  OAI221_X1 U19372 ( .B1(n17481), .B2(keyinput_228), .C1(n17794), .C2(
        keyinput_229), .A(n17480), .ZN(n17486) );
  AOI22_X1 U19373 ( .A1(P1_EBX_REG_9__SCAN_IN), .A2(keyinput_234), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_230), .ZN(n17482) );
  OAI221_X1 U19374 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(keyinput_234), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_230), .A(n17482), .ZN(n17485) );
  AOI22_X1 U19375 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_232), .B1(
        P1_EBX_REG_12__SCAN_IN), .B2(keyinput_231), .ZN(n17483) );
  OAI221_X1 U19376 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_232), .C1(
        P1_EBX_REG_12__SCAN_IN), .C2(keyinput_231), .A(n17483), .ZN(n17484) );
  NOR4_X1 U19377 ( .A1(n17487), .A2(n17486), .A3(n17485), .A4(n17484), .ZN(
        n17613) );
  AOI22_X1 U19378 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput_213), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(keyinput_214), .ZN(n17488) );
  OAI221_X1 U19379 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput_213), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput_214), .A(n17488), .ZN(n17593) );
  INV_X1 U19380 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n22192) );
  OAI22_X1 U19381 ( .A1(n22192), .A2(keyinput_201), .B1(keyinput_202), .B2(
        P1_REIP_REG_9__SCAN_IN), .ZN(n17489) );
  AOI221_X1 U19382 ( .B1(n22192), .B2(keyinput_201), .C1(
        P1_REIP_REG_9__SCAN_IN), .C2(keyinput_202), .A(n17489), .ZN(n17584) );
  OAI22_X1 U19383 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_192), .B1(
        keyinput_188), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n17490) );
  AOI221_X1 U19384 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_192), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_188), .A(n17490), .ZN(n17577)
         );
  XNOR2_X1 U19385 ( .A(n17643), .B(keyinput_187), .ZN(n17571) );
  INV_X1 U19386 ( .A(keyinput_186), .ZN(n17565) );
  INV_X1 U19387 ( .A(keyinput_180), .ZN(n17557) );
  AOI22_X1 U19388 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_171), 
        .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_172), .ZN(n17491) );
  OAI221_X1 U19389 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_171), 
        .C1(P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_172), .A(n17491), .ZN(
        n17549) );
  INV_X1 U19390 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n17548) );
  AOI22_X1 U19391 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_168), .B1(
        n22851), .B2(keyinput_169), .ZN(n17492) );
  OAI221_X1 U19392 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_168), .C1(
        n22851), .C2(keyinput_169), .A(n17492), .ZN(n17546) );
  INV_X1 U19393 ( .A(READY2), .ZN(n17494) );
  AOI22_X1 U19394 ( .A1(n17494), .A2(keyinput_165), .B1(n20701), .B2(
        keyinput_166), .ZN(n17493) );
  OAI221_X1 U19395 ( .B1(n17494), .B2(keyinput_165), .C1(n20701), .C2(
        keyinput_166), .A(n17493), .ZN(n17542) );
  INV_X1 U19396 ( .A(keyinput_154), .ZN(n17524) );
  INV_X1 U19397 ( .A(DATAI_9_), .ZN(n17496) );
  AOI22_X1 U19398 ( .A1(DATAI_8_), .A2(keyinput_152), .B1(n17496), .B2(
        keyinput_151), .ZN(n17495) );
  OAI221_X1 U19399 ( .B1(DATAI_8_), .B2(keyinput_152), .C1(n17496), .C2(
        keyinput_151), .A(n17495), .ZN(n17522) );
  INV_X1 U19400 ( .A(keyinput_150), .ZN(n17521) );
  INV_X1 U19401 ( .A(DATAI_10_), .ZN(n17684) );
  XOR2_X1 U19402 ( .A(DATAI_15_), .B(keyinput_145), .Z(n17520) );
  INV_X1 U19403 ( .A(keyinput_144), .ZN(n17514) );
  OAI22_X1 U19404 ( .A1(n17652), .A2(keyinput_134), .B1(n17651), .B2(
        keyinput_135), .ZN(n17497) );
  AOI221_X1 U19405 ( .B1(n17652), .B2(keyinput_134), .C1(keyinput_135), .C2(
        n17651), .A(n17497), .ZN(n17504) );
  INV_X1 U19406 ( .A(DATAI_24_), .ZN(n17502) );
  INV_X1 U19407 ( .A(DATAI_28_), .ZN(n17658) );
  INV_X1 U19408 ( .A(DATAI_30_), .ZN(n17654) );
  AOI22_X1 U19409 ( .A1(DATAI_29_), .A2(keyinput_131), .B1(n17654), .B2(
        keyinput_130), .ZN(n17498) );
  OAI221_X1 U19410 ( .B1(DATAI_29_), .B2(keyinput_131), .C1(n17654), .C2(
        keyinput_130), .A(n17498), .ZN(n17501) );
  OAI22_X1 U19411 ( .A1(DATAI_31_), .A2(keyinput_129), .B1(keyinput_128), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n17499) );
  AOI221_X1 U19412 ( .B1(DATAI_31_), .B2(keyinput_129), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_128), .A(n17499), .ZN(n17500) );
  AOI22_X1 U19413 ( .A1(n17504), .A2(n17503), .B1(DATAI_22_), .B2(keyinput_138), .ZN(n17505) );
  OAI21_X1 U19414 ( .B1(DATAI_22_), .B2(keyinput_138), .A(n17505), .ZN(n17512)
         );
  AOI22_X1 U19415 ( .A1(DATAI_23_), .A2(keyinput_137), .B1(DATAI_21_), .B2(
        keyinput_139), .ZN(n17506) );
  OAI221_X1 U19416 ( .B1(DATAI_23_), .B2(keyinput_137), .C1(DATAI_21_), .C2(
        keyinput_139), .A(n17506), .ZN(n17511) );
  OAI22_X1 U19417 ( .A1(n17665), .A2(keyinput_141), .B1(keyinput_140), .B2(
        DATAI_20_), .ZN(n17507) );
  AOI221_X1 U19418 ( .B1(n17665), .B2(keyinput_141), .C1(DATAI_20_), .C2(
        keyinput_140), .A(n17507), .ZN(n17510) );
  OAI22_X1 U19419 ( .A1(DATAI_17_), .A2(keyinput_143), .B1(DATAI_18_), .B2(
        keyinput_142), .ZN(n17508) );
  AOI221_X1 U19420 ( .B1(DATAI_17_), .B2(keyinput_143), .C1(keyinput_142), 
        .C2(DATAI_18_), .A(n17508), .ZN(n17509) );
  OAI211_X1 U19421 ( .C1(n17512), .C2(n17511), .A(n17510), .B(n17509), .ZN(
        n17513) );
  OAI221_X1 U19422 ( .B1(DATAI_16_), .B2(keyinput_144), .C1(n17673), .C2(
        n17514), .A(n17513), .ZN(n17519) );
  AOI22_X1 U19423 ( .A1(DATAI_13_), .A2(keyinput_147), .B1(DATAI_14_), .B2(
        keyinput_146), .ZN(n17515) );
  OAI221_X1 U19424 ( .B1(DATAI_13_), .B2(keyinput_147), .C1(DATAI_14_), .C2(
        keyinput_146), .A(n17515), .ZN(n17518) );
  AOI22_X1 U19425 ( .A1(DATAI_11_), .A2(keyinput_149), .B1(DATAI_12_), .B2(
        keyinput_148), .ZN(n17516) );
  OAI221_X1 U19426 ( .B1(DATAI_11_), .B2(keyinput_149), .C1(DATAI_12_), .C2(
        keyinput_148), .A(n17516), .ZN(n17517) );
  AOI221_X1 U19427 ( .B1(DATAI_6_), .B2(n17524), .C1(n17690), .C2(keyinput_154), .A(n17523), .ZN(n17531) );
  INV_X1 U19428 ( .A(DATAI_5_), .ZN(n17526) );
  AOI22_X1 U19429 ( .A1(n17527), .A2(keyinput_156), .B1(n17526), .B2(
        keyinput_155), .ZN(n17525) );
  OAI221_X1 U19430 ( .B1(n17527), .B2(keyinput_156), .C1(n17526), .C2(
        keyinput_155), .A(n17525), .ZN(n17530) );
  INV_X1 U19431 ( .A(DATAI_2_), .ZN(n17694) );
  OAI22_X1 U19432 ( .A1(n17694), .A2(keyinput_158), .B1(keyinput_157), .B2(
        DATAI_3_), .ZN(n17528) );
  AOI221_X1 U19433 ( .B1(n17694), .B2(keyinput_158), .C1(DATAI_3_), .C2(
        keyinput_157), .A(n17528), .ZN(n17529) );
  OAI21_X1 U19434 ( .B1(n17531), .B2(n17530), .A(n17529), .ZN(n17540) );
  OAI22_X1 U19435 ( .A1(n17533), .A2(keyinput_163), .B1(HOLD), .B2(
        keyinput_161), .ZN(n17532) );
  AOI221_X1 U19436 ( .B1(n17533), .B2(keyinput_163), .C1(keyinput_161), .C2(
        HOLD), .A(n17532), .ZN(n17536) );
  INV_X1 U19437 ( .A(NA), .ZN(n22378) );
  OAI22_X1 U19438 ( .A1(n22378), .A2(keyinput_162), .B1(keyinput_159), .B2(
        DATAI_1_), .ZN(n17534) );
  AOI221_X1 U19439 ( .B1(n22378), .B2(keyinput_162), .C1(DATAI_1_), .C2(
        keyinput_159), .A(n17534), .ZN(n17535) );
  OAI211_X1 U19440 ( .C1(DATAI_0_), .C2(keyinput_160), .A(n17536), .B(n17535), 
        .ZN(n17537) );
  AOI21_X1 U19441 ( .B1(DATAI_0_), .B2(keyinput_160), .A(n17537), .ZN(n17539)
         );
  NOR2_X1 U19442 ( .A1(READY1), .A2(keyinput_164), .ZN(n17538) );
  AOI221_X1 U19443 ( .B1(n17540), .B2(n17539), .C1(keyinput_164), .C2(READY1), 
        .A(n17538), .ZN(n17541) );
  OAI22_X1 U19444 ( .A1(keyinput_167), .A2(n17544), .B1(n17542), .B2(n17541), 
        .ZN(n17543) );
  AOI21_X1 U19445 ( .B1(keyinput_167), .B2(n17544), .A(n17543), .ZN(n17545) );
  OAI22_X1 U19446 ( .A1(keyinput_170), .A2(n17548), .B1(n17546), .B2(n17545), 
        .ZN(n17547) );
  AOI22_X1 U19447 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_176), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_174), .ZN(n17550) );
  OAI221_X1 U19448 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_176), 
        .C1(P1_FLUSH_REG_SCAN_IN), .C2(keyinput_174), .A(n17550), .ZN(n17555)
         );
  AOI22_X1 U19449 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_175), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_178), .ZN(n17551) );
  OAI221_X1 U19450 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_175), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_178), .A(n17551), .ZN(
        n17554) );
  AOI22_X1 U19451 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_177), .B1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_179), .ZN(n17552) );
  OAI221_X1 U19452 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_177), 
        .C1(P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_179), .A(n17552), .ZN(
        n17553) );
  AOI221_X1 U19453 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n17557), .C1(n20521), 
        .C2(keyinput_180), .A(n17556), .ZN(n17563) );
  XOR2_X1 U19454 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_181), .Z(n17562)
         );
  OAI22_X1 U19455 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_184), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_183), .ZN(n17558) );
  AOI221_X1 U19456 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_184), .C1(
        keyinput_183), .C2(P1_REIP_REG_28__SCAN_IN), .A(n17558), .ZN(n17561)
         );
  OAI22_X1 U19457 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_182), .B1(
        keyinput_185), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n17559) );
  AOI221_X1 U19458 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_182), .C1(
        P1_REIP_REG_26__SCAN_IN), .C2(keyinput_185), .A(n17559), .ZN(n17560)
         );
  OAI211_X1 U19459 ( .C1(n17563), .C2(n17562), .A(n17561), .B(n17560), .ZN(
        n17564) );
  OAI221_X1 U19460 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_186), .C1(
        n17734), .C2(n17565), .A(n17564), .ZN(n17570) );
  INV_X1 U19461 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20500) );
  AOI22_X1 U19462 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_191), .B1(
        n20500), .B2(keyinput_193), .ZN(n17566) );
  OAI221_X1 U19463 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_191), .C1(
        n20500), .C2(keyinput_193), .A(n17566), .ZN(n17569) );
  AOI22_X1 U19464 ( .A1(n17737), .A2(keyinput_189), .B1(n20504), .B2(
        keyinput_190), .ZN(n17567) );
  OAI221_X1 U19465 ( .B1(n17737), .B2(keyinput_189), .C1(n20504), .C2(
        keyinput_190), .A(n17567), .ZN(n17568) );
  INV_X1 U19466 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n17743) );
  AOI22_X1 U19467 ( .A1(n17743), .A2(keyinput_194), .B1(keyinput_196), .B2(
        n17744), .ZN(n17572) );
  OAI221_X1 U19468 ( .B1(n17743), .B2(keyinput_194), .C1(n17744), .C2(
        keyinput_196), .A(n17572), .ZN(n17576) );
  INV_X1 U19469 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U19470 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_197), .B1(
        n17574), .B2(keyinput_195), .ZN(n17573) );
  OAI221_X1 U19471 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_197), .C1(
        n17574), .C2(keyinput_195), .A(n17573), .ZN(n17575) );
  AOI22_X1 U19472 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(keyinput_200), .B1(
        n17751), .B2(keyinput_198), .ZN(n17578) );
  OAI221_X1 U19473 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(keyinput_200), .C1(
        n17751), .C2(keyinput_198), .A(n17578), .ZN(n17579) );
  XOR2_X1 U19474 ( .A(P1_REIP_REG_6__SCAN_IN), .B(keyinput_205), .Z(n17582) );
  AOI22_X1 U19475 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_203), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(keyinput_204), .ZN(n17580) );
  OAI221_X1 U19476 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_203), .C1(
        P1_REIP_REG_7__SCAN_IN), .C2(keyinput_204), .A(n17580), .ZN(n17581) );
  AOI211_X1 U19477 ( .C1(n17584), .C2(n17583), .A(n17582), .B(n17581), .ZN(
        n17589) );
  AOI22_X1 U19478 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_207), .B1(n22150), .B2(keyinput_206), .ZN(n17585) );
  OAI221_X1 U19479 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_207), .C1(
        n22150), .C2(keyinput_206), .A(n17585), .ZN(n17588) );
  OAI22_X1 U19480 ( .A1(n22124), .A2(keyinput_209), .B1(keyinput_208), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n17586) );
  AOI221_X1 U19481 ( .B1(n22124), .B2(keyinput_209), .C1(
        P1_REIP_REG_3__SCAN_IN), .C2(keyinput_208), .A(n17586), .ZN(n17587) );
  OAI22_X1 U19482 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(keyinput_210), .B1(
        keyinput_211), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n17590) );
  AOI221_X1 U19483 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(keyinput_210), .C1(
        P1_REIP_REG_0__SCAN_IN), .C2(keyinput_211), .A(n17590), .ZN(n17592) );
  NOR2_X1 U19484 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_212), .ZN(n17591)
         );
  OAI22_X1 U19485 ( .A1(n17596), .A2(keyinput_216), .B1(keyinput_217), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n17595) );
  AOI221_X1 U19486 ( .B1(n17596), .B2(keyinput_216), .C1(
        P1_EBX_REG_26__SCAN_IN), .C2(keyinput_217), .A(n17595), .ZN(n17602) );
  AOI22_X1 U19487 ( .A1(P1_EBX_REG_22__SCAN_IN), .A2(keyinput_221), .B1(n17598), .B2(keyinput_220), .ZN(n17597) );
  OAI221_X1 U19488 ( .B1(P1_EBX_REG_22__SCAN_IN), .B2(keyinput_221), .C1(
        n17598), .C2(keyinput_220), .A(n17597), .ZN(n17601) );
  AOI22_X1 U19489 ( .A1(P1_EBX_REG_24__SCAN_IN), .A2(keyinput_219), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_218), .ZN(n17599) );
  OAI221_X1 U19490 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(keyinput_219), .C1(
        P1_EBX_REG_25__SCAN_IN), .C2(keyinput_218), .A(n17599), .ZN(n17600) );
  AOI211_X1 U19491 ( .C1(n17603), .C2(n17602), .A(n17601), .B(n17600), .ZN(
        n17611) );
  AOI22_X1 U19492 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_222), .B1(n17605), .B2(keyinput_223), .ZN(n17604) );
  OAI221_X1 U19493 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_222), .C1(
        n17605), .C2(keyinput_223), .A(n17604), .ZN(n17610) );
  OAI22_X1 U19494 ( .A1(n22237), .A2(keyinput_227), .B1(keyinput_226), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n17606) );
  AOI221_X1 U19495 ( .B1(n22237), .B2(keyinput_227), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput_226), .A(n17606), .ZN(n17609) );
  OAI22_X1 U19496 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(keyinput_224), .B1(
        keyinput_225), .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n17607) );
  AOI221_X1 U19497 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput_224), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_225), .A(n17607), .ZN(n17608) );
  OAI211_X1 U19498 ( .C1(n17611), .C2(n17610), .A(n17609), .B(n17608), .ZN(
        n17612) );
  AOI22_X1 U19499 ( .A1(n17613), .A2(n17612), .B1(keyinput_235), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n17614) );
  OAI21_X1 U19500 ( .B1(keyinput_235), .B2(P1_EBX_REG_8__SCAN_IN), .A(n17614), 
        .ZN(n17615) );
  OAI221_X1 U19501 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n17616), .C1(n14246), 
        .C2(keyinput_236), .A(n17615), .ZN(n17626) );
  AOI22_X1 U19502 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_244), .B1(n22481), .B2(keyinput_245), .ZN(n17617) );
  OAI221_X1 U19503 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_244), .C1(
        n22481), .C2(keyinput_245), .A(n17617), .ZN(n17625) );
  AOI22_X1 U19504 ( .A1(n17805), .A2(keyinput_242), .B1(n14225), .B2(
        keyinput_243), .ZN(n17618) );
  OAI221_X1 U19505 ( .B1(n17805), .B2(keyinput_242), .C1(n14225), .C2(
        keyinput_243), .A(n17618), .ZN(n17622) );
  AOI22_X1 U19506 ( .A1(P1_EBX_REG_2__SCAN_IN), .A2(keyinput_241), .B1(n17620), 
        .B2(keyinput_240), .ZN(n17619) );
  OAI221_X1 U19507 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(keyinput_241), .C1(n17620), .C2(keyinput_240), .A(n17619), .ZN(n17621) );
  AOI211_X1 U19508 ( .C1(keyinput_239), .C2(P1_EBX_REG_4__SCAN_IN), .A(n17622), 
        .B(n17621), .ZN(n17623) );
  OAI21_X1 U19509 ( .B1(keyinput_239), .B2(P1_EBX_REG_4__SCAN_IN), .A(n17623), 
        .ZN(n17624) );
  AOI22_X1 U19510 ( .A1(n22450), .A2(keyinput_249), .B1(n22465), .B2(
        keyinput_247), .ZN(n17628) );
  OAI221_X1 U19511 ( .B1(n22450), .B2(keyinput_249), .C1(n22465), .C2(
        keyinput_247), .A(n17628), .ZN(n17631) );
  AOI22_X1 U19512 ( .A1(P1_EAX_REG_27__SCAN_IN), .A2(keyinput_248), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_246), .ZN(n17629) );
  OAI221_X1 U19513 ( .B1(P1_EAX_REG_27__SCAN_IN), .B2(keyinput_248), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_246), .A(n17629), .ZN(n17630) );
  AOI22_X1 U19514 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_250), .B1(n22436), .B2(keyinput_251), .ZN(n17632) );
  OAI221_X1 U19515 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_250), .C1(
        n22436), .C2(keyinput_251), .A(n17632), .ZN(n17635) );
  OAI22_X1 U19516 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(keyinput_252), .B1(
        keyinput_253), .B2(P1_EAX_REG_22__SCAN_IN), .ZN(n17633) );
  AOI221_X1 U19517 ( .B1(P1_EAX_REG_23__SCAN_IN), .B2(keyinput_252), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_253), .A(n17633), .ZN(n17634) );
  INV_X1 U19518 ( .A(keyinput_126), .ZN(n17824) );
  INV_X1 U19519 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n22154) );
  OAI22_X1 U19520 ( .A1(n22154), .A2(keyinput_109), .B1(n14238), .B2(
        keyinput_110), .ZN(n17636) );
  AOI221_X1 U19521 ( .B1(n22154), .B2(keyinput_109), .C1(keyinput_110), .C2(
        n14238), .A(n17636), .ZN(n17812) );
  INV_X1 U19522 ( .A(keyinput_108), .ZN(n17801) );
  OAI22_X1 U19523 ( .A1(n17638), .A2(keyinput_94), .B1(keyinput_95), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n17637) );
  AOI221_X1 U19524 ( .B1(n17638), .B2(keyinput_94), .C1(P1_EBX_REG_20__SCAN_IN), .C2(keyinput_95), .A(n17637), .ZN(n17787) );
  OAI22_X1 U19525 ( .A1(n17640), .A2(keyinput_85), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(keyinput_86), .ZN(n17639) );
  AOI221_X1 U19526 ( .B1(n17640), .B2(keyinput_85), .C1(keyinput_86), .C2(
        P1_EBX_REG_29__SCAN_IN), .A(n17639), .ZN(n17770) );
  OAI22_X1 U19527 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(keyinput_74), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(keyinput_73), .ZN(n17641) );
  AOI221_X1 U19528 ( .B1(P1_REIP_REG_9__SCAN_IN), .B2(keyinput_74), .C1(
        keyinput_73), .C2(P1_REIP_REG_10__SCAN_IN), .A(n17641), .ZN(n17758) );
  OAI22_X1 U19529 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(keyinput_64), .B1(
        keyinput_63), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n17642) );
  AOI221_X1 U19530 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(keyinput_64), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(keyinput_63), .A(n17642), .ZN(n17749) );
  XOR2_X1 U19531 ( .A(n17643), .B(keyinput_59), .Z(n17741) );
  INV_X1 U19532 ( .A(keyinput_58), .ZN(n17733) );
  INV_X1 U19533 ( .A(keyinput_52), .ZN(n17725) );
  INV_X1 U19534 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22328) );
  AOI22_X1 U19535 ( .A1(keyinput_44), .A2(P1_STATEBS16_REG_SCAN_IN), .B1(
        n22328), .B2(keyinput_43), .ZN(n17644) );
  OAI221_X1 U19536 ( .B1(keyinput_44), .B2(P1_STATEBS16_REG_SCAN_IN), .C1(
        n22328), .C2(keyinput_43), .A(n17644), .ZN(n17716) );
  INV_X1 U19537 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17646) );
  AOI22_X1 U19538 ( .A1(n22851), .A2(keyinput_41), .B1(keyinput_40), .B2(
        n17646), .ZN(n17645) );
  OAI221_X1 U19539 ( .B1(n22851), .B2(keyinput_41), .C1(n17646), .C2(
        keyinput_40), .A(n17645), .ZN(n17714) );
  AOI22_X1 U19540 ( .A1(READY2), .A2(keyinput_37), .B1(n20701), .B2(
        keyinput_38), .ZN(n17647) );
  OAI221_X1 U19541 ( .B1(READY2), .B2(keyinput_37), .C1(n20701), .C2(
        keyinput_38), .A(n17647), .ZN(n17711) );
  OAI22_X1 U19542 ( .A1(DATAI_5_), .A2(keyinput_27), .B1(DATAI_4_), .B2(
        keyinput_28), .ZN(n17648) );
  AOI221_X1 U19543 ( .B1(DATAI_5_), .B2(keyinput_27), .C1(keyinput_28), .C2(
        DATAI_4_), .A(n17648), .ZN(n17697) );
  AOI22_X1 U19544 ( .A1(DATAI_8_), .A2(keyinput_24), .B1(DATAI_9_), .B2(
        keyinput_23), .ZN(n17649) );
  OAI221_X1 U19545 ( .B1(DATAI_8_), .B2(keyinput_24), .C1(DATAI_9_), .C2(
        keyinput_23), .A(n17649), .ZN(n17688) );
  INV_X1 U19546 ( .A(keyinput_22), .ZN(n17685) );
  XOR2_X1 U19547 ( .A(DATAI_15_), .B(keyinput_17), .Z(n17683) );
  INV_X1 U19548 ( .A(keyinput_16), .ZN(n17674) );
  OAI22_X1 U19549 ( .A1(n17652), .A2(keyinput_6), .B1(n17651), .B2(keyinput_7), 
        .ZN(n17650) );
  AOI221_X1 U19550 ( .B1(n17652), .B2(keyinput_6), .C1(keyinput_7), .C2(n17651), .A(n17650), .ZN(n17660) );
  AOI22_X1 U19551 ( .A1(DATAI_29_), .A2(keyinput_3), .B1(n17654), .B2(
        keyinput_2), .ZN(n17653) );
  OAI221_X1 U19552 ( .B1(DATAI_29_), .B2(keyinput_3), .C1(n17654), .C2(
        keyinput_2), .A(n17653), .ZN(n17657) );
  OAI22_X1 U19553 ( .A1(DATAI_31_), .A2(keyinput_1), .B1(keyinput_0), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n17655) );
  AOI22_X1 U19554 ( .A1(n17660), .A2(n17659), .B1(DATAI_22_), .B2(keyinput_10), 
        .ZN(n17661) );
  OAI21_X1 U19555 ( .B1(DATAI_22_), .B2(keyinput_10), .A(n17661), .ZN(n17671)
         );
  AOI22_X1 U19556 ( .A1(keyinput_11), .A2(DATAI_21_), .B1(n17663), .B2(
        keyinput_9), .ZN(n17662) );
  OAI221_X1 U19557 ( .B1(keyinput_11), .B2(DATAI_21_), .C1(n17663), .C2(
        keyinput_9), .A(n17662), .ZN(n17670) );
  OAI22_X1 U19558 ( .A1(n17665), .A2(keyinput_13), .B1(n16199), .B2(
        keyinput_12), .ZN(n17664) );
  AOI221_X1 U19559 ( .B1(n17665), .B2(keyinput_13), .C1(keyinput_12), .C2(
        n16199), .A(n17664), .ZN(n17669) );
  OAI22_X1 U19560 ( .A1(n17667), .A2(keyinput_15), .B1(DATAI_18_), .B2(
        keyinput_14), .ZN(n17666) );
  AOI221_X1 U19561 ( .B1(n17667), .B2(keyinput_15), .C1(keyinput_14), .C2(
        DATAI_18_), .A(n17666), .ZN(n17668) );
  OAI211_X1 U19562 ( .C1(n17671), .C2(n17670), .A(n17669), .B(n17668), .ZN(
        n17672) );
  OAI221_X1 U19563 ( .B1(DATAI_16_), .B2(n17674), .C1(n17673), .C2(keyinput_16), .A(n17672), .ZN(n17682) );
  INV_X1 U19564 ( .A(DATAI_13_), .ZN(n17677) );
  INV_X1 U19565 ( .A(DATAI_14_), .ZN(n17676) );
  AOI22_X1 U19566 ( .A1(n17677), .A2(keyinput_19), .B1(n17676), .B2(
        keyinput_18), .ZN(n17675) );
  OAI221_X1 U19567 ( .B1(n17677), .B2(keyinput_19), .C1(n17676), .C2(
        keyinput_18), .A(n17675), .ZN(n17681) );
  INV_X1 U19568 ( .A(DATAI_11_), .ZN(n17679) );
  AOI22_X1 U19569 ( .A1(DATAI_12_), .A2(keyinput_20), .B1(n17679), .B2(
        keyinput_21), .ZN(n17678) );
  OAI221_X1 U19570 ( .B1(DATAI_12_), .B2(keyinput_20), .C1(n17679), .C2(
        keyinput_21), .A(n17678), .ZN(n17680) );
  INV_X1 U19571 ( .A(DATAI_7_), .ZN(n17687) );
  NAND2_X1 U19572 ( .A1(n17687), .A2(keyinput_25), .ZN(n17686) );
  INV_X1 U19573 ( .A(keyinput_26), .ZN(n17689) );
  AOI22_X1 U19574 ( .A1(keyinput_29), .A2(DATAI_3_), .B1(n17694), .B2(
        keyinput_30), .ZN(n17693) );
  OAI221_X1 U19575 ( .B1(keyinput_29), .B2(DATAI_3_), .C1(n17694), .C2(
        keyinput_30), .A(n17693), .ZN(n17695) );
  AOI21_X1 U19576 ( .B1(n17697), .B2(n17696), .A(n17695), .ZN(n17698) );
  INV_X1 U19577 ( .A(DATAI_1_), .ZN(n17700) );
  AOI22_X1 U19578 ( .A1(n22378), .A2(keyinput_34), .B1(keyinput_31), .B2(
        n17700), .ZN(n17699) );
  OAI221_X1 U19579 ( .B1(n22378), .B2(keyinput_34), .C1(n17700), .C2(
        keyinput_31), .A(n17699), .ZN(n17704) );
  INV_X1 U19580 ( .A(DATAI_0_), .ZN(n17702) );
  AOI22_X1 U19581 ( .A1(HOLD), .A2(keyinput_33), .B1(n17702), .B2(keyinput_32), 
        .ZN(n17701) );
  OAI221_X1 U19582 ( .B1(HOLD), .B2(keyinput_33), .C1(n17702), .C2(keyinput_32), .A(n17701), .ZN(n17703) );
  AOI211_X1 U19583 ( .C1(keyinput_35), .C2(BS16), .A(n17704), .B(n17703), .ZN(
        n17705) );
  OAI21_X1 U19584 ( .B1(keyinput_35), .B2(BS16), .A(n17705), .ZN(n17706) );
  INV_X1 U19585 ( .A(n17706), .ZN(n17708) );
  OAI22_X1 U19586 ( .A1(n17711), .A2(n17710), .B1(keyinput_39), .B2(
        P1_ADS_N_REG_SCAN_IN), .ZN(n17712) );
  AOI21_X1 U19587 ( .B1(keyinput_39), .B2(P1_ADS_N_REG_SCAN_IN), .A(n17712), 
        .ZN(n17713) );
  AOI22_X1 U19588 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_51), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_50), .ZN(n17718) );
  OAI221_X1 U19589 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_51), .C1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_50), .A(n17718), .ZN(
        n17723) );
  AOI22_X1 U19590 ( .A1(keyinput_47), .A2(P1_W_R_N_REG_SCAN_IN), .B1(n14721), 
        .B2(keyinput_46), .ZN(n17719) );
  OAI221_X1 U19591 ( .B1(keyinput_47), .B2(P1_W_R_N_REG_SCAN_IN), .C1(n14721), 
        .C2(keyinput_46), .A(n17719), .ZN(n17722) );
  INV_X1 U19592 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20542) );
  INV_X1 U19593 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20546) );
  AOI22_X1 U19594 ( .A1(n20542), .A2(keyinput_49), .B1(keyinput_48), .B2(
        n20546), .ZN(n17720) );
  OAI221_X1 U19595 ( .B1(n20542), .B2(keyinput_49), .C1(n20546), .C2(
        keyinput_48), .A(n17720), .ZN(n17721) );
  AOI221_X1 U19596 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n17725), .C1(n20521), 
        .C2(keyinput_52), .A(n17724), .ZN(n17731) );
  XOR2_X1 U19597 ( .A(P1_REIP_REG_30__SCAN_IN), .B(keyinput_53), .Z(n17730) );
  OAI22_X1 U19598 ( .A1(n20513), .A2(keyinput_56), .B1(keyinput_55), .B2(
        P1_REIP_REG_28__SCAN_IN), .ZN(n17726) );
  AOI221_X1 U19599 ( .B1(n20513), .B2(keyinput_56), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_55), .A(n17726), .ZN(n17729) );
  OAI22_X1 U19600 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_54), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .ZN(n17727) );
  AOI221_X1 U19601 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .C1(
        keyinput_57), .C2(P1_REIP_REG_26__SCAN_IN), .A(n17727), .ZN(n17728) );
  OAI211_X1 U19602 ( .C1(n17731), .C2(n17730), .A(n17729), .B(n17728), .ZN(
        n17732) );
  OAI221_X1 U19603 ( .B1(P1_REIP_REG_25__SCAN_IN), .B2(keyinput_58), .C1(
        n17734), .C2(n17733), .A(n17732), .ZN(n17740) );
  AOI22_X1 U19604 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(keyinput_60), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .ZN(n17735) );
  OAI221_X1 U19605 ( .B1(P1_REIP_REG_23__SCAN_IN), .B2(keyinput_60), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_62), .A(n17735), .ZN(n17739) );
  AOI22_X1 U19606 ( .A1(n17737), .A2(keyinput_61), .B1(n20500), .B2(
        keyinput_65), .ZN(n17736) );
  OAI221_X1 U19607 ( .B1(n17737), .B2(keyinput_61), .C1(n20500), .C2(
        keyinput_65), .A(n17736), .ZN(n17738) );
  AOI22_X1 U19608 ( .A1(n17744), .A2(keyinput_68), .B1(n17743), .B2(
        keyinput_66), .ZN(n17742) );
  OAI221_X1 U19609 ( .B1(n17744), .B2(keyinput_68), .C1(n17743), .C2(
        keyinput_66), .A(n17742), .ZN(n17748) );
  INV_X1 U19610 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n17746) );
  AOI22_X1 U19611 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_67), .B1(n17746), .B2(keyinput_69), .ZN(n17745) );
  OAI221_X1 U19612 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_67), .C1(
        n17746), .C2(keyinput_69), .A(n17745), .ZN(n17747) );
  AOI22_X1 U19613 ( .A1(n17751), .A2(keyinput_70), .B1(keyinput_72), .B2(
        n22211), .ZN(n17750) );
  OAI221_X1 U19614 ( .B1(n17751), .B2(keyinput_70), .C1(n22211), .C2(
        keyinput_72), .A(n17750), .ZN(n17752) );
  XNOR2_X1 U19615 ( .A(n17753), .B(keyinput_75), .ZN(n17756) );
  AOI22_X1 U19616 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(keyinput_76), .B1(
        P1_REIP_REG_6__SCAN_IN), .B2(keyinput_77), .ZN(n17754) );
  OAI221_X1 U19617 ( .B1(P1_REIP_REG_7__SCAN_IN), .B2(keyinput_76), .C1(
        P1_REIP_REG_6__SCAN_IN), .C2(keyinput_77), .A(n17754), .ZN(n17755) );
  AOI211_X1 U19618 ( .C1(n17758), .C2(n17757), .A(n17756), .B(n17755), .ZN(
        n17763) );
  AOI22_X1 U19619 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_79), .B1(n22150), 
        .B2(keyinput_78), .ZN(n17759) );
  OAI221_X1 U19620 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_79), .C1(n22150), .C2(keyinput_78), .A(n17759), .ZN(n17762) );
  OAI22_X1 U19621 ( .A1(n22124), .A2(keyinput_81), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(keyinput_80), .ZN(n17760) );
  AOI221_X1 U19622 ( .B1(n22124), .B2(keyinput_81), .C1(keyinput_80), .C2(
        P1_REIP_REG_3__SCAN_IN), .A(n17760), .ZN(n17761) );
  OAI21_X1 U19623 ( .B1(n17763), .B2(n17762), .A(n17761), .ZN(n17767) );
  INV_X1 U19624 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20547) );
  OAI22_X1 U19625 ( .A1(n14610), .A2(keyinput_82), .B1(n20547), .B2(
        keyinput_83), .ZN(n17764) );
  AOI221_X1 U19626 ( .B1(n14610), .B2(keyinput_82), .C1(keyinput_83), .C2(
        n20547), .A(n17764), .ZN(n17766) );
  AOI22_X1 U19627 ( .A1(n17770), .A2(n17769), .B1(keyinput_89), .B2(n17772), 
        .ZN(n17771) );
  OAI21_X1 U19628 ( .B1(keyinput_89), .B2(n17772), .A(n17771), .ZN(n17780) );
  AOI22_X1 U19629 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_88), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_87), .ZN(n17773) );
  OAI221_X1 U19630 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_88), .C1(
        P1_EBX_REG_28__SCAN_IN), .C2(keyinput_87), .A(n17773), .ZN(n17779) );
  OAI22_X1 U19631 ( .A1(n17775), .A2(keyinput_91), .B1(keyinput_90), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n17774) );
  AOI221_X1 U19632 ( .B1(n17775), .B2(keyinput_91), .C1(P1_EBX_REG_25__SCAN_IN), .C2(keyinput_90), .A(n17774), .ZN(n17778) );
  OAI22_X1 U19633 ( .A1(P1_EBX_REG_23__SCAN_IN), .A2(keyinput_92), .B1(
        keyinput_93), .B2(P1_EBX_REG_22__SCAN_IN), .ZN(n17776) );
  AOI221_X1 U19634 ( .B1(P1_EBX_REG_23__SCAN_IN), .B2(keyinput_92), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_93), .A(n17776), .ZN(n17777) );
  AOI22_X1 U19635 ( .A1(n22237), .A2(keyinput_99), .B1(n17782), .B2(
        keyinput_96), .ZN(n17781) );
  OAI221_X1 U19636 ( .B1(n22237), .B2(keyinput_99), .C1(n17782), .C2(
        keyinput_96), .A(n17781), .ZN(n17785) );
  AOI22_X1 U19637 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput_98), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(keyinput_97), .ZN(n17783) );
  OAI221_X1 U19638 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput_98), .C1(
        P1_EBX_REG_18__SCAN_IN), .C2(keyinput_97), .A(n17783), .ZN(n17784) );
  OAI22_X1 U19639 ( .A1(n17789), .A2(keyinput_102), .B1(keyinput_106), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n17788) );
  AOI221_X1 U19640 ( .B1(n17789), .B2(keyinput_102), .C1(P1_EBX_REG_9__SCAN_IN), .C2(keyinput_106), .A(n17788), .ZN(n17790) );
  OAI21_X1 U19641 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(keyinput_100), .A(n17790), 
        .ZN(n17791) );
  OAI22_X1 U19642 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_103), .B1(
        P1_EBX_REG_11__SCAN_IN), .B2(keyinput_104), .ZN(n17792) );
  AOI221_X1 U19643 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_103), .C1(
        keyinput_104), .C2(P1_EBX_REG_11__SCAN_IN), .A(n17792), .ZN(n17796) );
  OAI22_X1 U19644 ( .A1(n17794), .A2(keyinput_101), .B1(n22191), .B2(
        keyinput_105), .ZN(n17793) );
  AOI221_X1 U19645 ( .B1(n17794), .B2(keyinput_101), .C1(keyinput_105), .C2(
        n22191), .A(n17793), .ZN(n17795) );
  INV_X1 U19646 ( .A(keyinput_107), .ZN(n17797) );
  OAI221_X1 U19647 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n17801), .C1(n14246), 
        .C2(keyinput_108), .A(n17800), .ZN(n17811) );
  AOI22_X1 U19648 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_116), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(keyinput_117), .ZN(n17802) );
  OAI221_X1 U19649 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_116), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_117), .A(n17802), .ZN(n17810) );
  AOI22_X1 U19650 ( .A1(P1_EBX_REG_3__SCAN_IN), .A2(keyinput_112), .B1(
        P1_EBX_REG_4__SCAN_IN), .B2(keyinput_111), .ZN(n17803) );
  OAI221_X1 U19651 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(keyinput_112), .C1(
        P1_EBX_REG_4__SCAN_IN), .C2(keyinput_111), .A(n17803), .ZN(n17807) );
  AOI22_X1 U19652 ( .A1(P1_EBX_REG_0__SCAN_IN), .A2(keyinput_115), .B1(n17805), 
        .B2(keyinput_114), .ZN(n17804) );
  OAI221_X1 U19653 ( .B1(P1_EBX_REG_0__SCAN_IN), .B2(keyinput_115), .C1(n17805), .C2(keyinput_114), .A(n17804), .ZN(n17806) );
  AOI211_X1 U19654 ( .C1(keyinput_113), .C2(P1_EBX_REG_2__SCAN_IN), .A(n17807), 
        .B(n17806), .ZN(n17808) );
  OAI21_X1 U19655 ( .B1(keyinput_113), .B2(P1_EBX_REG_2__SCAN_IN), .A(n17808), 
        .ZN(n17809) );
  AOI211_X1 U19656 ( .C1(n17812), .C2(n17811), .A(n17810), .B(n17809), .ZN(
        n17817) );
  AOI22_X1 U19657 ( .A1(n22465), .A2(keyinput_119), .B1(keyinput_120), .B2(
        n22458), .ZN(n17813) );
  OAI221_X1 U19658 ( .B1(n22465), .B2(keyinput_119), .C1(n22458), .C2(
        keyinput_120), .A(n17813), .ZN(n17816) );
  AOI22_X1 U19659 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(keyinput_121), .B1(n22472), .B2(keyinput_118), .ZN(n17814) );
  OAI221_X1 U19660 ( .B1(P1_EAX_REG_26__SCAN_IN), .B2(keyinput_121), .C1(
        n22472), .C2(keyinput_118), .A(n17814), .ZN(n17815) );
  NOR3_X1 U19661 ( .A1(n17817), .A2(n17816), .A3(n17815), .ZN(n17822) );
  AOI22_X1 U19662 ( .A1(n22443), .A2(keyinput_122), .B1(keyinput_123), .B2(
        n22436), .ZN(n17818) );
  OAI221_X1 U19663 ( .B1(n22443), .B2(keyinput_122), .C1(n22436), .C2(
        keyinput_123), .A(n17818), .ZN(n17821) );
  OAI22_X1 U19664 ( .A1(n22430), .A2(keyinput_124), .B1(keyinput_125), .B2(
        P1_EAX_REG_22__SCAN_IN), .ZN(n17819) );
  AOI221_X1 U19665 ( .B1(n22430), .B2(keyinput_124), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput_125), .A(n17819), .ZN(n17820) );
  OAI21_X1 U19666 ( .B1(n17822), .B2(n17821), .A(n17820), .ZN(n17823) );
  OAI221_X1 U19667 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(n17824), .C1(n22420), 
        .C2(keyinput_126), .A(n17823), .ZN(n17826) );
  AOI21_X1 U19668 ( .B1(n17826), .B2(keyinput_127), .A(keyinput_255), .ZN(
        n17828) );
  INV_X1 U19669 ( .A(keyinput_127), .ZN(n17825) );
  AOI21_X1 U19670 ( .B1(n17826), .B2(n17825), .A(n22413), .ZN(n17827) );
  AOI22_X1 U19671 ( .A1(n22413), .A2(n17828), .B1(keyinput_255), .B2(n17827), 
        .ZN(n17829) );
  OAI22_X1 U19672 ( .A1(n17832), .A2(n22663), .B1(n17831), .B2(n22659), .ZN(
        n17836) );
  OAI22_X1 U19673 ( .A1(n17834), .A2(n22667), .B1(n22673), .B2(n17833), .ZN(
        n17835) );
  AOI211_X1 U19674 ( .C1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .C2(n17837), .A(
        n17836), .B(n17835), .ZN(n17838) );
  XNOR2_X1 U19675 ( .A(n17839), .B(n17838), .ZN(P1_U3099) );
  AOI22_X1 U19676 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n17840), .B1(n19012), 
        .B2(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17841) );
  INV_X1 U19677 ( .A(n17841), .ZN(P2_U2816) );
  AOI22_X1 U19678 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19124), .B1(n17862), 
        .B2(n17842), .ZN(n17848) );
  AOI222_X1 U19679 ( .A1(n17846), .A2(n17871), .B1(n17870), .B2(n17845), .C1(
        n17844), .C2(n17843), .ZN(n17847) );
  OAI211_X1 U19680 ( .C1(n17849), .C2(n17877), .A(n17848), .B(n17847), .ZN(
        P2_U3010) );
  AOI22_X1 U19681 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19124), .B1(n17862), 
        .B2(n19051), .ZN(n17859) );
  NOR2_X1 U19682 ( .A1(n17850), .A2(n17873), .ZN(n17857) );
  OAI22_X1 U19683 ( .A1(n17854), .A2(n17853), .B1(n17852), .B2(n17851), .ZN(
        n17855) );
  AOI21_X1 U19684 ( .B1(n17857), .B2(n17856), .A(n17855), .ZN(n17858) );
  OAI211_X1 U19685 ( .C1(n17860), .C2(n17877), .A(n17859), .B(n17858), .ZN(
        P2_U3008) );
  AOI22_X1 U19686 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19124), .B1(n17862), 
        .B2(n17861), .ZN(n17876) );
  OAI21_X1 U19687 ( .B1(n17865), .B2(n17864), .A(n17863), .ZN(n19303) );
  NAND2_X1 U19688 ( .A1(n17868), .A2(n17867), .ZN(n17869) );
  XNOR2_X1 U19689 ( .A(n17866), .B(n17869), .ZN(n19300) );
  AOI22_X1 U19690 ( .A1(n19300), .A2(n17871), .B1(n17870), .B2(n19297), .ZN(
        n17872) );
  OAI21_X1 U19691 ( .B1(n19303), .B2(n17873), .A(n17872), .ZN(n17874) );
  INV_X1 U19692 ( .A(n17874), .ZN(n17875) );
  OAI211_X1 U19693 ( .C1(n17878), .C2(n17877), .A(n17876), .B(n17875), .ZN(
        P2_U3006) );
  INV_X1 U19694 ( .A(n17901), .ZN(n17903) );
  INV_X1 U19695 ( .A(n17879), .ZN(n19013) );
  NAND3_X1 U19696 ( .A1(n17880), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n17881) );
  OAI21_X1 U19697 ( .B1(n19825), .B2(n19013), .A(n17881), .ZN(n17882) );
  AOI21_X1 U19698 ( .B1(n19987), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n17882), 
        .ZN(n17883) );
  OAI22_X1 U19699 ( .A1(n19987), .A2(n17901), .B1(n17903), .B2(n17883), .ZN(
        P2_U3605) );
  NAND2_X1 U19700 ( .A1(n19940), .A2(n17884), .ZN(n19959) );
  INV_X1 U19701 ( .A(n19959), .ZN(n17889) );
  NAND2_X1 U19702 ( .A1(n17885), .A2(n19992), .ZN(n17891) );
  NAND2_X1 U19703 ( .A1(n19311), .A2(n17891), .ZN(n17900) );
  INV_X1 U19704 ( .A(n17900), .ZN(n17887) );
  OAI22_X1 U19705 ( .A1(n19940), .A2(n17887), .B1(n17886), .B2(n19975), .ZN(
        n17888) );
  AOI21_X1 U19706 ( .B1(n19992), .B2(n17889), .A(n17888), .ZN(n17890) );
  AOI22_X1 U19707 ( .A1(n17903), .A2(n19871), .B1(n17890), .B2(n17901), .ZN(
        P2_U3603) );
  AOI21_X1 U19708 ( .B1(n19841), .B2(n17892), .A(n17891), .ZN(n17894) );
  OAI22_X1 U19709 ( .A1(n17892), .A2(n19311), .B1(n19026), .B2(n19975), .ZN(
        n17893) );
  NOR2_X1 U19710 ( .A1(n17894), .A2(n17893), .ZN(n17895) );
  AOI22_X1 U19711 ( .A1(n17903), .A2(n19985), .B1(n17895), .B2(n17901), .ZN(
        P2_U3604) );
  NOR2_X1 U19712 ( .A1(n17896), .A2(n19975), .ZN(n17899) );
  NAND2_X1 U19713 ( .A1(n19928), .A2(n19842), .ZN(n19910) );
  AOI211_X1 U19714 ( .C1(n19910), .C2(n19885), .A(n19841), .B(n15037), .ZN(
        n17898) );
  AOI211_X1 U19715 ( .C1(n19960), .C2(n17900), .A(n17899), .B(n17898), .ZN(
        n17902) );
  AOI22_X1 U19716 ( .A1(n17903), .A2(n19898), .B1(n17902), .B2(n17901), .ZN(
        P2_U3602) );
  NAND2_X1 U19717 ( .A1(n17904), .A2(n22311), .ZN(n17907) );
  OAI21_X1 U19718 ( .B1(n14423), .B2(n17053), .A(n17911), .ZN(n17905) );
  OAI21_X1 U19719 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17911), .A(n17905), 
        .ZN(n17906) );
  OAI221_X1 U19720 ( .B1(n17907), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17907), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17906), .ZN(P2_U2822) );
  INV_X1 U19721 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17910) );
  OAI221_X1 U19722 ( .B1(n17911), .B2(n17910), .C1(n17909), .C2(n17908), .A(
        n17907), .ZN(P2_U2823) );
  OAI22_X1 U19723 ( .A1(n22347), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17980), .ZN(n17912) );
  INV_X1 U19724 ( .A(n17912), .ZN(P2_U3611) );
  INV_X1 U19725 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17913) );
  AOI22_X1 U19726 ( .A1(n17980), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17913), 
        .B2(n22347), .ZN(P2_U3608) );
  AOI21_X1 U19727 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n22312), .ZN(n17914) );
  INV_X1 U19728 ( .A(n17914), .ZN(P2_U2815) );
  AOI22_X1 U19729 ( .A1(n17947), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17916) );
  OAI21_X1 U19730 ( .B1(n14081), .B2(n17949), .A(n17916), .ZN(P2_U2951) );
  INV_X1 U19731 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17918) );
  AOI22_X1 U19732 ( .A1(n17947), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17917) );
  OAI21_X1 U19733 ( .B1(n17918), .B2(n17949), .A(n17917), .ZN(P2_U2950) );
  INV_X1 U19734 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17920) );
  AOI22_X1 U19735 ( .A1(n17947), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17919) );
  OAI21_X1 U19736 ( .B1(n17920), .B2(n17949), .A(n17919), .ZN(P2_U2949) );
  INV_X1 U19737 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17922) );
  AOI22_X1 U19738 ( .A1(n17936), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17921) );
  OAI21_X1 U19739 ( .B1(n17922), .B2(n17949), .A(n17921), .ZN(P2_U2948) );
  INV_X1 U19740 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17924) );
  AOI22_X1 U19741 ( .A1(n17947), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17923) );
  OAI21_X1 U19742 ( .B1(n17924), .B2(n17949), .A(n17923), .ZN(P2_U2947) );
  INV_X1 U19743 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17926) );
  AOI22_X1 U19744 ( .A1(n17936), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17925) );
  OAI21_X1 U19745 ( .B1(n17926), .B2(n17949), .A(n17925), .ZN(P2_U2946) );
  AOI22_X1 U19746 ( .A1(n17936), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17927) );
  OAI21_X1 U19747 ( .B1(n17928), .B2(n17949), .A(n17927), .ZN(P2_U2945) );
  AOI22_X1 U19748 ( .A1(n17936), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17929) );
  OAI21_X1 U19749 ( .B1(n17930), .B2(n17949), .A(n17929), .ZN(P2_U2944) );
  AOI22_X1 U19750 ( .A1(n17936), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17931) );
  OAI21_X1 U19751 ( .B1(n17932), .B2(n17949), .A(n17931), .ZN(P2_U2943) );
  AOI22_X1 U19752 ( .A1(n17947), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17933) );
  OAI21_X1 U19753 ( .B1(n17934), .B2(n17949), .A(n17933), .ZN(P2_U2942) );
  AOI22_X1 U19754 ( .A1(n17936), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17937) );
  OAI21_X1 U19755 ( .B1(n17938), .B2(n17949), .A(n17937), .ZN(P2_U2941) );
  AOI22_X1 U19756 ( .A1(n17947), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17939) );
  OAI21_X1 U19757 ( .B1(n17940), .B2(n17949), .A(n17939), .ZN(P2_U2940) );
  AOI22_X1 U19758 ( .A1(n17947), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17941) );
  OAI21_X1 U19759 ( .B1(n17942), .B2(n17949), .A(n17941), .ZN(P2_U2939) );
  AOI22_X1 U19760 ( .A1(n17947), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17943) );
  OAI21_X1 U19761 ( .B1(n17944), .B2(n17949), .A(n17943), .ZN(P2_U2938) );
  AOI22_X1 U19762 ( .A1(n17947), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17945) );
  OAI21_X1 U19763 ( .B1(n17946), .B2(n17949), .A(n17945), .ZN(P2_U2937) );
  AOI22_X1 U19764 ( .A1(n17947), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17935), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17948) );
  OAI21_X1 U19765 ( .B1(n17950), .B2(n17949), .A(n17948), .ZN(P2_U2936) );
  INV_X1 U19766 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17951) );
  AOI22_X1 U19767 ( .A1(n17980), .A2(n17951), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n22347), .ZN(n17952) );
  OAI21_X1 U19768 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n22346), .A(n17952), 
        .ZN(P2_U2817) );
  NAND2_X1 U19769 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17980), .ZN(n17975) );
  OAI222_X1 U19770 ( .A1(n17975), .A2(n17053), .B1(n17953), .B2(n17980), .C1(
        n12060), .C2(n17977), .ZN(P2_U3212) );
  INV_X1 U19771 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17954) );
  OAI222_X1 U19772 ( .A1(n17977), .A2(n15268), .B1(n17954), .B2(n17980), .C1(
        n12060), .C2(n22351), .ZN(P2_U3213) );
  INV_X1 U19773 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n17955) );
  OAI222_X1 U19774 ( .A1(n17977), .A2(n14069), .B1(n17955), .B2(n17980), .C1(
        n15268), .C2(n22351), .ZN(P2_U3214) );
  INV_X1 U19775 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n17956) );
  OAI222_X1 U19776 ( .A1(n17977), .A2(n14106), .B1(n17956), .B2(n17980), .C1(
        n14069), .C2(n22351), .ZN(P2_U3215) );
  INV_X1 U19777 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n17957) );
  OAI222_X1 U19778 ( .A1(n17977), .A2(n19046), .B1(n17957), .B2(n17980), .C1(
        n14106), .C2(n22351), .ZN(P2_U3216) );
  INV_X1 U19779 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n17958) );
  OAI222_X1 U19780 ( .A1(n17977), .A2(n17044), .B1(n17958), .B2(n17980), .C1(
        n19046), .C2(n22351), .ZN(P2_U3217) );
  INV_X1 U19781 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n17959) );
  OAI222_X1 U19782 ( .A1(n17977), .A2(n14116), .B1(n17959), .B2(n17980), .C1(
        n17044), .C2(n22351), .ZN(P2_U3218) );
  INV_X1 U19783 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n17960) );
  OAI222_X1 U19784 ( .A1(n17977), .A2(n17961), .B1(n17960), .B2(n17980), .C1(
        n14116), .C2(n22351), .ZN(P2_U3219) );
  INV_X1 U19785 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20417) );
  OAI222_X1 U19786 ( .A1(n22351), .A2(n17961), .B1(n20417), .B2(n17980), .C1(
        n17962), .C2(n17977), .ZN(P2_U3220) );
  INV_X1 U19787 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20419) );
  OAI222_X1 U19788 ( .A1(n22351), .A2(n17962), .B1(n20419), .B2(n17980), .C1(
        n12472), .C2(n17977), .ZN(P2_U3221) );
  INV_X1 U19789 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20421) );
  OAI222_X1 U19790 ( .A1(n22351), .A2(n12472), .B1(n20421), .B2(n17980), .C1(
        n17963), .C2(n17977), .ZN(P2_U3222) );
  INV_X1 U19791 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20423) );
  OAI222_X1 U19792 ( .A1(n22351), .A2(n17963), .B1(n20423), .B2(n17980), .C1(
        n19084), .C2(n17977), .ZN(P2_U3223) );
  INV_X1 U19793 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20425) );
  OAI222_X1 U19794 ( .A1(n22351), .A2(n19084), .B1(n20425), .B2(n17980), .C1(
        n17964), .C2(n17977), .ZN(P2_U3224) );
  INV_X1 U19795 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20427) );
  OAI222_X1 U19796 ( .A1(n17975), .A2(n17964), .B1(n20427), .B2(n17980), .C1(
        n17965), .C2(n17977), .ZN(P2_U3225) );
  INV_X1 U19797 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20429) );
  OAI222_X1 U19798 ( .A1(n17975), .A2(n17965), .B1(n20429), .B2(n17980), .C1(
        n17966), .C2(n17977), .ZN(P2_U3226) );
  INV_X1 U19799 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20431) );
  OAI222_X1 U19800 ( .A1(n17975), .A2(n17966), .B1(n20431), .B2(n17980), .C1(
        n17967), .C2(n17977), .ZN(P2_U3227) );
  INV_X1 U19801 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20433) );
  OAI222_X1 U19802 ( .A1(n17975), .A2(n17967), .B1(n20433), .B2(n17980), .C1(
        n17968), .C2(n17977), .ZN(P2_U3228) );
  INV_X1 U19803 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20435) );
  OAI222_X1 U19804 ( .A1(n17977), .A2(n17969), .B1(n20435), .B2(n17980), .C1(
        n17968), .C2(n22351), .ZN(P2_U3229) );
  INV_X1 U19805 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20437) );
  OAI222_X1 U19806 ( .A1(n17975), .A2(n17969), .B1(n20437), .B2(n17980), .C1(
        n17970), .C2(n17977), .ZN(P2_U3230) );
  INV_X1 U19807 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20439) );
  OAI222_X1 U19808 ( .A1(n17977), .A2(n16901), .B1(n20439), .B2(n17980), .C1(
        n17970), .C2(n22351), .ZN(P2_U3231) );
  INV_X1 U19809 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20441) );
  OAI222_X1 U19810 ( .A1(n17977), .A2(n16882), .B1(n20441), .B2(n17980), .C1(
        n16901), .C2(n22351), .ZN(P2_U3232) );
  INV_X1 U19811 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20443) );
  OAI222_X1 U19812 ( .A1(n17977), .A2(n17971), .B1(n20443), .B2(n17980), .C1(
        n16882), .C2(n22351), .ZN(P2_U3233) );
  INV_X1 U19813 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20445) );
  OAI222_X1 U19814 ( .A1(n17977), .A2(n16862), .B1(n20445), .B2(n17980), .C1(
        n17971), .C2(n22351), .ZN(P2_U3234) );
  INV_X1 U19815 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20447) );
  OAI222_X1 U19816 ( .A1(n17977), .A2(n17972), .B1(n20447), .B2(n17980), .C1(
        n16862), .C2(n22351), .ZN(P2_U3235) );
  INV_X1 U19817 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20449) );
  OAI222_X1 U19818 ( .A1(n17975), .A2(n17972), .B1(n20449), .B2(n17980), .C1(
        n17973), .C2(n17977), .ZN(P2_U3236) );
  INV_X1 U19819 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20451) );
  OAI222_X1 U19820 ( .A1(n17977), .A2(n19207), .B1(n20451), .B2(n17980), .C1(
        n17973), .C2(n22351), .ZN(P2_U3237) );
  INV_X1 U19821 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20453) );
  OAI222_X1 U19822 ( .A1(n17975), .A2(n19207), .B1(n20453), .B2(n17980), .C1(
        n14159), .C2(n17977), .ZN(P2_U3238) );
  INV_X1 U19823 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20455) );
  OAI222_X1 U19824 ( .A1(n17975), .A2(n14159), .B1(n20455), .B2(n17980), .C1(
        n17974), .C2(n17977), .ZN(P2_U3239) );
  INV_X1 U19825 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20458) );
  OAI222_X1 U19826 ( .A1(n17975), .A2(n17974), .B1(n20458), .B2(n17980), .C1(
        n17976), .C2(n17977), .ZN(P2_U3240) );
  INV_X1 U19827 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20461) );
  OAI222_X1 U19828 ( .A1(n17977), .A2(n19255), .B1(n20461), .B2(n17980), .C1(
        n17976), .C2(n22351), .ZN(P2_U3241) );
  OAI22_X1 U19829 ( .A1(n22347), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17980), .ZN(n17978) );
  INV_X1 U19830 ( .A(n17978), .ZN(P2_U3588) );
  OAI22_X1 U19831 ( .A1(n22347), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17980), .ZN(n17979) );
  INV_X1 U19832 ( .A(n17979), .ZN(P2_U3587) );
  MUX2_X1 U19833 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n22347), .Z(P2_U3586) );
  OAI22_X1 U19834 ( .A1(n22347), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17980), .ZN(n17981) );
  INV_X1 U19835 ( .A(n17981), .ZN(P2_U3585) );
  INV_X1 U19836 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20796) );
  NOR3_X1 U19837 ( .A1(n17983), .A2(n21294), .A3(n17982), .ZN(n17984) );
  NOR2_X1 U19838 ( .A1(n21294), .A2(n18348), .ZN(n18351) );
  NAND4_X1 U19839 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .A4(n18351), .ZN(n17987) );
  NAND2_X1 U19840 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17989), .ZN(n18003) );
  INV_X1 U19841 ( .A(n18003), .ZN(n18012) );
  INV_X2 U19842 ( .A(n18352), .ZN(n18350) );
  AOI21_X1 U19843 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n18315), .A(n17989), .ZN(
        n17986) );
  INV_X1 U19844 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19569) );
  OAI22_X1 U19845 ( .A1(n18012), .A2(n17986), .B1(n19569), .B2(n18350), .ZN(
        P3_U2699) );
  INV_X1 U19846 ( .A(n17987), .ZN(n17991) );
  AOI21_X1 U19847 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n18315), .A(n17991), .ZN(
        n17988) );
  INV_X1 U19848 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19612) );
  OAI22_X1 U19849 ( .A1(n17989), .A2(n17988), .B1(n19612), .B2(n18350), .ZN(
        P3_U2700) );
  INV_X1 U19850 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18354) );
  INV_X1 U19851 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20771) );
  NOR2_X1 U19852 ( .A1(n18354), .A2(n20771), .ZN(n17990) );
  AOI21_X1 U19853 ( .B1(n17990), .B2(n18355), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17992) );
  INV_X1 U19854 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19655) );
  AOI221_X1 U19855 ( .B1(n17992), .B2(n18350), .C1(n19655), .C2(n18352), .A(
        n17991), .ZN(P3_U2701) );
  AOI22_X1 U19856 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17996) );
  AOI22_X1 U19857 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17995) );
  AOI22_X1 U19858 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17994) );
  AOI22_X1 U19859 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17993) );
  NAND4_X1 U19860 ( .A1(n17996), .A2(n17995), .A3(n17994), .A4(n17993), .ZN(
        n18002) );
  AOI22_X1 U19861 ( .A1(n18390), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18000) );
  AOI22_X1 U19862 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17999) );
  AOI22_X1 U19863 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17998) );
  AOI22_X1 U19864 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17997) );
  NAND4_X1 U19865 ( .A1(n18000), .A2(n17999), .A3(n17998), .A4(n17997), .ZN(
        n18001) );
  NOR2_X1 U19866 ( .A1(n18002), .A2(n18001), .ZN(n21366) );
  INV_X1 U19867 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20847) );
  NAND2_X1 U19868 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18014), .ZN(n18008) );
  NOR2_X1 U19869 ( .A1(n20847), .A2(n18008), .ZN(n18084) );
  NAND3_X1 U19870 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n18005) );
  NAND4_X1 U19871 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n18004) );
  NOR3_X1 U19872 ( .A1(n20796), .A2(n18005), .A3(n18004), .ZN(n18015) );
  NAND2_X1 U19873 ( .A1(n18355), .A2(n18015), .ZN(n18042) );
  INV_X1 U19874 ( .A(n18042), .ZN(n18112) );
  OAI21_X1 U19875 ( .B1(n18352), .B2(n18112), .A(P3_EBX_REG_8__SCAN_IN), .ZN(
        n18006) );
  OAI21_X1 U19876 ( .B1(n18084), .B2(P3_EBX_REG_8__SCAN_IN), .A(n18006), .ZN(
        n18007) );
  OAI21_X1 U19877 ( .B1(n21366), .B2(n18350), .A(n18007), .ZN(P3_U2695) );
  INV_X1 U19878 ( .A(n18008), .ZN(n18011) );
  AOI21_X1 U19879 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n18315), .A(n18011), .ZN(
        n18009) );
  OAI22_X1 U19880 ( .A1(n18112), .A2(n18009), .B1(n19447), .B2(n18350), .ZN(
        P3_U2696) );
  AOI21_X1 U19881 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18315), .A(n18014), .ZN(
        n18010) );
  INV_X1 U19882 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19488) );
  OAI22_X1 U19883 ( .A1(n18011), .A2(n18010), .B1(n19488), .B2(n18350), .ZN(
        P3_U2697) );
  AOI21_X1 U19884 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18315), .A(n18012), .ZN(
        n18013) );
  INV_X1 U19885 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19529) );
  OAI22_X1 U19886 ( .A1(n18014), .A2(n18013), .B1(n19529), .B2(n18350), .ZN(
        P3_U2698) );
  NAND4_X1 U19887 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n18043) );
  NAND3_X1 U19888 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .ZN(n18058) );
  NOR2_X1 U19889 ( .A1(n18043), .A2(n18058), .ZN(n18037) );
  AND3_X1 U19890 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18015), .A3(n18037), .ZN(
        n18126) );
  NAND2_X1 U19891 ( .A1(n18351), .A2(n18126), .ZN(n18038) );
  AOI22_X1 U19892 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18019) );
  AOI22_X1 U19893 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18018) );
  AOI22_X1 U19894 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18017) );
  AOI22_X1 U19895 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18016) );
  NAND4_X1 U19896 ( .A1(n18019), .A2(n18018), .A3(n18017), .A4(n18016), .ZN(
        n18025) );
  AOI22_X1 U19897 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U19898 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U19899 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U19900 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18020) );
  NAND4_X1 U19901 ( .A1(n18023), .A2(n18022), .A3(n18021), .A4(n18020), .ZN(
        n18024) );
  NOR2_X1 U19902 ( .A1(n18025), .A2(n18024), .ZN(n21348) );
  NAND3_X1 U19903 ( .A1(n18038), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n18350), 
        .ZN(n18026) );
  OAI221_X1 U19904 ( .B1(n18038), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n18315), 
        .C2(n21348), .A(n18026), .ZN(P3_U2687) );
  AOI22_X1 U19905 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18036) );
  AOI22_X1 U19906 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18035) );
  AOI22_X1 U19907 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18027) );
  OAI21_X1 U19908 ( .B1(n18086), .B2(n19447), .A(n18027), .ZN(n18033) );
  AOI22_X1 U19909 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18031) );
  AOI22_X1 U19910 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18030) );
  AOI22_X1 U19911 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18029) );
  AOI22_X1 U19912 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18028) );
  NAND4_X1 U19913 ( .A1(n18031), .A2(n18030), .A3(n18029), .A4(n18028), .ZN(
        n18032) );
  AOI211_X1 U19914 ( .C1(n18456), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n18033), .B(n18032), .ZN(n18034) );
  NAND3_X1 U19915 ( .A1(n18036), .A2(n18035), .A3(n18034), .ZN(n21357) );
  INV_X1 U19916 ( .A(n21357), .ZN(n18041) );
  AOI21_X1 U19917 ( .B1(n18112), .B2(n18037), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n18040) );
  NAND2_X1 U19918 ( .A1(n18315), .A2(n18038), .ZN(n18039) );
  OAI22_X1 U19919 ( .A1(n18041), .A2(n18350), .B1(n18040), .B2(n18039), .ZN(
        P3_U2688) );
  NOR2_X1 U19920 ( .A1(n18043), .A2(n18042), .ZN(n18099) );
  NAND2_X1 U19921 ( .A1(n21267), .A2(n18099), .ZN(n18057) );
  INV_X1 U19922 ( .A(n18057), .ZN(n18083) );
  AND3_X1 U19923 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n18083), .ZN(n18056) );
  AOI22_X1 U19924 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18350), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(n18083), .ZN(n18055) );
  AOI22_X1 U19925 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18053) );
  AOI22_X1 U19926 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18052) );
  AOI22_X1 U19927 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18044) );
  OAI21_X1 U19928 ( .B1(n18086), .B2(n19529), .A(n18044), .ZN(n18050) );
  AOI22_X1 U19929 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18048) );
  AOI22_X1 U19930 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18047) );
  AOI22_X1 U19931 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18046) );
  AOI22_X1 U19932 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18045) );
  NAND4_X1 U19933 ( .A1(n18048), .A2(n18047), .A3(n18046), .A4(n18045), .ZN(
        n18049) );
  AOI211_X1 U19934 ( .C1(n18181), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n18050), .B(n18049), .ZN(n18051) );
  NAND3_X1 U19935 ( .A1(n18053), .A2(n18052), .A3(n18051), .ZN(n21198) );
  INV_X1 U19936 ( .A(n21198), .ZN(n18054) );
  OAI22_X1 U19937 ( .A1(n18056), .A2(n18055), .B1(n18054), .B2(n18350), .ZN(
        P3_U2690) );
  AOI21_X1 U19938 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18315), .A(n18056), .ZN(
        n18071) );
  NOR2_X1 U19939 ( .A1(n18058), .A2(n18057), .ZN(n18070) );
  AOI22_X1 U19940 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18068) );
  AOI22_X1 U19941 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11152), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18067) );
  AOI22_X1 U19942 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18317), .B1(
        P3_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n20804), .ZN(n18059) );
  OAI21_X1 U19943 ( .B1(n19488), .B2(n18086), .A(n18059), .ZN(n18065) );
  AOI22_X1 U19944 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18063) );
  AOI22_X1 U19945 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n18462), .ZN(n18062) );
  AOI22_X1 U19946 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11128), .B1(
        P3_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n18434), .ZN(n18061) );
  AOI22_X1 U19947 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18421), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n18455), .ZN(n18060) );
  NAND4_X1 U19948 ( .A1(n18063), .A2(n18062), .A3(n18061), .A4(n18060), .ZN(
        n18064) );
  AOI211_X1 U19949 ( .C1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .C2(n18409), .A(
        n18065), .B(n18064), .ZN(n18066) );
  NAND3_X1 U19950 ( .A1(n18068), .A2(n18067), .A3(n18066), .ZN(n21351) );
  INV_X1 U19951 ( .A(n21351), .ZN(n18069) );
  OAI22_X1 U19952 ( .A1(n18071), .A2(n18070), .B1(n18069), .B2(n18315), .ZN(
        P3_U2689) );
  AOI22_X1 U19953 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U19954 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U19955 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U19956 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18072) );
  NAND4_X1 U19957 ( .A1(n18075), .A2(n18074), .A3(n18073), .A4(n18072), .ZN(
        n18081) );
  AOI22_X1 U19958 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18079) );
  AOI22_X1 U19959 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18078) );
  AOI22_X1 U19960 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18077) );
  AOI22_X1 U19961 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18076) );
  NAND4_X1 U19962 ( .A1(n18079), .A2(n18078), .A3(n18077), .A4(n18076), .ZN(
        n18080) );
  NOR2_X1 U19963 ( .A1(n18081), .A2(n18080), .ZN(n21203) );
  NOR3_X1 U19964 ( .A1(n18352), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n18083), .ZN(
        n18082) );
  AOI221_X1 U19965 ( .B1(n21203), .B2(n18352), .C1(n18083), .C2(
        P3_EBX_REG_12__SCAN_IN), .A(n18082), .ZN(P3_U2691) );
  AND3_X1 U19966 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n18084), .ZN(n18124) );
  AOI21_X1 U19967 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18315), .A(n18111), .ZN(
        n18098) );
  AOI22_X1 U19968 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U19969 ( .A1(n18434), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U19970 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18085) );
  OAI21_X1 U19971 ( .B1(n18086), .B2(n19612), .A(n18085), .ZN(n18093) );
  AOI22_X1 U19972 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18091) );
  AOI22_X1 U19973 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18090) );
  AOI22_X1 U19974 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18089) );
  AOI22_X1 U19975 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18088) );
  NAND4_X1 U19976 ( .A1(n18091), .A2(n18090), .A3(n18089), .A4(n18088), .ZN(
        n18092) );
  AOI211_X1 U19977 ( .C1(n18181), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n18093), .B(n18092), .ZN(n18094) );
  NAND3_X1 U19978 ( .A1(n18096), .A2(n18095), .A3(n18094), .ZN(n21206) );
  INV_X1 U19979 ( .A(n21206), .ZN(n18097) );
  OAI22_X1 U19980 ( .A1(n18099), .A2(n18098), .B1(n18097), .B2(n18350), .ZN(
        P3_U2692) );
  AOI21_X1 U19981 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18315), .A(n18124), .ZN(
        n18110) );
  AOI22_X1 U19982 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18103) );
  AOI22_X1 U19983 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18102) );
  AOI22_X1 U19984 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U19985 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18100) );
  NAND4_X1 U19986 ( .A1(n18103), .A2(n18102), .A3(n18101), .A4(n18100), .ZN(
        n18109) );
  AOI22_X1 U19987 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18107) );
  AOI22_X1 U19988 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18106) );
  AOI22_X1 U19989 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U19990 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18104) );
  NAND4_X1 U19991 ( .A1(n18107), .A2(n18106), .A3(n18105), .A4(n18104), .ZN(
        n18108) );
  NOR2_X1 U19992 ( .A1(n18109), .A2(n18108), .ZN(n21209) );
  OAI22_X1 U19993 ( .A1(n18111), .A2(n18110), .B1(n21209), .B2(n18315), .ZN(
        P3_U2693) );
  OAI221_X1 U19994 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(P3_EBX_REG_8__SCAN_IN), 
        .C1(P3_EBX_REG_9__SCAN_IN), .C2(n18112), .A(n18315), .ZN(n18123) );
  AOI22_X1 U19995 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18116) );
  AOI22_X1 U19996 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U19997 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U19998 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18113) );
  NAND4_X1 U19999 ( .A1(n18116), .A2(n18115), .A3(n18114), .A4(n18113), .ZN(
        n18122) );
  AOI22_X1 U20000 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18120) );
  AOI22_X1 U20001 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18119) );
  AOI22_X1 U20002 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18118) );
  AOI22_X1 U20003 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18117) );
  NAND4_X1 U20004 ( .A1(n18120), .A2(n18119), .A3(n18118), .A4(n18117), .ZN(
        n18121) );
  NOR2_X1 U20005 ( .A1(n18122), .A2(n18121), .ZN(n21215) );
  OAI22_X1 U20006 ( .A1(n18124), .A2(n18123), .B1(n21215), .B2(n18350), .ZN(
        P3_U2694) );
  INV_X1 U20007 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21144) );
  INV_X1 U20008 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n21104) );
  INV_X1 U20009 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n21093) );
  INV_X1 U20010 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n21044) );
  NOR3_X1 U20011 ( .A1(n21104), .A2(n21093), .A3(n21044), .ZN(n18125) );
  NAND4_X1 U20012 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n18125), .ZN(n18238) );
  NAND2_X1 U20013 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18127) );
  INV_X1 U20014 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n18314) );
  INV_X1 U20015 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20990) );
  NAND2_X1 U20016 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18126), .ZN(n18344) );
  NOR2_X1 U20017 ( .A1(n20990), .A2(n18344), .ZN(n18343) );
  NAND2_X1 U20018 ( .A1(n18355), .A2(n18343), .ZN(n18313) );
  NAND3_X1 U20019 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(P3_EBX_REG_19__SCAN_IN), 
        .A3(n18329), .ZN(n18226) );
  NOR4_X1 U20020 ( .A1(n21144), .A2(n18238), .A3(n18127), .A4(n18226), .ZN(
        n18224) );
  NAND2_X1 U20021 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n18224), .ZN(n18223) );
  INV_X1 U20022 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n21167) );
  INV_X1 U20023 ( .A(n18223), .ZN(n18128) );
  OAI33_X1 U20024 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18223), .A3(n21294), 
        .B1(n21167), .B2(n18352), .B3(n18128), .ZN(P3_U2672) );
  AOI22_X1 U20025 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18421), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18132) );
  AOI22_X1 U20026 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n20804), .ZN(n18131) );
  AOI22_X1 U20027 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18453), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U20028 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__6__SCAN_IN), .B2(n18455), .ZN(n18129) );
  NAND4_X1 U20029 ( .A1(n18132), .A2(n18131), .A3(n18130), .A4(n18129), .ZN(
        n18138) );
  AOI22_X1 U20030 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18136) );
  AOI22_X1 U20031 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11128), .B1(
        P3_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n18461), .ZN(n18135) );
  AOI22_X1 U20032 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18134) );
  AOI22_X1 U20033 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n18434), .ZN(n18133) );
  NAND4_X1 U20034 ( .A1(n18136), .A2(n18135), .A3(n18134), .A4(n18133), .ZN(
        n18137) );
  NOR2_X1 U20035 ( .A1(n18138), .A2(n18137), .ZN(n18244) );
  AOI22_X1 U20036 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18142) );
  AOI22_X1 U20037 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18141) );
  AOI22_X1 U20038 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U20039 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18139) );
  NAND4_X1 U20040 ( .A1(n18142), .A2(n18141), .A3(n18140), .A4(n18139), .ZN(
        n18148) );
  AOI22_X1 U20041 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18146) );
  AOI22_X1 U20042 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18145) );
  AOI22_X1 U20043 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18144) );
  AOI22_X1 U20044 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18143) );
  NAND4_X1 U20045 ( .A1(n18146), .A2(n18145), .A3(n18144), .A4(n18143), .ZN(
        n18147) );
  NOR2_X1 U20046 ( .A1(n18148), .A2(n18147), .ZN(n18239) );
  AOI22_X1 U20047 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18152) );
  AOI22_X1 U20048 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18151) );
  AOI22_X1 U20049 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18150) );
  AOI22_X1 U20050 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18149) );
  NAND4_X1 U20051 ( .A1(n18152), .A2(n18151), .A3(n18150), .A4(n18149), .ZN(
        n18159) );
  AOI22_X1 U20052 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U20053 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U20054 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U20055 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18154) );
  NAND4_X1 U20056 ( .A1(n18157), .A2(n18156), .A3(n18155), .A4(n18154), .ZN(
        n18158) );
  NOR2_X1 U20057 ( .A1(n18159), .A2(n18158), .ZN(n18261) );
  AOI22_X1 U20058 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18163) );
  AOI22_X1 U20059 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18162) );
  AOI22_X1 U20060 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18161) );
  AOI22_X1 U20061 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18160) );
  NAND4_X1 U20062 ( .A1(n18163), .A2(n18162), .A3(n18161), .A4(n18160), .ZN(
        n18169) );
  AOI22_X1 U20063 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18167) );
  AOI22_X1 U20064 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18166) );
  AOI22_X1 U20065 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18165) );
  AOI22_X1 U20066 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18164) );
  NAND4_X1 U20067 ( .A1(n18167), .A2(n18166), .A3(n18165), .A4(n18164), .ZN(
        n18168) );
  NOR2_X1 U20068 ( .A1(n18169), .A2(n18168), .ZN(n18271) );
  AOI22_X1 U20069 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U20070 ( .A1(n18462), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U20071 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18171) );
  AOI22_X1 U20072 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18170) );
  NAND4_X1 U20073 ( .A1(n18173), .A2(n18172), .A3(n18171), .A4(n18170), .ZN(
        n18179) );
  AOI22_X1 U20074 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U20075 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U20076 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18175) );
  AOI22_X1 U20077 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18379), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18174) );
  NAND4_X1 U20078 ( .A1(n18177), .A2(n18176), .A3(n18175), .A4(n18174), .ZN(
        n18178) );
  NOR2_X1 U20079 ( .A1(n18179), .A2(n18178), .ZN(n18272) );
  NOR2_X1 U20080 ( .A1(n18271), .A2(n18272), .ZN(n18270) );
  AOI22_X1 U20081 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U20082 ( .A1(n18434), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18189) );
  AOI22_X1 U20083 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n15716), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18180) );
  OAI21_X1 U20084 ( .B1(n18202), .B2(n19698), .A(n18180), .ZN(n18187) );
  AOI22_X1 U20085 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U20086 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18184) );
  AOI22_X1 U20087 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18181), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18183) );
  AOI22_X1 U20088 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18182) );
  NAND4_X1 U20089 ( .A1(n18185), .A2(n18184), .A3(n18183), .A4(n18182), .ZN(
        n18186) );
  AOI211_X1 U20090 ( .C1(n18414), .C2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n18187), .B(n18186), .ZN(n18188) );
  NAND3_X1 U20091 ( .A1(n18190), .A2(n18189), .A3(n18188), .ZN(n18266) );
  NAND2_X1 U20092 ( .A1(n18270), .A2(n18266), .ZN(n18265) );
  NOR2_X1 U20093 ( .A1(n18261), .A2(n18265), .ZN(n18260) );
  AOI22_X1 U20094 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18200) );
  AOI22_X1 U20095 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U20096 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18191) );
  OAI21_X1 U20097 ( .B1(n18202), .B2(n19612), .A(n18191), .ZN(n18197) );
  AOI22_X1 U20098 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18195) );
  AOI22_X1 U20099 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18194) );
  AOI22_X1 U20100 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18193) );
  AOI22_X1 U20101 ( .A1(n15725), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18192) );
  NAND4_X1 U20102 ( .A1(n18195), .A2(n18194), .A3(n18193), .A4(n18192), .ZN(
        n18196) );
  AOI211_X1 U20103 ( .C1(n18390), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18197), .B(n18196), .ZN(n18198) );
  NAND3_X1 U20104 ( .A1(n18200), .A2(n18199), .A3(n18198), .ZN(n18254) );
  NAND2_X1 U20105 ( .A1(n18260), .A2(n18254), .ZN(n18253) );
  NOR2_X1 U20106 ( .A1(n18239), .A2(n18253), .ZN(n18250) );
  AOI22_X1 U20107 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U20108 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18210) );
  AOI22_X1 U20109 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18201) );
  OAI21_X1 U20110 ( .B1(n18202), .B2(n19529), .A(n18201), .ZN(n18208) );
  AOI22_X1 U20111 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18206) );
  AOI22_X1 U20112 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18205) );
  AOI22_X1 U20113 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n18204) );
  AOI22_X1 U20114 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18203) );
  NAND4_X1 U20115 ( .A1(n18206), .A2(n18205), .A3(n18204), .A4(n18203), .ZN(
        n18207) );
  AOI211_X1 U20116 ( .C1(n18379), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n18208), .B(n18207), .ZN(n18209) );
  NAND3_X1 U20117 ( .A1(n18211), .A2(n18210), .A3(n18209), .ZN(n18249) );
  NAND2_X1 U20118 ( .A1(n18250), .A2(n18249), .ZN(n18248) );
  NOR2_X1 U20119 ( .A1(n18244), .A2(n18248), .ZN(n18243) );
  AOI22_X1 U20120 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U20121 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U20122 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18213) );
  AOI22_X1 U20123 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18212) );
  NAND4_X1 U20124 ( .A1(n18215), .A2(n18214), .A3(n18213), .A4(n18212), .ZN(
        n18221) );
  AOI22_X1 U20125 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18219) );
  AOI22_X1 U20126 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U20127 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18217) );
  AOI22_X1 U20128 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18216) );
  NAND4_X1 U20129 ( .A1(n18219), .A2(n18218), .A3(n18217), .A4(n18216), .ZN(
        n18220) );
  NOR2_X1 U20130 ( .A1(n18221), .A2(n18220), .ZN(n18222) );
  XOR2_X1 U20131 ( .A(n18243), .B(n18222), .Z(n21310) );
  OAI211_X1 U20132 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n18224), .A(n18223), .B(
        n18350), .ZN(n18225) );
  OAI21_X1 U20133 ( .B1(n21310), .B2(n18350), .A(n18225), .ZN(P3_U2673) );
  INV_X1 U20134 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n21014) );
  NAND2_X1 U20135 ( .A1(n21267), .A2(n18329), .ZN(n18328) );
  NOR2_X1 U20136 ( .A1(n21014), .A2(n18328), .ZN(n18300) );
  NAND2_X1 U20137 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18300), .ZN(n18256) );
  NAND2_X1 U20138 ( .A1(n18315), .A2(n18226), .ZN(n18301) );
  AOI22_X1 U20139 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n18230) );
  AOI22_X1 U20140 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18229) );
  AOI22_X1 U20141 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18228) );
  AOI22_X1 U20142 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n18227) );
  NAND4_X1 U20143 ( .A1(n18230), .A2(n18229), .A3(n18228), .A4(n18227), .ZN(
        n18236) );
  AOI22_X1 U20144 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18234) );
  AOI22_X1 U20145 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18233) );
  AOI22_X1 U20146 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U20147 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n18231) );
  NAND4_X1 U20148 ( .A1(n18234), .A2(n18233), .A3(n18232), .A4(n18231), .ZN(
        n18235) );
  NOR2_X1 U20149 ( .A1(n18236), .A2(n18235), .ZN(n21257) );
  OR2_X1 U20150 ( .A1(n21257), .A2(n18315), .ZN(n18237) );
  OAI221_X1 U20151 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18256), .C1(n21044), 
        .C2(n18301), .A(n18237), .ZN(P3_U2682) );
  NOR2_X1 U20152 ( .A1(n18256), .A2(n18238), .ZN(n18255) );
  INV_X1 U20153 ( .A(n18255), .ZN(n18242) );
  AOI21_X1 U20154 ( .B1(n18239), .B2(n18253), .A(n18250), .ZN(n21324) );
  INV_X1 U20155 ( .A(n21324), .ZN(n18241) );
  NAND3_X1 U20156 ( .A1(n18242), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18315), 
        .ZN(n18240) );
  OAI221_X1 U20157 ( .B1(n18242), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18315), 
        .C2(n18241), .A(n18240), .ZN(P3_U2676) );
  NAND3_X1 U20158 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n18255), .ZN(n18247) );
  AOI21_X1 U20159 ( .B1(n18244), .B2(n18248), .A(n18243), .ZN(n21316) );
  INV_X1 U20160 ( .A(n21316), .ZN(n18246) );
  NAND3_X1 U20161 ( .A1(n18247), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18350), 
        .ZN(n18245) );
  OAI221_X1 U20162 ( .B1(n18247), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18315), 
        .C2(n18246), .A(n18245), .ZN(P3_U2674) );
  INV_X1 U20163 ( .A(n18247), .ZN(n18252) );
  AOI22_X1 U20164 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18350), .B1(
        P3_EBX_REG_27__SCAN_IN), .B2(n18255), .ZN(n18251) );
  OAI21_X1 U20165 ( .B1(n18250), .B2(n18249), .A(n18248), .ZN(n21323) );
  OAI22_X1 U20166 ( .A1(n18252), .A2(n18251), .B1(n21323), .B2(n18350), .ZN(
        P3_U2675) );
  OAI21_X1 U20167 ( .B1(n18260), .B2(n18254), .A(n18253), .ZN(n21304) );
  NOR2_X1 U20168 ( .A1(n18255), .A2(n21104), .ZN(n18257) );
  INV_X1 U20169 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n21066) );
  NOR2_X1 U20170 ( .A1(n21044), .A2(n18256), .ZN(n18276) );
  NAND2_X1 U20171 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n18276), .ZN(n18269) );
  NOR2_X1 U20172 ( .A1(n21066), .A2(n18269), .ZN(n18275) );
  NAND2_X1 U20173 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n18275), .ZN(n18259) );
  NOR2_X1 U20174 ( .A1(n21093), .A2(n18259), .ZN(n18264) );
  AOI22_X1 U20175 ( .A1(n18257), .A2(n18350), .B1(n18264), .B2(n21104), .ZN(
        n18258) );
  OAI21_X1 U20176 ( .B1(n21304), .B2(n18350), .A(n18258), .ZN(P3_U2677) );
  INV_X1 U20177 ( .A(n18259), .ZN(n18268) );
  AOI21_X1 U20178 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18350), .A(n18268), .ZN(
        n18263) );
  AOI21_X1 U20179 ( .B1(n18261), .B2(n18265), .A(n18260), .ZN(n21290) );
  INV_X1 U20180 ( .A(n21290), .ZN(n18262) );
  OAI22_X1 U20181 ( .A1(n18264), .A2(n18263), .B1(n18262), .B2(n18350), .ZN(
        P3_U2678) );
  AOI21_X1 U20182 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18315), .A(n18275), .ZN(
        n18267) );
  OAI21_X1 U20183 ( .B1(n18270), .B2(n18266), .A(n18265), .ZN(n21334) );
  OAI22_X1 U20184 ( .A1(n18268), .A2(n18267), .B1(n21334), .B2(n18350), .ZN(
        P3_U2679) );
  INV_X1 U20185 ( .A(n18269), .ZN(n18289) );
  AOI21_X1 U20186 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18315), .A(n18289), .ZN(
        n18274) );
  AOI21_X1 U20187 ( .B1(n18272), .B2(n18271), .A(n18270), .ZN(n21335) );
  INV_X1 U20188 ( .A(n21335), .ZN(n18273) );
  OAI22_X1 U20189 ( .A1(n18275), .A2(n18274), .B1(n18273), .B2(n18315), .ZN(
        P3_U2680) );
  AOI21_X1 U20190 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18315), .A(n18276), .ZN(
        n18288) );
  AOI22_X1 U20191 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n11152), .B1(
        n18379), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18286) );
  AOI22_X1 U20192 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__6__SCAN_IN), .B2(n18434), .ZN(n18285) );
  AOI22_X1 U20193 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18277) );
  OAI21_X1 U20194 ( .B1(n11190), .B2(n19488), .A(n18277), .ZN(n18283) );
  AOI22_X1 U20195 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18421), .B1(
        P3_INSTQUEUE_REG_4__6__SCAN_IN), .B2(n11149), .ZN(n18281) );
  AOI22_X1 U20196 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18462), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n18455), .ZN(n18280) );
  AOI22_X1 U20197 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n11127), .ZN(n18279) );
  AOI22_X1 U20198 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18453), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n20804), .ZN(n18278) );
  NAND4_X1 U20199 ( .A1(n18281), .A2(n18280), .A3(n18279), .A4(n18278), .ZN(
        n18282) );
  AOI211_X1 U20200 ( .C1(n11130), .C2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n18283), .B(n18282), .ZN(n18284) );
  NAND3_X1 U20201 ( .A1(n18286), .A2(n18285), .A3(n18284), .ZN(n21266) );
  INV_X1 U20202 ( .A(n21266), .ZN(n18287) );
  OAI22_X1 U20203 ( .A1(n18289), .A2(n18288), .B1(n18287), .B2(n18350), .ZN(
        P3_U2681) );
  AOI22_X1 U20204 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U20205 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18292) );
  AOI22_X1 U20206 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18291) );
  AOI22_X1 U20207 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18290) );
  NAND4_X1 U20208 ( .A1(n18293), .A2(n18292), .A3(n18291), .A4(n18290), .ZN(
        n18299) );
  AOI22_X1 U20209 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18297) );
  AOI22_X1 U20210 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18296) );
  AOI22_X1 U20211 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18295) );
  AOI22_X1 U20212 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18294) );
  NAND4_X1 U20213 ( .A1(n18297), .A2(n18296), .A3(n18295), .A4(n18294), .ZN(
        n18298) );
  NOR2_X1 U20214 ( .A1(n18299), .A2(n18298), .ZN(n21262) );
  NOR2_X1 U20215 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18300), .ZN(n18302) );
  OAI22_X1 U20216 ( .A1(n21262), .A2(n18350), .B1(n18302), .B2(n18301), .ZN(
        P3_U2683) );
  AOI22_X1 U20217 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U20218 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U20219 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18303) );
  OAI21_X1 U20220 ( .B1(n11190), .B2(n19655), .A(n18303), .ZN(n18309) );
  AOI22_X1 U20221 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18307) );
  AOI22_X1 U20222 ( .A1(n18462), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18306) );
  AOI22_X1 U20223 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18305) );
  AOI22_X1 U20224 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18304) );
  NAND4_X1 U20225 ( .A1(n18307), .A2(n18306), .A3(n18305), .A4(n18304), .ZN(
        n18308) );
  AOI211_X1 U20226 ( .C1(n11130), .C2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A(
        n18309), .B(n18308), .ZN(n18310) );
  NAND3_X1 U20227 ( .A1(n18312), .A2(n18311), .A3(n18310), .ZN(n21280) );
  AOI21_X1 U20228 ( .B1(n18314), .B2(n18313), .A(n18329), .ZN(n18316) );
  MUX2_X1 U20229 ( .A(n21280), .B(n18316), .S(n18315), .Z(P3_U2685) );
  AOI22_X1 U20230 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18321) );
  AOI22_X1 U20231 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18320) );
  AOI22_X1 U20232 ( .A1(n15725), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18317), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18319) );
  AOI22_X1 U20233 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18318) );
  NAND4_X1 U20234 ( .A1(n18321), .A2(n18320), .A3(n18319), .A4(n18318), .ZN(
        n18327) );
  AOI22_X1 U20235 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18325) );
  AOI22_X1 U20236 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18324) );
  AOI22_X1 U20237 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n18323) );
  AOI22_X1 U20238 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18322) );
  NAND4_X1 U20239 ( .A1(n18325), .A2(n18324), .A3(n18323), .A4(n18322), .ZN(
        n18326) );
  NOR2_X1 U20240 ( .A1(n18327), .A2(n18326), .ZN(n21279) );
  INV_X1 U20241 ( .A(n18328), .ZN(n18331) );
  NAND2_X1 U20242 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n18329), .ZN(n18330) );
  OAI21_X1 U20243 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n18331), .A(n18330), .ZN(
        n18332) );
  AOI22_X1 U20244 ( .A1(n18352), .A2(n21279), .B1(n18332), .B2(n18350), .ZN(
        P3_U2684) );
  AOI22_X1 U20245 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U20246 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18335) );
  AOI22_X1 U20247 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18334) );
  AOI22_X1 U20248 ( .A1(n18317), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18333) );
  NAND4_X1 U20249 ( .A1(n18336), .A2(n18335), .A3(n18334), .A4(n18333), .ZN(
        n18342) );
  AOI22_X1 U20250 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18340) );
  AOI22_X1 U20251 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18339) );
  AOI22_X1 U20252 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18338) );
  AOI22_X1 U20253 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18337) );
  NAND4_X1 U20254 ( .A1(n18340), .A2(n18339), .A3(n18338), .A4(n18337), .ZN(
        n18341) );
  NOR2_X1 U20255 ( .A1(n18342), .A2(n18341), .ZN(n21289) );
  AOI21_X1 U20256 ( .B1(n20990), .B2(n18344), .A(n18343), .ZN(n18345) );
  AOI22_X1 U20257 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18348), .B1(n18351), 
        .B2(n18345), .ZN(n18346) );
  OAI21_X1 U20258 ( .B1(n21289), .B2(n18350), .A(n18346), .ZN(P3_U2686) );
  NAND2_X1 U20259 ( .A1(n18354), .A2(n20771), .ZN(n20776) );
  OAI21_X1 U20260 ( .B1(n20771), .B2(n18354), .A(n20776), .ZN(n18347) );
  INV_X1 U20261 ( .A(n18347), .ZN(n20768) );
  AOI22_X1 U20262 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n18348), .B1(n20768), .B2(
        n18351), .ZN(n18349) );
  OAI21_X1 U20263 ( .B1(n19698), .B2(n18350), .A(n18349), .ZN(P3_U2702) );
  AOI22_X1 U20264 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18352), .B1(
        n18351), .B2(n18354), .ZN(n18353) );
  OAI21_X1 U20265 ( .B1(n18355), .B2(n18354), .A(n18353), .ZN(P3_U2703) );
  INV_X1 U20266 ( .A(n18522), .ZN(n18357) );
  OAI21_X1 U20267 ( .B1(n21874), .B2(n20712), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n18356) );
  OAI21_X1 U20268 ( .B1(n18357), .B2(n21936), .A(n18356), .ZN(P3_U2634) );
  INV_X1 U20269 ( .A(n18358), .ZN(n18364) );
  INV_X1 U20270 ( .A(n18359), .ZN(n18360) );
  OAI21_X1 U20271 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n18361), .A(n18360), .ZN(
        n21934) );
  INV_X1 U20272 ( .A(n20707), .ZN(n18362) );
  OAI21_X1 U20273 ( .B1(n18362), .B2(n18364), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18363) );
  OAI221_X1 U20274 ( .B1(n18364), .B2(n21934), .C1(n18364), .C2(n19364), .A(
        n18363), .ZN(P3_U2863) );
  AOI22_X1 U20275 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18374) );
  AOI22_X1 U20276 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18373) );
  AOI22_X1 U20277 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18365) );
  OAI21_X1 U20278 ( .B1(n11184), .B2(n19447), .A(n18365), .ZN(n18371) );
  AOI22_X1 U20279 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18369) );
  AOI22_X1 U20280 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n18368) );
  AOI22_X1 U20281 ( .A1(n15715), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n18367) );
  AOI22_X1 U20282 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18366) );
  NAND4_X1 U20283 ( .A1(n18369), .A2(n18368), .A3(n18367), .A4(n18366), .ZN(
        n18370) );
  AOI211_X1 U20284 ( .C1(n18453), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n18371), .B(n18370), .ZN(n18372) );
  AOI22_X1 U20285 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18461), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18378) );
  AOI22_X1 U20286 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18455), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18377) );
  AOI22_X1 U20287 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18423), .B1(
        P3_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n11126), .ZN(n18376) );
  AOI22_X1 U20288 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20804), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18375) );
  NAND4_X1 U20289 ( .A1(n18378), .A2(n18377), .A3(n18376), .A4(n18375), .ZN(
        n18385) );
  AOI22_X1 U20290 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18379), .B1(
        P3_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n18421), .ZN(n18383) );
  AOI22_X1 U20291 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18382) );
  AOI22_X1 U20292 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18381) );
  AOI22_X1 U20293 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18380) );
  NAND4_X1 U20294 ( .A1(n18383), .A2(n18382), .A3(n18381), .A4(n18380), .ZN(
        n18384) );
  AOI22_X1 U20295 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18389) );
  AOI22_X1 U20296 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18388) );
  AOI22_X1 U20297 ( .A1(n18181), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18387) );
  AOI22_X1 U20298 ( .A1(n18423), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18386) );
  NAND4_X1 U20299 ( .A1(n18389), .A2(n18388), .A3(n18387), .A4(n18386), .ZN(
        n18396) );
  AOI22_X1 U20300 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18390), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18394) );
  AOI22_X1 U20301 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18393) );
  AOI22_X1 U20302 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U20303 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18391) );
  NAND4_X1 U20304 ( .A1(n18394), .A2(n18393), .A3(n18392), .A4(n18391), .ZN(
        n18395) );
  AOI22_X1 U20305 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n18407), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U20306 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18399) );
  AOI22_X1 U20307 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18398) );
  AOI22_X1 U20308 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18397) );
  NAND4_X1 U20309 ( .A1(n18400), .A2(n18399), .A3(n18398), .A4(n18397), .ZN(
        n18406) );
  AOI22_X1 U20310 ( .A1(n11132), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n15713), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n18404) );
  AOI22_X1 U20311 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18403) );
  AOI22_X1 U20312 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18461), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18402) );
  AOI22_X1 U20313 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18401) );
  NAND4_X1 U20314 ( .A1(n18404), .A2(n18403), .A3(n18402), .A4(n18401), .ZN(
        n18405) );
  AOI22_X1 U20315 ( .A1(n11128), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18407), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U20316 ( .A1(n15713), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U20317 ( .A1(n18409), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11127), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18411) );
  AOI22_X1 U20318 ( .A1(n15725), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18410) );
  NAND4_X1 U20319 ( .A1(n18413), .A2(n18412), .A3(n18411), .A4(n18410), .ZN(
        n18420) );
  AOI22_X1 U20320 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18418) );
  AOI22_X1 U20321 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11131), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18417) );
  AOI22_X1 U20322 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18416) );
  AOI22_X1 U20323 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n18415) );
  NAND4_X1 U20324 ( .A1(n18418), .A2(n18417), .A3(n18416), .A4(n18415), .ZN(
        n18419) );
  NOR2_X2 U20325 ( .A1(n18420), .A2(n18419), .ZN(n21374) );
  NOR2_X2 U20326 ( .A1(n21248), .A2(n21374), .ZN(n18495) );
  AOI22_X1 U20327 ( .A1(n18379), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18432) );
  AOI22_X1 U20328 ( .A1(n18421), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18431) );
  AOI22_X1 U20329 ( .A1(n18455), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18422) );
  OAI21_X1 U20330 ( .B1(n11184), .B2(n19612), .A(n18422), .ZN(n18429) );
  AOI22_X1 U20331 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11152), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18427) );
  AOI22_X1 U20332 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18426) );
  AOI22_X1 U20333 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18425) );
  AOI22_X1 U20334 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18423), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18424) );
  NAND4_X1 U20335 ( .A1(n18427), .A2(n18426), .A3(n18425), .A4(n18424), .ZN(
        n18428) );
  AOI211_X1 U20336 ( .C1(n18453), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n18429), .B(n18428), .ZN(n18430) );
  NAND3_X1 U20337 ( .A1(n18432), .A2(n18431), .A3(n18430), .ZN(n21237) );
  NAND2_X1 U20338 ( .A1(n18495), .A2(n21237), .ZN(n18449) );
  AOI22_X1 U20339 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n18414), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n18445) );
  AOI22_X1 U20340 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18444) );
  AOI22_X1 U20341 ( .A1(n18453), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11126), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18433) );
  OAI21_X1 U20342 ( .B1(n11184), .B2(n19529), .A(n18433), .ZN(n18442) );
  AOI22_X1 U20343 ( .A1(n15715), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18440) );
  AOI22_X1 U20344 ( .A1(n11149), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18439) );
  AOI22_X1 U20345 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18435), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18438) );
  AOI22_X1 U20346 ( .A1(n18436), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n18437) );
  NAND4_X1 U20347 ( .A1(n18440), .A2(n18439), .A3(n18438), .A4(n18437), .ZN(
        n18441) );
  AOI211_X1 U20348 ( .C1(n18423), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n18442), .B(n18441), .ZN(n18443) );
  NAND3_X1 U20349 ( .A1(n18445), .A2(n18444), .A3(n18443), .ZN(n21227) );
  NAND2_X1 U20350 ( .A1(n18448), .A2(n21227), .ZN(n18447) );
  AOI21_X1 U20351 ( .B1(n21728), .B2(n18446), .A(n18721), .ZN(n18481) );
  XOR2_X1 U20352 ( .A(n21223), .B(n18447), .Z(n18479) );
  XOR2_X1 U20353 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n18479), .Z(
        n18843) );
  XOR2_X1 U20354 ( .A(n21227), .B(n18448), .Z(n18475) );
  XOR2_X1 U20355 ( .A(n21231), .B(n18449), .Z(n18473) );
  XOR2_X1 U20356 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n18473), .Z(
        n18868) );
  AND2_X1 U20357 ( .A1(n21248), .A2(n21374), .ZN(n18450) );
  NAND2_X1 U20358 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18451), .ZN(
        n18470) );
  NAND2_X1 U20359 ( .A1(n21374), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18469) );
  INV_X1 U20360 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21481) );
  XNOR2_X1 U20361 ( .A(n21374), .B(n21481), .ZN(n18901) );
  AOI22_X1 U20362 ( .A1(n11132), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11149), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18460) );
  AOI22_X1 U20363 ( .A1(n18454), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18453), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18459) );
  AOI22_X1 U20364 ( .A1(n11127), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20804), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18458) );
  AOI22_X1 U20365 ( .A1(n18456), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18455), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18457) );
  NAND4_X1 U20366 ( .A1(n18460), .A2(n18459), .A3(n18458), .A4(n18457), .ZN(
        n18468) );
  AOI22_X1 U20367 ( .A1(n11130), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18434), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18466) );
  AOI22_X1 U20368 ( .A1(n18461), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11128), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18465) );
  AOI22_X1 U20369 ( .A1(n18414), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n18462), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U20370 ( .A1(n11152), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18421), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18463) );
  NAND4_X1 U20371 ( .A1(n18466), .A2(n18465), .A3(n18464), .A4(n18463), .ZN(
        n18467) );
  INV_X1 U20372 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21472) );
  NAND2_X1 U20373 ( .A1(n18901), .A2(n18908), .ZN(n18900) );
  NAND2_X1 U20374 ( .A1(n18469), .A2(n18900), .ZN(n18894) );
  NAND2_X1 U20375 ( .A1(n18895), .A2(n18894), .ZN(n18893) );
  NAND2_X1 U20376 ( .A1(n18470), .A2(n18893), .ZN(n18471) );
  NAND2_X1 U20377 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18471), .ZN(
        n18472) );
  INV_X1 U20378 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21507) );
  XNOR2_X1 U20379 ( .A(n21507), .B(n18471), .ZN(n18884) );
  XOR2_X1 U20380 ( .A(n21237), .B(n18495), .Z(n18883) );
  NAND2_X1 U20381 ( .A1(n18884), .A2(n18883), .ZN(n18882) );
  NAND2_X1 U20382 ( .A1(n18472), .A2(n18882), .ZN(n18867) );
  NAND2_X1 U20383 ( .A1(n18868), .A2(n18867), .ZN(n18866) );
  NAND2_X1 U20384 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18473), .ZN(
        n18474) );
  NAND2_X1 U20385 ( .A1(n18475), .A2(n18477), .ZN(n18478) );
  NAND2_X1 U20386 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18854), .ZN(
        n18853) );
  NAND2_X1 U20387 ( .A1(n18478), .A2(n18853), .ZN(n18842) );
  NAND2_X1 U20388 ( .A1(n18843), .A2(n18842), .ZN(n18841) );
  NAND2_X1 U20389 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18479), .ZN(
        n18480) );
  NAND2_X2 U20390 ( .A1(n18841), .A2(n18480), .ZN(n18548) );
  NAND2_X1 U20391 ( .A1(n18481), .A2(n18548), .ZN(n18483) );
  OAI21_X1 U20392 ( .B1(n18486), .B2(n18485), .A(n18484), .ZN(n21882) );
  NOR2_X1 U20393 ( .A1(n19657), .A2(n18488), .ZN(n21394) );
  NOR2_X1 U20394 ( .A1(n21395), .A2(n21394), .ZN(n21384) );
  INV_X1 U20395 ( .A(n18489), .ZN(n21415) );
  OR2_X2 U20396 ( .A1(n19657), .A2(n21940), .ZN(n18914) );
  OAI21_X1 U20397 ( .B1(n21374), .B2(n18909), .A(n21248), .ZN(n18493) );
  NAND2_X1 U20398 ( .A1(n18493), .A2(n21237), .ZN(n18503) );
  NOR2_X1 U20399 ( .A1(n21231), .A2(n18503), .ZN(n18492) );
  NAND2_X1 U20400 ( .A1(n18492), .A2(n21227), .ZN(n18508) );
  NOR2_X1 U20401 ( .A1(n21223), .A2(n18508), .ZN(n18512) );
  NAND2_X1 U20402 ( .A1(n18512), .A2(n21450), .ZN(n18513) );
  XOR2_X1 U20403 ( .A(n21227), .B(n18492), .Z(n18505) );
  XNOR2_X1 U20404 ( .A(n21237), .B(n18494), .ZN(n18500) );
  AND2_X1 U20405 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18500), .ZN(
        n18501) );
  INV_X1 U20406 ( .A(n18909), .ZN(n21375) );
  INV_X1 U20407 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21492) );
  NOR2_X1 U20408 ( .A1(n18496), .A2(n21492), .ZN(n18499) );
  NOR2_X1 U20409 ( .A1(n21374), .A2(n21472), .ZN(n18498) );
  NAND3_X1 U20410 ( .A1(n18909), .A2(n21374), .A3(n21472), .ZN(n18497) );
  OAI221_X1 U20411 ( .B1(n18498), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18909), .C2(n21374), .A(n18497), .ZN(n18891) );
  NOR2_X1 U20412 ( .A1(n18499), .A2(n18890), .ZN(n18881) );
  XOR2_X1 U20413 ( .A(n21507), .B(n18500), .Z(n18880) );
  NOR2_X1 U20414 ( .A1(n18881), .A2(n18880), .ZN(n18879) );
  INV_X1 U20415 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21506) );
  NOR2_X1 U20416 ( .A1(n18502), .A2(n21506), .ZN(n18504) );
  XNOR2_X1 U20417 ( .A(n21231), .B(n18503), .ZN(n18870) );
  INV_X1 U20418 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18506) );
  XOR2_X1 U20419 ( .A(n18506), .B(n18505), .Z(n18856) );
  XNOR2_X1 U20420 ( .A(n21223), .B(n18508), .ZN(n18510) );
  NOR2_X1 U20421 ( .A1(n18509), .A2(n18510), .ZN(n18511) );
  INV_X1 U20422 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21448) );
  XNOR2_X1 U20423 ( .A(n18510), .B(n18509), .ZN(n18846) );
  XOR2_X1 U20424 ( .A(n21450), .B(n18512), .Z(n18515) );
  NOR2_X1 U20425 ( .A1(n18513), .A2(n18517), .ZN(n18519) );
  INV_X1 U20426 ( .A(n18513), .ZN(n18518) );
  NAND2_X1 U20427 ( .A1(n18515), .A2(n18514), .ZN(n18836) );
  INV_X1 U20428 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21548) );
  OAI22_X2 U20429 ( .A1(n21563), .A2(n18830), .B1(n18915), .B2(n21562), .ZN(
        n18787) );
  INV_X1 U20430 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21596) );
  INV_X1 U20431 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18590) );
  NOR2_X1 U20432 ( .A1(n21869), .A2(n21850), .ZN(n21561) );
  NAND3_X1 U20433 ( .A1(n21561), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18572) );
  NOR2_X1 U20434 ( .A1(n18590), .A2(n18572), .ZN(n21605) );
  INV_X1 U20435 ( .A(n21605), .ZN(n18520) );
  NOR2_X1 U20436 ( .A1(n21596), .A2(n18520), .ZN(n21612) );
  NAND2_X1 U20437 ( .A1(n21612), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n21817) );
  NAND2_X1 U20438 ( .A1(n18787), .A2(n21458), .ZN(n18594) );
  INV_X1 U20439 ( .A(n18594), .ZN(n18757) );
  INV_X1 U20440 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21833) );
  INV_X1 U20441 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21816) );
  NOR2_X1 U20442 ( .A1(n21833), .A2(n21816), .ZN(n21807) );
  INV_X1 U20443 ( .A(n21807), .ZN(n18533) );
  AOI22_X1 U20444 ( .A1(n21622), .A2(n11144), .B1(n21604), .B2(n18779), .ZN(
        n18521) );
  INV_X1 U20445 ( .A(n18521), .ZN(n18565) );
  AOI21_X1 U20446 ( .B1(n18757), .B2(n18533), .A(n18565), .ZN(n18764) );
  INV_X1 U20447 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18537) );
  NAND2_X1 U20448 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18582) );
  NAND2_X1 U20449 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18557) );
  NOR2_X1 U20450 ( .A1(n20979), .A2(n11315), .ZN(n18760) );
  AOI21_X1 U20451 ( .B1(n18568), .B2(n20979), .A(n18886), .ZN(n18767) );
  OAI21_X1 U20452 ( .B1(n18760), .B2(n18910), .A(n18767), .ZN(n18543) );
  AOI21_X1 U20453 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18697), .A(
        n19704), .ZN(n18570) );
  NOR3_X1 U20454 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18570), .A3(
        n20979), .ZN(n18544) );
  NAND2_X2 U20455 ( .A1(n21936), .A2(n18522), .ZN(n21822) );
  INV_X1 U20456 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21821) );
  NOR2_X1 U20457 ( .A1(n18541), .A2(n11315), .ZN(n18540) );
  INV_X1 U20458 ( .A(n18540), .ZN(n21011) );
  OAI21_X1 U20459 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18760), .A(
        n21011), .ZN(n20996) );
  OAI22_X1 U20460 ( .A1(n21822), .A2(n21821), .B1(n18759), .B2(n20996), .ZN(
        n18524) );
  AOI211_X1 U20461 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18543), .A(
        n18544), .B(n18524), .ZN(n18535) );
  NAND2_X1 U20462 ( .A1(n21741), .A2(n18537), .ZN(n18538) );
  INV_X1 U20463 ( .A(n18538), .ZN(n18616) );
  AOI21_X1 U20464 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18721), .A(
        n18616), .ZN(n18532) );
  NOR2_X1 U20465 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18794) );
  INV_X1 U20466 ( .A(n18794), .ZN(n18573) );
  NOR3_X1 U20467 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n18573), .ZN(n18588) );
  NAND2_X1 U20468 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21741), .ZN(
        n18525) );
  AOI22_X1 U20469 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n21741), .B1(
        n18721), .B2(n21548), .ZN(n18818) );
  NAND2_X1 U20470 ( .A1(n18525), .A2(n18816), .ZN(n18791) );
  NAND2_X1 U20471 ( .A1(n18791), .A2(n21458), .ZN(n18530) );
  NAND2_X1 U20472 ( .A1(n21741), .A2(n18755), .ZN(n18644) );
  INV_X1 U20473 ( .A(n18529), .ZN(n18531) );
  NAND2_X1 U20474 ( .A1(n18531), .A2(n18530), .ZN(n18643) );
  NAND2_X1 U20475 ( .A1(n21807), .A2(n18643), .ZN(n18536) );
  NAND2_X1 U20476 ( .A1(n18644), .A2(n18536), .ZN(n18601) );
  XNOR2_X1 U20477 ( .A(n18532), .B(n18601), .ZN(n21819) );
  NOR2_X1 U20478 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18533), .ZN(
        n21818) );
  AOI22_X1 U20479 ( .A1(n18812), .A2(n21819), .B1(n18757), .B2(n21818), .ZN(
        n18534) );
  OAI211_X1 U20480 ( .C1(n18764), .C2(n18537), .A(n18535), .B(n18534), .ZN(
        P3_U2812) );
  INV_X1 U20481 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21787) );
  NOR3_X1 U20482 ( .A1(n21741), .A2(n18537), .A3(n18536), .ZN(n18615) );
  NOR2_X1 U20483 ( .A1(n18538), .A2(n18601), .ZN(n18605) );
  NOR2_X1 U20484 ( .A1(n18615), .A2(n18605), .ZN(n18539) );
  XNOR2_X1 U20485 ( .A(n21787), .B(n18539), .ZN(n21791) );
  NAND2_X1 U20486 ( .A1(n21807), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n21449) );
  NOR2_X1 U20487 ( .A1(n21449), .A2(n18594), .ZN(n18625) );
  INV_X1 U20488 ( .A(n21449), .ZN(n21459) );
  NAND2_X1 U20489 ( .A1(n21459), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n21453) );
  NOR2_X1 U20490 ( .A1(n21604), .A2(n21453), .ZN(n21786) );
  NOR2_X1 U20491 ( .A1(n21622), .A2(n21453), .ZN(n21776) );
  OAI22_X1 U20492 ( .A1(n21786), .A2(n18830), .B1(n21776), .B2(n18915), .ZN(
        n18626) );
  OAI22_X1 U20493 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18540), .B1(
        n11315), .B2(n18620), .ZN(n21013) );
  NOR3_X1 U20494 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18570), .A3(
        n18541), .ZN(n18542) );
  AOI221_X1 U20495 ( .B1(n18544), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(
        n18543), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18542), .ZN(
        n18545) );
  INV_X2 U20496 ( .A(n21822), .ZN(n21866) );
  NAND2_X1 U20497 ( .A1(n21866), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21788) );
  OAI211_X1 U20498 ( .C1(n21013), .C2(n18759), .A(n18545), .B(n21788), .ZN(
        n18546) );
  AOI221_X1 U20499 ( .B1(n18625), .B2(n21787), .C1(n18626), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n18546), .ZN(n18547) );
  OAI21_X1 U20500 ( .B1(n21791), .B2(n18829), .A(n18547), .ZN(P3_U2811) );
  INV_X1 U20501 ( .A(n18552), .ZN(n18553) );
  NAND2_X1 U20502 ( .A1(n18553), .A2(n18715), .ZN(n18559) );
  INV_X1 U20503 ( .A(n18572), .ZN(n21572) );
  INV_X1 U20504 ( .A(n18548), .ZN(n18549) );
  NAND2_X1 U20505 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n21559) );
  NOR3_X1 U20506 ( .A1(n18549), .A2(n21741), .A3(n21559), .ZN(n18801) );
  NAND3_X1 U20507 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21572), .A3(
        n18801), .ZN(n18770) );
  NAND3_X1 U20508 ( .A1(n18588), .A2(n18802), .A3(n18590), .ZN(n18771) );
  AOI22_X1 U20509 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18770), .B1(
        n18771), .B2(n21596), .ZN(n18551) );
  XOR2_X1 U20510 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18551), .Z(
        n21621) );
  INV_X1 U20511 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20954) );
  NOR2_X1 U20512 ( .A1(n21822), .A2(n20954), .ZN(n21619) );
  INV_X1 U20513 ( .A(n18910), .ZN(n18672) );
  NOR2_X1 U20514 ( .A1(n18552), .A2(n11315), .ZN(n18773) );
  INV_X1 U20515 ( .A(n18773), .ZN(n20950) );
  OAI21_X1 U20516 ( .B1(n18553), .B2(n18873), .A(n18911), .ZN(n18774) );
  AOI21_X1 U20517 ( .B1(n18672), .B2(n20950), .A(n18774), .ZN(n18561) );
  INV_X1 U20518 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20962) );
  NAND2_X1 U20519 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18773), .ZN(
        n20963) );
  OAI21_X1 U20520 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18773), .A(
        n20963), .ZN(n20953) );
  OAI22_X1 U20521 ( .A1(n18561), .A2(n20962), .B1(n18759), .B2(n20953), .ZN(
        n18554) );
  AOI211_X1 U20522 ( .C1(n18812), .C2(n21621), .A(n21619), .B(n18554), .ZN(
        n18556) );
  OAI221_X1 U20523 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21612), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18787), .A(n18565), .ZN(
        n18555) );
  OAI211_X1 U20524 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18559), .A(
        n18556), .B(n18555), .ZN(P3_U2815) );
  INV_X1 U20525 ( .A(n18759), .ZN(n18739) );
  INV_X1 U20526 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18560) );
  AND2_X1 U20527 ( .A1(n20981), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18762) );
  AOI21_X1 U20528 ( .B1(n18560), .B2(n20963), .A(n18762), .ZN(n20965) );
  INV_X1 U20529 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n21837) );
  NOR2_X1 U20530 ( .A1(n21822), .A2(n21837), .ZN(n18563) );
  OAI21_X1 U20531 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18557), .ZN(n18558) );
  OAI22_X1 U20532 ( .A1(n18561), .A2(n18560), .B1(n18559), .B2(n18558), .ZN(
        n18562) );
  AOI211_X1 U20533 ( .C1(n18739), .C2(n20965), .A(n18563), .B(n18562), .ZN(
        n18567) );
  AOI22_X1 U20534 ( .A1(n18721), .A2(n21833), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n21741), .ZN(n18564) );
  XOR2_X1 U20535 ( .A(n18643), .B(n18564), .Z(n21835) );
  AOI22_X1 U20536 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18565), .B1(
        n18812), .B2(n21835), .ZN(n18566) );
  OAI211_X1 U20537 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n18594), .A(
        n18567), .B(n18566), .ZN(P3_U2814) );
  NOR2_X1 U20538 ( .A1(n20913), .A2(n11315), .ZN(n18780) );
  AOI21_X1 U20539 ( .B1(n18568), .B2(n20913), .A(n18672), .ZN(n18569) );
  OAI21_X1 U20540 ( .B1(n18780), .B2(n18569), .A(n18911), .ZN(n18587) );
  OR2_X1 U20541 ( .A1(n20913), .A2(n18570), .ZN(n18584) );
  NAND2_X1 U20542 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18780), .ZN(
        n18580) );
  OAI21_X1 U20543 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18780), .A(
        n18580), .ZN(n20916) );
  OAI22_X1 U20544 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18584), .B1(
        n20916), .B2(n18759), .ZN(n18571) );
  AOI21_X1 U20545 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18587), .A(
        n18571), .ZN(n18579) );
  NOR2_X1 U20546 ( .A1(n21562), .A2(n18572), .ZN(n21577) );
  NOR2_X1 U20547 ( .A1(n21563), .A2(n18572), .ZN(n21576) );
  OAI22_X1 U20548 ( .A1(n21577), .A2(n18915), .B1(n21576), .B2(n18830), .ZN(
        n18591) );
  INV_X1 U20549 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21592) );
  AND2_X1 U20550 ( .A1(n21561), .A2(n18801), .ZN(n18575) );
  NOR2_X1 U20551 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18573), .ZN(
        n18574) );
  AOI22_X1 U20552 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18575), .B1(
        n18574), .B2(n18802), .ZN(n18576) );
  XOR2_X1 U20553 ( .A(n21592), .B(n18576), .Z(n21585) );
  AOI22_X1 U20554 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18591), .B1(
        n18812), .B2(n21585), .ZN(n18578) );
  NAND2_X1 U20555 ( .A1(n21866), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n21587) );
  INV_X1 U20556 ( .A(n21561), .ZN(n21567) );
  INV_X1 U20557 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21566) );
  NOR2_X1 U20558 ( .A1(n21567), .A2(n21566), .ZN(n21581) );
  NAND3_X1 U20559 ( .A1(n21581), .A2(n21592), .A3(n18787), .ZN(n18577) );
  NAND4_X1 U20560 ( .A1(n18579), .A2(n18578), .A3(n21587), .A4(n18577), .ZN(
        P3_U2818) );
  INV_X1 U20561 ( .A(n18787), .ZN(n18815) );
  NAND2_X1 U20562 ( .A1(n21572), .A2(n18590), .ZN(n21846) );
  INV_X1 U20563 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18999) );
  NOR2_X1 U20564 ( .A1(n21822), .A2(n18999), .ZN(n18586) );
  INV_X1 U20565 ( .A(n18580), .ZN(n18581) );
  NAND2_X1 U20566 ( .A1(n11258), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20937) );
  OAI21_X1 U20567 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18581), .A(
        n20937), .ZN(n20935) );
  OAI21_X1 U20568 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18582), .ZN(n18583) );
  OAI22_X1 U20569 ( .A1(n18759), .A2(n20935), .B1(n18584), .B2(n18583), .ZN(
        n18585) );
  AOI211_X1 U20570 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18587), .A(
        n18586), .B(n18585), .ZN(n18593) );
  AOI22_X1 U20571 ( .A1(n21572), .A2(n18801), .B1(n18588), .B2(n18802), .ZN(
        n18589) );
  XOR2_X1 U20572 ( .A(n18590), .B(n18589), .Z(n21839) );
  AOI22_X1 U20573 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18591), .B1(
        n18812), .B2(n21839), .ZN(n18592) );
  OAI211_X1 U20574 ( .C1(n18815), .C2(n21846), .A(n18593), .B(n18592), .ZN(
        P3_U2817) );
  NAND2_X1 U20575 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21460) );
  INV_X1 U20576 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21634) );
  NOR2_X1 U20577 ( .A1(n21460), .A2(n21634), .ZN(n21629) );
  NAND2_X1 U20578 ( .A1(n21459), .A2(n21629), .ZN(n21630) );
  NOR2_X1 U20579 ( .A1(n18620), .A2(n11315), .ZN(n18622) );
  OAI22_X1 U20580 ( .A1(n18597), .A2(n18873), .B1(n18622), .B2(n18910), .ZN(
        n18595) );
  NOR2_X1 U20581 ( .A1(n18886), .A2(n18595), .ZN(n18618) );
  OAI21_X1 U20582 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18758), .A(
        n18618), .ZN(n18611) );
  INV_X1 U20583 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18596) );
  INV_X1 U20584 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n21040) );
  NAND2_X1 U20585 ( .A1(n18597), .A2(n18715), .ZN(n18609) );
  AOI221_X1 U20586 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n18596), .C2(n21040), .A(
        n18609), .ZN(n18600) );
  INV_X1 U20587 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21058) );
  NAND2_X1 U20588 ( .A1(n18597), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18621) );
  NOR2_X1 U20589 ( .A1(n21040), .A2(n18621), .ZN(n18598) );
  OAI22_X1 U20590 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18598), .B1(
        n11315), .B2(n18631), .ZN(n21053) );
  OAI22_X1 U20591 ( .A1(n21822), .A2(n21058), .B1(n18759), .B2(n21053), .ZN(
        n18599) );
  AOI211_X1 U20592 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n18611), .A(
        n18600), .B(n18599), .ZN(n18604) );
  OAI22_X1 U20593 ( .A1(n21456), .A2(n18915), .B1(n21752), .B2(n18830), .ZN(
        n18612) );
  NOR2_X1 U20594 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18606) );
  NAND3_X1 U20595 ( .A1(n18616), .A2(n18606), .A3(n21634), .ZN(n18637) );
  NAND3_X1 U20596 ( .A1(n21629), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18601), .ZN(n18647) );
  INV_X1 U20597 ( .A(n18644), .ZN(n18602) );
  AOI21_X1 U20598 ( .B1(n18637), .B2(n18647), .A(n18602), .ZN(n18638) );
  XOR2_X1 U20599 ( .A(n18638), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n21637) );
  AOI22_X1 U20600 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18612), .B1(
        n18812), .B2(n21637), .ZN(n18603) );
  OAI211_X1 U20601 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18708), .A(
        n18604), .B(n18603), .ZN(P3_U2808) );
  INV_X1 U20602 ( .A(n21460), .ZN(n18607) );
  AOI22_X1 U20603 ( .A1(n18607), .A2(n18615), .B1(n18606), .B2(n18605), .ZN(
        n18608) );
  XOR2_X1 U20604 ( .A(n18608), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n21466) );
  INV_X1 U20605 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n21032) );
  NOR2_X1 U20606 ( .A1(n21822), .A2(n21032), .ZN(n21463) );
  XNOR2_X1 U20607 ( .A(n21040), .B(n18621), .ZN(n21036) );
  OAI22_X1 U20608 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18609), .B1(
        n21036), .B2(n18759), .ZN(n18610) );
  AOI211_X1 U20609 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n18611), .A(
        n21463), .B(n18610), .ZN(n18614) );
  NOR2_X1 U20610 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n21460), .ZN(
        n21464) );
  AOI22_X1 U20611 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18612), .B1(
        n21464), .B2(n18625), .ZN(n18613) );
  OAI211_X1 U20612 ( .C1(n21466), .C2(n18829), .A(n18614), .B(n18613), .ZN(
        P3_U2809) );
  OAI221_X1 U20613 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18616), 
        .C1(n21787), .C2(n18615), .A(n18644), .ZN(n18617) );
  XOR2_X1 U20614 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n18617), .Z(
        n21792) );
  AOI221_X1 U20615 ( .B1(n18620), .B2(n18619), .C1(n19703), .C2(n18619), .A(
        n18618), .ZN(n18624) );
  OAI21_X1 U20616 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18622), .A(
        n18621), .ZN(n21028) );
  AOI21_X1 U20617 ( .B1(n18759), .B2(n18758), .A(n21028), .ZN(n18623) );
  AOI211_X1 U20618 ( .C1(P3_REIP_REG_20__SCAN_IN), .C2(n21866), .A(n18624), 
        .B(n18623), .ZN(n18628) );
  NOR2_X1 U20619 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n21787), .ZN(
        n21793) );
  AOI22_X1 U20620 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18626), .B1(
        n18625), .B2(n21793), .ZN(n18627) );
  OAI211_X1 U20621 ( .C1(n18829), .C2(n21792), .A(n18628), .B(n18627), .ZN(
        P3_U2810) );
  INV_X1 U20622 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21641) );
  INV_X1 U20623 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21766) );
  NOR2_X1 U20624 ( .A1(n21641), .A2(n21766), .ZN(n21753) );
  AOI21_X1 U20625 ( .B1(n21753), .B2(n21752), .A(n18830), .ZN(n18635) );
  NOR2_X1 U20626 ( .A1(n21758), .A2(n18915), .ZN(n18629) );
  AOI22_X1 U20627 ( .A1(n21752), .A2(n18635), .B1(n21456), .B2(n18629), .ZN(
        n18642) );
  INV_X1 U20628 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21061) );
  NOR2_X1 U20629 ( .A1(n18631), .A2(n11315), .ZN(n18632) );
  OAI22_X1 U20630 ( .A1(n18651), .A2(n19703), .B1(n18632), .B2(n18910), .ZN(
        n18630) );
  NOR2_X1 U20631 ( .A1(n18886), .A2(n18630), .ZN(n18649) );
  AOI221_X1 U20632 ( .B1(n18631), .B2(n21061), .C1(n19703), .C2(n21061), .A(
        n18649), .ZN(n18634) );
  NAND2_X1 U20633 ( .A1(n18651), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18661) );
  OAI21_X1 U20634 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18632), .A(
        n18661), .ZN(n21064) );
  AOI21_X1 U20635 ( .B1(n18759), .B2(n18758), .A(n21064), .ZN(n18633) );
  AOI211_X1 U20636 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n21866), .A(n18634), 
        .B(n18633), .ZN(n18641) );
  INV_X1 U20637 ( .A(n18635), .ZN(n18636) );
  OAI21_X1 U20638 ( .B1(n21758), .B2(n18915), .A(n18636), .ZN(n18668) );
  NOR2_X1 U20639 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18637), .ZN(
        n18645) );
  OAI221_X1 U20640 ( .B1(n18645), .B2(n18721), .C1(n18645), .C2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n18638), .ZN(n18639) );
  XOR2_X1 U20641 ( .A(n21766), .B(n18639), .Z(n21763) );
  AOI22_X1 U20642 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18668), .B1(
        n18812), .B2(n21763), .ZN(n18640) );
  OAI211_X1 U20643 ( .C1(n18642), .C2(n21641), .A(n18641), .B(n18640), .ZN(
        P3_U2807) );
  INV_X1 U20644 ( .A(n21630), .ZN(n21643) );
  OAI221_X1 U20645 ( .B1(n18646), .B2(n18645), .C1(n18646), .C2(n21766), .A(
        n18644), .ZN(n18660) );
  INV_X1 U20646 ( .A(n21753), .ZN(n21768) );
  OAI21_X1 U20647 ( .B1(n21741), .B2(n18706), .A(n18705), .ZN(n18648) );
  XOR2_X1 U20648 ( .A(n18648), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n21649) );
  OAI21_X1 U20649 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18758), .A(
        n18649), .ZN(n18665) );
  INV_X1 U20650 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18650) );
  INV_X1 U20651 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n21078) );
  NAND2_X1 U20652 ( .A1(n18651), .A2(n18715), .ZN(n18662) );
  AOI221_X1 U20653 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n18650), .C2(n21078), .A(
        n18662), .ZN(n18654) );
  INV_X1 U20654 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n21099) );
  NOR2_X1 U20655 ( .A1(n21078), .A2(n18661), .ZN(n18652) );
  OAI22_X1 U20656 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18652), .B1(
        n11315), .B2(n18698), .ZN(n21092) );
  OAI22_X1 U20657 ( .A1(n21822), .A2(n21099), .B1(n18759), .B2(n21092), .ZN(
        n18653) );
  AOI211_X1 U20658 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n18665), .A(
        n18654), .B(n18653), .ZN(n18658) );
  NAND3_X1 U20659 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21752), .A3(
        n21753), .ZN(n18655) );
  INV_X1 U20660 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21654) );
  XOR2_X1 U20661 ( .A(n18655), .B(n21654), .Z(n21646) );
  NAND2_X1 U20662 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21758), .ZN(
        n18656) );
  XOR2_X1 U20663 ( .A(n21654), .B(n18656), .Z(n21647) );
  AOI22_X1 U20664 ( .A1(n18779), .A2(n21646), .B1(n11144), .B2(n21647), .ZN(
        n18657) );
  OAI211_X1 U20665 ( .C1(n18829), .C2(n21649), .A(n18658), .B(n18657), .ZN(
        P3_U2805) );
  AOI21_X1 U20666 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18660), .A(
        n18659), .ZN(n21775) );
  INV_X1 U20667 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n21087) );
  NOR2_X1 U20668 ( .A1(n21822), .A2(n21087), .ZN(n18664) );
  XNOR2_X1 U20669 ( .A(n21078), .B(n18661), .ZN(n21082) );
  OAI22_X1 U20670 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18662), .B1(
        n21082), .B2(n18759), .ZN(n18663) );
  AOI211_X1 U20671 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n18665), .A(
        n18664), .B(n18663), .ZN(n18670) );
  NOR2_X1 U20672 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21768), .ZN(
        n18666) );
  AOI22_X1 U20673 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18668), .B1(
        n18667), .B2(n18666), .ZN(n18669) );
  OAI211_X1 U20674 ( .C1(n21775), .C2(n18829), .A(n18670), .B(n18669), .ZN(
        P3_U2806) );
  INV_X1 U20675 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n21105) );
  NOR2_X2 U20676 ( .A1(n18698), .A2(n21105), .ZN(n18687) );
  NAND2_X1 U20677 ( .A1(n18671), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18688) );
  NOR2_X1 U20678 ( .A1(n18743), .A2(n11315), .ZN(n18741) );
  AOI21_X1 U20679 ( .B1(n11314), .B2(n18688), .A(n18741), .ZN(n21129) );
  AND3_X1 U20680 ( .A1(n11314), .A2(n18715), .A3(n18671), .ZN(n18676) );
  OAI21_X1 U20681 ( .B1(n18698), .B2(n11315), .A(n18672), .ZN(n18673) );
  OAI211_X1 U20682 ( .C1(n18687), .C2(n18873), .A(n18673), .B(n18911), .ZN(
        n18704) );
  AOI21_X1 U20683 ( .B1(n18697), .B2(n21105), .A(n18704), .ZN(n18696) );
  INV_X1 U20684 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18695) );
  NAND3_X1 U20685 ( .A1(n18687), .A2(n18695), .A3(n18715), .ZN(n18690) );
  NAND2_X1 U20686 ( .A1(n21866), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n18674) );
  OAI221_X1 U20687 ( .B1(n11314), .B2(n18696), .C1(n11314), .C2(n18690), .A(
        n18674), .ZN(n18675) );
  AOI211_X1 U20688 ( .C1(n18739), .C2(n21129), .A(n18676), .B(n18675), .ZN(
        n18684) );
  NAND2_X1 U20689 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21753), .ZN(
        n21655) );
  INV_X1 U20690 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18711) );
  NOR3_X1 U20691 ( .A1(n21655), .A2(n18711), .A3(n21654), .ZN(n21689) );
  NAND2_X1 U20692 ( .A1(n21689), .A2(n21752), .ZN(n21681) );
  AOI22_X1 U20693 ( .A1(n11144), .A2(n21666), .B1(n18779), .B2(n21681), .ZN(
        n18712) );
  NAND2_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18712), .ZN(
        n18692) );
  OAI211_X1 U20695 ( .C1(n18779), .C2(n11144), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18692), .ZN(n18683) );
  INV_X1 U20696 ( .A(n21689), .ZN(n21678) );
  NOR2_X1 U20697 ( .A1(n21678), .A2(n18708), .ZN(n18734) );
  NAND3_X1 U20698 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18734), .A3(
        n21743), .ZN(n18682) );
  NOR2_X1 U20699 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18721), .ZN(
        n18718) );
  AOI21_X1 U20700 ( .B1(n18721), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n18718), .ZN(n21747) );
  AOI21_X1 U20701 ( .B1(n18711), .B2(n21654), .A(n18721), .ZN(n18677) );
  INV_X1 U20702 ( .A(n18677), .ZN(n18678) );
  INV_X1 U20703 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21738) );
  NAND2_X1 U20704 ( .A1(n18679), .A2(n21738), .ZN(n21748) );
  INV_X1 U20705 ( .A(n21748), .ZN(n18719) );
  NOR2_X1 U20706 ( .A1(n18679), .A2(n21738), .ZN(n18720) );
  NOR2_X1 U20707 ( .A1(n18719), .A2(n18720), .ZN(n18686) );
  OAI211_X1 U20708 ( .C1(n21747), .C2(n18680), .A(n18812), .B(n21727), .ZN(
        n18681) );
  NAND4_X1 U20709 ( .A1(n18684), .A2(n18683), .A3(n18682), .A4(n18681), .ZN(
        P3_U2802) );
  OAI21_X1 U20710 ( .B1(n18721), .B2(n18686), .A(n18685), .ZN(n21674) );
  NAND2_X1 U20711 ( .A1(n18687), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18699) );
  INV_X1 U20712 ( .A(n18699), .ZN(n18689) );
  OAI21_X1 U20713 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n18689), .A(
        n18688), .ZN(n21120) );
  NAND2_X1 U20714 ( .A1(n21866), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21675) );
  OAI211_X1 U20715 ( .C1(n18759), .C2(n21120), .A(n18690), .B(n21675), .ZN(
        n18691) );
  AOI21_X1 U20716 ( .B1(n18812), .B2(n21674), .A(n18691), .ZN(n18694) );
  OAI21_X1 U20717 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18734), .A(
        n18692), .ZN(n18693) );
  OAI211_X1 U20718 ( .C1(n18696), .C2(n18695), .A(n18694), .B(n18693), .ZN(
        P3_U2803) );
  OAI21_X1 U20719 ( .B1(n18698), .B2(n19703), .A(n21105), .ZN(n18703) );
  NOR2_X1 U20720 ( .A1(n18698), .A2(n11315), .ZN(n18700) );
  OAI21_X1 U20721 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18700), .A(
        n18699), .ZN(n21109) );
  AOI21_X1 U20722 ( .B1(n18759), .B2(n18758), .A(n21109), .ZN(n18702) );
  NAND2_X1 U20723 ( .A1(n21866), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n21662) );
  INV_X1 U20724 ( .A(n21662), .ZN(n18701) );
  AOI211_X1 U20725 ( .C1(n18704), .C2(n18703), .A(n18702), .B(n18701), .ZN(
        n18710) );
  OAI221_X1 U20726 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n21741), 
        .C1(n21654), .C2(n18706), .A(n18705), .ZN(n18707) );
  XOR2_X1 U20727 ( .A(n18711), .B(n18707), .Z(n21661) );
  OAI211_X1 U20728 ( .C1(n18712), .C2(n18711), .A(n18710), .B(n18709), .ZN(
        P3_U2804) );
  INV_X1 U20729 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21388) );
  NAND2_X1 U20730 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21713) );
  NOR2_X1 U20731 ( .A1(n21743), .A2(n21738), .ZN(n21688) );
  INV_X1 U20732 ( .A(n21688), .ZN(n21677) );
  NOR2_X1 U20733 ( .A1(n21677), .A2(n21681), .ZN(n21734) );
  INV_X1 U20734 ( .A(n21734), .ZN(n18754) );
  OR2_X1 U20735 ( .A1(n21713), .A2(n18754), .ZN(n18713) );
  XNOR2_X1 U20736 ( .A(n21388), .B(n18713), .ZN(n21716) );
  INV_X1 U20737 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21169) );
  INV_X1 U20738 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n18714) );
  INV_X1 U20739 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19001) );
  NOR2_X1 U20740 ( .A1(n21822), .A2(n19001), .ZN(n21720) );
  NAND2_X1 U20741 ( .A1(n11244), .A2(n18715), .ZN(n18731) );
  XNOR2_X1 U20742 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18716) );
  NOR2_X1 U20743 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18758), .ZN(
        n18738) );
  OR2_X1 U20744 ( .A1(n19703), .A2(n11244), .ZN(n18742) );
  OAI211_X1 U20745 ( .C1(n18741), .C2(n18910), .A(n18911), .B(n18742), .ZN(
        n18746) );
  NOR2_X1 U20746 ( .A1(n18738), .A2(n18746), .ZN(n18730) );
  OAI22_X1 U20747 ( .A1(n18731), .A2(n18716), .B1(n18730), .B2(n21169), .ZN(
        n18717) );
  AOI211_X1 U20748 ( .C1(n21155), .C2(n18739), .A(n21720), .B(n18717), .ZN(
        n18725) );
  NAND2_X1 U20749 ( .A1(n18719), .A2(n18718), .ZN(n18747) );
  INV_X1 U20750 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21692) );
  NAND3_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18721), .A3(
        n18720), .ZN(n21731) );
  INV_X1 U20752 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21706) );
  OAI33_X1 U20753 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n18747), .B1(n21692), .B2(
        n21731), .B3(n21706), .ZN(n18722) );
  XNOR2_X1 U20754 ( .A(n21388), .B(n18722), .ZN(n21723) );
  OR2_X1 U20755 ( .A1(n21677), .A2(n21666), .ZN(n21729) );
  NOR2_X1 U20756 ( .A1(n21729), .A2(n21713), .ZN(n18723) );
  XNOR2_X1 U20757 ( .A(n21388), .B(n18723), .ZN(n21721) );
  AOI22_X1 U20758 ( .A1(n18812), .A2(n21723), .B1(n11144), .B2(n21721), .ZN(
        n18724) );
  OAI211_X1 U20759 ( .C1(n21716), .C2(n18830), .A(n18725), .B(n18724), .ZN(
        P3_U2799) );
  AOI22_X1 U20760 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n21731), .B1(
        n18747), .B2(n21692), .ZN(n18726) );
  XOR2_X1 U20761 ( .A(n21706), .B(n18726), .Z(n21712) );
  NOR2_X1 U20762 ( .A1(n21677), .A2(n21692), .ZN(n18735) );
  INV_X1 U20763 ( .A(n18735), .ZN(n21703) );
  OAI21_X1 U20764 ( .B1(n21681), .B2(n21703), .A(n18779), .ZN(n18753) );
  OAI21_X1 U20765 ( .B1(n21682), .B2(n18915), .A(n18753), .ZN(n18750) );
  INV_X1 U20766 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n18729) );
  OAI21_X1 U20767 ( .B1(n18728), .B2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n18727), .ZN(n21178) );
  OAI22_X1 U20768 ( .A1(n18730), .A2(n18729), .B1(n18759), .B2(n21178), .ZN(
        n18733) );
  INV_X1 U20769 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21166) );
  OAI22_X1 U20770 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18731), .B1(
        n21822), .B2(n21166), .ZN(n18732) );
  AOI211_X1 U20771 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18750), .A(
        n18733), .B(n18732), .ZN(n18737) );
  NAND3_X1 U20772 ( .A1(n18735), .A2(n18734), .A3(n21706), .ZN(n18736) );
  OAI211_X1 U20773 ( .C1(n21712), .C2(n18829), .A(n18737), .B(n18736), .ZN(
        P3_U2800) );
  INV_X1 U20774 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21153) );
  NOR2_X1 U20775 ( .A1(n21822), .A2(n21153), .ZN(n21696) );
  NOR2_X1 U20776 ( .A1(n18739), .A2(n18738), .ZN(n18744) );
  OAI21_X1 U20777 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18741), .A(
        n18740), .ZN(n21150) );
  OAI22_X1 U20778 ( .A1(n18744), .A2(n21150), .B1(n18743), .B2(n18742), .ZN(
        n18745) );
  AOI211_X1 U20779 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n18746), .A(
        n21696), .B(n18745), .ZN(n18752) );
  NAND2_X1 U20780 ( .A1(n18747), .A2(n21731), .ZN(n18748) );
  XOR2_X1 U20781 ( .A(n18748), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n21697) );
  OAI21_X1 U20782 ( .B1(n21729), .B2(n18915), .A(n21692), .ZN(n18749) );
  AOI22_X1 U20783 ( .A1(n18812), .A2(n21697), .B1(n18750), .B2(n18749), .ZN(
        n18751) );
  OAI211_X1 U20784 ( .C1(n18754), .C2(n18753), .A(n18752), .B(n18751), .ZN(
        P3_U2801) );
  AOI21_X1 U20785 ( .B1(n20981), .B2(n19704), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18768) );
  OAI21_X1 U20786 ( .B1(n18756), .B2(n21816), .A(n18755), .ZN(n21825) );
  AOI21_X1 U20787 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18757), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18763) );
  INV_X1 U20788 ( .A(n18760), .ZN(n18761) );
  OAI21_X1 U20789 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n18762), .A(
        n18761), .ZN(n20984) );
  OAI22_X1 U20790 ( .A1(n18764), .A2(n18763), .B1(n18896), .B2(n20984), .ZN(
        n18765) );
  AOI21_X1 U20791 ( .B1(n18812), .B2(n21825), .A(n18765), .ZN(n18766) );
  NAND2_X1 U20792 ( .A1(n21866), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21828) );
  OAI211_X1 U20793 ( .C1(n18768), .C2(n18767), .A(n18766), .B(n21828), .ZN(
        P3_U2813) );
  OAI21_X1 U20794 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n11212), .A(
        n21618), .ZN(n21597) );
  AOI21_X1 U20795 ( .B1(n21596), .B2(n18769), .A(n21616), .ZN(n21595) );
  NAND2_X1 U20796 ( .A1(n18771), .A2(n18770), .ZN(n18772) );
  XOR2_X1 U20797 ( .A(n18772), .B(n21596), .Z(n21598) );
  AOI21_X1 U20798 ( .B1(n11311), .B2(n20937), .A(n18773), .ZN(n20939) );
  INV_X1 U20799 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20942) );
  NOR2_X1 U20800 ( .A1(n21822), .A2(n20942), .ZN(n21600) );
  AOI21_X1 U20801 ( .B1(n20939), .B2(n18904), .A(n21600), .ZN(n18776) );
  OAI221_X1 U20802 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11258), .C1(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19704), .A(n18774), .ZN(
        n18775) );
  OAI211_X1 U20803 ( .C1(n21598), .C2(n18829), .A(n18776), .B(n18775), .ZN(
        n18777) );
  AOI21_X1 U20804 ( .B1(n18779), .B2(n21595), .A(n18777), .ZN(n18778) );
  OAI21_X1 U20805 ( .B1(n18915), .B2(n21597), .A(n18778), .ZN(P3_U2816) );
  AOI22_X1 U20806 ( .A1(n11144), .A2(n21562), .B1(n18779), .B2(n21563), .ZN(
        n18814) );
  NAND2_X1 U20807 ( .A1(n18911), .A2(n18873), .ZN(n18905) );
  INV_X1 U20808 ( .A(n18905), .ZN(n18805) );
  AOI21_X1 U20809 ( .B1(n19704), .B2(n18782), .A(n18805), .ZN(n18796) );
  INV_X1 U20810 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20899) );
  NOR2_X1 U20811 ( .A1(n21822), .A2(n20899), .ZN(n18784) );
  NAND2_X1 U20812 ( .A1(n18782), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20901) );
  AOI21_X1 U20813 ( .B1(n11310), .B2(n20901), .A(n18780), .ZN(n18781) );
  INV_X1 U20814 ( .A(n18781), .ZN(n20904) );
  NAND2_X1 U20815 ( .A1(n18782), .A2(n19704), .ZN(n18795) );
  OAI22_X1 U20816 ( .A1(n18896), .A2(n20904), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18795), .ZN(n18783) );
  AOI211_X1 U20817 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18796), .A(
        n18784), .B(n18783), .ZN(n18789) );
  AOI22_X1 U20818 ( .A1(n21561), .A2(n18801), .B1(n18794), .B2(n18802), .ZN(
        n18785) );
  XOR2_X1 U20819 ( .A(n21566), .B(n18785), .Z(n21560) );
  NAND2_X1 U20820 ( .A1(n21561), .A2(n21566), .ZN(n21571) );
  OAI21_X1 U20821 ( .B1(n21561), .B2(n21566), .A(n21571), .ZN(n18786) );
  AOI22_X1 U20822 ( .A1(n18812), .A2(n21560), .B1(n18787), .B2(n18786), .ZN(
        n18788) );
  OAI211_X1 U20823 ( .C1(n18814), .C2(n21566), .A(n18789), .B(n18788), .ZN(
        P3_U2819) );
  AOI21_X1 U20824 ( .B1(n21741), .B2(n21869), .A(n18801), .ZN(n18790) );
  AOI21_X1 U20825 ( .B1(n21869), .B2(n18791), .A(n18790), .ZN(n18793) );
  AOI221_X1 U20826 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18801), .C1(
        n21869), .C2(n18802), .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18792) );
  AOI21_X1 U20827 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18793), .A(
        n18792), .ZN(n21854) );
  NOR3_X1 U20828 ( .A1(n21561), .A2(n18794), .A3(n18815), .ZN(n18799) );
  NAND3_X1 U20829 ( .A1(n18807), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20884) );
  INV_X1 U20830 ( .A(n20884), .ZN(n18808) );
  OAI21_X1 U20831 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18808), .A(
        n20901), .ZN(n20886) );
  INV_X1 U20832 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20871) );
  NAND4_X1 U20833 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(n11159), .A4(n19704), .ZN(
        n18806) );
  NOR2_X1 U20834 ( .A1(n20871), .A2(n18806), .ZN(n18804) );
  AOI22_X1 U20835 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18796), .B1(
        n18804), .B2(n18795), .ZN(n18797) );
  NAND2_X1 U20836 ( .A1(n21866), .A2(P3_REIP_REG_10__SCAN_IN), .ZN(n21855) );
  OAI211_X1 U20837 ( .C1(n18896), .C2(n20886), .A(n18797), .B(n21855), .ZN(
        n18798) );
  AOI211_X1 U20838 ( .C1(n21854), .C2(n18812), .A(n18799), .B(n18798), .ZN(
        n18800) );
  OAI21_X1 U20839 ( .B1(n18814), .B2(n21850), .A(n18800), .ZN(P3_U2820) );
  NOR2_X1 U20840 ( .A1(n18802), .A2(n18801), .ZN(n18803) );
  XOR2_X1 U20841 ( .A(n18803), .B(n21869), .Z(n21864) );
  AOI211_X1 U20842 ( .C1(n18806), .C2(n20871), .A(n18805), .B(n18804), .ZN(
        n18811) );
  NAND2_X1 U20843 ( .A1(n18807), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18821) );
  AOI21_X1 U20844 ( .B1(n20871), .B2(n18821), .A(n18808), .ZN(n18809) );
  INV_X1 U20845 ( .A(n18809), .ZN(n20878) );
  INV_X1 U20846 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n20888) );
  OAI22_X1 U20847 ( .A1(n18896), .A2(n20878), .B1(n21822), .B2(n20888), .ZN(
        n18810) );
  AOI211_X1 U20848 ( .C1(n18812), .C2(n21864), .A(n18811), .B(n18810), .ZN(
        n18813) );
  OAI221_X1 U20849 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18815), .C1(
        n21869), .C2(n18814), .A(n18813), .ZN(P3_U2821) );
  OAI21_X1 U20850 ( .B1(n18818), .B2(n18817), .A(n18816), .ZN(n21552) );
  INV_X1 U20851 ( .A(n21552), .ZN(n21554) );
  AOI21_X1 U20852 ( .B1(n18820), .B2(n21548), .A(n18819), .ZN(n21553) );
  NAND2_X1 U20853 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n11159), .ZN(
        n18822) );
  NOR2_X1 U20854 ( .A1(n11315), .A2(n18822), .ZN(n20862) );
  OAI21_X1 U20855 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20862), .A(
        n18821), .ZN(n20863) );
  OAI21_X1 U20856 ( .B1(n11159), .B2(n18873), .A(n18911), .ZN(n18838) );
  AOI22_X1 U20857 ( .A1(n21866), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18838), .ZN(n18826) );
  INV_X1 U20858 ( .A(n18822), .ZN(n18824) );
  NAND2_X1 U20859 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18823) );
  OAI211_X1 U20860 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18824), .A(
        n19704), .B(n18823), .ZN(n18825) );
  OAI211_X1 U20861 ( .C1(n18896), .C2(n20863), .A(n18826), .B(n18825), .ZN(
        n18827) );
  AOI21_X1 U20862 ( .B1(n11144), .B2(n21553), .A(n18827), .ZN(n18828) );
  OAI221_X1 U20863 ( .B1(n21554), .B2(n18830), .C1(n21552), .C2(n18829), .A(
        n18828), .ZN(P3_U2822) );
  OAI21_X1 U20864 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18832), .A(
        n18831), .ZN(n21546) );
  INV_X1 U20865 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20851) );
  NAND2_X1 U20866 ( .A1(n11159), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18847) );
  AOI21_X1 U20867 ( .B1(n20851), .B2(n18847), .A(n20862), .ZN(n20843) );
  NAND2_X1 U20868 ( .A1(n11159), .A2(n19704), .ZN(n18833) );
  INV_X1 U20869 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n21541) );
  OAI22_X1 U20870 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18833), .B1(
        n21822), .B2(n21541), .ZN(n18834) );
  AOI21_X1 U20871 ( .B1(n20843), .B2(n18904), .A(n18834), .ZN(n18840) );
  NAND2_X1 U20872 ( .A1(n18836), .A2(n18835), .ZN(n18837) );
  XOR2_X1 U20873 ( .A(n18837), .B(n11322), .Z(n21544) );
  AOI22_X1 U20874 ( .A1(n11144), .A2(n21544), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18838), .ZN(n18839) );
  OAI211_X1 U20875 ( .C1(n18914), .C2(n21546), .A(n18840), .B(n18839), .ZN(
        P3_U2823) );
  OAI21_X1 U20876 ( .B1(n18843), .B2(n18842), .A(n18841), .ZN(n21534) );
  NOR2_X1 U20877 ( .A1(n18848), .A2(n19703), .ZN(n18844) );
  AOI22_X1 U20878 ( .A1(n21866), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18844), 
        .B2(n18849), .ZN(n18852) );
  AOI21_X1 U20879 ( .B1(n21448), .B2(n18846), .A(n18845), .ZN(n21531) );
  NOR2_X1 U20880 ( .A1(n18848), .A2(n11315), .ZN(n18859) );
  OAI21_X1 U20881 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18859), .A(
        n18847), .ZN(n20837) );
  OAI21_X1 U20882 ( .B1(n19703), .B2(n18848), .A(n18905), .ZN(n18862) );
  OAI22_X1 U20883 ( .A1(n18896), .A2(n20837), .B1(n18849), .B2(n18862), .ZN(
        n18850) );
  AOI21_X1 U20884 ( .B1(n11144), .B2(n21531), .A(n18850), .ZN(n18851) );
  OAI211_X1 U20885 ( .C1(n18914), .C2(n21534), .A(n18852), .B(n18851), .ZN(
        P3_U2824) );
  OAI21_X1 U20886 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18854), .A(
        n18853), .ZN(n21526) );
  AOI21_X1 U20887 ( .B1(n18857), .B2(n18856), .A(n18855), .ZN(n21523) );
  NOR2_X1 U20888 ( .A1(n18858), .A2(n11315), .ZN(n20818) );
  INV_X1 U20889 ( .A(n18859), .ZN(n18860) );
  OAI21_X1 U20890 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20818), .A(
        n18860), .ZN(n20819) );
  AOI21_X1 U20891 ( .B1(n18861), .B2(n18911), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18863) );
  OAI22_X1 U20892 ( .A1(n18896), .A2(n20819), .B1(n18863), .B2(n18862), .ZN(
        n18864) );
  AOI21_X1 U20893 ( .B1(n11144), .B2(n21523), .A(n18864), .ZN(n18865) );
  NAND2_X1 U20894 ( .A1(n21866), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n21524) );
  OAI211_X1 U20895 ( .C1(n18914), .C2(n21526), .A(n18865), .B(n21524), .ZN(
        P3_U2825) );
  OAI21_X1 U20896 ( .B1(n18868), .B2(n18867), .A(n18866), .ZN(n21515) );
  AOI21_X1 U20897 ( .B1(n18871), .B2(n18870), .A(n18869), .ZN(n21508) );
  INV_X1 U20898 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20816) );
  NOR2_X1 U20899 ( .A1(n21822), .A2(n20816), .ZN(n21513) );
  INV_X1 U20900 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20813) );
  AND3_X1 U20901 ( .A1(n20813), .A2(n18874), .A3(n19704), .ZN(n18872) );
  AOI211_X1 U20902 ( .C1(n11144), .C2(n21508), .A(n21513), .B(n18872), .ZN(
        n18876) );
  OAI21_X1 U20903 ( .B1(n18874), .B2(n18873), .A(n18911), .ZN(n18887) );
  NAND2_X1 U20904 ( .A1(n18874), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18877) );
  AOI21_X1 U20905 ( .B1(n20813), .B2(n18877), .A(n20818), .ZN(n20812) );
  AOI22_X1 U20906 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18887), .B1(
        n20812), .B2(n18904), .ZN(n18875) );
  OAI211_X1 U20907 ( .C1(n18914), .C2(n21515), .A(n18876), .B(n18875), .ZN(
        P3_U2826) );
  NOR2_X1 U20908 ( .A1(n20782), .A2(n11315), .ZN(n18878) );
  OAI21_X1 U20909 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18878), .A(
        n18877), .ZN(n20790) );
  AOI21_X1 U20910 ( .B1(n18881), .B2(n18880), .A(n18879), .ZN(n21502) );
  INV_X1 U20911 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n20793) );
  OAI21_X1 U20912 ( .B1(n18884), .B2(n18883), .A(n18882), .ZN(n21499) );
  OAI22_X1 U20913 ( .A1(n21822), .A2(n20793), .B1(n18914), .B2(n21499), .ZN(
        n18885) );
  AOI21_X1 U20914 ( .B1(n11144), .B2(n21502), .A(n18885), .ZN(n18889) );
  NOR2_X1 U20915 ( .A1(n18886), .A2(n20782), .ZN(n18899) );
  OAI21_X1 U20916 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18899), .A(
        n18887), .ZN(n18888) );
  OAI211_X1 U20917 ( .C1(n18896), .C2(n20790), .A(n18889), .B(n18888), .ZN(
        P3_U2827) );
  AOI21_X1 U20918 ( .B1(n18892), .B2(n18891), .A(n18890), .ZN(n21490) );
  INV_X1 U20919 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18990) );
  NOR2_X1 U20920 ( .A1(n21822), .A2(n18990), .ZN(n21489) );
  AOI22_X1 U20921 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n11315), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20782), .ZN(n20785) );
  OAI21_X1 U20922 ( .B1(n18895), .B2(n18894), .A(n18893), .ZN(n21485) );
  OAI22_X1 U20923 ( .A1(n18896), .A2(n20785), .B1(n18914), .B2(n21485), .ZN(
        n18897) );
  AOI211_X1 U20924 ( .C1(n11144), .C2(n21490), .A(n21489), .B(n18897), .ZN(
        n18898) );
  OAI221_X1 U20925 ( .B1(n18899), .B2(n20782), .C1(n18899), .C2(n19703), .A(
        n18898), .ZN(P3_U2828) );
  OAI21_X1 U20926 ( .B1(n18901), .B2(n18908), .A(n18900), .ZN(n21475) );
  NAND2_X1 U20927 ( .A1(n21472), .A2(n18909), .ZN(n18902) );
  XNOR2_X1 U20928 ( .A(n18902), .B(n18901), .ZN(n21476) );
  AOI22_X1 U20929 ( .A1(n21866), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n11144), 
        .B2(n21476), .ZN(n18907) );
  AOI22_X1 U20930 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18905), .B1(
        n18904), .B2(n11315), .ZN(n18906) );
  OAI211_X1 U20931 ( .C1(n18914), .C2(n21475), .A(n18907), .B(n18906), .ZN(
        P3_U2829) );
  AOI21_X1 U20932 ( .B1(n18909), .B2(n21472), .A(n18908), .ZN(n21471) );
  INV_X1 U20933 ( .A(n21471), .ZN(n21470) );
  NAND3_X1 U20934 ( .A1(n21389), .A2(n18911), .A3(n18910), .ZN(n18912) );
  AOI22_X1 U20935 ( .A1(n21866), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18912), .ZN(n18913) );
  OAI221_X1 U20936 ( .B1(n21471), .B2(n18915), .C1(n21470), .C2(n18914), .A(
        n18913), .ZN(P3_U2830) );
  NOR2_X1 U20937 ( .A1(n19363), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19402) );
  NOR2_X1 U20938 ( .A1(n21903), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19385) );
  INV_X1 U20939 ( .A(n19385), .ZN(n19393) );
  NOR2_X1 U20940 ( .A1(n21900), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19412) );
  INV_X1 U20941 ( .A(n19412), .ZN(n19411) );
  NAND2_X1 U20942 ( .A1(n19393), .A2(n19411), .ZN(n18916) );
  AOI22_X1 U20943 ( .A1(n19402), .A2(n18918), .B1(n18917), .B2(n18916), .ZN(
        n18919) );
  OAI21_X1 U20944 ( .B1(n18920), .B2(n21903), .A(n18919), .ZN(P3_U2866) );
  INV_X1 U20945 ( .A(n19389), .ZN(n19408) );
  OAI21_X1 U20946 ( .B1(n18921), .B2(n19408), .A(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18922) );
  OAI21_X1 U20947 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18923), .A(
        n18922), .ZN(P3_U2864) );
  NOR4_X1 U20948 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18927) );
  NOR4_X1 U20949 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18926) );
  NOR4_X1 U20950 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18925) );
  NOR4_X1 U20951 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18924) );
  NAND4_X1 U20952 ( .A1(n18927), .A2(n18926), .A3(n18925), .A4(n18924), .ZN(
        n18933) );
  NOR4_X1 U20953 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18931) );
  AOI211_X1 U20954 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18930) );
  NOR4_X1 U20955 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18929) );
  NOR4_X1 U20956 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18928) );
  NAND4_X1 U20957 ( .A1(n18931), .A2(n18930), .A3(n18929), .A4(n18928), .ZN(
        n18932) );
  NOR2_X1 U20958 ( .A1(n18933), .A2(n18932), .ZN(n18946) );
  INV_X1 U20959 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18935) );
  OAI21_X1 U20960 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18946), .ZN(n18934) );
  OAI21_X1 U20961 ( .B1(n18946), .B2(n18935), .A(n18934), .ZN(P3_U3293) );
  INV_X1 U20962 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18938) );
  AOI21_X1 U20963 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18936) );
  INV_X1 U20964 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18942) );
  OAI221_X1 U20965 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18936), .C1(n18942), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18946), .ZN(n18937) );
  OAI21_X1 U20966 ( .B1(n18946), .B2(n18938), .A(n18937), .ZN(P3_U3292) );
  INV_X1 U20967 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18940) );
  NOR3_X1 U20968 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18941) );
  OAI21_X1 U20969 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18941), .A(n18946), .ZN(
        n18939) );
  OAI21_X1 U20970 ( .B1(n18946), .B2(n18940), .A(n18939), .ZN(P3_U2638) );
  INV_X1 U20971 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22316) );
  AOI21_X1 U20972 ( .B1(n18942), .B2(n22316), .A(n18941), .ZN(n18945) );
  INV_X1 U20973 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18944) );
  INV_X1 U20974 ( .A(n18946), .ZN(n18943) );
  AOI22_X1 U20975 ( .A1(n18946), .A2(n18945), .B1(n18944), .B2(n18943), .ZN(
        P3_U2639) );
  INV_X1 U20976 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19008) );
  AOI22_X1 U20977 ( .A1(n22323), .A2(n18947), .B1(n19008), .B2(n19006), .ZN(
        P3_U3297) );
  OAI22_X1 U20978 ( .A1(n19006), .A2(n18948), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n22323), .ZN(n18949) );
  INV_X1 U20979 ( .A(n18949), .ZN(P3_U3294) );
  AOI21_X1 U20980 ( .B1(n22377), .B2(n22320), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18950) );
  AOI22_X1 U20981 ( .A1(n22323), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18950), 
        .B2(n19006), .ZN(P3_U2635) );
  INV_X1 U20982 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n21380) );
  AOI22_X1 U20983 ( .A1(n21871), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18951) );
  OAI21_X1 U20984 ( .B1(n21380), .B2(n18967), .A(n18951), .ZN(P3_U2767) );
  INV_X1 U20985 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n21367) );
  AOI22_X1 U20986 ( .A1(n21871), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18952) );
  OAI21_X1 U20987 ( .B1(n21367), .B2(n18967), .A(n18952), .ZN(P3_U2766) );
  INV_X1 U20988 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n21244) );
  AOI22_X1 U20989 ( .A1(n21871), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18953) );
  OAI21_X1 U20990 ( .B1(n21244), .B2(n18967), .A(n18953), .ZN(P3_U2765) );
  INV_X1 U20991 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n21235) );
  AOI22_X1 U20992 ( .A1(n21871), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18954) );
  OAI21_X1 U20993 ( .B1(n21235), .B2(n18967), .A(n18954), .ZN(P3_U2764) );
  INV_X1 U20994 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n21219) );
  AOI22_X1 U20995 ( .A1(n21871), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18955) );
  OAI21_X1 U20996 ( .B1(n21219), .B2(n18967), .A(n18955), .ZN(P3_U2763) );
  INV_X1 U20997 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20747) );
  AOI22_X1 U20998 ( .A1(n21871), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18956) );
  OAI21_X1 U20999 ( .B1(n20747), .B2(n18967), .A(n18956), .ZN(P3_U2762) );
  INV_X1 U21000 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20749) );
  AOI22_X1 U21001 ( .A1(n21871), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18957) );
  OAI21_X1 U21002 ( .B1(n20749), .B2(n18967), .A(n18957), .ZN(P3_U2761) );
  INV_X1 U21003 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n21195) );
  AOI22_X1 U21004 ( .A1(n21871), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18958) );
  OAI21_X1 U21005 ( .B1(n21195), .B2(n18967), .A(n18958), .ZN(P3_U2760) );
  INV_X1 U21006 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n21252) );
  AOI22_X1 U21007 ( .A1(n21871), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18959) );
  OAI21_X1 U21008 ( .B1(n21252), .B2(n18967), .A(n18959), .ZN(P3_U2759) );
  INV_X1 U21009 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n21213) );
  AOI22_X1 U21010 ( .A1(n18977), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18960) );
  OAI21_X1 U21011 ( .B1(n21213), .B2(n18967), .A(n18960), .ZN(P3_U2758) );
  INV_X1 U21012 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n20755) );
  AOI22_X1 U21013 ( .A1(n18977), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18961) );
  OAI21_X1 U21014 ( .B1(n20755), .B2(n18967), .A(n18961), .ZN(P3_U2757) );
  INV_X1 U21015 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n21251) );
  AOI22_X1 U21016 ( .A1(n18977), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18962) );
  OAI21_X1 U21017 ( .B1(n21251), .B2(n18967), .A(n18962), .ZN(P3_U2756) );
  INV_X1 U21018 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20758) );
  AOI22_X1 U21019 ( .A1(n18977), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18963) );
  OAI21_X1 U21020 ( .B1(n20758), .B2(n18967), .A(n18963), .ZN(P3_U2755) );
  INV_X1 U21021 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n21253) );
  AOI22_X1 U21022 ( .A1(n18977), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18964) );
  OAI21_X1 U21023 ( .B1(n21253), .B2(n18967), .A(n18964), .ZN(P3_U2754) );
  INV_X1 U21024 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n21353) );
  AOI22_X1 U21025 ( .A1(n18977), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18965) );
  OAI21_X1 U21026 ( .B1(n21353), .B2(n18967), .A(n18965), .ZN(P3_U2753) );
  INV_X1 U21027 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21360) );
  AOI22_X1 U21028 ( .A1(n18977), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18966) );
  OAI21_X1 U21029 ( .B1(n21360), .B2(n18967), .A(n18966), .ZN(P3_U2752) );
  INV_X1 U21030 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n20716) );
  NAND2_X1 U21031 ( .A1(n18968), .A2(n11367), .ZN(n18987) );
  AOI22_X1 U21032 ( .A1(n18977), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18969) );
  OAI21_X1 U21033 ( .B1(n20716), .B2(n18987), .A(n18969), .ZN(P3_U2751) );
  INV_X1 U21034 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U21035 ( .A1(n18977), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18970) );
  OAI21_X1 U21036 ( .B1(n20718), .B2(n18987), .A(n18970), .ZN(P3_U2750) );
  INV_X1 U21037 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20720) );
  AOI22_X1 U21038 ( .A1(n18977), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18971) );
  OAI21_X1 U21039 ( .B1(n20720), .B2(n18987), .A(n18971), .ZN(P3_U2749) );
  INV_X1 U21040 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U21041 ( .A1(n21871), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18972) );
  OAI21_X1 U21042 ( .B1(n20722), .B2(n18987), .A(n18972), .ZN(P3_U2748) );
  INV_X1 U21043 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n21265) );
  AOI22_X1 U21044 ( .A1(n21871), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18973) );
  OAI21_X1 U21045 ( .B1(n21265), .B2(n18987), .A(n18973), .ZN(P3_U2747) );
  INV_X1 U21046 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n21291) );
  AOI22_X1 U21047 ( .A1(n21871), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18974) );
  OAI21_X1 U21048 ( .B1(n21291), .B2(n18987), .A(n18974), .ZN(P3_U2746) );
  INV_X1 U21049 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n21292) );
  AOI22_X1 U21050 ( .A1(n21871), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18975) );
  OAI21_X1 U21051 ( .B1(n21292), .B2(n18987), .A(n18975), .ZN(P3_U2745) );
  INV_X1 U21052 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n20727) );
  AOI22_X1 U21053 ( .A1(n21871), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18976) );
  OAI21_X1 U21054 ( .B1(n20727), .B2(n18987), .A(n18976), .ZN(P3_U2744) );
  INV_X1 U21055 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n20729) );
  AOI22_X1 U21056 ( .A1(n18977), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18978) );
  OAI21_X1 U21057 ( .B1(n20729), .B2(n18987), .A(n18978), .ZN(P3_U2743) );
  INV_X1 U21058 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U21059 ( .A1(n21871), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18979), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18980) );
  OAI21_X1 U21060 ( .B1(n20731), .B2(n18987), .A(n18980), .ZN(P3_U2742) );
  INV_X1 U21061 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n21300) );
  AOI22_X1 U21062 ( .A1(n21871), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18981) );
  OAI21_X1 U21063 ( .B1(n21300), .B2(n18987), .A(n18981), .ZN(P3_U2741) );
  INV_X1 U21064 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U21065 ( .A1(n21871), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18982) );
  OAI21_X1 U21066 ( .B1(n20735), .B2(n18987), .A(n18982), .ZN(P3_U2740) );
  INV_X1 U21067 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U21068 ( .A1(n21871), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18983) );
  OAI21_X1 U21069 ( .B1(n20737), .B2(n18987), .A(n18983), .ZN(P3_U2739) );
  INV_X1 U21070 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n21312) );
  AOI22_X1 U21071 ( .A1(n21871), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18984) );
  OAI21_X1 U21072 ( .B1(n21312), .B2(n18987), .A(n18984), .ZN(P3_U2738) );
  INV_X1 U21073 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U21074 ( .A1(n21871), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18985), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18986) );
  OAI21_X1 U21075 ( .B1(n20740), .B2(n18987), .A(n18986), .ZN(P3_U2737) );
  AOI21_X1 U21076 ( .B1(n19006), .B2(P3_ADS_N_REG_SCAN_IN), .A(n22317), .ZN(
        n18988) );
  INV_X1 U21077 ( .A(n18988), .ZN(P3_U2633) );
  NOR2_X1 U21078 ( .A1(n19006), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n22371) );
  INV_X2 U21079 ( .A(n22371), .ZN(n19002) );
  AOI22_X1 U21080 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n19006), .ZN(n18989) );
  OAI21_X1 U21081 ( .B1(n18990), .B2(n19002), .A(n18989), .ZN(P3_U3032) );
  AOI22_X1 U21082 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n19006), .ZN(n18991) );
  OAI21_X1 U21083 ( .B1(n20793), .B2(n19002), .A(n18991), .ZN(P3_U3033) );
  AOI22_X1 U21084 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n19006), .ZN(n18992) );
  OAI21_X1 U21085 ( .B1(n20816), .B2(n19002), .A(n18992), .ZN(P3_U3034) );
  INV_X1 U21086 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U21087 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n19006), .ZN(n18993) );
  OAI21_X1 U21088 ( .B1(n20822), .B2(n19002), .A(n18993), .ZN(P3_U3035) );
  INV_X1 U21089 ( .A(n18997), .ZN(n19000) );
  AOI22_X1 U21090 ( .A1(n22371), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n19006), .ZN(n18994) );
  OAI21_X1 U21091 ( .B1(n19000), .B2(n20822), .A(n18994), .ZN(P3_U3036) );
  AOI22_X1 U21092 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_5__SCAN_IN), .B2(n19006), .ZN(n18995) );
  OAI21_X1 U21093 ( .B1(n21541), .B2(n19002), .A(n18995), .ZN(P3_U3037) );
  AOI22_X1 U21094 ( .A1(n22371), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_ADDRESS_REG_6__SCAN_IN), .B2(n19006), .ZN(n18996) );
  OAI21_X1 U21095 ( .B1(n19000), .B2(n21541), .A(n18996), .ZN(P3_U3038) );
  AOI22_X1 U21096 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n18997), .B1(
        P3_ADDRESS_REG_7__SCAN_IN), .B2(n19006), .ZN(n18998) );
  OAI21_X1 U21097 ( .B1(n20888), .B2(n19002), .A(n18998), .ZN(P3_U3039) );
  INV_X1 U21098 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20897) );
  INV_X1 U21099 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20418) );
  OAI222_X1 U21100 ( .A1(n19002), .A2(n20897), .B1(n20418), .B2(n22323), .C1(
        n20888), .C2(n19000), .ZN(P3_U3040) );
  INV_X1 U21101 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n20420) );
  OAI222_X1 U21102 ( .A1(n19002), .A2(n20899), .B1(n20420), .B2(n22323), .C1(
        n20897), .C2(n19000), .ZN(P3_U3041) );
  INV_X1 U21103 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20925) );
  INV_X1 U21104 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n20422) );
  OAI222_X1 U21105 ( .A1(n19002), .A2(n20925), .B1(n20422), .B2(n22323), .C1(
        n20899), .C2(n19000), .ZN(P3_U3042) );
  INV_X1 U21106 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n20424) );
  OAI222_X1 U21107 ( .A1(n19002), .A2(n18999), .B1(n20424), .B2(n22323), .C1(
        n20925), .C2(n19000), .ZN(P3_U3043) );
  INV_X1 U21108 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n20426) );
  OAI222_X1 U21109 ( .A1(n19002), .A2(n20942), .B1(n20426), .B2(n22323), .C1(
        n18999), .C2(n19000), .ZN(P3_U3044) );
  INV_X1 U21110 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20428) );
  OAI222_X1 U21111 ( .A1(n19002), .A2(n20954), .B1(n20428), .B2(n22323), .C1(
        n20942), .C2(n19000), .ZN(P3_U3045) );
  INV_X1 U21112 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n20430) );
  OAI222_X1 U21113 ( .A1(n19002), .A2(n21837), .B1(n20430), .B2(n22323), .C1(
        n20954), .C2(n19000), .ZN(P3_U3046) );
  INV_X1 U21114 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20985) );
  INV_X1 U21115 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n20432) );
  OAI222_X1 U21116 ( .A1(n19002), .A2(n20985), .B1(n20432), .B2(n22323), .C1(
        n21837), .C2(n19000), .ZN(P3_U3047) );
  INV_X1 U21117 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n20434) );
  OAI222_X1 U21118 ( .A1(n19002), .A2(n21821), .B1(n20434), .B2(n22323), .C1(
        n20985), .C2(n19000), .ZN(P3_U3048) );
  INV_X1 U21119 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n21006) );
  INV_X1 U21120 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n20436) );
  OAI222_X1 U21121 ( .A1(n19002), .A2(n21006), .B1(n20436), .B2(n22323), .C1(
        n21821), .C2(n19000), .ZN(P3_U3049) );
  INV_X1 U21122 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n21801) );
  INV_X1 U21123 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n20438) );
  OAI222_X1 U21124 ( .A1(n19002), .A2(n21801), .B1(n20438), .B2(n22323), .C1(
        n21006), .C2(n19000), .ZN(P3_U3050) );
  INV_X1 U21125 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n20440) );
  OAI222_X1 U21126 ( .A1(n19002), .A2(n21032), .B1(n20440), .B2(n22323), .C1(
        n21801), .C2(n19000), .ZN(P3_U3051) );
  INV_X1 U21127 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n20442) );
  OAI222_X1 U21128 ( .A1(n19002), .A2(n21058), .B1(n20442), .B2(n22323), .C1(
        n21032), .C2(n19000), .ZN(P3_U3052) );
  INV_X1 U21129 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n21068) );
  INV_X1 U21130 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n20444) );
  OAI222_X1 U21131 ( .A1(n19002), .A2(n21068), .B1(n20444), .B2(n22323), .C1(
        n21058), .C2(n19000), .ZN(P3_U3053) );
  INV_X1 U21132 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20446) );
  OAI222_X1 U21133 ( .A1(n19002), .A2(n21087), .B1(n20446), .B2(n22323), .C1(
        n21068), .C2(n19000), .ZN(P3_U3054) );
  INV_X1 U21134 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20448) );
  OAI222_X1 U21135 ( .A1(n21087), .A2(n19000), .B1(n20448), .B2(n22323), .C1(
        n21099), .C2(n19002), .ZN(P3_U3055) );
  INV_X1 U21136 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n21100) );
  INV_X1 U21137 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n20450) );
  OAI222_X1 U21138 ( .A1(n19002), .A2(n21100), .B1(n20450), .B2(n22323), .C1(
        n21099), .C2(n19000), .ZN(P3_U3056) );
  INV_X1 U21139 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20452) );
  INV_X1 U21140 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n21117) );
  OAI222_X1 U21141 ( .A1(n21100), .A2(n19000), .B1(n20452), .B2(n22323), .C1(
        n21117), .C2(n19002), .ZN(P3_U3057) );
  INV_X1 U21142 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21750) );
  INV_X1 U21143 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n20454) );
  OAI222_X1 U21144 ( .A1(n19002), .A2(n21750), .B1(n20454), .B2(n22323), .C1(
        n21117), .C2(n19000), .ZN(P3_U3058) );
  INV_X1 U21145 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n20456) );
  OAI222_X1 U21146 ( .A1(n21750), .A2(n19000), .B1(n20456), .B2(n22323), .C1(
        n21153), .C2(n19002), .ZN(P3_U3059) );
  INV_X1 U21147 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n20459) );
  OAI222_X1 U21148 ( .A1(n19002), .A2(n21166), .B1(n20459), .B2(n22323), .C1(
        n21153), .C2(n19000), .ZN(P3_U3060) );
  INV_X1 U21149 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n20462) );
  OAI222_X1 U21150 ( .A1(n19002), .A2(n19001), .B1(n20462), .B2(n22323), .C1(
        n21166), .C2(n19000), .ZN(P3_U3061) );
  OAI22_X1 U21151 ( .A1(n19006), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n22323), .ZN(n19003) );
  INV_X1 U21152 ( .A(n19003), .ZN(P3_U3277) );
  OAI22_X1 U21153 ( .A1(n19006), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n22323), .ZN(n19004) );
  INV_X1 U21154 ( .A(n19004), .ZN(P3_U3276) );
  OAI22_X1 U21155 ( .A1(n19006), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n22323), .ZN(n19005) );
  INV_X1 U21156 ( .A(n19005), .ZN(P3_U3275) );
  OAI22_X1 U21157 ( .A1(n19006), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n22323), .ZN(n19007) );
  INV_X1 U21158 ( .A(n19007), .ZN(P3_U3274) );
  NOR4_X1 U21159 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n19010)
         );
  NOR4_X1 U21160 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n19008), .ZN(n19009) );
  INV_X2 U21161 ( .A(n19699), .ZN(U215) );
  NAND3_X1 U21162 ( .A1(n19010), .A2(n19009), .A3(U215), .ZN(U213) );
  NAND4_X1 U21163 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .A3(n19322), .A4(n22349), .ZN(n19011) );
  OAI211_X1 U21164 ( .C1(n19014), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        n19023) );
  INV_X1 U21165 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22355) );
  NOR2_X1 U21166 ( .A1(n22359), .A2(n19903), .ZN(n19015) );
  NOR2_X1 U21167 ( .A1(n19016), .A2(n19015), .ZN(n19021) );
  AOI21_X1 U21168 ( .B1(n22356), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n11295), 
        .ZN(n19019) );
  MUX2_X1 U21169 ( .A(n19019), .B(n19018), .S(n19017), .Z(n19020) );
  OAI21_X1 U21170 ( .B1(n19021), .B2(n19020), .A(n19023), .ZN(n19022) );
  OAI21_X1 U21171 ( .B1(n19023), .B2(n22355), .A(n19022), .ZN(P2_U3610) );
  INV_X1 U21172 ( .A(n19086), .ZN(n19122) );
  AOI22_X1 U21173 ( .A1(n11121), .A2(P2_EBX_REG_1__SCAN_IN), .B1(n19239), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21174 ( .B1(n19215), .B2(n19025), .A(n19024), .ZN(n19028) );
  OAI22_X1 U21175 ( .A1(n19268), .A2(n19026), .B1(n19256), .B2(n17053), .ZN(
        n19027) );
  AOI211_X1 U21176 ( .C1(n19251), .C2(n19029), .A(n19028), .B(n19027), .ZN(
        n19033) );
  AOI22_X1 U21177 ( .A1(n19031), .A2(n19244), .B1(n19030), .B2(n19842), .ZN(
        n19032) );
  OAI211_X1 U21178 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19122), .A(
        n19033), .B(n19032), .ZN(P2_U2854) );
  OAI21_X1 U21179 ( .B1(n12445), .B2(n19210), .A(n19294), .ZN(n19036) );
  OAI22_X1 U21180 ( .A1(n19034), .A2(n19215), .B1(n11561), .B2(n19208), .ZN(
        n19035) );
  AOI211_X1 U21181 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19237), .A(n19036), .B(
        n19035), .ZN(n19043) );
  NOR2_X1 U21182 ( .A1(n15794), .A2(n19037), .ZN(n19039) );
  XNOR2_X1 U21183 ( .A(n19039), .B(n19038), .ZN(n19041) );
  AOI22_X1 U21184 ( .A1(n19041), .A2(n19244), .B1(n19251), .B2(n19040), .ZN(
        n19042) );
  OAI211_X1 U21185 ( .C1(n19268), .C2(n20070), .A(n19043), .B(n19042), .ZN(
        P2_U2850) );
  OAI21_X1 U21186 ( .B1(n19044), .B2(n19210), .A(n19294), .ZN(n19048) );
  OAI22_X1 U21187 ( .A1(n19256), .A2(n19046), .B1(n19045), .B2(n19215), .ZN(
        n19047) );
  AOI211_X1 U21188 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19239), .A(
        n19048), .B(n19047), .ZN(n19055) );
  NAND2_X1 U21189 ( .A1(n15795), .A2(n19049), .ZN(n19050) );
  XNOR2_X1 U21190 ( .A(n19051), .B(n19050), .ZN(n19053) );
  AOI22_X1 U21191 ( .A1(n19053), .A2(n19244), .B1(n19251), .B2(n19052), .ZN(
        n19054) );
  OAI211_X1 U21192 ( .C1(n19268), .C2(n19056), .A(n19055), .B(n19054), .ZN(
        P2_U2849) );
  NAND2_X1 U21193 ( .A1(n15795), .A2(n19057), .ZN(n19059) );
  XNOR2_X1 U21194 ( .A(n19059), .B(n19058), .ZN(n19068) );
  INV_X1 U21195 ( .A(n19814), .ZN(n19062) );
  AOI22_X1 U21196 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19239), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19237), .ZN(n19060) );
  OAI211_X1 U21197 ( .C1(n19210), .C2(n11907), .A(n19060), .B(n19294), .ZN(
        n19061) );
  AOI21_X1 U21198 ( .B1(n19241), .B2(n19062), .A(n19061), .ZN(n19063) );
  OAI21_X1 U21199 ( .B1(n19064), .B2(n19166), .A(n19063), .ZN(n19065) );
  AOI21_X1 U21200 ( .B1(n19066), .B2(n19261), .A(n19065), .ZN(n19067) );
  OAI21_X1 U21201 ( .B1(n19068), .B2(n19316), .A(n19067), .ZN(P2_U2845) );
  INV_X1 U21202 ( .A(n19069), .ZN(n19076) );
  INV_X1 U21203 ( .A(n19070), .ZN(n19074) );
  AOI22_X1 U21204 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19237), .ZN(n19071) );
  OAI211_X1 U21205 ( .C1(n19072), .C2(n19208), .A(n19294), .B(n19071), .ZN(
        n19073) );
  AOI21_X1 U21206 ( .B1(n19241), .B2(n19074), .A(n19073), .ZN(n19075) );
  OAI21_X1 U21207 ( .B1(n19076), .B2(n19166), .A(n19075), .ZN(n19077) );
  AOI21_X1 U21208 ( .B1(n19078), .B2(n19261), .A(n19077), .ZN(n19082) );
  OAI211_X1 U21209 ( .C1(n19080), .C2(n19083), .A(n19265), .B(n19079), .ZN(
        n19081) );
  OAI211_X1 U21210 ( .C1(n19122), .C2(n19083), .A(n19082), .B(n19081), .ZN(
        P2_U2844) );
  OAI22_X1 U21211 ( .A1(n11908), .A2(n19210), .B1(n19084), .B2(n19256), .ZN(
        n19085) );
  AOI211_X1 U21212 ( .C1(n19087), .C2(n19086), .A(n19124), .B(n19085), .ZN(
        n19098) );
  AOI22_X1 U21213 ( .A1(n19088), .A2(n19261), .B1(n19239), .B2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n19097) );
  OAI22_X1 U21214 ( .A1(n19090), .A2(n19166), .B1(n19089), .B2(n19268), .ZN(
        n19091) );
  INV_X1 U21215 ( .A(n19091), .ZN(n19096) );
  OAI21_X1 U21216 ( .B1(n19094), .B2(n19093), .A(n19092), .ZN(n19095) );
  NAND4_X1 U21217 ( .A1(n19098), .A2(n19097), .A3(n19096), .A4(n19095), .ZN(
        P2_U2842) );
  NAND2_X1 U21218 ( .A1(n15795), .A2(n19099), .ZN(n19101) );
  XNOR2_X1 U21219 ( .A(n19101), .B(n19100), .ZN(n19110) );
  AOI22_X1 U21220 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19239), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19237), .ZN(n19102) );
  OAI211_X1 U21221 ( .C1(n19210), .C2(n12487), .A(n19102), .B(n19294), .ZN(
        n19103) );
  AOI21_X1 U21222 ( .B1(n19104), .B2(n19241), .A(n19103), .ZN(n19105) );
  OAI21_X1 U21223 ( .B1(n19106), .B2(n19166), .A(n19105), .ZN(n19107) );
  AOI21_X1 U21224 ( .B1(n19108), .B2(n19261), .A(n19107), .ZN(n19109) );
  OAI21_X1 U21225 ( .B1(n19110), .B2(n19316), .A(n19109), .ZN(P2_U2839) );
  AOI22_X1 U21226 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19237), .ZN(n19115) );
  AOI22_X1 U21227 ( .A1(n19111), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n19114) );
  OAI211_X1 U21228 ( .C1(n19112), .C2(n19123), .A(n19244), .B(n19131), .ZN(
        n19113) );
  AND4_X1 U21229 ( .A1(n19115), .A2(n19114), .A3(n19294), .A4(n19113), .ZN(
        n19121) );
  INV_X1 U21230 ( .A(n19116), .ZN(n19117) );
  OAI22_X1 U21231 ( .A1(n19118), .A2(n19166), .B1(n19117), .B2(n19268), .ZN(
        n19119) );
  INV_X1 U21232 ( .A(n19119), .ZN(n19120) );
  OAI211_X1 U21233 ( .C1(n19123), .C2(n19122), .A(n19121), .B(n19120), .ZN(
        P2_U2838) );
  AOI21_X1 U21234 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n11121), .A(n19124), .ZN(
        n19125) );
  OAI21_X1 U21235 ( .B1(n11550), .B2(n19208), .A(n19125), .ZN(n19126) );
  AOI21_X1 U21236 ( .B1(n19237), .B2(P2_REIP_REG_18__SCAN_IN), .A(n19126), 
        .ZN(n19127) );
  OAI21_X1 U21237 ( .B1(n19128), .B2(n19166), .A(n19127), .ZN(n19133) );
  AOI211_X1 U21238 ( .C1(n19131), .C2(n19130), .A(n19316), .B(n19129), .ZN(
        n19132) );
  AOI211_X1 U21239 ( .C1(n19261), .C2(n19134), .A(n19133), .B(n19132), .ZN(
        n19135) );
  OAI21_X1 U21240 ( .B1(n19136), .B2(n19268), .A(n19135), .ZN(P2_U2837) );
  INV_X1 U21241 ( .A(n19137), .ZN(n19139) );
  AOI22_X1 U21242 ( .A1(n19139), .A2(n19251), .B1(n19241), .B2(n19138), .ZN(
        n19150) );
  AOI211_X1 U21243 ( .C1(n19142), .C2(n19141), .A(n19316), .B(n19140), .ZN(
        n19145) );
  AOI22_X1 U21244 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19239), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19237), .ZN(n19143) );
  NAND2_X1 U21245 ( .A1(n19294), .A2(n19143), .ZN(n19144) );
  NOR2_X1 U21246 ( .A1(n19145), .A2(n19144), .ZN(n19146) );
  OAI21_X1 U21247 ( .B1(n19210), .B2(n12497), .A(n19146), .ZN(n19147) );
  AOI21_X1 U21248 ( .B1(n19148), .B2(n19261), .A(n19147), .ZN(n19149) );
  NAND2_X1 U21249 ( .A1(n19150), .A2(n19149), .ZN(P2_U2836) );
  AOI22_X1 U21250 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19237), .ZN(n19159) );
  AOI22_X1 U21251 ( .A1(n19151), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n19158) );
  AOI22_X1 U21252 ( .A1(n19152), .A2(n19227), .B1(n20019), .B2(n19241), .ZN(
        n19157) );
  AOI21_X1 U21253 ( .B1(n19154), .B2(n11239), .A(n19153), .ZN(n19155) );
  NAND2_X1 U21254 ( .A1(n19244), .A2(n19155), .ZN(n19156) );
  NAND4_X1 U21255 ( .A1(n19159), .A2(n19158), .A3(n19157), .A4(n19156), .ZN(
        P2_U2833) );
  AOI211_X1 U21256 ( .C1(n19162), .C2(n19161), .A(n19160), .B(n19316), .ZN(
        n19163) );
  INV_X1 U21257 ( .A(n19163), .ZN(n19172) );
  AOI22_X1 U21258 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19237), .ZN(n19171) );
  AOI22_X1 U21259 ( .A1(n19164), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n19170) );
  OAI22_X1 U21260 ( .A1(n19167), .A2(n19166), .B1(n19165), .B2(n19268), .ZN(
        n19168) );
  INV_X1 U21261 ( .A(n19168), .ZN(n19169) );
  NAND4_X1 U21262 ( .A1(n19172), .A2(n19171), .A3(n19170), .A4(n19169), .ZN(
        P2_U2832) );
  AOI22_X1 U21263 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19237), .ZN(n19184) );
  AOI22_X1 U21264 ( .A1(n19173), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n19183) );
  INV_X1 U21265 ( .A(n19174), .ZN(n19175) );
  AOI22_X1 U21266 ( .A1(n19176), .A2(n19227), .B1(n19175), .B2(n19241), .ZN(
        n19182) );
  INV_X1 U21267 ( .A(n19179), .ZN(n19177) );
  OAI221_X1 U21268 ( .B1(n19180), .B2(n19179), .C1(n19178), .C2(n19177), .A(
        n19244), .ZN(n19181) );
  NAND4_X1 U21269 ( .A1(n19184), .A2(n19183), .A3(n19182), .A4(n19181), .ZN(
        P2_U2831) );
  AOI22_X1 U21270 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n11121), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19237), .ZN(n19196) );
  AOI22_X1 U21271 ( .A1(n19185), .A2(n19261), .B1(n19253), .B2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n19195) );
  INV_X1 U21272 ( .A(n19186), .ZN(n19189) );
  INV_X1 U21273 ( .A(n19187), .ZN(n19188) );
  AOI22_X1 U21274 ( .A1(n19189), .A2(n19251), .B1(n19241), .B2(n19188), .ZN(
        n19194) );
  OAI211_X1 U21275 ( .C1(n19192), .C2(n19191), .A(n19244), .B(n19190), .ZN(
        n19193) );
  NAND4_X1 U21276 ( .A1(n19196), .A2(n19195), .A3(n19194), .A4(n19193), .ZN(
        P2_U2830) );
  AOI22_X1 U21277 ( .A1(n19197), .A2(n19261), .B1(P2_EBX_REG_26__SCAN_IN), 
        .B2(n11121), .ZN(n19206) );
  AOI22_X1 U21278 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19239), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19237), .ZN(n19205) );
  AOI22_X1 U21279 ( .A1(n19199), .A2(n19227), .B1(n19198), .B2(n19241), .ZN(
        n19204) );
  OAI211_X1 U21280 ( .C1(n19202), .C2(n19201), .A(n19244), .B(n19200), .ZN(
        n19203) );
  NAND4_X1 U21281 ( .A1(n19206), .A2(n19205), .A3(n19204), .A4(n19203), .ZN(
        P2_U2829) );
  OAI22_X1 U21282 ( .A1(n19209), .A2(n19208), .B1(n19207), .B2(n19256), .ZN(
        n19212) );
  NOR2_X1 U21283 ( .A1(n19210), .A2(n12522), .ZN(n19211) );
  AOI211_X1 U21284 ( .C1(n19213), .C2(n19251), .A(n19212), .B(n19211), .ZN(
        n19214) );
  OAI21_X1 U21285 ( .B1(n19216), .B2(n19215), .A(n19214), .ZN(n19217) );
  INV_X1 U21286 ( .A(n19217), .ZN(n19222) );
  OAI211_X1 U21287 ( .C1(n19220), .C2(n19219), .A(n19244), .B(n19218), .ZN(
        n19221) );
  OAI211_X1 U21288 ( .C1(n19268), .C2(n19223), .A(n19222), .B(n19221), .ZN(
        P2_U2828) );
  AOI22_X1 U21289 ( .A1(n19224), .A2(n19261), .B1(n19237), .B2(
        P2_REIP_REG_28__SCAN_IN), .ZN(n19235) );
  AOI22_X1 U21290 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n11121), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19239), .ZN(n19234) );
  INV_X1 U21291 ( .A(n19225), .ZN(n19226) );
  AOI22_X1 U21292 ( .A1(n19228), .A2(n19227), .B1(n19226), .B2(n19241), .ZN(
        n19233) );
  OAI211_X1 U21293 ( .C1(n19231), .C2(n19230), .A(n19244), .B(n19229), .ZN(
        n19232) );
  NAND4_X1 U21294 ( .A1(n19235), .A2(n19234), .A3(n19233), .A4(n19232), .ZN(
        P2_U2827) );
  INV_X1 U21295 ( .A(n19236), .ZN(n19238) );
  AOI22_X1 U21296 ( .A1(n19238), .A2(n19261), .B1(n19237), .B2(
        P2_REIP_REG_29__SCAN_IN), .ZN(n19250) );
  AOI22_X1 U21297 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n11121), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19239), .ZN(n19249) );
  AOI22_X1 U21298 ( .A1(n19242), .A2(n19251), .B1(n19241), .B2(n19240), .ZN(
        n19248) );
  OAI211_X1 U21299 ( .C1(n19246), .C2(n19245), .A(n19244), .B(n19243), .ZN(
        n19247) );
  NAND4_X1 U21300 ( .A1(n19250), .A2(n19249), .A3(n19248), .A4(n19247), .ZN(
        P2_U2826) );
  AOI22_X1 U21301 ( .A1(n11121), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19253), .ZN(n19257) );
  AND2_X1 U21302 ( .A1(n19257), .A2(n11720), .ZN(n19258) );
  AOI21_X1 U21303 ( .B1(n19262), .B2(n19261), .A(n19260), .ZN(n19267) );
  NAND3_X1 U21304 ( .A1(n19265), .A2(n19264), .A3(n19263), .ZN(n19266) );
  OAI211_X1 U21305 ( .C1(n19269), .C2(n19268), .A(n19267), .B(n19266), .ZN(
        P2_U2824) );
  NAND3_X1 U21306 ( .A1(n19274), .A2(n19271), .A3(n19270), .ZN(n19272) );
  OAI21_X1 U21307 ( .B1(n19274), .B2(n19273), .A(n19272), .ZN(P2_U3595) );
  INV_X1 U21308 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19278) );
  OR2_X1 U21309 ( .A1(n19275), .A2(n19278), .ZN(n19284) );
  AOI22_X1 U21310 ( .A1(n19299), .A2(n19277), .B1(n19298), .B2(n19276), .ZN(
        n19283) );
  NAND2_X1 U21311 ( .A1(n19279), .A2(n19278), .ZN(n19282) );
  NAND2_X1 U21312 ( .A1(n19292), .A2(n19280), .ZN(n19281) );
  AND4_X1 U21313 ( .A1(n19284), .A2(n19283), .A3(n19282), .A4(n19281), .ZN(
        n19286) );
  OAI211_X1 U21314 ( .C1(n19287), .C2(n19302), .A(n19286), .B(n19285), .ZN(
        P2_U3046) );
  AOI211_X1 U21315 ( .C1(n19307), .C2(n19290), .A(n19289), .B(n19288), .ZN(
        n19296) );
  NAND2_X1 U21316 ( .A1(n19292), .A2(n19291), .ZN(n19293) );
  OAI21_X1 U21317 ( .B1(n14116), .B2(n19294), .A(n19293), .ZN(n19295) );
  NOR2_X1 U21318 ( .A1(n19296), .A2(n19295), .ZN(n19306) );
  AOI22_X1 U21319 ( .A1(n19300), .A2(n19299), .B1(n19298), .B2(n19297), .ZN(
        n19301) );
  OAI21_X1 U21320 ( .B1(n19303), .B2(n19302), .A(n19301), .ZN(n19304) );
  INV_X1 U21321 ( .A(n19304), .ZN(n19305) );
  OAI211_X1 U21322 ( .C1(n19308), .C2(n19307), .A(n19306), .B(n19305), .ZN(
        P2_U3038) );
  NAND2_X1 U21323 ( .A1(n19321), .A2(n19309), .ZN(n19326) );
  OAI21_X1 U21324 ( .B1(n19311), .B2(n19310), .A(n19332), .ZN(n19315) );
  NAND2_X1 U21325 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n22359), .ZN(n19312) );
  AOI21_X1 U21326 ( .B1(n19313), .B2(n19326), .A(n19312), .ZN(n19314) );
  AOI21_X1 U21327 ( .B1(n19326), .B2(n19315), .A(n19314), .ZN(n19317) );
  NAND2_X1 U21328 ( .A1(n19317), .A2(n19316), .ZN(P2_U3177) );
  INV_X1 U21329 ( .A(n19318), .ZN(n19331) );
  OAI21_X1 U21330 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19320), .A(n19319), 
        .ZN(n19327) );
  AOI21_X1 U21331 ( .B1(n22359), .B2(n19903), .A(n19321), .ZN(n19323) );
  OAI22_X1 U21332 ( .A1(n19324), .A2(n19332), .B1(n19323), .B2(n19322), .ZN(
        n19325) );
  AOI221_X1 U21333 ( .B1(n22349), .B2(n19327), .C1(n19326), .C2(n19327), .A(
        n19325), .ZN(n19329) );
  OAI211_X1 U21334 ( .C1(n19331), .C2(n19330), .A(n19329), .B(n19328), .ZN(
        P2_U3176) );
  NOR2_X1 U21335 ( .A1(n19333), .A2(n19332), .ZN(n19336) );
  MUX2_X1 U21336 ( .A(P2_MORE_REG_SCAN_IN), .B(n19334), .S(n19336), .Z(
        P2_U3609) );
  OAI21_X1 U21337 ( .B1(n19336), .B2(n12377), .A(n19335), .ZN(P2_U2819) );
  INV_X1 U21338 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20698) );
  INV_X1 U21339 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19362) );
  AOI22_X1 U21340 ( .A1(n19699), .A2(n20698), .B1(n19362), .B2(U215), .ZN(U282) );
  OAI22_X1 U21341 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19699), .ZN(n19337) );
  INV_X1 U21342 ( .A(n19337), .ZN(U281) );
  OAI22_X1 U21343 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19699), .ZN(n19338) );
  INV_X1 U21344 ( .A(n19338), .ZN(U280) );
  OAI22_X1 U21345 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19699), .ZN(n19339) );
  INV_X1 U21346 ( .A(n19339), .ZN(U279) );
  OAI22_X1 U21347 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19699), .ZN(n19340) );
  INV_X1 U21348 ( .A(n19340), .ZN(U278) );
  OAI22_X1 U21349 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19699), .ZN(n19341) );
  INV_X1 U21350 ( .A(n19341), .ZN(U277) );
  OAI22_X1 U21351 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19699), .ZN(n19342) );
  INV_X1 U21352 ( .A(n19342), .ZN(U276) );
  OAI22_X1 U21353 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19699), .ZN(n19343) );
  INV_X1 U21354 ( .A(n19343), .ZN(U275) );
  OAI22_X1 U21355 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19699), .ZN(n19344) );
  INV_X1 U21356 ( .A(n19344), .ZN(U274) );
  OAI22_X1 U21357 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19699), .ZN(n19345) );
  INV_X1 U21358 ( .A(n19345), .ZN(U273) );
  OAI22_X1 U21359 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19699), .ZN(n19346) );
  INV_X1 U21360 ( .A(n19346), .ZN(U272) );
  OAI22_X1 U21361 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19699), .ZN(n19347) );
  INV_X1 U21362 ( .A(n19347), .ZN(U271) );
  OAI22_X1 U21363 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19360), .ZN(n19348) );
  INV_X1 U21364 ( .A(n19348), .ZN(U270) );
  OAI22_X1 U21365 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19699), .ZN(n19349) );
  INV_X1 U21366 ( .A(n19349), .ZN(U269) );
  OAI22_X1 U21367 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19360), .ZN(n19350) );
  INV_X1 U21368 ( .A(n19350), .ZN(U268) );
  OAI22_X1 U21369 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19699), .ZN(n19351) );
  INV_X1 U21370 ( .A(n19351), .ZN(U267) );
  OAI22_X1 U21371 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19360), .ZN(n19352) );
  INV_X1 U21372 ( .A(n19352), .ZN(U266) );
  OAI22_X1 U21373 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19699), .ZN(n19353) );
  INV_X1 U21374 ( .A(n19353), .ZN(U265) );
  OAI22_X1 U21375 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19360), .ZN(n19354) );
  INV_X1 U21376 ( .A(n19354), .ZN(U264) );
  OAI22_X1 U21377 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n19360), .ZN(n19355) );
  INV_X1 U21378 ( .A(n19355), .ZN(U263) );
  OAI22_X1 U21379 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n19360), .ZN(n19356) );
  INV_X1 U21380 ( .A(n19356), .ZN(U262) );
  OAI22_X1 U21381 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n19360), .ZN(n19357) );
  INV_X1 U21382 ( .A(n19357), .ZN(U261) );
  OAI22_X1 U21383 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n19360), .ZN(n19358) );
  INV_X1 U21384 ( .A(n19358), .ZN(U260) );
  OAI22_X1 U21385 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n19360), .ZN(n19359) );
  INV_X1 U21386 ( .A(n19359), .ZN(U259) );
  OAI22_X1 U21387 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19360), .ZN(n19361) );
  INV_X1 U21388 ( .A(n19361), .ZN(U258) );
  NAND3_X1 U21389 ( .A1(n21895), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19373) );
  NOR2_X2 U21390 ( .A1(n19373), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19723) );
  INV_X1 U21391 ( .A(n19723), .ZN(n19660) );
  NOR2_X2 U21392 ( .A1(n19362), .A2(n19703), .ZN(n19442) );
  INV_X1 U21393 ( .A(n19442), .ZN(n19383) );
  INV_X1 U21394 ( .A(n19373), .ZN(n19365) );
  NAND2_X1 U21395 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19365), .ZN(
        n19712) );
  NAND2_X1 U21396 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19704), .ZN(n19436) );
  INV_X1 U21397 ( .A(n19436), .ZN(n19443) );
  NOR2_X1 U21398 ( .A1(n21923), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n20766) );
  INV_X1 U21399 ( .A(n20766), .ZN(n21916) );
  NOR2_X1 U21400 ( .A1(n21903), .A2(n19363), .ZN(n19433) );
  AND2_X1 U21401 ( .A1(n21916), .A2(n19433), .ZN(n19706) );
  INV_X1 U21402 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n21222) );
  NOR2_X2 U21403 ( .A1(n21222), .A2(n19571), .ZN(n19441) );
  AOI22_X1 U21404 ( .A1(n19797), .A2(n19443), .B1(n19706), .B2(n19441), .ZN(
        n19369) );
  NAND2_X1 U21405 ( .A1(n19364), .A2(n19705), .ZN(n19374) );
  INV_X1 U21406 ( .A(n19374), .ZN(n19404) );
  AOI22_X1 U21407 ( .A1(n19704), .A2(n19365), .B1(n19433), .B2(n19404), .ZN(
        n19709) );
  NAND2_X1 U21408 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19433), .ZN(
        n19793) );
  INV_X1 U21409 ( .A(n19793), .ZN(n19781) );
  NOR2_X1 U21410 ( .A1(n19367), .A2(n19366), .ZN(n19449) );
  NAND2_X1 U21411 ( .A1(n21294), .A2(n19449), .ZN(n19428) );
  INV_X1 U21412 ( .A(n19428), .ZN(n19444) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19444), .ZN(n19368) );
  OAI211_X1 U21414 ( .C1(n19660), .C2(n19383), .A(n19369), .B(n19368), .ZN(
        P3_U2995) );
  NAND2_X1 U21415 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19385), .ZN(
        n19384) );
  NOR2_X2 U21416 ( .A1(n21892), .A2(n19384), .ZN(n19729) );
  INV_X1 U21417 ( .A(n19729), .ZN(n19717) );
  NAND2_X1 U21418 ( .A1(n21892), .A2(n19433), .ZN(n19805) );
  INV_X1 U21419 ( .A(n19805), .ZN(n19788) );
  NOR2_X1 U21420 ( .A1(n19797), .A2(n19788), .ZN(n19439) );
  NOR2_X1 U21421 ( .A1(n20766), .A2(n19439), .ZN(n19713) );
  AOI22_X1 U21422 ( .A1(n19723), .A2(n19443), .B1(n19441), .B2(n19713), .ZN(
        n19372) );
  NOR2_X1 U21423 ( .A1(n19723), .A2(n19729), .ZN(n19379) );
  OAI21_X1 U21424 ( .B1(n19379), .B2(n19389), .A(n19439), .ZN(n19370) );
  OAI211_X1 U21425 ( .C1(n19788), .C2(n21923), .A(n19705), .B(n19370), .ZN(
        n19714) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19714), .B1(
        n19444), .B2(n19788), .ZN(n19371) );
  OAI211_X1 U21427 ( .C1(n19383), .C2(n19717), .A(n19372), .B(n19371), .ZN(
        P3_U2987) );
  NOR2_X2 U21428 ( .A1(n19384), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19734) );
  INV_X1 U21429 ( .A(n19734), .ZN(n19727) );
  NOR2_X1 U21430 ( .A1(n20766), .A2(n19373), .ZN(n19718) );
  AOI22_X1 U21431 ( .A1(n19443), .A2(n19729), .B1(n19441), .B2(n19718), .ZN(
        n19378) );
  INV_X1 U21432 ( .A(n19384), .ZN(n19376) );
  NOR2_X1 U21433 ( .A1(n21900), .A2(n21903), .ZN(n19375) );
  NOR2_X1 U21434 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19374), .ZN(
        n19432) );
  AOI22_X1 U21435 ( .A1(n19704), .A2(n19376), .B1(n19375), .B2(n19432), .ZN(
        n19719) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19719), .B1(
        n19444), .B2(n19797), .ZN(n19377) );
  OAI211_X1 U21437 ( .C1(n19383), .C2(n19727), .A(n19378), .B(n19377), .ZN(
        P3_U2979) );
  NAND2_X1 U21438 ( .A1(n21895), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19397) );
  NOR2_X2 U21439 ( .A1(n19393), .A2(n19397), .ZN(n19740) );
  INV_X1 U21440 ( .A(n19740), .ZN(n19583) );
  NOR2_X1 U21441 ( .A1(n20766), .A2(n19379), .ZN(n19722) );
  AOI22_X1 U21442 ( .A1(n19443), .A2(n19734), .B1(n19441), .B2(n19722), .ZN(
        n19382) );
  NOR2_X1 U21443 ( .A1(n19734), .A2(n19740), .ZN(n19388) );
  OAI21_X1 U21444 ( .B1(n21923), .B2(n21892), .A(n19705), .ZN(n19438) );
  OAI22_X1 U21445 ( .A1(n19703), .A2(n19388), .B1(n19438), .B2(n19379), .ZN(
        n19380) );
  INV_X1 U21446 ( .A(n19380), .ZN(n19724) );
  AOI22_X1 U21447 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19444), .ZN(n19381) );
  OAI211_X1 U21448 ( .C1(n19383), .C2(n19583), .A(n19382), .B(n19381), .ZN(
        P3_U2971) );
  NAND2_X1 U21449 ( .A1(n21895), .A2(n21892), .ZN(n21897) );
  NOR2_X2 U21450 ( .A1(n21897), .A2(n19393), .ZN(n19746) );
  NOR2_X1 U21451 ( .A1(n20766), .A2(n19384), .ZN(n19728) );
  AOI22_X1 U21452 ( .A1(n19442), .A2(n19746), .B1(n19441), .B2(n19728), .ZN(
        n19387) );
  OAI211_X1 U21453 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n19704), .A(
        n19404), .B(n19385), .ZN(n19730) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19730), .B1(
        n19444), .B2(n19729), .ZN(n19386) );
  OAI211_X1 U21455 ( .C1(n19436), .C2(n19583), .A(n19387), .B(n19386), .ZN(
        P3_U2963) );
  NAND2_X1 U21456 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19402), .ZN(
        n19629) );
  NOR2_X1 U21457 ( .A1(n20766), .A2(n19388), .ZN(n19733) );
  AOI22_X1 U21458 ( .A1(n19442), .A2(n19752), .B1(n19441), .B2(n19733), .ZN(
        n19392) );
  NAND2_X1 U21459 ( .A1(n19738), .A2(n19629), .ZN(n19399) );
  INV_X1 U21460 ( .A(n19399), .ZN(n19398) );
  OAI21_X1 U21461 ( .B1(n19398), .B2(n19389), .A(n19388), .ZN(n19390) );
  OAI211_X1 U21462 ( .C1(n19734), .C2(n21923), .A(n19705), .B(n19390), .ZN(
        n19735) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19735), .B1(
        n19444), .B2(n19734), .ZN(n19391) );
  OAI211_X1 U21464 ( .C1(n19436), .C2(n19738), .A(n19392), .B(n19391), .ZN(
        P3_U2955) );
  NAND2_X1 U21465 ( .A1(n21892), .A2(n19402), .ZN(n19744) );
  INV_X1 U21466 ( .A(n19744), .ZN(n19757) );
  NAND2_X1 U21467 ( .A1(n21895), .A2(n21916), .ZN(n19430) );
  NOR2_X1 U21468 ( .A1(n19393), .A2(n19430), .ZN(n19739) );
  AOI22_X1 U21469 ( .A1(n19442), .A2(n19757), .B1(n19441), .B2(n19739), .ZN(
        n19396) );
  NOR2_X1 U21470 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19393), .ZN(
        n19394) );
  AOI22_X1 U21471 ( .A1(n19704), .A2(n19402), .B1(n19404), .B2(n19394), .ZN(
        n19741) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19741), .B1(
        n19443), .B2(n19752), .ZN(n19395) );
  OAI211_X1 U21473 ( .C1(n19428), .C2(n19583), .A(n19396), .B(n19395), .ZN(
        P3_U2947) );
  INV_X1 U21474 ( .A(n19397), .ZN(n19415) );
  NAND2_X1 U21475 ( .A1(n19415), .A2(n19412), .ZN(n19755) );
  INV_X1 U21476 ( .A(n19755), .ZN(n19762) );
  NOR2_X1 U21477 ( .A1(n20766), .A2(n19398), .ZN(n19745) );
  AOI22_X1 U21478 ( .A1(n19442), .A2(n19762), .B1(n19441), .B2(n19745), .ZN(
        n19401) );
  NAND2_X1 U21479 ( .A1(n19744), .A2(n19755), .ZN(n19407) );
  INV_X1 U21480 ( .A(n19438), .ZN(n19425) );
  AOI22_X1 U21481 ( .A1(n19704), .A2(n19407), .B1(n19425), .B2(n19399), .ZN(
        n19747) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19747), .B1(
        n19443), .B2(n19757), .ZN(n19400) );
  OAI211_X1 U21483 ( .C1(n19428), .C2(n19738), .A(n19401), .B(n19400), .ZN(
        P3_U2939) );
  NOR2_X2 U21484 ( .A1(n21897), .A2(n19411), .ZN(n19768) );
  INV_X1 U21485 ( .A(n19402), .ZN(n19403) );
  NOR2_X1 U21486 ( .A1(n20766), .A2(n19403), .ZN(n19750) );
  AOI22_X1 U21487 ( .A1(n19442), .A2(n19768), .B1(n19441), .B2(n19750), .ZN(
        n19406) );
  NAND3_X1 U21488 ( .A1(n19412), .A2(n19404), .A3(n19421), .ZN(n19751) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19751), .B1(
        n19444), .B2(n19752), .ZN(n19405) );
  OAI211_X1 U21490 ( .C1(n19436), .C2(n19755), .A(n19406), .B(n19405), .ZN(
        P3_U2931) );
  NAND2_X1 U21491 ( .A1(n21900), .A2(n21903), .ZN(n19429) );
  NOR2_X1 U21492 ( .A1(n21895), .A2(n19429), .ZN(n19419) );
  NAND2_X1 U21493 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19419), .ZN(
        n19766) );
  INV_X1 U21494 ( .A(n19766), .ZN(n19776) );
  AND2_X1 U21495 ( .A1(n21916), .A2(n19407), .ZN(n19756) );
  AOI22_X1 U21496 ( .A1(n19442), .A2(n19776), .B1(n19441), .B2(n19756), .ZN(
        n19410) );
  AOI21_X1 U21497 ( .B1(n19679), .B2(n19766), .A(n19438), .ZN(n19416) );
  AOI22_X1 U21498 ( .A1(n19408), .A2(n19416), .B1(n19425), .B2(n19407), .ZN(
        n19758) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19758), .B1(
        n19443), .B2(n19768), .ZN(n19409) );
  OAI211_X1 U21500 ( .C1(n19428), .C2(n19744), .A(n19410), .B(n19409), .ZN(
        P3_U2923) );
  NAND2_X1 U21501 ( .A1(n21892), .A2(n19419), .ZN(n19772) );
  NOR2_X1 U21502 ( .A1(n19430), .A2(n19411), .ZN(n19761) );
  AOI22_X1 U21503 ( .A1(n19442), .A2(n19782), .B1(n19441), .B2(n19761), .ZN(
        n19414) );
  AOI22_X1 U21504 ( .A1(n19704), .A2(n19419), .B1(n19432), .B2(n19412), .ZN(
        n19763) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19763), .B1(
        n19444), .B2(n19762), .ZN(n19413) );
  OAI211_X1 U21506 ( .C1(n19436), .C2(n19766), .A(n19414), .B(n19413), .ZN(
        P3_U2915) );
  INV_X1 U21507 ( .A(n19429), .ZN(n19431) );
  NAND2_X1 U21508 ( .A1(n19415), .A2(n19431), .ZN(n19642) );
  INV_X1 U21509 ( .A(n19642), .ZN(n19789) );
  AOI21_X1 U21510 ( .B1(n19679), .B2(n19766), .A(n20766), .ZN(n19767) );
  AOI22_X1 U21511 ( .A1(n19442), .A2(n19789), .B1(n19441), .B2(n19767), .ZN(
        n19418) );
  NAND2_X1 U21512 ( .A1(n19772), .A2(n19642), .ZN(n19424) );
  AOI21_X1 U21513 ( .B1(n19704), .B2(n19424), .A(n19416), .ZN(n19769) );
  AOI22_X1 U21514 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19769), .B1(
        n19443), .B2(n19782), .ZN(n19417) );
  OAI211_X1 U21515 ( .C1(n19428), .C2(n19679), .A(n19418), .B(n19417), .ZN(
        P3_U2907) );
  AND2_X1 U21516 ( .A1(n21916), .A2(n19419), .ZN(n19773) );
  AOI22_X1 U21517 ( .A1(n19443), .A2(n19789), .B1(n19441), .B2(n19773), .ZN(
        n19423) );
  OAI21_X1 U21518 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19429), .A(n19766), 
        .ZN(n19420) );
  NAND3_X1 U21519 ( .A1(n19705), .A2(n19421), .A3(n19420), .ZN(n19774) );
  NOR2_X2 U21520 ( .A1(n21897), .A2(n19429), .ZN(n19800) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19774), .B1(
        n19442), .B2(n19800), .ZN(n19422) );
  OAI211_X1 U21522 ( .C1(n19428), .C2(n19766), .A(n19423), .B(n19422), .ZN(
        P3_U2899) );
  AND2_X1 U21523 ( .A1(n21916), .A2(n19424), .ZN(n19780) );
  AOI22_X1 U21524 ( .A1(n19443), .A2(n19800), .B1(n19441), .B2(n19780), .ZN(
        n19427) );
  INV_X1 U21525 ( .A(n19800), .ZN(n19786) );
  NAND2_X1 U21526 ( .A1(n19793), .A2(n19786), .ZN(n19437) );
  AOI22_X1 U21527 ( .A1(n19704), .A2(n19437), .B1(n19425), .B2(n19424), .ZN(
        n19783) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19783), .B1(
        n19442), .B2(n19781), .ZN(n19426) );
  OAI211_X1 U21529 ( .C1(n19428), .C2(n19772), .A(n19427), .B(n19426), .ZN(
        P3_U2891) );
  NOR2_X1 U21530 ( .A1(n19430), .A2(n19429), .ZN(n19787) );
  AOI22_X1 U21531 ( .A1(n19442), .A2(n19788), .B1(n19441), .B2(n19787), .ZN(
        n19435) );
  AOI22_X1 U21532 ( .A1(n19704), .A2(n19433), .B1(n19432), .B2(n19431), .ZN(
        n19790) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19790), .B1(
        n19444), .B2(n19789), .ZN(n19434) );
  OAI211_X1 U21534 ( .C1(n19793), .C2(n19436), .A(n19435), .B(n19434), .ZN(
        P3_U2883) );
  INV_X1 U21535 ( .A(n19437), .ZN(n19440) );
  OAI22_X1 U21536 ( .A1(n19439), .A2(n19703), .B1(n19440), .B2(n19438), .ZN(
        n19798) );
  NOR2_X1 U21537 ( .A1(n20766), .A2(n19440), .ZN(n19795) );
  AOI22_X1 U21538 ( .A1(n19442), .A2(n19797), .B1(n19441), .B2(n19795), .ZN(
        n19446) );
  AOI22_X1 U21539 ( .A1(n19444), .A2(n19800), .B1(n19443), .B2(n19788), .ZN(
        n19445) );
  OAI211_X1 U21540 ( .C1(n19447), .C2(n19798), .A(n19446), .B(n19445), .ZN(
        P3_U2875) );
  OAI22_X1 U21541 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19699), .ZN(n19448) );
  INV_X1 U21542 ( .A(n19448), .ZN(U257) );
  INV_X1 U21543 ( .A(n19449), .ZN(n19707) );
  NOR2_X1 U21544 ( .A1(n19707), .A2(n21433), .ZN(n19484) );
  INV_X1 U21545 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19450) );
  NOR2_X2 U21546 ( .A1(n19450), .A2(n19703), .ZN(n19483) );
  INV_X1 U21547 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n21226) );
  NOR2_X2 U21548 ( .A1(n21226), .A2(n19571), .ZN(n19482) );
  AOI22_X1 U21549 ( .A1(n19723), .A2(n19483), .B1(n19706), .B2(n19482), .ZN(
        n19452) );
  AOI22_X1 U21550 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19709), .B1(
        n19797), .B2(n19485), .ZN(n19451) );
  OAI211_X1 U21551 ( .C1(n19793), .C2(n19481), .A(n19452), .B(n19451), .ZN(
        P3_U2994) );
  AOI22_X1 U21552 ( .A1(n19723), .A2(n19485), .B1(n19713), .B2(n19482), .ZN(
        n19454) );
  AOI22_X1 U21553 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19714), .B1(
        n19729), .B2(n19483), .ZN(n19453) );
  OAI211_X1 U21554 ( .C1(n19805), .C2(n19481), .A(n19454), .B(n19453), .ZN(
        P3_U2986) );
  AOI22_X1 U21555 ( .A1(n19734), .A2(n19483), .B1(n19718), .B2(n19482), .ZN(
        n19456) );
  AOI22_X1 U21556 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19719), .B1(
        n19729), .B2(n19485), .ZN(n19455) );
  OAI211_X1 U21557 ( .C1(n19712), .C2(n19481), .A(n19456), .B(n19455), .ZN(
        P3_U2978) );
  AOI22_X1 U21558 ( .A1(n19740), .A2(n19483), .B1(n19722), .B2(n19482), .ZN(
        n19458) );
  AOI22_X1 U21559 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19724), .B1(
        n19734), .B2(n19485), .ZN(n19457) );
  OAI211_X1 U21560 ( .C1(n19660), .C2(n19481), .A(n19458), .B(n19457), .ZN(
        P3_U2970) );
  AOI22_X1 U21561 ( .A1(n19728), .A2(n19482), .B1(n19746), .B2(n19483), .ZN(
        n19460) );
  AOI22_X1 U21562 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19730), .B1(
        n19740), .B2(n19485), .ZN(n19459) );
  OAI211_X1 U21563 ( .C1(n19717), .C2(n19481), .A(n19460), .B(n19459), .ZN(
        P3_U2962) );
  AOI22_X1 U21564 ( .A1(n19746), .A2(n19485), .B1(n19733), .B2(n19482), .ZN(
        n19462) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19735), .B1(
        n19752), .B2(n19483), .ZN(n19461) );
  OAI211_X1 U21566 ( .C1(n19727), .C2(n19481), .A(n19462), .B(n19461), .ZN(
        P3_U2954) );
  AOI22_X1 U21567 ( .A1(n19752), .A2(n19485), .B1(n19739), .B2(n19482), .ZN(
        n19464) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19741), .B1(
        n19757), .B2(n19483), .ZN(n19463) );
  OAI211_X1 U21569 ( .C1(n19583), .C2(n19481), .A(n19464), .B(n19463), .ZN(
        P3_U2946) );
  AOI22_X1 U21570 ( .A1(n19757), .A2(n19485), .B1(n19745), .B2(n19482), .ZN(
        n19466) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19747), .B1(
        n19762), .B2(n19483), .ZN(n19465) );
  OAI211_X1 U21572 ( .C1(n19738), .C2(n19481), .A(n19466), .B(n19465), .ZN(
        P3_U2938) );
  AOI22_X1 U21573 ( .A1(n19762), .A2(n19485), .B1(n19750), .B2(n19482), .ZN(
        n19468) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19751), .B1(
        n19768), .B2(n19483), .ZN(n19467) );
  OAI211_X1 U21575 ( .C1(n19629), .C2(n19481), .A(n19468), .B(n19467), .ZN(
        P3_U2930) );
  AOI22_X1 U21576 ( .A1(n19768), .A2(n19485), .B1(n19756), .B2(n19482), .ZN(
        n19470) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19758), .B1(
        n19776), .B2(n19483), .ZN(n19469) );
  OAI211_X1 U21578 ( .C1(n19744), .C2(n19481), .A(n19470), .B(n19469), .ZN(
        P3_U2922) );
  AOI22_X1 U21579 ( .A1(n19782), .A2(n19483), .B1(n19761), .B2(n19482), .ZN(
        n19472) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19763), .B1(
        n19776), .B2(n19485), .ZN(n19471) );
  OAI211_X1 U21581 ( .C1(n19755), .C2(n19481), .A(n19472), .B(n19471), .ZN(
        P3_U2914) );
  AOI22_X1 U21582 ( .A1(n19782), .A2(n19485), .B1(n19767), .B2(n19482), .ZN(
        n19474) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19769), .B1(
        n19789), .B2(n19483), .ZN(n19473) );
  OAI211_X1 U21584 ( .C1(n19679), .C2(n19481), .A(n19474), .B(n19473), .ZN(
        P3_U2906) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19482), .ZN(n19476) );
  AOI22_X1 U21586 ( .A1(n19789), .A2(n19485), .B1(n19800), .B2(n19483), .ZN(
        n19475) );
  OAI211_X1 U21587 ( .C1(n19766), .C2(n19481), .A(n19476), .B(n19475), .ZN(
        P3_U2898) );
  AOI22_X1 U21588 ( .A1(n19781), .A2(n19483), .B1(n19780), .B2(n19482), .ZN(
        n19478) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19783), .B1(
        n19800), .B2(n19485), .ZN(n19477) );
  OAI211_X1 U21590 ( .C1(n19772), .C2(n19481), .A(n19478), .B(n19477), .ZN(
        P3_U2890) );
  AOI22_X1 U21591 ( .A1(n19781), .A2(n19485), .B1(n19787), .B2(n19482), .ZN(
        n19480) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19790), .B1(
        n19788), .B2(n19483), .ZN(n19479) );
  OAI211_X1 U21593 ( .C1(n19642), .C2(n19481), .A(n19480), .B(n19479), .ZN(
        P3_U2882) );
  AOI22_X1 U21594 ( .A1(n19797), .A2(n19483), .B1(n19795), .B2(n19482), .ZN(
        n19487) );
  AOI22_X1 U21595 ( .A1(n19788), .A2(n19485), .B1(n19800), .B2(n19484), .ZN(
        n19486) );
  OAI211_X1 U21596 ( .C1(n19488), .C2(n19798), .A(n19487), .B(n19486), .ZN(
        P3_U2874) );
  OAI22_X1 U21597 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19699), .ZN(n19489) );
  INV_X1 U21598 ( .A(n19489), .ZN(U256) );
  INV_X1 U21599 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n21256) );
  NOR2_X1 U21600 ( .A1(n21256), .A2(n19703), .ZN(n19526) );
  INV_X1 U21601 ( .A(n19526), .ZN(n19519) );
  NAND2_X1 U21602 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19704), .ZN(n19522) );
  INV_X1 U21603 ( .A(n19522), .ZN(n19524) );
  AND2_X1 U21604 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n19705), .ZN(n19523) );
  AOI22_X1 U21605 ( .A1(n19723), .A2(n19524), .B1(n19706), .B2(n19523), .ZN(
        n19492) );
  NOR2_X2 U21606 ( .A1(n19490), .A2(n19707), .ZN(n19525) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19525), .ZN(n19491) );
  OAI211_X1 U21608 ( .C1(n19712), .C2(n19519), .A(n19492), .B(n19491), .ZN(
        P3_U2993) );
  AOI22_X1 U21609 ( .A1(n19729), .A2(n19524), .B1(n19713), .B2(n19523), .ZN(
        n19494) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19525), .ZN(n19493) );
  OAI211_X1 U21611 ( .C1(n19660), .C2(n19519), .A(n19494), .B(n19493), .ZN(
        P3_U2985) );
  AOI22_X1 U21612 ( .A1(n19729), .A2(n19526), .B1(n19718), .B2(n19523), .ZN(
        n19496) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19525), .ZN(n19495) );
  OAI211_X1 U21614 ( .C1(n19727), .C2(n19522), .A(n19496), .B(n19495), .ZN(
        P3_U2977) );
  AOI22_X1 U21615 ( .A1(n19740), .A2(n19524), .B1(n19722), .B2(n19523), .ZN(
        n19498) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19525), .ZN(n19497) );
  OAI211_X1 U21617 ( .C1(n19727), .C2(n19519), .A(n19498), .B(n19497), .ZN(
        P3_U2969) );
  AOI22_X1 U21618 ( .A1(n19728), .A2(n19523), .B1(n19746), .B2(n19524), .ZN(
        n19500) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19525), .ZN(n19499) );
  OAI211_X1 U21620 ( .C1(n19583), .C2(n19519), .A(n19500), .B(n19499), .ZN(
        P3_U2961) );
  AOI22_X1 U21621 ( .A1(n19752), .A2(n19524), .B1(n19733), .B2(n19523), .ZN(
        n19502) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19525), .ZN(n19501) );
  OAI211_X1 U21623 ( .C1(n19738), .C2(n19519), .A(n19502), .B(n19501), .ZN(
        P3_U2953) );
  AOI22_X1 U21624 ( .A1(n19752), .A2(n19526), .B1(n19739), .B2(n19523), .ZN(
        n19504) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19525), .ZN(n19503) );
  OAI211_X1 U21626 ( .C1(n19744), .C2(n19522), .A(n19504), .B(n19503), .ZN(
        P3_U2945) );
  AOI22_X1 U21627 ( .A1(n19762), .A2(n19524), .B1(n19745), .B2(n19523), .ZN(
        n19506) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19525), .ZN(n19505) );
  OAI211_X1 U21629 ( .C1(n19744), .C2(n19519), .A(n19506), .B(n19505), .ZN(
        P3_U2937) );
  AOI22_X1 U21630 ( .A1(n19762), .A2(n19526), .B1(n19750), .B2(n19523), .ZN(
        n19508) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19751), .B1(
        n19752), .B2(n19525), .ZN(n19507) );
  OAI211_X1 U21632 ( .C1(n19679), .C2(n19522), .A(n19508), .B(n19507), .ZN(
        P3_U2929) );
  AOI22_X1 U21633 ( .A1(n19776), .A2(n19524), .B1(n19756), .B2(n19523), .ZN(
        n19510) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19525), .ZN(n19509) );
  OAI211_X1 U21635 ( .C1(n19679), .C2(n19519), .A(n19510), .B(n19509), .ZN(
        P3_U2921) );
  AOI22_X1 U21636 ( .A1(n19782), .A2(n19524), .B1(n19761), .B2(n19523), .ZN(
        n19512) );
  AOI22_X1 U21637 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19525), .ZN(n19511) );
  OAI211_X1 U21638 ( .C1(n19766), .C2(n19519), .A(n19512), .B(n19511), .ZN(
        P3_U2913) );
  AOI22_X1 U21639 ( .A1(n19789), .A2(n19524), .B1(n19767), .B2(n19523), .ZN(
        n19514) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19525), .ZN(n19513) );
  OAI211_X1 U21641 ( .C1(n19772), .C2(n19519), .A(n19514), .B(n19513), .ZN(
        P3_U2905) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19523), .ZN(n19516) );
  AOI22_X1 U21643 ( .A1(n19776), .A2(n19525), .B1(n19789), .B2(n19526), .ZN(
        n19515) );
  OAI211_X1 U21644 ( .C1(n19786), .C2(n19522), .A(n19516), .B(n19515), .ZN(
        P3_U2897) );
  AOI22_X1 U21645 ( .A1(n19781), .A2(n19524), .B1(n19780), .B2(n19523), .ZN(
        n19518) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19525), .ZN(n19517) );
  OAI211_X1 U21647 ( .C1(n19786), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P3_U2889) );
  AOI22_X1 U21648 ( .A1(n19781), .A2(n19526), .B1(n19787), .B2(n19523), .ZN(
        n19521) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19525), .ZN(n19520) );
  OAI211_X1 U21650 ( .C1(n19805), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P3_U2881) );
  AOI22_X1 U21651 ( .A1(n19797), .A2(n19524), .B1(n19795), .B2(n19523), .ZN(
        n19528) );
  AOI22_X1 U21652 ( .A1(n19788), .A2(n19526), .B1(n19800), .B2(n19525), .ZN(
        n19527) );
  OAI211_X1 U21653 ( .C1(n19529), .C2(n19798), .A(n19528), .B(n19527), .ZN(
        P3_U2873) );
  OAI22_X1 U21654 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19699), .ZN(n19530) );
  INV_X1 U21655 ( .A(n19530), .ZN(U255) );
  NAND2_X1 U21656 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19704), .ZN(n19562) );
  NAND2_X1 U21657 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n19704), .ZN(n19557) );
  INV_X1 U21658 ( .A(n19557), .ZN(n19564) );
  INV_X1 U21659 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n21234) );
  NOR2_X2 U21660 ( .A1(n21234), .A2(n19571), .ZN(n19563) );
  AOI22_X1 U21661 ( .A1(n19797), .A2(n19564), .B1(n19706), .B2(n19563), .ZN(
        n19532) );
  NOR2_X2 U21662 ( .A1(n21442), .A2(n19707), .ZN(n19565) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19565), .ZN(n19531) );
  OAI211_X1 U21664 ( .C1(n19660), .C2(n19562), .A(n19532), .B(n19531), .ZN(
        P3_U2992) );
  AOI22_X1 U21665 ( .A1(n19723), .A2(n19564), .B1(n19713), .B2(n19563), .ZN(
        n19534) );
  AOI22_X1 U21666 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19565), .ZN(n19533) );
  OAI211_X1 U21667 ( .C1(n19717), .C2(n19562), .A(n19534), .B(n19533), .ZN(
        P3_U2984) );
  AOI22_X1 U21668 ( .A1(n19729), .A2(n19564), .B1(n19718), .B2(n19563), .ZN(
        n19536) );
  AOI22_X1 U21669 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19565), .ZN(n19535) );
  OAI211_X1 U21670 ( .C1(n19727), .C2(n19562), .A(n19536), .B(n19535), .ZN(
        P3_U2976) );
  INV_X1 U21671 ( .A(n19562), .ZN(n19566) );
  AOI22_X1 U21672 ( .A1(n19740), .A2(n19566), .B1(n19722), .B2(n19563), .ZN(
        n19538) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19565), .ZN(n19537) );
  OAI211_X1 U21674 ( .C1(n19727), .C2(n19557), .A(n19538), .B(n19537), .ZN(
        P3_U2968) );
  AOI22_X1 U21675 ( .A1(n19728), .A2(n19563), .B1(n19746), .B2(n19566), .ZN(
        n19540) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19565), .ZN(n19539) );
  OAI211_X1 U21677 ( .C1(n19583), .C2(n19557), .A(n19540), .B(n19539), .ZN(
        P3_U2960) );
  AOI22_X1 U21678 ( .A1(n19746), .A2(n19564), .B1(n19733), .B2(n19563), .ZN(
        n19542) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19565), .ZN(n19541) );
  OAI211_X1 U21680 ( .C1(n19629), .C2(n19562), .A(n19542), .B(n19541), .ZN(
        P3_U2952) );
  AOI22_X1 U21681 ( .A1(n19752), .A2(n19564), .B1(n19739), .B2(n19563), .ZN(
        n19544) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19565), .ZN(n19543) );
  OAI211_X1 U21683 ( .C1(n19744), .C2(n19562), .A(n19544), .B(n19543), .ZN(
        P3_U2944) );
  AOI22_X1 U21684 ( .A1(n19757), .A2(n19564), .B1(n19745), .B2(n19563), .ZN(
        n19546) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19565), .ZN(n19545) );
  OAI211_X1 U21686 ( .C1(n19755), .C2(n19562), .A(n19546), .B(n19545), .ZN(
        P3_U2936) );
  AOI22_X1 U21687 ( .A1(n19762), .A2(n19564), .B1(n19750), .B2(n19563), .ZN(
        n19548) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19751), .B1(
        n19752), .B2(n19565), .ZN(n19547) );
  OAI211_X1 U21689 ( .C1(n19679), .C2(n19562), .A(n19548), .B(n19547), .ZN(
        P3_U2928) );
  AOI22_X1 U21690 ( .A1(n19768), .A2(n19564), .B1(n19756), .B2(n19563), .ZN(
        n19550) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19565), .ZN(n19549) );
  OAI211_X1 U21692 ( .C1(n19766), .C2(n19562), .A(n19550), .B(n19549), .ZN(
        P3_U2920) );
  AOI22_X1 U21693 ( .A1(n19782), .A2(n19566), .B1(n19761), .B2(n19563), .ZN(
        n19552) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19565), .ZN(n19551) );
  OAI211_X1 U21695 ( .C1(n19766), .C2(n19557), .A(n19552), .B(n19551), .ZN(
        P3_U2912) );
  AOI22_X1 U21696 ( .A1(n19782), .A2(n19564), .B1(n19767), .B2(n19563), .ZN(
        n19554) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19565), .ZN(n19553) );
  OAI211_X1 U21698 ( .C1(n19642), .C2(n19562), .A(n19554), .B(n19553), .ZN(
        P3_U2904) );
  AOI22_X1 U21699 ( .A1(n19800), .A2(n19566), .B1(n19773), .B2(n19563), .ZN(
        n19556) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19774), .B1(
        n19776), .B2(n19565), .ZN(n19555) );
  OAI211_X1 U21701 ( .C1(n19642), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P3_U2896) );
  AOI22_X1 U21702 ( .A1(n19800), .A2(n19564), .B1(n19780), .B2(n19563), .ZN(
        n19559) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19565), .ZN(n19558) );
  OAI211_X1 U21704 ( .C1(n19793), .C2(n19562), .A(n19559), .B(n19558), .ZN(
        P3_U2888) );
  AOI22_X1 U21705 ( .A1(n19781), .A2(n19564), .B1(n19787), .B2(n19563), .ZN(
        n19561) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19565), .ZN(n19560) );
  OAI211_X1 U21707 ( .C1(n19805), .C2(n19562), .A(n19561), .B(n19560), .ZN(
        P3_U2880) );
  AOI22_X1 U21708 ( .A1(n19788), .A2(n19564), .B1(n19795), .B2(n19563), .ZN(
        n19568) );
  AOI22_X1 U21709 ( .A1(n19797), .A2(n19566), .B1(n19800), .B2(n19565), .ZN(
        n19567) );
  OAI211_X1 U21710 ( .C1(n19569), .C2(n19798), .A(n19568), .B(n19567), .ZN(
        P3_U2872) );
  OAI22_X1 U21711 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19699), .ZN(n19570) );
  INV_X1 U21712 ( .A(n19570), .ZN(U254) );
  INV_X1 U21713 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n21329) );
  NOR2_X1 U21714 ( .A1(n21329), .A2(n19703), .ZN(n19607) );
  NAND2_X1 U21715 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19704), .ZN(n19605) );
  INV_X1 U21716 ( .A(n19605), .ZN(n19609) );
  INV_X1 U21717 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n21242) );
  NOR2_X2 U21718 ( .A1(n21242), .A2(n19571), .ZN(n19606) );
  AOI22_X1 U21719 ( .A1(n19797), .A2(n19609), .B1(n19706), .B2(n19606), .ZN(
        n19574) );
  NOR2_X2 U21720 ( .A1(n19572), .A2(n19707), .ZN(n19608) );
  AOI22_X1 U21721 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19608), .ZN(n19573) );
  OAI211_X1 U21722 ( .C1(n19660), .C2(n19602), .A(n19574), .B(n19573), .ZN(
        P3_U2991) );
  AOI22_X1 U21723 ( .A1(n19723), .A2(n19609), .B1(n19713), .B2(n19606), .ZN(
        n19576) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19608), .ZN(n19575) );
  OAI211_X1 U21725 ( .C1(n19717), .C2(n19602), .A(n19576), .B(n19575), .ZN(
        P3_U2983) );
  AOI22_X1 U21726 ( .A1(n19729), .A2(n19609), .B1(n19718), .B2(n19606), .ZN(
        n19578) );
  AOI22_X1 U21727 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19608), .ZN(n19577) );
  OAI211_X1 U21728 ( .C1(n19727), .C2(n19602), .A(n19578), .B(n19577), .ZN(
        P3_U2975) );
  AOI22_X1 U21729 ( .A1(n19734), .A2(n19609), .B1(n19722), .B2(n19606), .ZN(
        n19580) );
  AOI22_X1 U21730 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19608), .ZN(n19579) );
  OAI211_X1 U21731 ( .C1(n19583), .C2(n19602), .A(n19580), .B(n19579), .ZN(
        P3_U2967) );
  AOI22_X1 U21732 ( .A1(n19728), .A2(n19606), .B1(n19746), .B2(n19607), .ZN(
        n19582) );
  AOI22_X1 U21733 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19608), .ZN(n19581) );
  OAI211_X1 U21734 ( .C1(n19583), .C2(n19605), .A(n19582), .B(n19581), .ZN(
        P3_U2959) );
  AOI22_X1 U21735 ( .A1(n19746), .A2(n19609), .B1(n19733), .B2(n19606), .ZN(
        n19585) );
  AOI22_X1 U21736 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19608), .ZN(n19584) );
  OAI211_X1 U21737 ( .C1(n19629), .C2(n19602), .A(n19585), .B(n19584), .ZN(
        P3_U2951) );
  AOI22_X1 U21738 ( .A1(n19752), .A2(n19609), .B1(n19739), .B2(n19606), .ZN(
        n19587) );
  AOI22_X1 U21739 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19608), .ZN(n19586) );
  OAI211_X1 U21740 ( .C1(n19744), .C2(n19602), .A(n19587), .B(n19586), .ZN(
        P3_U2943) );
  AOI22_X1 U21741 ( .A1(n19757), .A2(n19609), .B1(n19745), .B2(n19606), .ZN(
        n19589) );
  AOI22_X1 U21742 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19608), .ZN(n19588) );
  OAI211_X1 U21743 ( .C1(n19755), .C2(n19602), .A(n19589), .B(n19588), .ZN(
        P3_U2935) );
  AOI22_X1 U21744 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19751), .B1(
        n19750), .B2(n19606), .ZN(n19591) );
  AOI22_X1 U21745 ( .A1(n19752), .A2(n19608), .B1(n19768), .B2(n19607), .ZN(
        n19590) );
  OAI211_X1 U21746 ( .C1(n19755), .C2(n19605), .A(n19591), .B(n19590), .ZN(
        P3_U2927) );
  AOI22_X1 U21747 ( .A1(n19776), .A2(n19607), .B1(n19756), .B2(n19606), .ZN(
        n19593) );
  AOI22_X1 U21748 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19608), .ZN(n19592) );
  OAI211_X1 U21749 ( .C1(n19679), .C2(n19605), .A(n19593), .B(n19592), .ZN(
        P3_U2919) );
  AOI22_X1 U21750 ( .A1(n19776), .A2(n19609), .B1(n19761), .B2(n19606), .ZN(
        n19595) );
  AOI22_X1 U21751 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19608), .ZN(n19594) );
  OAI211_X1 U21752 ( .C1(n19772), .C2(n19602), .A(n19595), .B(n19594), .ZN(
        P3_U2911) );
  AOI22_X1 U21753 ( .A1(n19782), .A2(n19609), .B1(n19767), .B2(n19606), .ZN(
        n19597) );
  AOI22_X1 U21754 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19608), .ZN(n19596) );
  OAI211_X1 U21755 ( .C1(n19642), .C2(n19602), .A(n19597), .B(n19596), .ZN(
        P3_U2903) );
  AOI22_X1 U21756 ( .A1(n19800), .A2(n19607), .B1(n19773), .B2(n19606), .ZN(
        n19599) );
  AOI22_X1 U21757 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19774), .B1(
        n19776), .B2(n19608), .ZN(n19598) );
  OAI211_X1 U21758 ( .C1(n19642), .C2(n19605), .A(n19599), .B(n19598), .ZN(
        P3_U2895) );
  AOI22_X1 U21759 ( .A1(n19800), .A2(n19609), .B1(n19780), .B2(n19606), .ZN(
        n19601) );
  AOI22_X1 U21760 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19608), .ZN(n19600) );
  OAI211_X1 U21761 ( .C1(n19793), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P3_U2887) );
  AOI22_X1 U21762 ( .A1(n19788), .A2(n19607), .B1(n19787), .B2(n19606), .ZN(
        n19604) );
  AOI22_X1 U21763 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19608), .ZN(n19603) );
  OAI211_X1 U21764 ( .C1(n19793), .C2(n19605), .A(n19604), .B(n19603), .ZN(
        P3_U2879) );
  AOI22_X1 U21765 ( .A1(n19797), .A2(n19607), .B1(n19795), .B2(n19606), .ZN(
        n19611) );
  AOI22_X1 U21766 ( .A1(n19788), .A2(n19609), .B1(n19800), .B2(n19608), .ZN(
        n19610) );
  OAI211_X1 U21767 ( .C1(n19612), .C2(n19798), .A(n19611), .B(n19610), .ZN(
        P3_U2871) );
  OAI22_X1 U21768 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19699), .ZN(n19613) );
  INV_X1 U21769 ( .A(n19613), .ZN(U253) );
  INV_X1 U21770 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19614) );
  NOR2_X1 U21771 ( .A1(n19614), .A2(n19703), .ZN(n19650) );
  INV_X1 U21772 ( .A(n19650), .ZN(n19648) );
  NAND2_X1 U21773 ( .A1(n19704), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19645) );
  INV_X1 U21774 ( .A(n19645), .ZN(n19652) );
  AND2_X1 U21775 ( .A1(n19705), .A2(BUF2_REG_2__SCAN_IN), .ZN(n19649) );
  AOI22_X1 U21776 ( .A1(n19797), .A2(n19652), .B1(n19706), .B2(n19649), .ZN(
        n19616) );
  NOR2_X2 U21777 ( .A1(n21434), .A2(n19707), .ZN(n19651) );
  AOI22_X1 U21778 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19651), .ZN(n19615) );
  OAI211_X1 U21779 ( .C1(n19660), .C2(n19648), .A(n19616), .B(n19615), .ZN(
        P3_U2990) );
  AOI22_X1 U21780 ( .A1(n19729), .A2(n19650), .B1(n19713), .B2(n19649), .ZN(
        n19618) );
  AOI22_X1 U21781 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19651), .ZN(n19617) );
  OAI211_X1 U21782 ( .C1(n19660), .C2(n19645), .A(n19618), .B(n19617), .ZN(
        P3_U2982) );
  AOI22_X1 U21783 ( .A1(n19729), .A2(n19652), .B1(n19718), .B2(n19649), .ZN(
        n19620) );
  AOI22_X1 U21784 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19651), .ZN(n19619) );
  OAI211_X1 U21785 ( .C1(n19727), .C2(n19648), .A(n19620), .B(n19619), .ZN(
        P3_U2974) );
  AOI22_X1 U21786 ( .A1(n19740), .A2(n19650), .B1(n19722), .B2(n19649), .ZN(
        n19622) );
  AOI22_X1 U21787 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19651), .ZN(n19621) );
  OAI211_X1 U21788 ( .C1(n19727), .C2(n19645), .A(n19622), .B(n19621), .ZN(
        P3_U2966) );
  AOI22_X1 U21789 ( .A1(n19740), .A2(n19652), .B1(n19728), .B2(n19649), .ZN(
        n19624) );
  AOI22_X1 U21790 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19651), .ZN(n19623) );
  OAI211_X1 U21791 ( .C1(n19738), .C2(n19648), .A(n19624), .B(n19623), .ZN(
        P3_U2958) );
  AOI22_X1 U21792 ( .A1(n19746), .A2(n19652), .B1(n19733), .B2(n19649), .ZN(
        n19626) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19651), .ZN(n19625) );
  OAI211_X1 U21794 ( .C1(n19629), .C2(n19648), .A(n19626), .B(n19625), .ZN(
        P3_U2950) );
  AOI22_X1 U21795 ( .A1(n19739), .A2(n19649), .B1(n19757), .B2(n19650), .ZN(
        n19628) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19651), .ZN(n19627) );
  OAI211_X1 U21797 ( .C1(n19629), .C2(n19645), .A(n19628), .B(n19627), .ZN(
        P3_U2942) );
  AOI22_X1 U21798 ( .A1(n19762), .A2(n19650), .B1(n19745), .B2(n19649), .ZN(
        n19631) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19651), .ZN(n19630) );
  OAI211_X1 U21800 ( .C1(n19744), .C2(n19645), .A(n19631), .B(n19630), .ZN(
        P3_U2934) );
  AOI22_X1 U21801 ( .A1(n19762), .A2(n19652), .B1(n19750), .B2(n19649), .ZN(
        n19633) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19751), .B1(
        n19752), .B2(n19651), .ZN(n19632) );
  OAI211_X1 U21803 ( .C1(n19679), .C2(n19648), .A(n19633), .B(n19632), .ZN(
        P3_U2926) );
  AOI22_X1 U21804 ( .A1(n19768), .A2(n19652), .B1(n19756), .B2(n19649), .ZN(
        n19635) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19651), .ZN(n19634) );
  OAI211_X1 U21806 ( .C1(n19766), .C2(n19648), .A(n19635), .B(n19634), .ZN(
        P3_U2918) );
  AOI22_X1 U21807 ( .A1(n19782), .A2(n19650), .B1(n19761), .B2(n19649), .ZN(
        n19637) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19651), .ZN(n19636) );
  OAI211_X1 U21809 ( .C1(n19766), .C2(n19645), .A(n19637), .B(n19636), .ZN(
        P3_U2910) );
  AOI22_X1 U21810 ( .A1(n19782), .A2(n19652), .B1(n19767), .B2(n19649), .ZN(
        n19639) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19651), .ZN(n19638) );
  OAI211_X1 U21812 ( .C1(n19642), .C2(n19648), .A(n19639), .B(n19638), .ZN(
        P3_U2902) );
  AOI22_X1 U21813 ( .A1(n19800), .A2(n19650), .B1(n19773), .B2(n19649), .ZN(
        n19641) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19774), .B1(
        n19776), .B2(n19651), .ZN(n19640) );
  OAI211_X1 U21815 ( .C1(n19642), .C2(n19645), .A(n19641), .B(n19640), .ZN(
        P3_U2894) );
  AOI22_X1 U21816 ( .A1(n19781), .A2(n19650), .B1(n19780), .B2(n19649), .ZN(
        n19644) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19651), .ZN(n19643) );
  OAI211_X1 U21818 ( .C1(n19786), .C2(n19645), .A(n19644), .B(n19643), .ZN(
        P3_U2886) );
  AOI22_X1 U21819 ( .A1(n19781), .A2(n19652), .B1(n19787), .B2(n19649), .ZN(
        n19647) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19651), .ZN(n19646) );
  OAI211_X1 U21821 ( .C1(n19805), .C2(n19648), .A(n19647), .B(n19646), .ZN(
        P3_U2878) );
  AOI22_X1 U21822 ( .A1(n19797), .A2(n19650), .B1(n19795), .B2(n19649), .ZN(
        n19654) );
  AOI22_X1 U21823 ( .A1(n19788), .A2(n19652), .B1(n19800), .B2(n19651), .ZN(
        n19653) );
  OAI211_X1 U21824 ( .C1(n19655), .C2(n19798), .A(n19654), .B(n19653), .ZN(
        P3_U2870) );
  OAI22_X1 U21825 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19699), .ZN(n19656) );
  INV_X1 U21826 ( .A(n19656), .ZN(U252) );
  INV_X1 U21827 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n21298) );
  NOR2_X1 U21828 ( .A1(n21298), .A2(n19703), .ZN(n19693) );
  INV_X1 U21829 ( .A(n19693), .ZN(n19691) );
  NAND2_X1 U21830 ( .A1(n19704), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19688) );
  INV_X1 U21831 ( .A(n19688), .ZN(n19695) );
  AND2_X1 U21832 ( .A1(n19705), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19692) );
  AOI22_X1 U21833 ( .A1(n19797), .A2(n19695), .B1(n19706), .B2(n19692), .ZN(
        n19659) );
  NOR2_X2 U21834 ( .A1(n19657), .A2(n19707), .ZN(n19694) );
  AOI22_X1 U21835 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19694), .ZN(n19658) );
  OAI211_X1 U21836 ( .C1(n19660), .C2(n19691), .A(n19659), .B(n19658), .ZN(
        P3_U2989) );
  AOI22_X1 U21837 ( .A1(n19723), .A2(n19695), .B1(n19713), .B2(n19692), .ZN(
        n19662) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19694), .ZN(n19661) );
  OAI211_X1 U21839 ( .C1(n19717), .C2(n19691), .A(n19662), .B(n19661), .ZN(
        P3_U2981) );
  AOI22_X1 U21840 ( .A1(n19734), .A2(n19693), .B1(n19718), .B2(n19692), .ZN(
        n19664) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19694), .ZN(n19663) );
  OAI211_X1 U21842 ( .C1(n19717), .C2(n19688), .A(n19664), .B(n19663), .ZN(
        P3_U2973) );
  AOI22_X1 U21843 ( .A1(n19740), .A2(n19693), .B1(n19722), .B2(n19692), .ZN(
        n19666) );
  AOI22_X1 U21844 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19694), .ZN(n19665) );
  OAI211_X1 U21845 ( .C1(n19727), .C2(n19688), .A(n19666), .B(n19665), .ZN(
        P3_U2965) );
  AOI22_X1 U21846 ( .A1(n19740), .A2(n19695), .B1(n19728), .B2(n19692), .ZN(
        n19668) );
  AOI22_X1 U21847 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19694), .ZN(n19667) );
  OAI211_X1 U21848 ( .C1(n19738), .C2(n19691), .A(n19668), .B(n19667), .ZN(
        P3_U2957) );
  AOI22_X1 U21849 ( .A1(n19752), .A2(n19693), .B1(n19733), .B2(n19692), .ZN(
        n19670) );
  AOI22_X1 U21850 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19694), .ZN(n19669) );
  OAI211_X1 U21851 ( .C1(n19738), .C2(n19688), .A(n19670), .B(n19669), .ZN(
        P3_U2949) );
  AOI22_X1 U21852 ( .A1(n19752), .A2(n19695), .B1(n19739), .B2(n19692), .ZN(
        n19672) );
  AOI22_X1 U21853 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19694), .ZN(n19671) );
  OAI211_X1 U21854 ( .C1(n19744), .C2(n19691), .A(n19672), .B(n19671), .ZN(
        P3_U2941) );
  AOI22_X1 U21855 ( .A1(n19762), .A2(n19693), .B1(n19745), .B2(n19692), .ZN(
        n19674) );
  AOI22_X1 U21856 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19694), .ZN(n19673) );
  OAI211_X1 U21857 ( .C1(n19744), .C2(n19688), .A(n19674), .B(n19673), .ZN(
        P3_U2933) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19751), .B1(
        n19750), .B2(n19692), .ZN(n19676) );
  AOI22_X1 U21859 ( .A1(n19752), .A2(n19694), .B1(n19768), .B2(n19693), .ZN(
        n19675) );
  OAI211_X1 U21860 ( .C1(n19755), .C2(n19688), .A(n19676), .B(n19675), .ZN(
        P3_U2925) );
  AOI22_X1 U21861 ( .A1(n19776), .A2(n19693), .B1(n19756), .B2(n19692), .ZN(
        n19678) );
  AOI22_X1 U21862 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19694), .ZN(n19677) );
  OAI211_X1 U21863 ( .C1(n19679), .C2(n19688), .A(n19678), .B(n19677), .ZN(
        P3_U2917) );
  AOI22_X1 U21864 ( .A1(n19776), .A2(n19695), .B1(n19761), .B2(n19692), .ZN(
        n19681) );
  AOI22_X1 U21865 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19694), .ZN(n19680) );
  OAI211_X1 U21866 ( .C1(n19772), .C2(n19691), .A(n19681), .B(n19680), .ZN(
        P3_U2909) );
  AOI22_X1 U21867 ( .A1(n19789), .A2(n19693), .B1(n19767), .B2(n19692), .ZN(
        n19683) );
  AOI22_X1 U21868 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19694), .ZN(n19682) );
  OAI211_X1 U21869 ( .C1(n19772), .C2(n19688), .A(n19683), .B(n19682), .ZN(
        P3_U2901) );
  AOI22_X1 U21870 ( .A1(n19789), .A2(n19695), .B1(n19773), .B2(n19692), .ZN(
        n19685) );
  AOI22_X1 U21871 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19774), .B1(
        n19776), .B2(n19694), .ZN(n19684) );
  OAI211_X1 U21872 ( .C1(n19786), .C2(n19691), .A(n19685), .B(n19684), .ZN(
        P3_U2893) );
  AOI22_X1 U21873 ( .A1(n19781), .A2(n19693), .B1(n19780), .B2(n19692), .ZN(
        n19687) );
  AOI22_X1 U21874 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19694), .ZN(n19686) );
  OAI211_X1 U21875 ( .C1(n19786), .C2(n19688), .A(n19687), .B(n19686), .ZN(
        P3_U2885) );
  AOI22_X1 U21876 ( .A1(n19781), .A2(n19695), .B1(n19787), .B2(n19692), .ZN(
        n19690) );
  AOI22_X1 U21877 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19694), .ZN(n19689) );
  OAI211_X1 U21878 ( .C1(n19805), .C2(n19691), .A(n19690), .B(n19689), .ZN(
        P3_U2877) );
  AOI22_X1 U21879 ( .A1(n19797), .A2(n19693), .B1(n19795), .B2(n19692), .ZN(
        n19697) );
  AOI22_X1 U21880 ( .A1(n19788), .A2(n19695), .B1(n19800), .B2(n19694), .ZN(
        n19696) );
  OAI211_X1 U21881 ( .C1(n19698), .C2(n19798), .A(n19697), .B(n19696), .ZN(
        P3_U2869) );
  OAI22_X1 U21882 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19699), .ZN(n19701) );
  INV_X1 U21883 ( .A(n19701), .ZN(U251) );
  INV_X1 U21884 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19702) );
  NOR2_X1 U21885 ( .A1(n19703), .A2(n19702), .ZN(n19775) );
  INV_X1 U21886 ( .A(n19775), .ZN(n19804) );
  NAND2_X1 U21887 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19704), .ZN(n19779) );
  INV_X1 U21888 ( .A(n19779), .ZN(n19796) );
  AND2_X1 U21889 ( .A1(n19705), .A2(BUF2_REG_0__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U21890 ( .A1(n19723), .A2(n19796), .B1(n19706), .B2(n19794), .ZN(
        n19711) );
  NOR2_X2 U21891 ( .A1(n19708), .A2(n19707), .ZN(n19799) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19709), .B1(
        n19781), .B2(n19799), .ZN(n19710) );
  OAI211_X1 U21893 ( .C1(n19712), .C2(n19804), .A(n19711), .B(n19710), .ZN(
        P3_U2988) );
  AOI22_X1 U21894 ( .A1(n19723), .A2(n19775), .B1(n19713), .B2(n19794), .ZN(
        n19716) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19714), .B1(
        n19788), .B2(n19799), .ZN(n19715) );
  OAI211_X1 U21896 ( .C1(n19717), .C2(n19779), .A(n19716), .B(n19715), .ZN(
        P3_U2980) );
  AOI22_X1 U21897 ( .A1(n19729), .A2(n19775), .B1(n19718), .B2(n19794), .ZN(
        n19721) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19719), .B1(
        n19797), .B2(n19799), .ZN(n19720) );
  OAI211_X1 U21899 ( .C1(n19727), .C2(n19779), .A(n19721), .B(n19720), .ZN(
        P3_U2972) );
  AOI22_X1 U21900 ( .A1(n19740), .A2(n19796), .B1(n19722), .B2(n19794), .ZN(
        n19726) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19724), .B1(
        n19723), .B2(n19799), .ZN(n19725) );
  OAI211_X1 U21902 ( .C1(n19727), .C2(n19804), .A(n19726), .B(n19725), .ZN(
        P3_U2964) );
  AOI22_X1 U21903 ( .A1(n19740), .A2(n19775), .B1(n19728), .B2(n19794), .ZN(
        n19732) );
  AOI22_X1 U21904 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19730), .B1(
        n19729), .B2(n19799), .ZN(n19731) );
  OAI211_X1 U21905 ( .C1(n19738), .C2(n19779), .A(n19732), .B(n19731), .ZN(
        P3_U2956) );
  AOI22_X1 U21906 ( .A1(n19752), .A2(n19796), .B1(n19733), .B2(n19794), .ZN(
        n19737) );
  AOI22_X1 U21907 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19735), .B1(
        n19734), .B2(n19799), .ZN(n19736) );
  OAI211_X1 U21908 ( .C1(n19738), .C2(n19804), .A(n19737), .B(n19736), .ZN(
        P3_U2948) );
  AOI22_X1 U21909 ( .A1(n19752), .A2(n19775), .B1(n19739), .B2(n19794), .ZN(
        n19743) );
  AOI22_X1 U21910 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19741), .B1(
        n19740), .B2(n19799), .ZN(n19742) );
  OAI211_X1 U21911 ( .C1(n19744), .C2(n19779), .A(n19743), .B(n19742), .ZN(
        P3_U2940) );
  AOI22_X1 U21912 ( .A1(n19757), .A2(n19775), .B1(n19745), .B2(n19794), .ZN(
        n19749) );
  AOI22_X1 U21913 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19799), .ZN(n19748) );
  OAI211_X1 U21914 ( .C1(n19755), .C2(n19779), .A(n19749), .B(n19748), .ZN(
        P3_U2932) );
  AOI22_X1 U21915 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19751), .B1(
        n19750), .B2(n19794), .ZN(n19754) );
  AOI22_X1 U21916 ( .A1(n19752), .A2(n19799), .B1(n19768), .B2(n19796), .ZN(
        n19753) );
  OAI211_X1 U21917 ( .C1(n19755), .C2(n19804), .A(n19754), .B(n19753), .ZN(
        P3_U2924) );
  AOI22_X1 U21918 ( .A1(n19768), .A2(n19775), .B1(n19756), .B2(n19794), .ZN(
        n19760) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19758), .B1(
        n19757), .B2(n19799), .ZN(n19759) );
  OAI211_X1 U21920 ( .C1(n19766), .C2(n19779), .A(n19760), .B(n19759), .ZN(
        P3_U2916) );
  AOI22_X1 U21921 ( .A1(n19782), .A2(n19796), .B1(n19761), .B2(n19794), .ZN(
        n19765) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19763), .B1(
        n19762), .B2(n19799), .ZN(n19764) );
  OAI211_X1 U21923 ( .C1(n19766), .C2(n19804), .A(n19765), .B(n19764), .ZN(
        P3_U2908) );
  AOI22_X1 U21924 ( .A1(n19789), .A2(n19796), .B1(n19767), .B2(n19794), .ZN(
        n19771) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19769), .B1(
        n19768), .B2(n19799), .ZN(n19770) );
  OAI211_X1 U21926 ( .C1(n19772), .C2(n19804), .A(n19771), .B(n19770), .ZN(
        P3_U2900) );
  AOI22_X1 U21927 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19774), .B1(
        n19773), .B2(n19794), .ZN(n19778) );
  AOI22_X1 U21928 ( .A1(n19776), .A2(n19799), .B1(n19789), .B2(n19775), .ZN(
        n19777) );
  OAI211_X1 U21929 ( .C1(n19786), .C2(n19779), .A(n19778), .B(n19777), .ZN(
        P3_U2892) );
  AOI22_X1 U21930 ( .A1(n19781), .A2(n19796), .B1(n19780), .B2(n19794), .ZN(
        n19785) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19783), .B1(
        n19782), .B2(n19799), .ZN(n19784) );
  OAI211_X1 U21932 ( .C1(n19786), .C2(n19804), .A(n19785), .B(n19784), .ZN(
        P3_U2884) );
  AOI22_X1 U21933 ( .A1(n19788), .A2(n19796), .B1(n19787), .B2(n19794), .ZN(
        n19792) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19790), .B1(
        n19789), .B2(n19799), .ZN(n19791) );
  OAI211_X1 U21935 ( .C1(n19793), .C2(n19804), .A(n19792), .B(n19791), .ZN(
        P3_U2876) );
  AOI22_X1 U21936 ( .A1(n19797), .A2(n19796), .B1(n19795), .B2(n19794), .ZN(
        n19803) );
  INV_X1 U21937 ( .A(n19798), .ZN(n19801) );
  AOI22_X1 U21938 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19801), .B1(
        n19800), .B2(n19799), .ZN(n19802) );
  OAI211_X1 U21939 ( .C1(n19805), .C2(n19804), .A(n19803), .B(n19802), .ZN(
        P3_U2868) );
  AOI22_X1 U21940 ( .A1(n20064), .A2(n19806), .B1(n20111), .B2(
        P2_EAX_REG_14__SCAN_IN), .ZN(n19807) );
  OAI21_X1 U21941 ( .B1(n20071), .B2(n19808), .A(n19807), .ZN(P2_U2905) );
  AOI22_X1 U21942 ( .A1(n20064), .A2(n19809), .B1(n20111), .B2(
        P2_EAX_REG_12__SCAN_IN), .ZN(n19810) );
  OAI21_X1 U21943 ( .B1(n20071), .B2(n19811), .A(n19810), .ZN(P2_U2907) );
  AOI22_X1 U21944 ( .A1(n20064), .A2(n19812), .B1(n20111), .B2(
        P2_EAX_REG_10__SCAN_IN), .ZN(n19813) );
  OAI21_X1 U21945 ( .B1(n20071), .B2(n19814), .A(n19813), .ZN(P2_U2909) );
  AOI22_X1 U21946 ( .A1(n20064), .A2(n19815), .B1(n20111), .B2(
        P2_EAX_REG_9__SCAN_IN), .ZN(n19816) );
  OAI21_X1 U21947 ( .B1(n20071), .B2(n19817), .A(n19816), .ZN(P2_U2910) );
  NOR2_X2 U21948 ( .A1(n12011), .A2(n20293), .ZN(n20002) );
  AOI22_X1 U21949 ( .A1(n20296), .A2(n19819), .B1(n20295), .B2(n20002), .ZN(
        n19823) );
  INV_X1 U21950 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20681) );
  INV_X1 U21951 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n21340) );
  OAI22_X1 U21952 ( .A1(n20681), .A2(n19821), .B1(n21340), .B2(n19820), .ZN(
        n19981) );
  AOI22_X1 U21953 ( .A1(n20285), .A2(n19981), .B1(n20299), .B2(n20003), .ZN(
        n19822) );
  OAI211_X1 U21954 ( .C1(n20210), .C2(n19824), .A(n19823), .B(n19822), .ZN(
        P2_U3175) );
  INV_X1 U21955 ( .A(n19981), .ZN(n20017) );
  NOR2_X1 U21956 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19826), .ZN(
        n20303) );
  AOI22_X1 U21957 ( .A1(n20003), .A2(n20304), .B1(n20002), .B2(n20303), .ZN(
        n19835) );
  AOI21_X1 U21958 ( .B1(n20316), .B2(n20309), .A(n19841), .ZN(n19827) );
  NOR2_X1 U21959 ( .A1(n19827), .A2(n15037), .ZN(n19831) );
  NAND3_X1 U21960 ( .A1(n19985), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19851) );
  NOR2_X1 U21961 ( .A1(n19987), .A2(n19851), .ZN(n20310) );
  INV_X1 U21962 ( .A(n20310), .ZN(n19840) );
  INV_X1 U21963 ( .A(n19962), .ZN(n20006) );
  AOI21_X1 U21964 ( .B1(n11145), .B2(n20006), .A(n20005), .ZN(n19829) );
  AOI21_X1 U21965 ( .B1(n19831), .B2(n19840), .A(n19829), .ZN(n19830) );
  OAI21_X1 U21966 ( .B1(n20303), .B2(n20310), .A(n19831), .ZN(n19833) );
  OAI21_X1 U21967 ( .B1(n11145), .B2(n20303), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19832) );
  NAND2_X1 U21968 ( .A1(n19833), .A2(n19832), .ZN(n20305) );
  AOI22_X1 U21969 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20306), .B1(
        n19819), .B2(n20305), .ZN(n19834) );
  OAI211_X1 U21970 ( .C1(n20017), .C2(n20309), .A(n19835), .B(n19834), .ZN(
        P2_U3167) );
  OAI21_X1 U21971 ( .B1(n19838), .B2(n20310), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19837) );
  OAI21_X1 U21972 ( .B1(n19851), .B2(n15037), .A(n19837), .ZN(n20311) );
  AOI22_X1 U21973 ( .A1(n20311), .A2(n19819), .B1(n20002), .B2(n20310), .ZN(
        n19847) );
  NOR2_X1 U21974 ( .A1(n20310), .A2(n19838), .ZN(n19839) );
  AOI211_X1 U21975 ( .C1(n19962), .C2(n19840), .A(n20291), .B(n19839), .ZN(
        n19845) );
  OR2_X1 U21976 ( .A1(n19842), .A2(n19841), .ZN(n19990) );
  OAI21_X1 U21977 ( .B1(n19843), .B2(n19990), .A(n19851), .ZN(n19844) );
  OAI21_X1 U21978 ( .B1(n19845), .B2(n20005), .A(n19844), .ZN(n20313) );
  AOI22_X1 U21979 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20313), .B1(
        n20304), .B2(n19981), .ZN(n19846) );
  OAI211_X1 U21980 ( .C1(n19984), .C2(n20323), .A(n19847), .B(n19846), .ZN(
        P2_U3159) );
  INV_X1 U21981 ( .A(n19848), .ZN(n19854) );
  INV_X1 U21982 ( .A(n19849), .ZN(n19850) );
  NAND2_X1 U21983 ( .A1(n19850), .A2(n19972), .ZN(n19945) );
  NOR2_X1 U21984 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19851), .ZN(
        n20317) );
  OAI21_X1 U21985 ( .B1(n19852), .B2(n20317), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19853) );
  OAI21_X1 U21986 ( .B1(n19854), .B2(n19945), .A(n19853), .ZN(n20318) );
  AOI22_X1 U21987 ( .A1(n20318), .A2(n19819), .B1(n20002), .B2(n20317), .ZN(
        n19861) );
  OAI21_X1 U21988 ( .B1(n20319), .B2(n20312), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19856) );
  OAI21_X1 U21989 ( .B1(n19945), .B2(n19898), .A(n19856), .ZN(n19859) );
  INV_X1 U21990 ( .A(n20317), .ZN(n19857) );
  OAI211_X1 U21991 ( .C1(n12182), .C2(n19962), .A(n19857), .B(n15037), .ZN(
        n19858) );
  NAND3_X1 U21992 ( .A1(n19859), .A2(n19858), .A3(n20009), .ZN(n20320) );
  AOI22_X1 U21993 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n20003), .B2(n20319), .ZN(n19860) );
  OAI211_X1 U21994 ( .C1(n20017), .C2(n20323), .A(n19861), .B(n19860), .ZN(
        P2_U3151) );
  NAND3_X1 U21995 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19871), .ZN(n19872) );
  INV_X1 U21996 ( .A(n12174), .ZN(n19863) );
  NOR2_X1 U21997 ( .A1(n19987), .A2(n19872), .ZN(n20324) );
  OAI21_X1 U21998 ( .B1(n19863), .B2(n20324), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19862) );
  OAI21_X1 U21999 ( .B1(n19872), .B2(n15037), .A(n19862), .ZN(n20325) );
  AOI22_X1 U22000 ( .A1(n20325), .A2(n19819), .B1(n20002), .B2(n20324), .ZN(
        n19868) );
  AOI211_X1 U22001 ( .C1(n19863), .C2(n20006), .A(n19992), .B(n20324), .ZN(
        n19864) );
  NOR2_X1 U22002 ( .A1(n20291), .A2(n19864), .ZN(n19866) );
  OAI21_X1 U22003 ( .B1(n19941), .B2(n19959), .A(n19872), .ZN(n19865) );
  NAND2_X1 U22004 ( .A1(n19866), .A2(n19865), .ZN(n20326) );
  AOI22_X1 U22005 ( .A1(n20003), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n19867) );
  OAI211_X1 U22006 ( .C1(n20017), .C2(n20329), .A(n19868), .B(n19867), .ZN(
        P2_U3143) );
  INV_X1 U22007 ( .A(n20331), .ZN(n19869) );
  NAND2_X1 U22008 ( .A1(n20262), .A2(n19869), .ZN(n19870) );
  AOI21_X1 U22009 ( .B1(n19870), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n15037), 
        .ZN(n19877) );
  NAND3_X1 U22010 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19985), .A3(
        n19871), .ZN(n19895) );
  NOR2_X1 U22011 ( .A1(n19987), .A2(n19895), .ZN(n20337) );
  NOR2_X1 U22012 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19872), .ZN(
        n20330) );
  NOR2_X1 U22013 ( .A1(n20337), .A2(n20330), .ZN(n19880) );
  INV_X1 U22014 ( .A(n20005), .ZN(n19876) );
  NOR2_X1 U22015 ( .A1(n19873), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22016 ( .B1(n19874), .B2(n20330), .A(n20009), .ZN(n19875) );
  INV_X1 U22017 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U22018 ( .A1(n20331), .A2(n19981), .B1(n20002), .B2(n20330), .ZN(
        n19883) );
  INV_X1 U22019 ( .A(n19877), .ZN(n19881) );
  OAI21_X1 U22020 ( .B1(n19878), .B2(n20330), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19879) );
  AOI22_X1 U22021 ( .A1(n19819), .A2(n20332), .B1(n20338), .B2(n20003), .ZN(
        n19882) );
  OAI211_X1 U22022 ( .C1(n20336), .C2(n19884), .A(n19883), .B(n19882), .ZN(
        P2_U3135) );
  AOI22_X1 U22023 ( .A1(n20338), .A2(n19981), .B1(n20337), .B2(n20002), .ZN(
        n19894) );
  OAI21_X1 U22024 ( .B1(n19885), .B2(n19990), .A(n19992), .ZN(n19892) );
  INV_X1 U22025 ( .A(n19895), .ZN(n19889) );
  INV_X1 U22026 ( .A(n20337), .ZN(n19887) );
  INV_X1 U22027 ( .A(n12177), .ZN(n19890) );
  NOR2_X1 U22028 ( .A1(n20337), .A2(n19890), .ZN(n19886) );
  AOI211_X1 U22029 ( .C1(n19962), .C2(n19887), .A(n20291), .B(n19886), .ZN(
        n19888) );
  OAI22_X1 U22030 ( .A1(n19892), .A2(n19889), .B1(n20005), .B2(n19888), .ZN(
        n20340) );
  OAI21_X1 U22031 ( .B1(n19890), .B2(n20337), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19891) );
  AOI22_X1 U22032 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20340), .B1(
        n19819), .B2(n20339), .ZN(n19893) );
  OAI211_X1 U22033 ( .C1(n19984), .C2(n20343), .A(n19894), .B(n19893), .ZN(
        P2_U3127) );
  NOR2_X1 U22034 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19895), .ZN(
        n20344) );
  AOI22_X1 U22035 ( .A1(n20345), .A2(n19981), .B1(n20002), .B2(n20344), .ZN(
        n19908) );
  INV_X1 U22036 ( .A(n20356), .ZN(n19896) );
  NOR2_X1 U22037 ( .A1(n20345), .A2(n19896), .ZN(n19897) );
  OAI21_X1 U22038 ( .B1(n19897), .B2(n19841), .A(n19992), .ZN(n19906) );
  NAND2_X1 U22039 ( .A1(n19898), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19943) );
  NOR2_X1 U22040 ( .A1(n19958), .A2(n19943), .ZN(n20350) );
  NOR2_X1 U22041 ( .A1(n20344), .A2(n20350), .ZN(n19904) );
  INV_X1 U22042 ( .A(n19904), .ZN(n19901) );
  INV_X1 U22043 ( .A(n20344), .ZN(n19899) );
  OAI211_X1 U22044 ( .C1(n12181), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n15037), 
        .B(n19899), .ZN(n19900) );
  OAI211_X1 U22045 ( .C1(n19906), .C2(n19901), .A(n20009), .B(n19900), .ZN(
        n20347) );
  OAI21_X1 U22046 ( .B1(n19902), .B2(n20344), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19905) );
  AOI22_X1 U22047 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20347), .B1(
        n19819), .B2(n20346), .ZN(n19907) );
  OAI211_X1 U22048 ( .C1(n19984), .C2(n20356), .A(n19908), .B(n19907), .ZN(
        P2_U3119) );
  OR2_X1 U22049 ( .A1(n19985), .A2(n19943), .ZN(n19918) );
  OAI21_X1 U22050 ( .B1(n19911), .B2(n20350), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19909) );
  OAI21_X1 U22051 ( .B1(n19918), .B2(n15037), .A(n19909), .ZN(n20351) );
  AOI22_X1 U22052 ( .A1(n20351), .A2(n19819), .B1(n20350), .B2(n20002), .ZN(
        n19917) );
  OAI21_X1 U22053 ( .B1(n19910), .B2(n19841), .A(n19918), .ZN(n19915) );
  INV_X1 U22054 ( .A(n19911), .ZN(n19913) );
  INV_X1 U22055 ( .A(n20350), .ZN(n19912) );
  OAI211_X1 U22056 ( .C1(n19913), .C2(n19962), .A(n15037), .B(n19912), .ZN(
        n19914) );
  NAND3_X1 U22057 ( .A1(n19915), .A2(n20009), .A3(n19914), .ZN(n20353) );
  AOI22_X1 U22058 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20003), .ZN(n19916) );
  OAI211_X1 U22059 ( .C1(n20017), .C2(n20356), .A(n19917), .B(n19916), .ZN(
        P2_U3111) );
  OR2_X1 U22060 ( .A1(n19972), .A2(n19943), .ZN(n19921) );
  NOR2_X1 U22061 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19918), .ZN(
        n20357) );
  OAI21_X1 U22062 ( .B1(n12189), .B2(n20357), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19919) );
  OAI21_X1 U22063 ( .B1(n15037), .B2(n19921), .A(n19919), .ZN(n20358) );
  AOI22_X1 U22064 ( .A1(n20358), .A2(n19819), .B1(n20002), .B2(n20357), .ZN(
        n19926) );
  AOI211_X1 U22065 ( .C1(n12189), .C2(n20006), .A(n19992), .B(n20357), .ZN(
        n19924) );
  OAI221_X1 U22066 ( .B1(n19841), .B2(n20369), .C1(n19841), .C2(n20363), .A(
        n19921), .ZN(n19922) );
  NAND2_X1 U22067 ( .A1(n20009), .A2(n19922), .ZN(n19923) );
  AOI22_X1 U22068 ( .A1(n20003), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n20359), .ZN(n19925) );
  OAI211_X1 U22069 ( .C1(n20017), .C2(n20363), .A(n19926), .B(n19925), .ZN(
        P2_U3103) );
  NOR2_X1 U22070 ( .A1(n19943), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19934) );
  INV_X1 U22071 ( .A(n19934), .ZN(n19936) );
  NOR2_X1 U22072 ( .A1(n19987), .A2(n19936), .ZN(n20364) );
  AOI22_X1 U22073 ( .A1(n20360), .A2(n19981), .B1(n20002), .B2(n20364), .ZN(
        n19939) );
  OAI21_X1 U22074 ( .B1(n19929), .B2(n19990), .A(n19992), .ZN(n19937) );
  INV_X1 U22075 ( .A(n19930), .ZN(n19932) );
  OAI21_X1 U22076 ( .B1(n19992), .B2(n20364), .A(n20009), .ZN(n19931) );
  OAI21_X1 U22077 ( .B1(n19932), .B2(n19962), .A(n19931), .ZN(n19933) );
  OAI21_X1 U22078 ( .B1(n19937), .B2(n19934), .A(n19933), .ZN(n20366) );
  OAI21_X1 U22079 ( .B1(n19930), .B2(n20364), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19935) );
  OAI21_X1 U22080 ( .B1(n19937), .B2(n19936), .A(n19935), .ZN(n20365) );
  AOI22_X1 U22081 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20366), .B1(
        n19819), .B2(n20365), .ZN(n19938) );
  OAI211_X1 U22082 ( .C1(n19984), .C2(n20232), .A(n19939), .B(n19938), .ZN(
        P2_U3095) );
  NOR3_X2 U22083 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19943), .ZN(n20370) );
  AOI22_X1 U22084 ( .A1(n20371), .A2(n19981), .B1(n20002), .B2(n20370), .ZN(
        n19955) );
  NOR2_X1 U22085 ( .A1(n20371), .A2(n20273), .ZN(n19944) );
  OAI21_X1 U22086 ( .B1(n19944), .B2(n19841), .A(n19992), .ZN(n19953) );
  NOR2_X1 U22087 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19945), .ZN(
        n19949) );
  INV_X1 U22088 ( .A(n19950), .ZN(n19947) );
  INV_X1 U22089 ( .A(n20370), .ZN(n19946) );
  OAI211_X1 U22090 ( .C1(n19947), .C2(n19962), .A(n19946), .B(n15037), .ZN(
        n19948) );
  OAI211_X1 U22091 ( .C1(n19953), .C2(n19949), .A(n20009), .B(n19948), .ZN(
        n20373) );
  INV_X1 U22092 ( .A(n19949), .ZN(n19952) );
  OAI21_X1 U22093 ( .B1(n19950), .B2(n20370), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19951) );
  AOI22_X1 U22094 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20373), .B1(
        n19819), .B2(n20372), .ZN(n19954) );
  OAI211_X1 U22095 ( .C1(n19984), .C2(n20381), .A(n19955), .B(n19954), .ZN(
        P2_U3087) );
  INV_X1 U22096 ( .A(n19956), .ZN(n19957) );
  NOR2_X1 U22097 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19986) );
  INV_X1 U22098 ( .A(n19986), .ZN(n20001) );
  NOR2_X1 U22099 ( .A1(n19958), .A2(n20001), .ZN(n20376) );
  AOI22_X1 U22100 ( .A1(n20273), .A2(n19981), .B1(n20002), .B2(n20376), .ZN(
        n19970) );
  OAI21_X1 U22101 ( .B1(n19960), .B2(n19959), .A(n19992), .ZN(n19968) );
  NAND2_X1 U22102 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19986), .ZN(
        n19967) );
  INV_X1 U22103 ( .A(n19967), .ZN(n19965) );
  INV_X1 U22104 ( .A(n12187), .ZN(n19963) );
  OAI21_X1 U22105 ( .B1(n19992), .B2(n20376), .A(n20009), .ZN(n19961) );
  OAI21_X1 U22106 ( .B1(n19963), .B2(n19962), .A(n19961), .ZN(n19964) );
  OAI21_X1 U22107 ( .B1(n19968), .B2(n19965), .A(n19964), .ZN(n20378) );
  OAI21_X1 U22108 ( .B1(n12187), .B2(n20376), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19966) );
  OAI21_X1 U22109 ( .B1(n19968), .B2(n19967), .A(n19966), .ZN(n20377) );
  AOI22_X1 U22110 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20378), .B1(
        n19819), .B2(n20377), .ZN(n19969) );
  OAI211_X1 U22111 ( .C1(n19984), .C2(n20276), .A(n19970), .B(n19969), .ZN(
        P2_U3079) );
  NOR3_X2 U22112 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19985), .A3(
        n20001), .ZN(n20382) );
  OAI21_X1 U22113 ( .B1(n19976), .B2(n20382), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19974) );
  INV_X1 U22114 ( .A(n19972), .ZN(n19973) );
  NAND3_X1 U22115 ( .A1(n19973), .A2(n19992), .A3(n19986), .ZN(n19977) );
  NAND2_X1 U22116 ( .A1(n19974), .A2(n19977), .ZN(n20383) );
  AOI22_X1 U22117 ( .A1(n20383), .A2(n19819), .B1(n20002), .B2(n20382), .ZN(
        n19983) );
  AOI211_X1 U22118 ( .C1(n20394), .C2(n20276), .A(n15037), .B(n19841), .ZN(
        n19980) );
  AOI21_X1 U22119 ( .B1(n19976), .B2(n19975), .A(n20382), .ZN(n19978) );
  OAI21_X1 U22120 ( .B1(n19978), .B2(n19992), .A(n19977), .ZN(n19979) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n19981), .ZN(n19982) );
  OAI211_X1 U22122 ( .C1(n19984), .C2(n20394), .A(n19983), .B(n19982), .ZN(
        P2_U3071) );
  NAND2_X1 U22123 ( .A1(n19986), .A2(n19985), .ZN(n19989) );
  NOR2_X1 U22124 ( .A1(n19987), .A2(n19989), .ZN(n20388) );
  OAI21_X1 U22125 ( .B1(n19993), .B2(n20388), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19988) );
  OAI21_X1 U22126 ( .B1(n19989), .B2(n15037), .A(n19988), .ZN(n20389) );
  AOI22_X1 U22127 ( .A1(n20389), .A2(n19819), .B1(n20002), .B2(n20388), .ZN(
        n20000) );
  INV_X1 U22128 ( .A(n19998), .ZN(n19991) );
  OAI21_X1 U22129 ( .B1(n19991), .B2(n19990), .A(n19989), .ZN(n19996) );
  AOI211_X1 U22130 ( .C1(n19993), .C2(n20006), .A(n19992), .B(n20388), .ZN(
        n19994) );
  NOR2_X1 U22131 ( .A1(n20291), .A2(n19994), .ZN(n19995) );
  NAND2_X1 U22132 ( .A1(n19996), .A2(n19995), .ZN(n20391) );
  AOI22_X1 U22133 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n20003), .B2(n20398), .ZN(n19999) );
  OAI211_X1 U22134 ( .C1(n20017), .C2(n20394), .A(n20000), .B(n19999), .ZN(
        P2_U3063) );
  NOR3_X2 U22135 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n20001), .ZN(n20397) );
  AOI22_X1 U22136 ( .A1(n20003), .A2(n20285), .B1(n20002), .B2(n20397), .ZN(
        n20016) );
  AOI21_X1 U22137 ( .B1(n20405), .B2(n20289), .A(n19841), .ZN(n20004) );
  NOR2_X1 U22138 ( .A1(n20004), .A2(n15037), .ZN(n20011) );
  AOI21_X1 U22139 ( .B1(n20012), .B2(n20006), .A(n20005), .ZN(n20007) );
  AOI21_X1 U22140 ( .B1(n20011), .B2(n20008), .A(n20007), .ZN(n20010) );
  OAI21_X1 U22141 ( .B1(n20295), .B2(n20397), .A(n20011), .ZN(n20014) );
  OAI21_X1 U22142 ( .B1(n20012), .B2(n20397), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20013) );
  NAND2_X1 U22143 ( .A1(n20014), .A2(n20013), .ZN(n20401) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n19819), .ZN(n20015) );
  OAI211_X1 U22145 ( .C1(n20017), .C2(n20289), .A(n20016), .B(n20015), .ZN(
        P2_U3055) );
  INV_X1 U22146 ( .A(n20024), .ZN(n20018) );
  AOI22_X1 U22147 ( .A1(n20113), .A2(n20018), .B1(n20111), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n20023) );
  AOI22_X1 U22148 ( .A1(n20115), .A2(BUF1_REG_22__SCAN_IN), .B1(n20114), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n20022) );
  AOI22_X1 U22149 ( .A1(n20020), .A2(n20119), .B1(n20117), .B2(n20019), .ZN(
        n20021) );
  NAND3_X1 U22150 ( .A1(n20023), .A2(n20022), .A3(n20021), .ZN(P2_U2897) );
  NOR2_X2 U22151 ( .A1(n12013), .A2(n20293), .ZN(n20058) );
  AOI22_X1 U22152 ( .A1(n20296), .A2(n20025), .B1(n20295), .B2(n20058), .ZN(
        n20027) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20300), .B1(
        n20285), .B2(n20052), .ZN(n20026) );
  OAI211_X1 U22154 ( .C1(n20055), .C2(n20309), .A(n20027), .B(n20026), .ZN(
        P2_U3174) );
  AOI22_X1 U22155 ( .A1(n20052), .A2(n20299), .B1(n20058), .B2(n20303), .ZN(
        n20029) );
  AOI22_X1 U22156 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20306), .B1(
        n20025), .B2(n20305), .ZN(n20028) );
  OAI211_X1 U22157 ( .C1(n20055), .C2(n20316), .A(n20029), .B(n20028), .ZN(
        P2_U3166) );
  AOI22_X1 U22158 ( .A1(n20311), .A2(n20025), .B1(n20058), .B2(n20310), .ZN(
        n20031) );
  AOI22_X1 U22159 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20059), .ZN(n20030) );
  OAI211_X1 U22160 ( .C1(n20062), .C2(n20316), .A(n20031), .B(n20030), .ZN(
        P2_U3158) );
  AOI22_X1 U22161 ( .A1(n20318), .A2(n20025), .B1(n20058), .B2(n20317), .ZN(
        n20033) );
  AOI22_X1 U22162 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n20319), .B2(n20059), .ZN(n20032) );
  OAI211_X1 U22163 ( .C1(n20062), .C2(n20323), .A(n20033), .B(n20032), .ZN(
        P2_U3150) );
  AOI22_X1 U22164 ( .A1(n20325), .A2(n20025), .B1(n20058), .B2(n20324), .ZN(
        n20035) );
  AOI22_X1 U22165 ( .A1(n20059), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20034) );
  OAI211_X1 U22166 ( .C1(n20062), .C2(n20329), .A(n20035), .B(n20034), .ZN(
        P2_U3142) );
  AOI22_X1 U22167 ( .A1(n20052), .A2(n20331), .B1(n20058), .B2(n20330), .ZN(
        n20037) );
  AOI22_X1 U22168 ( .A1(n20025), .A2(n20332), .B1(n20338), .B2(n20059), .ZN(
        n20036) );
  OAI211_X1 U22169 ( .C1(n20336), .C2(n12249), .A(n20037), .B(n20036), .ZN(
        P2_U3134) );
  AOI22_X1 U22170 ( .A1(n20059), .A2(n20345), .B1(n20337), .B2(n20058), .ZN(
        n20039) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20340), .B1(
        n20025), .B2(n20339), .ZN(n20038) );
  OAI211_X1 U22172 ( .C1(n20062), .C2(n20262), .A(n20039), .B(n20038), .ZN(
        P2_U3126) );
  AOI22_X1 U22173 ( .A1(n20052), .A2(n20345), .B1(n20058), .B2(n20344), .ZN(
        n20041) );
  AOI22_X1 U22174 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20347), .B1(
        n20025), .B2(n20346), .ZN(n20040) );
  OAI211_X1 U22175 ( .C1(n20055), .C2(n20356), .A(n20041), .B(n20040), .ZN(
        P2_U3118) );
  AOI22_X1 U22176 ( .A1(n20351), .A2(n20025), .B1(n20350), .B2(n20058), .ZN(
        n20043) );
  AOI22_X1 U22177 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20059), .ZN(n20042) );
  OAI211_X1 U22178 ( .C1(n20062), .C2(n20356), .A(n20043), .B(n20042), .ZN(
        P2_U3110) );
  AOI22_X1 U22179 ( .A1(n20358), .A2(n20025), .B1(n20058), .B2(n20357), .ZN(
        n20045) );
  AOI22_X1 U22180 ( .A1(n20059), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n20359), .ZN(n20044) );
  OAI211_X1 U22181 ( .C1(n20062), .C2(n20363), .A(n20045), .B(n20044), .ZN(
        P2_U3102) );
  AOI22_X1 U22182 ( .A1(n20052), .A2(n20360), .B1(n20364), .B2(n20058), .ZN(
        n20047) );
  AOI22_X1 U22183 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20366), .B1(
        n20025), .B2(n20365), .ZN(n20046) );
  OAI211_X1 U22184 ( .C1(n20055), .C2(n20232), .A(n20047), .B(n20046), .ZN(
        P2_U3094) );
  AOI22_X1 U22185 ( .A1(n20052), .A2(n20371), .B1(n20058), .B2(n20370), .ZN(
        n20049) );
  AOI22_X1 U22186 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20373), .B1(
        n20025), .B2(n20372), .ZN(n20048) );
  OAI211_X1 U22187 ( .C1(n20055), .C2(n20381), .A(n20049), .B(n20048), .ZN(
        P2_U3086) );
  AOI22_X1 U22188 ( .A1(n20052), .A2(n20273), .B1(n20058), .B2(n20376), .ZN(
        n20051) );
  AOI22_X1 U22189 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20378), .B1(
        n20025), .B2(n20377), .ZN(n20050) );
  OAI211_X1 U22190 ( .C1(n20055), .C2(n20276), .A(n20051), .B(n20050), .ZN(
        P2_U3078) );
  AOI22_X1 U22191 ( .A1(n20383), .A2(n20025), .B1(n20058), .B2(n20382), .ZN(
        n20054) );
  AOI22_X1 U22192 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20052), .ZN(n20053) );
  OAI211_X1 U22193 ( .C1(n20055), .C2(n20394), .A(n20054), .B(n20053), .ZN(
        P2_U3070) );
  AOI22_X1 U22194 ( .A1(n20389), .A2(n20025), .B1(n20058), .B2(n20388), .ZN(
        n20057) );
  AOI22_X1 U22195 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n20059), .B2(n20398), .ZN(n20056) );
  OAI211_X1 U22196 ( .C1(n20062), .C2(n20394), .A(n20057), .B(n20056), .ZN(
        P2_U3062) );
  AOI22_X1 U22197 ( .A1(n20059), .A2(n20285), .B1(n20058), .B2(n20397), .ZN(
        n20061) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20025), .ZN(n20060) );
  OAI211_X1 U22199 ( .C1(n20062), .C2(n20289), .A(n20061), .B(n20060), .ZN(
        P2_U3054) );
  AOI22_X1 U22200 ( .A1(n20064), .A2(n20063), .B1(n20111), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n20069) );
  OR3_X1 U22201 ( .A1(n20067), .A2(n20066), .A3(n20065), .ZN(n20068) );
  OAI211_X1 U22202 ( .C1(n20071), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P2_U2914) );
  AOI22_X1 U22203 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20297), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n20298), .ZN(n20110) );
  NOR2_X2 U22204 ( .A1(n15857), .A2(n20293), .ZN(n20106) );
  AOI22_X1 U22205 ( .A1(n20296), .A2(n20073), .B1(n20295), .B2(n20106), .ZN(
        n20075) );
  AOI22_X1 U22206 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20300), .B1(
        n20285), .B2(n20107), .ZN(n20074) );
  OAI211_X1 U22207 ( .C1(n20110), .C2(n20309), .A(n20075), .B(n20074), .ZN(
        P2_U3173) );
  AOI22_X1 U22208 ( .A1(n20102), .A2(n20304), .B1(n20106), .B2(n20303), .ZN(
        n20077) );
  AOI22_X1 U22209 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20306), .B1(
        n20073), .B2(n20305), .ZN(n20076) );
  OAI211_X1 U22210 ( .C1(n20105), .C2(n20309), .A(n20077), .B(n20076), .ZN(
        P2_U3165) );
  AOI22_X1 U22211 ( .A1(n20311), .A2(n20073), .B1(n20106), .B2(n20310), .ZN(
        n20079) );
  AOI22_X1 U22212 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20102), .ZN(n20078) );
  OAI211_X1 U22213 ( .C1(n20105), .C2(n20316), .A(n20079), .B(n20078), .ZN(
        P2_U3157) );
  AOI22_X1 U22214 ( .A1(n20318), .A2(n20073), .B1(n20106), .B2(n20317), .ZN(
        n20081) );
  AOI22_X1 U22215 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n20319), .B2(n20102), .ZN(n20080) );
  OAI211_X1 U22216 ( .C1(n20105), .C2(n20323), .A(n20081), .B(n20080), .ZN(
        P2_U3149) );
  AOI22_X1 U22217 ( .A1(n20325), .A2(n20073), .B1(n20106), .B2(n20324), .ZN(
        n20083) );
  AOI22_X1 U22218 ( .A1(n20102), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n20082) );
  OAI211_X1 U22219 ( .C1(n20105), .C2(n20329), .A(n20083), .B(n20082), .ZN(
        P2_U3141) );
  AOI22_X1 U22220 ( .A1(n20107), .A2(n20331), .B1(n20106), .B2(n20330), .ZN(
        n20085) );
  AOI22_X1 U22221 ( .A1(n20073), .A2(n20332), .B1(n20338), .B2(n20102), .ZN(
        n20084) );
  OAI211_X1 U22222 ( .C1(n20336), .C2(n12191), .A(n20085), .B(n20084), .ZN(
        P2_U3133) );
  AOI22_X1 U22223 ( .A1(n20102), .A2(n20345), .B1(n20337), .B2(n20106), .ZN(
        n20087) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20340), .B1(
        n20073), .B2(n20339), .ZN(n20086) );
  OAI211_X1 U22225 ( .C1(n20105), .C2(n20262), .A(n20087), .B(n20086), .ZN(
        P2_U3125) );
  AOI22_X1 U22226 ( .A1(n20107), .A2(n20345), .B1(n20106), .B2(n20344), .ZN(
        n20089) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20347), .B1(
        n20073), .B2(n20346), .ZN(n20088) );
  OAI211_X1 U22228 ( .C1(n20110), .C2(n20356), .A(n20089), .B(n20088), .ZN(
        P2_U3117) );
  AOI22_X1 U22229 ( .A1(n20351), .A2(n20073), .B1(n20350), .B2(n20106), .ZN(
        n20091) );
  AOI22_X1 U22230 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20102), .ZN(n20090) );
  OAI211_X1 U22231 ( .C1(n20105), .C2(n20356), .A(n20091), .B(n20090), .ZN(
        P2_U3109) );
  AOI22_X1 U22232 ( .A1(n20358), .A2(n20073), .B1(n20106), .B2(n20357), .ZN(
        n20093) );
  AOI22_X1 U22233 ( .A1(n20102), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n20359), .ZN(n20092) );
  OAI211_X1 U22234 ( .C1(n20105), .C2(n20363), .A(n20093), .B(n20092), .ZN(
        P2_U3101) );
  AOI22_X1 U22235 ( .A1(n20107), .A2(n20360), .B1(n20364), .B2(n20106), .ZN(
        n20095) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20366), .B1(
        n20073), .B2(n20365), .ZN(n20094) );
  OAI211_X1 U22237 ( .C1(n20110), .C2(n20232), .A(n20095), .B(n20094), .ZN(
        P2_U3093) );
  AOI22_X1 U22238 ( .A1(n20107), .A2(n20371), .B1(n20106), .B2(n20370), .ZN(
        n20097) );
  AOI22_X1 U22239 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20373), .B1(
        n20073), .B2(n20372), .ZN(n20096) );
  OAI211_X1 U22240 ( .C1(n20110), .C2(n20381), .A(n20097), .B(n20096), .ZN(
        P2_U3085) );
  AOI22_X1 U22241 ( .A1(n20102), .A2(n20384), .B1(n20106), .B2(n20376), .ZN(
        n20099) );
  AOI22_X1 U22242 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20378), .B1(
        n20073), .B2(n20377), .ZN(n20098) );
  OAI211_X1 U22243 ( .C1(n20105), .C2(n20381), .A(n20099), .B(n20098), .ZN(
        P2_U3077) );
  AOI22_X1 U22244 ( .A1(n20383), .A2(n20073), .B1(n20106), .B2(n20382), .ZN(
        n20101) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20107), .ZN(n20100) );
  OAI211_X1 U22246 ( .C1(n20110), .C2(n20394), .A(n20101), .B(n20100), .ZN(
        P2_U3069) );
  AOI22_X1 U22247 ( .A1(n20389), .A2(n20073), .B1(n20106), .B2(n20388), .ZN(
        n20104) );
  AOI22_X1 U22248 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n20102), .B2(n20398), .ZN(n20103) );
  OAI211_X1 U22249 ( .C1(n20105), .C2(n20394), .A(n20104), .B(n20103), .ZN(
        P2_U3061) );
  AOI22_X1 U22250 ( .A1(n20107), .A2(n20398), .B1(n20106), .B2(n20397), .ZN(
        n20109) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20073), .ZN(n20108) );
  OAI211_X1 U22252 ( .C1(n20110), .C2(n20405), .A(n20109), .B(n20108), .ZN(
        P2_U3053) );
  AOI22_X1 U22253 ( .A1(n20113), .A2(n20112), .B1(n20111), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n20123) );
  AOI22_X1 U22254 ( .A1(n20115), .A2(BUF1_REG_20__SCAN_IN), .B1(n20114), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n20122) );
  INV_X1 U22255 ( .A(n20116), .ZN(n20118) );
  AOI22_X1 U22256 ( .A1(n20120), .A2(n20119), .B1(n20118), .B2(n20117), .ZN(
        n20121) );
  NAND3_X1 U22257 ( .A1(n20123), .A2(n20122), .A3(n20121), .ZN(P2_U2899) );
  NOR2_X2 U22258 ( .A1(n20124), .A2(n20291), .ZN(n20161) );
  NOR2_X2 U22259 ( .A1(n20125), .A2(n20293), .ZN(n20159) );
  AOI22_X1 U22260 ( .A1(n20296), .A2(n20161), .B1(n20295), .B2(n20159), .ZN(
        n20127) );
  AOI22_X1 U22261 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20297), .ZN(n20164) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20155), .ZN(n20126) );
  OAI211_X1 U22263 ( .C1(n20158), .C2(n20405), .A(n20127), .B(n20126), .ZN(
        P2_U3172) );
  AOI22_X1 U22264 ( .A1(n20155), .A2(n20304), .B1(n20159), .B2(n20303), .ZN(
        n20129) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20306), .B1(
        n20161), .B2(n20305), .ZN(n20128) );
  OAI211_X1 U22266 ( .C1(n20158), .C2(n20309), .A(n20129), .B(n20128), .ZN(
        P2_U3164) );
  AOI22_X1 U22267 ( .A1(n20311), .A2(n20161), .B1(n20159), .B2(n20310), .ZN(
        n20131) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20313), .B1(
        n20304), .B2(n20160), .ZN(n20130) );
  OAI211_X1 U22269 ( .C1(n20164), .C2(n20323), .A(n20131), .B(n20130), .ZN(
        P2_U3156) );
  AOI22_X1 U22270 ( .A1(n20318), .A2(n20161), .B1(n20159), .B2(n20317), .ZN(
        n20133) );
  AOI22_X1 U22271 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n20319), .B2(n20155), .ZN(n20132) );
  OAI211_X1 U22272 ( .C1(n20158), .C2(n20323), .A(n20133), .B(n20132), .ZN(
        P2_U3148) );
  AOI22_X1 U22273 ( .A1(n20325), .A2(n20161), .B1(n20159), .B2(n20324), .ZN(
        n20135) );
  AOI22_X1 U22274 ( .A1(n20155), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20134) );
  OAI211_X1 U22275 ( .C1(n20158), .C2(n20329), .A(n20135), .B(n20134), .ZN(
        P2_U3140) );
  INV_X1 U22276 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n20138) );
  AOI22_X1 U22277 ( .A1(n20155), .A2(n20338), .B1(n20159), .B2(n20330), .ZN(
        n20137) );
  AOI22_X1 U22278 ( .A1(n20161), .A2(n20332), .B1(n20331), .B2(n20160), .ZN(
        n20136) );
  OAI211_X1 U22279 ( .C1(n20336), .C2(n20138), .A(n20137), .B(n20136), .ZN(
        P2_U3132) );
  AOI22_X1 U22280 ( .A1(n20160), .A2(n20338), .B1(n20337), .B2(n20159), .ZN(
        n20140) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20340), .B1(
        n20161), .B2(n20339), .ZN(n20139) );
  OAI211_X1 U22282 ( .C1(n20164), .C2(n20343), .A(n20140), .B(n20139), .ZN(
        P2_U3124) );
  AOI22_X1 U22283 ( .A1(n20160), .A2(n20345), .B1(n20159), .B2(n20344), .ZN(
        n20142) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20347), .B1(
        n20161), .B2(n20346), .ZN(n20141) );
  OAI211_X1 U22285 ( .C1(n20164), .C2(n20356), .A(n20142), .B(n20141), .ZN(
        P2_U3116) );
  AOI22_X1 U22286 ( .A1(n20351), .A2(n20161), .B1(n20350), .B2(n20159), .ZN(
        n20144) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20155), .ZN(n20143) );
  OAI211_X1 U22288 ( .C1(n20158), .C2(n20356), .A(n20144), .B(n20143), .ZN(
        P2_U3108) );
  AOI22_X1 U22289 ( .A1(n20358), .A2(n20161), .B1(n20159), .B2(n20357), .ZN(
        n20146) );
  AOI22_X1 U22290 ( .A1(n20155), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n20359), .ZN(n20145) );
  OAI211_X1 U22291 ( .C1(n20158), .C2(n20363), .A(n20146), .B(n20145), .ZN(
        P2_U3100) );
  AOI22_X1 U22292 ( .A1(n20155), .A2(n20371), .B1(n20364), .B2(n20159), .ZN(
        n20148) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20366), .B1(
        n20161), .B2(n20365), .ZN(n20147) );
  OAI211_X1 U22294 ( .C1(n20158), .C2(n20369), .A(n20148), .B(n20147), .ZN(
        P2_U3092) );
  AOI22_X1 U22295 ( .A1(n20160), .A2(n20371), .B1(n20159), .B2(n20370), .ZN(
        n20150) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20373), .B1(
        n20161), .B2(n20372), .ZN(n20149) );
  OAI211_X1 U22297 ( .C1(n20164), .C2(n20381), .A(n20150), .B(n20149), .ZN(
        P2_U3084) );
  AOI22_X1 U22298 ( .A1(n20155), .A2(n20384), .B1(n20159), .B2(n20376), .ZN(
        n20152) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20378), .B1(
        n20161), .B2(n20377), .ZN(n20151) );
  OAI211_X1 U22300 ( .C1(n20158), .C2(n20381), .A(n20152), .B(n20151), .ZN(
        P2_U3076) );
  AOI22_X1 U22301 ( .A1(n20383), .A2(n20161), .B1(n20159), .B2(n20382), .ZN(
        n20154) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20160), .ZN(n20153) );
  OAI211_X1 U22303 ( .C1(n20164), .C2(n20394), .A(n20154), .B(n20153), .ZN(
        P2_U3068) );
  AOI22_X1 U22304 ( .A1(n20389), .A2(n20161), .B1(n20159), .B2(n20388), .ZN(
        n20157) );
  AOI22_X1 U22305 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n20155), .B2(n20398), .ZN(n20156) );
  OAI211_X1 U22306 ( .C1(n20158), .C2(n20394), .A(n20157), .B(n20156), .ZN(
        P2_U3060) );
  AOI22_X1 U22307 ( .A1(n20160), .A2(n20398), .B1(n20397), .B2(n20159), .ZN(
        n20163) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20161), .ZN(n20162) );
  OAI211_X1 U22309 ( .C1(n20164), .C2(n20405), .A(n20163), .B(n20162), .ZN(
        P2_U3052) );
  NOR2_X2 U22310 ( .A1(n20165), .A2(n20291), .ZN(n20201) );
  NOR2_X2 U22311 ( .A1(n20166), .A2(n20293), .ZN(n20199) );
  AOI22_X1 U22312 ( .A1(n20296), .A2(n20201), .B1(n20295), .B2(n20199), .ZN(
        n20168) );
  AOI22_X1 U22313 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20297), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20298), .ZN(n20196) );
  AOI22_X1 U22314 ( .A1(n20285), .A2(n20193), .B1(n20299), .B2(n20200), .ZN(
        n20167) );
  OAI211_X1 U22315 ( .C1(n20210), .C2(n12122), .A(n20168), .B(n20167), .ZN(
        P2_U3171) );
  AOI22_X1 U22316 ( .A1(n20193), .A2(n20299), .B1(n20199), .B2(n20303), .ZN(
        n20170) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20306), .B1(
        n20201), .B2(n20305), .ZN(n20169) );
  OAI211_X1 U22318 ( .C1(n20196), .C2(n20316), .A(n20170), .B(n20169), .ZN(
        P2_U3163) );
  AOI22_X1 U22319 ( .A1(n20311), .A2(n20201), .B1(n20199), .B2(n20310), .ZN(
        n20172) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20313), .B1(
        n20304), .B2(n20193), .ZN(n20171) );
  OAI211_X1 U22321 ( .C1(n20196), .C2(n20323), .A(n20172), .B(n20171), .ZN(
        P2_U3155) );
  AOI22_X1 U22322 ( .A1(n20318), .A2(n20201), .B1(n20199), .B2(n20317), .ZN(
        n20174) );
  AOI22_X1 U22323 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n20319), .B2(n20200), .ZN(n20173) );
  OAI211_X1 U22324 ( .C1(n20204), .C2(n20323), .A(n20174), .B(n20173), .ZN(
        P2_U3147) );
  AOI22_X1 U22325 ( .A1(n20325), .A2(n20201), .B1(n20199), .B2(n20324), .ZN(
        n20176) );
  AOI22_X1 U22326 ( .A1(n20200), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n20175) );
  OAI211_X1 U22327 ( .C1(n20204), .C2(n20329), .A(n20176), .B(n20175), .ZN(
        P2_U3139) );
  AOI22_X1 U22328 ( .A1(n20200), .A2(n20338), .B1(n20199), .B2(n20330), .ZN(
        n20178) );
  AOI22_X1 U22329 ( .A1(n20201), .A2(n20332), .B1(n20331), .B2(n20193), .ZN(
        n20177) );
  OAI211_X1 U22330 ( .C1(n20336), .C2(n12100), .A(n20178), .B(n20177), .ZN(
        P2_U3131) );
  AOI22_X1 U22331 ( .A1(n20193), .A2(n20338), .B1(n20337), .B2(n20199), .ZN(
        n20180) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20340), .B1(
        n20201), .B2(n20339), .ZN(n20179) );
  OAI211_X1 U22333 ( .C1(n20196), .C2(n20343), .A(n20180), .B(n20179), .ZN(
        P2_U3123) );
  AOI22_X1 U22334 ( .A1(n20193), .A2(n20345), .B1(n20199), .B2(n20344), .ZN(
        n20182) );
  AOI22_X1 U22335 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20347), .B1(
        n20201), .B2(n20346), .ZN(n20181) );
  OAI211_X1 U22336 ( .C1(n20196), .C2(n20356), .A(n20182), .B(n20181), .ZN(
        P2_U3115) );
  AOI22_X1 U22337 ( .A1(n20351), .A2(n20201), .B1(n20350), .B2(n20199), .ZN(
        n20184) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20200), .ZN(n20183) );
  OAI211_X1 U22339 ( .C1(n20204), .C2(n20356), .A(n20184), .B(n20183), .ZN(
        P2_U3107) );
  AOI22_X1 U22340 ( .A1(n20358), .A2(n20201), .B1(n20199), .B2(n20357), .ZN(
        n20186) );
  AOI22_X1 U22341 ( .A1(n20200), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n20359), .ZN(n20185) );
  OAI211_X1 U22342 ( .C1(n20204), .C2(n20363), .A(n20186), .B(n20185), .ZN(
        P2_U3099) );
  AOI22_X1 U22343 ( .A1(n20200), .A2(n20371), .B1(n20364), .B2(n20199), .ZN(
        n20188) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20366), .B1(
        n20201), .B2(n20365), .ZN(n20187) );
  OAI211_X1 U22345 ( .C1(n20204), .C2(n20369), .A(n20188), .B(n20187), .ZN(
        P2_U3091) );
  AOI22_X1 U22346 ( .A1(n20193), .A2(n20371), .B1(n20370), .B2(n20199), .ZN(
        n20190) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20373), .B1(
        n20201), .B2(n20372), .ZN(n20189) );
  OAI211_X1 U22348 ( .C1(n20196), .C2(n20381), .A(n20190), .B(n20189), .ZN(
        P2_U3083) );
  AOI22_X1 U22349 ( .A1(n20200), .A2(n20384), .B1(n20376), .B2(n20199), .ZN(
        n20192) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20378), .B1(
        n20201), .B2(n20377), .ZN(n20191) );
  OAI211_X1 U22351 ( .C1(n20204), .C2(n20381), .A(n20192), .B(n20191), .ZN(
        P2_U3075) );
  AOI22_X1 U22352 ( .A1(n20383), .A2(n20201), .B1(n20199), .B2(n20382), .ZN(
        n20195) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20193), .ZN(n20194) );
  OAI211_X1 U22354 ( .C1(n20196), .C2(n20394), .A(n20195), .B(n20194), .ZN(
        P2_U3067) );
  AOI22_X1 U22355 ( .A1(n20389), .A2(n20201), .B1(n20199), .B2(n20388), .ZN(
        n20198) );
  AOI22_X1 U22356 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n20200), .B2(n20398), .ZN(n20197) );
  OAI211_X1 U22357 ( .C1(n20204), .C2(n20394), .A(n20198), .B(n20197), .ZN(
        P2_U3059) );
  AOI22_X1 U22358 ( .A1(n20200), .A2(n20285), .B1(n20397), .B2(n20199), .ZN(
        n20203) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20201), .ZN(n20202) );
  OAI211_X1 U22360 ( .C1(n20204), .C2(n20289), .A(n20203), .B(n20202), .ZN(
        P2_U3051) );
  INV_X1 U22361 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20209) );
  NOR2_X2 U22362 ( .A1(n20205), .A2(n20291), .ZN(n20245) );
  NOR2_X2 U22363 ( .A1(n20206), .A2(n20293), .ZN(n20243) );
  AOI22_X1 U22364 ( .A1(n20296), .A2(n20245), .B1(n20295), .B2(n20243), .ZN(
        n20208) );
  AOI22_X1 U22365 ( .A1(n20285), .A2(n20237), .B1(n20299), .B2(n20244), .ZN(
        n20207) );
  OAI211_X1 U22366 ( .C1(n20210), .C2(n20209), .A(n20208), .B(n20207), .ZN(
        P2_U3170) );
  AOI22_X1 U22367 ( .A1(n20237), .A2(n20299), .B1(n20243), .B2(n20303), .ZN(
        n20212) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20306), .B1(
        n20245), .B2(n20305), .ZN(n20211) );
  OAI211_X1 U22369 ( .C1(n20240), .C2(n20316), .A(n20212), .B(n20211), .ZN(
        P2_U3162) );
  AOI22_X1 U22370 ( .A1(n20311), .A2(n20245), .B1(n20243), .B2(n20310), .ZN(
        n20214) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20313), .B1(
        n20304), .B2(n20237), .ZN(n20213) );
  OAI211_X1 U22372 ( .C1(n20240), .C2(n20323), .A(n20214), .B(n20213), .ZN(
        P2_U3154) );
  AOI22_X1 U22373 ( .A1(n20318), .A2(n20245), .B1(n20243), .B2(n20317), .ZN(
        n20216) );
  AOI22_X1 U22374 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n20319), .B2(n20244), .ZN(n20215) );
  OAI211_X1 U22375 ( .C1(n20248), .C2(n20323), .A(n20216), .B(n20215), .ZN(
        P2_U3146) );
  AOI22_X1 U22376 ( .A1(n20325), .A2(n20245), .B1(n20243), .B2(n20324), .ZN(
        n20218) );
  AOI22_X1 U22377 ( .A1(n20244), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n20217) );
  OAI211_X1 U22378 ( .C1(n20248), .C2(n20329), .A(n20218), .B(n20217), .ZN(
        P2_U3138) );
  INV_X1 U22379 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20221) );
  AOI22_X1 U22380 ( .A1(n20237), .A2(n20331), .B1(n20243), .B2(n20330), .ZN(
        n20220) );
  AOI22_X1 U22381 ( .A1(n20245), .A2(n20332), .B1(n20338), .B2(n20244), .ZN(
        n20219) );
  OAI211_X1 U22382 ( .C1(n20336), .C2(n20221), .A(n20220), .B(n20219), .ZN(
        P2_U3130) );
  AOI22_X1 U22383 ( .A1(n20237), .A2(n20338), .B1(n20337), .B2(n20243), .ZN(
        n20223) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20340), .B1(
        n20245), .B2(n20339), .ZN(n20222) );
  OAI211_X1 U22385 ( .C1(n20240), .C2(n20343), .A(n20223), .B(n20222), .ZN(
        P2_U3122) );
  AOI22_X1 U22386 ( .A1(n20237), .A2(n20345), .B1(n20243), .B2(n20344), .ZN(
        n20225) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20347), .B1(
        n20245), .B2(n20346), .ZN(n20224) );
  OAI211_X1 U22388 ( .C1(n20240), .C2(n20356), .A(n20225), .B(n20224), .ZN(
        P2_U3114) );
  AOI22_X1 U22389 ( .A1(n20351), .A2(n20245), .B1(n20350), .B2(n20243), .ZN(
        n20227) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20244), .ZN(n20226) );
  OAI211_X1 U22391 ( .C1(n20248), .C2(n20356), .A(n20227), .B(n20226), .ZN(
        P2_U3106) );
  AOI22_X1 U22392 ( .A1(n20358), .A2(n20245), .B1(n20243), .B2(n20357), .ZN(
        n20229) );
  AOI22_X1 U22393 ( .A1(n20244), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n20359), .ZN(n20228) );
  OAI211_X1 U22394 ( .C1(n20248), .C2(n20363), .A(n20229), .B(n20228), .ZN(
        P2_U3098) );
  AOI22_X1 U22395 ( .A1(n20237), .A2(n20360), .B1(n20364), .B2(n20243), .ZN(
        n20231) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20366), .B1(
        n20245), .B2(n20365), .ZN(n20230) );
  OAI211_X1 U22397 ( .C1(n20240), .C2(n20232), .A(n20231), .B(n20230), .ZN(
        P2_U3090) );
  AOI22_X1 U22398 ( .A1(n20237), .A2(n20371), .B1(n20243), .B2(n20370), .ZN(
        n20234) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20373), .B1(
        n20245), .B2(n20372), .ZN(n20233) );
  OAI211_X1 U22400 ( .C1(n20240), .C2(n20381), .A(n20234), .B(n20233), .ZN(
        P2_U3082) );
  AOI22_X1 U22401 ( .A1(n20244), .A2(n20384), .B1(n20243), .B2(n20376), .ZN(
        n20236) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20378), .B1(
        n20245), .B2(n20377), .ZN(n20235) );
  OAI211_X1 U22403 ( .C1(n20248), .C2(n20381), .A(n20236), .B(n20235), .ZN(
        P2_U3074) );
  AOI22_X1 U22404 ( .A1(n20383), .A2(n20245), .B1(n20243), .B2(n20382), .ZN(
        n20239) );
  AOI22_X1 U22405 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20237), .ZN(n20238) );
  OAI211_X1 U22406 ( .C1(n20240), .C2(n20394), .A(n20239), .B(n20238), .ZN(
        P2_U3066) );
  AOI22_X1 U22407 ( .A1(n20389), .A2(n20245), .B1(n20243), .B2(n20388), .ZN(
        n20242) );
  AOI22_X1 U22408 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n20244), .B2(n20398), .ZN(n20241) );
  OAI211_X1 U22409 ( .C1(n20248), .C2(n20394), .A(n20242), .B(n20241), .ZN(
        P2_U3058) );
  AOI22_X1 U22410 ( .A1(n20244), .A2(n20285), .B1(n20243), .B2(n20397), .ZN(
        n20247) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20245), .ZN(n20246) );
  OAI211_X1 U22412 ( .C1(n20248), .C2(n20289), .A(n20247), .B(n20246), .ZN(
        P2_U3050) );
  AOI22_X1 U22413 ( .A1(n20304), .A2(n20284), .B1(n20283), .B2(n20303), .ZN(
        n20250) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20306), .B1(
        n20286), .B2(n20305), .ZN(n20249) );
  OAI211_X1 U22415 ( .C1(n20290), .C2(n20309), .A(n20250), .B(n20249), .ZN(
        P2_U3161) );
  AOI22_X1 U22416 ( .A1(n20311), .A2(n20286), .B1(n20283), .B2(n20310), .ZN(
        n20252) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20313), .B1(
        n20304), .B2(n20277), .ZN(n20251) );
  OAI211_X1 U22418 ( .C1(n20280), .C2(n20323), .A(n20252), .B(n20251), .ZN(
        P2_U3153) );
  AOI22_X1 U22419 ( .A1(n20318), .A2(n20286), .B1(n20283), .B2(n20317), .ZN(
        n20254) );
  AOI22_X1 U22420 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n20319), .B2(n20284), .ZN(n20253) );
  OAI211_X1 U22421 ( .C1(n20290), .C2(n20323), .A(n20254), .B(n20253), .ZN(
        P2_U3145) );
  AOI22_X1 U22422 ( .A1(n20325), .A2(n20286), .B1(n20283), .B2(n20324), .ZN(
        n20256) );
  AOI22_X1 U22423 ( .A1(n20284), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n20255) );
  OAI211_X1 U22424 ( .C1(n20290), .C2(n20329), .A(n20256), .B(n20255), .ZN(
        P2_U3137) );
  INV_X1 U22425 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20259) );
  AOI22_X1 U22426 ( .A1(n20277), .A2(n20331), .B1(n20283), .B2(n20330), .ZN(
        n20258) );
  AOI22_X1 U22427 ( .A1(n20286), .A2(n20332), .B1(n20338), .B2(n20284), .ZN(
        n20257) );
  OAI211_X1 U22428 ( .C1(n20336), .C2(n20259), .A(n20258), .B(n20257), .ZN(
        P2_U3129) );
  AOI22_X1 U22429 ( .A1(n20284), .A2(n20345), .B1(n20283), .B2(n20337), .ZN(
        n20261) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20340), .B1(
        n20286), .B2(n20339), .ZN(n20260) );
  OAI211_X1 U22431 ( .C1(n20290), .C2(n20262), .A(n20261), .B(n20260), .ZN(
        P2_U3121) );
  AOI22_X1 U22432 ( .A1(n20277), .A2(n20345), .B1(n20283), .B2(n20344), .ZN(
        n20264) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20347), .B1(
        n20286), .B2(n20346), .ZN(n20263) );
  OAI211_X1 U22434 ( .C1(n20280), .C2(n20356), .A(n20264), .B(n20263), .ZN(
        P2_U3113) );
  AOI22_X1 U22435 ( .A1(n20351), .A2(n20286), .B1(n20283), .B2(n20350), .ZN(
        n20266) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20284), .ZN(n20265) );
  OAI211_X1 U22437 ( .C1(n20290), .C2(n20356), .A(n20266), .B(n20265), .ZN(
        P2_U3105) );
  AOI22_X1 U22438 ( .A1(n20358), .A2(n20286), .B1(n20283), .B2(n20357), .ZN(
        n20268) );
  AOI22_X1 U22439 ( .A1(n20284), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n20359), .ZN(n20267) );
  OAI211_X1 U22440 ( .C1(n20290), .C2(n20363), .A(n20268), .B(n20267), .ZN(
        P2_U3097) );
  AOI22_X1 U22441 ( .A1(n20284), .A2(n20371), .B1(n20283), .B2(n20364), .ZN(
        n20270) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20366), .B1(
        n20286), .B2(n20365), .ZN(n20269) );
  OAI211_X1 U22443 ( .C1(n20290), .C2(n20369), .A(n20270), .B(n20269), .ZN(
        P2_U3089) );
  AOI22_X1 U22444 ( .A1(n20277), .A2(n20371), .B1(n20283), .B2(n20370), .ZN(
        n20272) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20373), .B1(
        n20286), .B2(n20372), .ZN(n20271) );
  OAI211_X1 U22446 ( .C1(n20280), .C2(n20381), .A(n20272), .B(n20271), .ZN(
        P2_U3081) );
  AOI22_X1 U22447 ( .A1(n20277), .A2(n20273), .B1(n20283), .B2(n20376), .ZN(
        n20275) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20378), .B1(
        n20286), .B2(n20377), .ZN(n20274) );
  OAI211_X1 U22449 ( .C1(n20280), .C2(n20276), .A(n20275), .B(n20274), .ZN(
        P2_U3073) );
  AOI22_X1 U22450 ( .A1(n20383), .A2(n20286), .B1(n20283), .B2(n20382), .ZN(
        n20279) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20277), .ZN(n20278) );
  OAI211_X1 U22452 ( .C1(n20280), .C2(n20394), .A(n20279), .B(n20278), .ZN(
        P2_U3065) );
  AOI22_X1 U22453 ( .A1(n20389), .A2(n20286), .B1(n20283), .B2(n20388), .ZN(
        n20282) );
  AOI22_X1 U22454 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n20284), .B2(n20398), .ZN(n20281) );
  OAI211_X1 U22455 ( .C1(n20290), .C2(n20394), .A(n20282), .B(n20281), .ZN(
        P2_U3057) );
  AOI22_X1 U22456 ( .A1(n20285), .A2(n20284), .B1(n20283), .B2(n20397), .ZN(
        n20288) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20286), .ZN(n20287) );
  OAI211_X1 U22458 ( .C1(n20290), .C2(n20289), .A(n20288), .B(n20287), .ZN(
        P2_U3049) );
  NOR2_X2 U22459 ( .A1(n20292), .A2(n20291), .ZN(n20400) );
  AOI22_X1 U22460 ( .A1(n20296), .A2(n20400), .B1(n20295), .B2(n11125), .ZN(
        n20302) );
  AOI22_X1 U22461 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20298), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20297), .ZN(n20406) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20300), .B1(
        n20299), .B2(n20390), .ZN(n20301) );
  OAI211_X1 U22463 ( .C1(n20395), .C2(n20405), .A(n20302), .B(n20301), .ZN(
        P2_U3168) );
  AOI22_X1 U22464 ( .A1(n20304), .A2(n20390), .B1(n11125), .B2(n20303), .ZN(
        n20308) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20306), .B1(
        n20400), .B2(n20305), .ZN(n20307) );
  OAI211_X1 U22466 ( .C1(n20395), .C2(n20309), .A(n20308), .B(n20307), .ZN(
        P2_U3160) );
  AOI22_X1 U22467 ( .A1(n20311), .A2(n20400), .B1(n11125), .B2(n20310), .ZN(
        n20315) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20313), .B1(
        n20312), .B2(n20390), .ZN(n20314) );
  OAI211_X1 U22469 ( .C1(n20395), .C2(n20316), .A(n20315), .B(n20314), .ZN(
        P2_U3152) );
  AOI22_X1 U22470 ( .A1(n20318), .A2(n20400), .B1(n11125), .B2(n20317), .ZN(
        n20322) );
  AOI22_X1 U22471 ( .A1(n20320), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n20319), .B2(n20390), .ZN(n20321) );
  OAI211_X1 U22472 ( .C1(n20395), .C2(n20323), .A(n20322), .B(n20321), .ZN(
        P2_U3144) );
  AOI22_X1 U22473 ( .A1(n20325), .A2(n20400), .B1(n11125), .B2(n20324), .ZN(
        n20328) );
  AOI22_X1 U22474 ( .A1(n20390), .A2(n20331), .B1(n20326), .B2(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20327) );
  OAI211_X1 U22475 ( .C1(n20395), .C2(n20329), .A(n20328), .B(n20327), .ZN(
        P2_U3136) );
  INV_X1 U22476 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n20335) );
  INV_X1 U22477 ( .A(n20395), .ZN(n20399) );
  AOI22_X1 U22478 ( .A1(n20399), .A2(n20331), .B1(n11125), .B2(n20330), .ZN(
        n20334) );
  AOI22_X1 U22479 ( .A1(n20400), .A2(n20332), .B1(n20338), .B2(n20390), .ZN(
        n20333) );
  OAI211_X1 U22480 ( .C1(n20336), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P2_U3128) );
  AOI22_X1 U22481 ( .A1(n20399), .A2(n20338), .B1(n20337), .B2(n11125), .ZN(
        n20342) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20340), .B1(
        n20400), .B2(n20339), .ZN(n20341) );
  OAI211_X1 U22483 ( .C1(n20406), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P2_U3120) );
  AOI22_X1 U22484 ( .A1(n20399), .A2(n20345), .B1(n11125), .B2(n20344), .ZN(
        n20349) );
  AOI22_X1 U22485 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20347), .B1(
        n20400), .B2(n20346), .ZN(n20348) );
  OAI211_X1 U22486 ( .C1(n20406), .C2(n20356), .A(n20349), .B(n20348), .ZN(
        P2_U3112) );
  AOI22_X1 U22487 ( .A1(n20351), .A2(n20400), .B1(n20350), .B2(n11125), .ZN(
        n20355) );
  AOI22_X1 U22488 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20353), .B1(
        n20352), .B2(n20390), .ZN(n20354) );
  OAI211_X1 U22489 ( .C1(n20395), .C2(n20356), .A(n20355), .B(n20354), .ZN(
        P2_U3104) );
  AOI22_X1 U22490 ( .A1(n20358), .A2(n20400), .B1(n11125), .B2(n20357), .ZN(
        n20362) );
  AOI22_X1 U22491 ( .A1(n20390), .A2(n20360), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n20359), .ZN(n20361) );
  OAI211_X1 U22492 ( .C1(n20395), .C2(n20363), .A(n20362), .B(n20361), .ZN(
        P2_U3096) );
  AOI22_X1 U22493 ( .A1(n20390), .A2(n20371), .B1(n20364), .B2(n11125), .ZN(
        n20368) );
  AOI22_X1 U22494 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20366), .B1(
        n20400), .B2(n20365), .ZN(n20367) );
  OAI211_X1 U22495 ( .C1(n20395), .C2(n20369), .A(n20368), .B(n20367), .ZN(
        P2_U3088) );
  AOI22_X1 U22496 ( .A1(n20399), .A2(n20371), .B1(n11125), .B2(n20370), .ZN(
        n20375) );
  AOI22_X1 U22497 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20373), .B1(
        n20400), .B2(n20372), .ZN(n20374) );
  OAI211_X1 U22498 ( .C1(n20406), .C2(n20381), .A(n20375), .B(n20374), .ZN(
        P2_U3080) );
  AOI22_X1 U22499 ( .A1(n20390), .A2(n20384), .B1(n11125), .B2(n20376), .ZN(
        n20380) );
  AOI22_X1 U22500 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20378), .B1(
        n20400), .B2(n20377), .ZN(n20379) );
  OAI211_X1 U22501 ( .C1(n20395), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P2_U3072) );
  AOI22_X1 U22502 ( .A1(n20383), .A2(n20400), .B1(n11125), .B2(n20382), .ZN(
        n20387) );
  AOI22_X1 U22503 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20385), .B1(
        n20384), .B2(n20399), .ZN(n20386) );
  OAI211_X1 U22504 ( .C1(n20406), .C2(n20394), .A(n20387), .B(n20386), .ZN(
        P2_U3064) );
  AOI22_X1 U22505 ( .A1(n20389), .A2(n20400), .B1(n11125), .B2(n20388), .ZN(
        n20393) );
  AOI22_X1 U22506 ( .A1(n20391), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n20390), .B2(n20398), .ZN(n20392) );
  OAI211_X1 U22507 ( .C1(n20395), .C2(n20394), .A(n20393), .B(n20392), .ZN(
        P2_U3056) );
  AOI22_X1 U22508 ( .A1(n20399), .A2(n20398), .B1(n20397), .B2(n11125), .ZN(
        n20404) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20402), .B1(
        n20401), .B2(n20400), .ZN(n20403) );
  OAI211_X1 U22510 ( .C1(n20406), .C2(n20405), .A(n20404), .B(n20403), .ZN(
        P2_U3048) );
  INV_X1 U22511 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20700) );
  INV_X1 U22512 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n20407) );
  AOI222_X1 U22513 ( .A1(n20698), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n20700), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n20407), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n20408) );
  OAI22_X1 U22514 ( .A1(n20457), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n20460), .ZN(n20409) );
  INV_X1 U22515 ( .A(n20409), .ZN(U376) );
  OAI22_X1 U22516 ( .A1(n20457), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n20460), .ZN(n20410) );
  INV_X1 U22517 ( .A(n20410), .ZN(U365) );
  OAI22_X1 U22518 ( .A1(n20457), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n20460), .ZN(n20411) );
  INV_X1 U22519 ( .A(n20411), .ZN(U354) );
  OAI22_X1 U22520 ( .A1(n20457), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n20408), .ZN(n20412) );
  INV_X1 U22521 ( .A(n20412), .ZN(U353) );
  OAI22_X1 U22522 ( .A1(n20457), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n20460), .ZN(n20413) );
  INV_X1 U22523 ( .A(n20413), .ZN(U352) );
  OAI22_X1 U22524 ( .A1(n20457), .A2(P3_ADDRESS_REG_5__SCAN_IN), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(n20460), .ZN(n20414) );
  INV_X1 U22525 ( .A(n20414), .ZN(U351) );
  INV_X2 U22526 ( .A(n20457), .ZN(n20460) );
  OAI22_X1 U22527 ( .A1(n20457), .A2(P3_ADDRESS_REG_6__SCAN_IN), .B1(
        P2_ADDRESS_REG_6__SCAN_IN), .B2(n20460), .ZN(n20415) );
  INV_X1 U22528 ( .A(n20415), .ZN(U350) );
  OAI22_X1 U22529 ( .A1(n20457), .A2(P3_ADDRESS_REG_7__SCAN_IN), .B1(
        P2_ADDRESS_REG_7__SCAN_IN), .B2(n20460), .ZN(n20416) );
  INV_X1 U22530 ( .A(n20416), .ZN(U349) );
  AOI22_X1 U22531 ( .A1(n20460), .A2(n20418), .B1(n20417), .B2(n20457), .ZN(
        U348) );
  AOI22_X1 U22532 ( .A1(n20460), .A2(n20420), .B1(n20419), .B2(n20457), .ZN(
        U347) );
  AOI22_X1 U22533 ( .A1(n20460), .A2(n20422), .B1(n20421), .B2(n20457), .ZN(
        U375) );
  AOI22_X1 U22534 ( .A1(n20460), .A2(n20424), .B1(n20423), .B2(n20457), .ZN(
        U374) );
  AOI22_X1 U22535 ( .A1(n20460), .A2(n20426), .B1(n20425), .B2(n20457), .ZN(
        U373) );
  AOI22_X1 U22536 ( .A1(n20460), .A2(n20428), .B1(n20427), .B2(n20457), .ZN(
        U372) );
  AOI22_X1 U22537 ( .A1(n20460), .A2(n20430), .B1(n20429), .B2(n20457), .ZN(
        U371) );
  AOI22_X1 U22538 ( .A1(n20460), .A2(n20432), .B1(n20431), .B2(n20457), .ZN(
        U370) );
  AOI22_X1 U22539 ( .A1(n20460), .A2(n20434), .B1(n20433), .B2(n20457), .ZN(
        U369) );
  AOI22_X1 U22540 ( .A1(n20460), .A2(n20436), .B1(n20435), .B2(n20457), .ZN(
        U368) );
  AOI22_X1 U22541 ( .A1(n20460), .A2(n20438), .B1(n20437), .B2(n20457), .ZN(
        U367) );
  AOI22_X1 U22542 ( .A1(n20460), .A2(n20440), .B1(n20439), .B2(n20457), .ZN(
        U366) );
  AOI22_X1 U22543 ( .A1(n20460), .A2(n20442), .B1(n20441), .B2(n20457), .ZN(
        U364) );
  AOI22_X1 U22544 ( .A1(n20460), .A2(n20444), .B1(n20443), .B2(n20457), .ZN(
        U363) );
  AOI22_X1 U22545 ( .A1(n20460), .A2(n20446), .B1(n20445), .B2(n20457), .ZN(
        U362) );
  AOI22_X1 U22546 ( .A1(n20460), .A2(n20448), .B1(n20447), .B2(n20457), .ZN(
        U361) );
  AOI22_X1 U22547 ( .A1(n20460), .A2(n20450), .B1(n20449), .B2(n20457), .ZN(
        U360) );
  AOI22_X1 U22548 ( .A1(n20408), .A2(n20452), .B1(n20451), .B2(n20457), .ZN(
        U359) );
  AOI22_X1 U22549 ( .A1(n20460), .A2(n20454), .B1(n20453), .B2(n20457), .ZN(
        U358) );
  AOI22_X1 U22550 ( .A1(n20460), .A2(n20456), .B1(n20455), .B2(n20457), .ZN(
        U357) );
  AOI22_X1 U22551 ( .A1(n20460), .A2(n20459), .B1(n20458), .B2(n20457), .ZN(
        U356) );
  AOI22_X1 U22552 ( .A1(n20408), .A2(n20462), .B1(n20461), .B2(n20457), .ZN(
        U355) );
  AOI22_X1 U22553 ( .A1(n21945), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20464) );
  OAI21_X1 U22554 ( .B1(n22391), .B2(n20481), .A(n20464), .ZN(P1_U2936) );
  AOI22_X1 U22555 ( .A1(n21945), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20465) );
  OAI21_X1 U22556 ( .B1(n22397), .B2(n20481), .A(n20465), .ZN(P1_U2935) );
  AOI22_X1 U22557 ( .A1(n21945), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20466) );
  OAI21_X1 U22558 ( .B1(n22403), .B2(n20481), .A(n20466), .ZN(P1_U2934) );
  AOI22_X1 U22559 ( .A1(n21945), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20467) );
  OAI21_X1 U22560 ( .B1(n22409), .B2(n20481), .A(n20467), .ZN(P1_U2933) );
  INV_X1 U22561 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n22417) );
  AOI22_X1 U22562 ( .A1(n21945), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20468) );
  OAI21_X1 U22563 ( .B1(n22417), .B2(n20481), .A(n20468), .ZN(P1_U2932) );
  AOI22_X1 U22564 ( .A1(n21945), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20469) );
  OAI21_X1 U22565 ( .B1(n13399), .B2(n20481), .A(n20469), .ZN(P1_U2931) );
  AOI22_X1 U22566 ( .A1(n21945), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20470) );
  OAI21_X1 U22567 ( .B1(n15299), .B2(n20481), .A(n20470), .ZN(P1_U2930) );
  AOI22_X1 U22568 ( .A1(n21945), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20471) );
  OAI21_X1 U22569 ( .B1(n13411), .B2(n20481), .A(n20471), .ZN(P1_U2929) );
  INV_X1 U22570 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n22439) );
  AOI22_X1 U22571 ( .A1(n21945), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20472) );
  OAI21_X1 U22572 ( .B1(n22439), .B2(n20481), .A(n20472), .ZN(P1_U2928) );
  INV_X1 U22573 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n22446) );
  AOI22_X1 U22574 ( .A1(n21945), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20473) );
  OAI21_X1 U22575 ( .B1(n22446), .B2(n20481), .A(n20473), .ZN(P1_U2927) );
  INV_X1 U22576 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n22453) );
  AOI22_X1 U22577 ( .A1(n21945), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20475) );
  OAI21_X1 U22578 ( .B1(n22453), .B2(n20481), .A(n20475), .ZN(P1_U2926) );
  INV_X1 U22579 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n22461) );
  AOI22_X1 U22580 ( .A1(n21945), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20476) );
  OAI21_X1 U22581 ( .B1(n22461), .B2(n20481), .A(n20476), .ZN(P1_U2925) );
  INV_X1 U22582 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n22468) );
  AOI22_X1 U22583 ( .A1(n21945), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20477) );
  OAI21_X1 U22584 ( .B1(n22468), .B2(n20481), .A(n20477), .ZN(P1_U2924) );
  INV_X1 U22585 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n22475) );
  AOI22_X1 U22586 ( .A1(n21945), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20478) );
  OAI21_X1 U22587 ( .B1(n22475), .B2(n20481), .A(n20478), .ZN(P1_U2923) );
  INV_X1 U22588 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n22485) );
  AOI22_X1 U22589 ( .A1(n21945), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20479) );
  OAI21_X1 U22590 ( .B1(n22485), .B2(n20481), .A(n20479), .ZN(P1_U2922) );
  AOI22_X1 U22591 ( .A1(n21945), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n20474), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20480) );
  OAI21_X1 U22592 ( .B1(n14497), .B2(n20481), .A(n20480), .ZN(P1_U2921) );
  OR2_X1 U22593 ( .A1(n22850), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20520) );
  INV_X1 U22594 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n22335) );
  NOR2_X1 U22595 ( .A1(n22335), .A2(n22850), .ZN(n20510) );
  OAI222_X1 U22596 ( .A1(n20520), .A2(n22124), .B1(n20482), .B2(n22853), .C1(
        n14610), .C2(n22331), .ZN(P1_U3197) );
  INV_X1 U22597 ( .A(n22331), .ZN(n20518) );
  AOI222_X1 U22598 ( .A1(n20515), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_2__SCAN_IN), 
        .C2(n20518), .ZN(n20483) );
  INV_X1 U22599 ( .A(n20483), .ZN(P1_U3198) );
  INV_X1 U22600 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n22123) );
  AOI22_X1 U22601 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n22850), .ZN(n20484) );
  OAI21_X1 U22602 ( .B1(n22123), .B2(n22331), .A(n20484), .ZN(P1_U3199) );
  AOI22_X1 U22603 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20518), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n22850), .ZN(n20485) );
  OAI21_X1 U22604 ( .B1(n22150), .B2(n20520), .A(n20485), .ZN(P1_U3200) );
  AOI22_X1 U22605 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n22850), .ZN(n20486) );
  OAI21_X1 U22606 ( .B1(n22150), .B2(n22331), .A(n20486), .ZN(P1_U3201) );
  AOI22_X1 U22607 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20518), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n22850), .ZN(n20487) );
  OAI21_X1 U22608 ( .B1(n22173), .B2(n20520), .A(n20487), .ZN(P1_U3202) );
  AOI222_X1 U22609 ( .A1(n20515), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20518), .ZN(n20488) );
  INV_X1 U22610 ( .A(n20488), .ZN(P1_U3203) );
  AOI222_X1 U22611 ( .A1(n20515), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20518), .ZN(n20489) );
  INV_X1 U22612 ( .A(n20489), .ZN(P1_U3204) );
  AOI222_X1 U22613 ( .A1(n20515), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20518), .ZN(n20490) );
  INV_X1 U22614 ( .A(n20490), .ZN(P1_U3205) );
  AOI222_X1 U22615 ( .A1(n20515), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20510), .ZN(n20491) );
  INV_X1 U22616 ( .A(n20491), .ZN(P1_U3206) );
  AOI222_X1 U22617 ( .A1(n20515), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20510), .ZN(n20492) );
  INV_X1 U22618 ( .A(n20492), .ZN(P1_U3207) );
  AOI222_X1 U22619 ( .A1(n20518), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20515), .ZN(n20493) );
  INV_X1 U22620 ( .A(n20493), .ZN(P1_U3208) );
  AOI222_X1 U22621 ( .A1(n20518), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20515), .ZN(n20494) );
  INV_X1 U22622 ( .A(n20494), .ZN(P1_U3209) );
  AOI222_X1 U22623 ( .A1(n20515), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20510), .ZN(n20495) );
  INV_X1 U22624 ( .A(n20495), .ZN(P1_U3210) );
  AOI222_X1 U22625 ( .A1(n20518), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20515), .ZN(n20496) );
  INV_X1 U22626 ( .A(n20496), .ZN(P1_U3211) );
  AOI222_X1 U22627 ( .A1(n20518), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20515), .ZN(n20497) );
  INV_X1 U22628 ( .A(n20497), .ZN(P1_U3212) );
  AOI222_X1 U22629 ( .A1(n20515), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20510), .ZN(n20498) );
  INV_X1 U22630 ( .A(n20498), .ZN(P1_U3213) );
  AOI22_X1 U22631 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n22850), .ZN(n20499) );
  OAI21_X1 U22632 ( .B1(n20500), .B2(n22331), .A(n20499), .ZN(P1_U3214) );
  INV_X1 U22633 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20502) );
  AOI22_X1 U22634 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n22850), .ZN(n20501) );
  OAI21_X1 U22635 ( .B1(n20502), .B2(n22331), .A(n20501), .ZN(P1_U3215) );
  AOI22_X1 U22636 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n20518), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n22850), .ZN(n20503) );
  OAI21_X1 U22637 ( .B1(n20504), .B2(n20520), .A(n20503), .ZN(P1_U3216) );
  AOI222_X1 U22638 ( .A1(n20515), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20510), .ZN(n20505) );
  INV_X1 U22639 ( .A(n20505), .ZN(P1_U3217) );
  AOI222_X1 U22640 ( .A1(n20515), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20510), .ZN(n20506) );
  INV_X1 U22641 ( .A(n20506), .ZN(P1_U3218) );
  AOI222_X1 U22642 ( .A1(n20515), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20518), .ZN(n20507) );
  INV_X1 U22643 ( .A(n20507), .ZN(P1_U3219) );
  AOI222_X1 U22644 ( .A1(n20515), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20510), .ZN(n20508) );
  INV_X1 U22645 ( .A(n20508), .ZN(P1_U3220) );
  AOI222_X1 U22646 ( .A1(n20515), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20518), .ZN(n20509) );
  INV_X1 U22647 ( .A(n20509), .ZN(P1_U3221) );
  AOI222_X1 U22648 ( .A1(n20515), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n22850), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20510), .ZN(n20511) );
  INV_X1 U22649 ( .A(n20511), .ZN(P1_U3222) );
  AOI22_X1 U22650 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n22850), .ZN(n20512) );
  OAI21_X1 U22651 ( .B1(n20513), .B2(n22331), .A(n20512), .ZN(P1_U3223) );
  AOI22_X1 U22652 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n20518), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n22850), .ZN(n20514) );
  OAI21_X1 U22653 ( .B1(n20517), .B2(n20520), .A(n20514), .ZN(P1_U3224) );
  AOI22_X1 U22654 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20515), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n22850), .ZN(n20516) );
  OAI21_X1 U22655 ( .B1(n20517), .B2(n22331), .A(n20516), .ZN(P1_U3225) );
  AOI22_X1 U22656 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20518), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n22850), .ZN(n20519) );
  OAI21_X1 U22657 ( .B1(n20521), .B2(n20520), .A(n20519), .ZN(P1_U3226) );
  OAI22_X1 U22658 ( .A1(n22850), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22853), .ZN(n20522) );
  INV_X1 U22659 ( .A(n20522), .ZN(P1_U3458) );
  NOR2_X1 U22660 ( .A1(P1_DATAWIDTH_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20523) );
  NAND2_X1 U22661 ( .A1(n20523), .A2(n20547), .ZN(n20543) );
  OAI21_X1 U22662 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20543), .ZN(n20534) );
  NOR4_X1 U22663 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20527) );
  NOR4_X1 U22664 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20526) );
  NOR4_X1 U22665 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20525) );
  NOR4_X1 U22666 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20524) );
  NAND4_X1 U22667 ( .A1(n20527), .A2(n20526), .A3(n20525), .A4(n20524), .ZN(
        n20533) );
  NOR4_X1 U22668 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20531) );
  AOI211_X1 U22669 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20530) );
  NOR4_X1 U22670 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20529) );
  NOR4_X1 U22671 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n20528) );
  NAND4_X1 U22672 ( .A1(n20531), .A2(n20530), .A3(n20529), .A4(n20528), .ZN(
        n20532) );
  OR2_X1 U22673 ( .A1(n20533), .A2(n20532), .ZN(n20545) );
  MUX2_X1 U22674 ( .A(n20534), .B(P1_BYTEENABLE_REG_3__SCAN_IN), .S(n20545), 
        .Z(P1_U2808) );
  OAI22_X1 U22675 ( .A1(n22850), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22853), .ZN(n20535) );
  INV_X1 U22676 ( .A(n20535), .ZN(P1_U3459) );
  NAND2_X1 U22677 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20540) );
  INV_X1 U22678 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n22307) );
  NOR2_X1 U22679 ( .A1(n20545), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20548) );
  OAI211_X1 U22680 ( .C1(n20536), .C2(n20547), .A(n22307), .B(n20548), .ZN(
        n20537) );
  INV_X1 U22681 ( .A(n20537), .ZN(n20538) );
  AOI21_X1 U22682 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n20545), .A(n20538), 
        .ZN(n20539) );
  OAI21_X1 U22683 ( .B1(n20540), .B2(n20545), .A(n20539), .ZN(P1_U3481) );
  OAI22_X1 U22684 ( .A1(n22850), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22853), .ZN(n20541) );
  INV_X1 U22685 ( .A(n20541), .ZN(P1_U3460) );
  AOI22_X1 U22686 ( .A1(n20548), .A2(n20543), .B1(n20542), .B2(n20545), .ZN(
        P1_U2807) );
  OAI22_X1 U22687 ( .A1(n22850), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22853), .ZN(n20544) );
  INV_X1 U22688 ( .A(n20544), .ZN(P1_U3461) );
  AOI22_X1 U22689 ( .A1(n20548), .A2(n20547), .B1(n20546), .B2(n20545), .ZN(
        P1_U3482) );
  INV_X1 U22690 ( .A(n20549), .ZN(n20550) );
  AOI21_X1 U22691 ( .B1(n20552), .B2(n20551), .A(n20550), .ZN(n22156) );
  AOI22_X1 U22692 ( .A1(n22159), .A2(n14221), .B1(n20572), .B2(n22156), .ZN(
        n20553) );
  OAI21_X1 U22693 ( .B1(n20574), .B2(n22154), .A(n20553), .ZN(P1_U2866) );
  AOI21_X1 U22694 ( .B1(n20556), .B2(n20555), .A(n20554), .ZN(n22213) );
  AOI22_X1 U22695 ( .A1(n22220), .A2(n14221), .B1(n20572), .B2(n22213), .ZN(
        n20557) );
  OAI21_X1 U22696 ( .B1(n20574), .B2(n20558), .A(n20557), .ZN(P1_U2860) );
  OR2_X1 U22697 ( .A1(n20560), .A2(n20559), .ZN(n20561) );
  AND2_X1 U22698 ( .A1(n20562), .A2(n20561), .ZN(n22189) );
  INV_X1 U22699 ( .A(n22189), .ZN(n20563) );
  OAI22_X1 U22700 ( .A1(n22195), .A2(n16146), .B1(n16143), .B2(n20563), .ZN(
        n20564) );
  INV_X1 U22701 ( .A(n20564), .ZN(n20565) );
  OAI21_X1 U22702 ( .B1(n20574), .B2(n22191), .A(n20565), .ZN(P1_U2862) );
  XNOR2_X1 U22703 ( .A(n20567), .B(n20566), .ZN(n22254) );
  AOI22_X1 U22704 ( .A1(n22257), .A2(n14221), .B1(n20572), .B2(n22254), .ZN(
        n20568) );
  OAI21_X1 U22705 ( .B1(n20574), .B2(n22248), .A(n20568), .ZN(P1_U2855) );
  INV_X1 U22706 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n22129) );
  AOI21_X1 U22707 ( .B1(n20571), .B2(n20570), .A(n20569), .ZN(n22126) );
  AOI22_X1 U22708 ( .A1(n22136), .A2(n14221), .B1(n20572), .B2(n22126), .ZN(
        n20573) );
  OAI21_X1 U22709 ( .B1(n20574), .B2(n22129), .A(n20573), .ZN(P1_U2868) );
  AOI22_X1 U22710 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20580) );
  OAI21_X1 U22711 ( .B1(n20577), .B2(n20576), .A(n20575), .ZN(n20578) );
  INV_X1 U22712 ( .A(n20578), .ZN(n21983) );
  AOI22_X1 U22713 ( .A1(n20595), .A2(n21983), .B1(n22136), .B2(n20614), .ZN(
        n20579) );
  OAI211_X1 U22714 ( .C1(n20634), .C2(n22138), .A(n20580), .B(n20579), .ZN(
        P1_U2995) );
  AOI22_X1 U22715 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n20586) );
  OAI21_X1 U22716 ( .B1(n20583), .B2(n20582), .A(n20581), .ZN(n20584) );
  INV_X1 U22717 ( .A(n20584), .ZN(n22001) );
  AOI22_X1 U22718 ( .A1(n20595), .A2(n22001), .B1(n22148), .B2(n20614), .ZN(
        n20585) );
  OAI211_X1 U22719 ( .C1(n20634), .C2(n22141), .A(n20586), .B(n20585), .ZN(
        P1_U2994) );
  AOI22_X1 U22720 ( .A1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n20592) );
  NAND2_X1 U22721 ( .A1(n20588), .A2(n20587), .ZN(n20589) );
  NAND2_X1 U22722 ( .A1(n20590), .A2(n20589), .ZN(n21996) );
  AOI22_X1 U22723 ( .A1(n21996), .A2(n20595), .B1(n22159), .B2(n20614), .ZN(
        n20591) );
  OAI211_X1 U22724 ( .C1(n20634), .C2(n22157), .A(n20592), .B(n20591), .ZN(
        P1_U2993) );
  AOI22_X1 U22725 ( .A1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n20597) );
  AOI21_X1 U22726 ( .B1(n20594), .B2(n20593), .A(n11210), .ZN(n22016) );
  AOI22_X1 U22727 ( .A1(n22016), .A2(n20595), .B1(n20614), .B2(n22171), .ZN(
        n20596) );
  OAI211_X1 U22728 ( .C1(n20634), .C2(n22165), .A(n20597), .B(n20596), .ZN(
        P1_U2992) );
  INV_X1 U22729 ( .A(n20604), .ZN(n20598) );
  MUX2_X1 U22730 ( .A(n20620), .B(n20598), .S(n20617), .Z(n20599) );
  NAND2_X1 U22731 ( .A1(n20599), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n20605) );
  OAI21_X1 U22732 ( .B1(n20599), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n20605), .ZN(n22043) );
  AOI22_X1 U22733 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n20602) );
  OAI22_X1 U22734 ( .A1(n22195), .A2(n20630), .B1(n22194), .B2(n20634), .ZN(
        n20600) );
  INV_X1 U22735 ( .A(n20600), .ZN(n20601) );
  OAI211_X1 U22736 ( .C1(n22280), .C2(n22043), .A(n20602), .B(n20601), .ZN(
        P1_U2989) );
  NOR2_X1 U22737 ( .A1(n22044), .A2(n22211), .ZN(n22059) );
  NOR2_X1 U22738 ( .A1(n20604), .A2(n20603), .ZN(n20606) );
  MUX2_X1 U22739 ( .A(n20603), .B(n20606), .S(n20605), .Z(n20607) );
  OAI22_X1 U22740 ( .A1(n22065), .A2(n22280), .B1(n20634), .B2(n22206), .ZN(
        n20608) );
  OAI21_X1 U22741 ( .B1(n20630), .B2(n22205), .A(n20609), .ZN(P1_U2988) );
  OAI21_X1 U22742 ( .B1(n20612), .B2(n20611), .A(n20610), .ZN(n20613) );
  INV_X1 U22743 ( .A(n20613), .ZN(n22058) );
  AOI22_X1 U22744 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n20616) );
  AOI22_X1 U22745 ( .A1(n20625), .A2(n22221), .B1(n20614), .B2(n22220), .ZN(
        n20615) );
  OAI211_X1 U22746 ( .C1(n22058), .C2(n22280), .A(n20616), .B(n20615), .ZN(
        P1_U2987) );
  NOR2_X1 U22747 ( .A1(n20617), .A2(n22078), .ZN(n20623) );
  OAI21_X1 U22748 ( .B1(n20620), .B2(n20619), .A(n20618), .ZN(n20621) );
  MUX2_X1 U22749 ( .A(n20623), .B(n20622), .S(n20621), .Z(n20624) );
  XOR2_X1 U22750 ( .A(n14281), .B(n20624), .Z(n22085) );
  AOI22_X1 U22751 ( .A1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n20627) );
  AOI22_X1 U22752 ( .A1(n22257), .A2(n20614), .B1(n22252), .B2(n20625), .ZN(
        n20626) );
  OAI211_X1 U22753 ( .C1(n22085), .C2(n22280), .A(n20627), .B(n20626), .ZN(
        P1_U2982) );
  AOI22_X1 U22754 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n20628), .B1(
        n22108), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n20633) );
  OAI22_X1 U22755 ( .A1(n22269), .A2(n20630), .B1(n20629), .B2(n22280), .ZN(
        n20631) );
  INV_X1 U22756 ( .A(n20631), .ZN(n20632) );
  OAI211_X1 U22757 ( .C1(n20634), .C2(n22266), .A(n20633), .B(n20632), .ZN(
        P1_U2980) );
  OAI21_X1 U22758 ( .B1(n20635), .B2(n22303), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20636) );
  OAI21_X1 U22759 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20637), .A(n20636), 
        .ZN(P1_U2803) );
  AOI21_X1 U22760 ( .B1(n22335), .B2(n22343), .A(P1_D_C_N_REG_SCAN_IN), .ZN(
        n20638) );
  AOI22_X1 U22761 ( .A1(n22853), .A2(P1_CODEFETCH_REG_SCAN_IN), .B1(n20638), 
        .B2(n22850), .ZN(P1_U2804) );
  INV_X1 U22762 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20641) );
  INV_X2 U22763 ( .A(U212), .ZN(n20682) );
  AOI22_X1 U22764 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n20695), .ZN(n20640) );
  OAI21_X1 U22765 ( .B1(n20641), .B2(n20680), .A(n20640), .ZN(U247) );
  AOI22_X1 U22766 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20695), .ZN(n20642) );
  OAI21_X1 U22767 ( .B1(n14743), .B2(n20680), .A(n20642), .ZN(U246) );
  AOI22_X1 U22768 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n20695), .ZN(n20643) );
  OAI21_X1 U22769 ( .B1(n14664), .B2(n20680), .A(n20643), .ZN(U245) );
  AOI22_X1 U22770 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20695), .ZN(n20644) );
  OAI21_X1 U22771 ( .B1(n14775), .B2(n20680), .A(n20644), .ZN(U244) );
  INV_X1 U22772 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U22773 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n20695), .ZN(n20645) );
  OAI21_X1 U22774 ( .B1(n20646), .B2(n20680), .A(n20645), .ZN(U243) );
  AOI22_X1 U22775 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20695), .ZN(n20647) );
  OAI21_X1 U22776 ( .B1(n14822), .B2(n20680), .A(n20647), .ZN(U242) );
  INV_X1 U22777 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20649) );
  AOI22_X1 U22778 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20695), .ZN(n20648) );
  OAI21_X1 U22779 ( .B1(n20649), .B2(n20680), .A(n20648), .ZN(U241) );
  AOI22_X1 U22780 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20695), .ZN(n20650) );
  OAI21_X1 U22781 ( .B1(n14786), .B2(n20680), .A(n20650), .ZN(U240) );
  AOI22_X1 U22782 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n20695), .ZN(n20651) );
  OAI21_X1 U22783 ( .B1(n15301), .B2(n20680), .A(n20651), .ZN(U239) );
  AOI22_X1 U22784 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20695), .ZN(n20652) );
  OAI21_X1 U22785 ( .B1(n20653), .B2(n20680), .A(n20652), .ZN(U238) );
  AOI22_X1 U22786 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n20695), .ZN(n20654) );
  OAI21_X1 U22787 ( .B1(n20655), .B2(n20680), .A(n20654), .ZN(U237) );
  AOI22_X1 U22788 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20695), .ZN(n20656) );
  OAI21_X1 U22789 ( .B1(n20657), .B2(n20680), .A(n20656), .ZN(U236) );
  AOI22_X1 U22790 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20695), .ZN(n20658) );
  OAI21_X1 U22791 ( .B1(n20659), .B2(n20680), .A(n20658), .ZN(U235) );
  AOI22_X1 U22792 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20695), .ZN(n20660) );
  OAI21_X1 U22793 ( .B1(n20661), .B2(n20680), .A(n20660), .ZN(U234) );
  INV_X1 U22794 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n20663) );
  AOI22_X1 U22795 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20695), .ZN(n20662) );
  OAI21_X1 U22796 ( .B1(n20663), .B2(n20680), .A(n20662), .ZN(U233) );
  AOI22_X1 U22797 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20695), .ZN(n20664) );
  OAI21_X1 U22798 ( .B1(n14494), .B2(n20680), .A(n20664), .ZN(U232) );
  INV_X1 U22799 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20666) );
  AOI22_X1 U22800 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n20695), .ZN(n20665) );
  OAI21_X1 U22801 ( .B1(n20666), .B2(n20680), .A(n20665), .ZN(U231) );
  INV_X1 U22802 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20668) );
  AOI22_X1 U22803 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n20695), .ZN(n20667) );
  OAI21_X1 U22804 ( .B1(n20668), .B2(n20680), .A(n20667), .ZN(U230) );
  INV_X1 U22805 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20670) );
  AOI22_X1 U22806 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20695), .ZN(n20669) );
  OAI21_X1 U22807 ( .B1(n20670), .B2(n20680), .A(n20669), .ZN(U229) );
  INV_X1 U22808 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20672) );
  AOI22_X1 U22809 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n20695), .ZN(n20671) );
  OAI21_X1 U22810 ( .B1(n20672), .B2(n20680), .A(n20671), .ZN(U228) );
  INV_X1 U22811 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20674) );
  AOI22_X1 U22812 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n20695), .ZN(n20673) );
  OAI21_X1 U22813 ( .B1(n20674), .B2(n20680), .A(n20673), .ZN(U227) );
  INV_X1 U22814 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20676) );
  AOI22_X1 U22815 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n20695), .ZN(n20675) );
  OAI21_X1 U22816 ( .B1(n20676), .B2(n20680), .A(n20675), .ZN(U226) );
  INV_X1 U22817 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20678) );
  AOI22_X1 U22818 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n20695), .ZN(n20677) );
  OAI21_X1 U22819 ( .B1(n20678), .B2(n20680), .A(n20677), .ZN(U225) );
  AOI22_X1 U22820 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n20695), .ZN(n20679) );
  OAI21_X1 U22821 ( .B1(n20681), .B2(n20680), .A(n20679), .ZN(U224) );
  INV_X1 U22822 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20684) );
  AOI22_X1 U22823 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n20695), .ZN(n20683) );
  OAI21_X1 U22824 ( .B1(n20684), .B2(n20680), .A(n20683), .ZN(U223) );
  INV_X1 U22825 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20686) );
  AOI22_X1 U22826 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n20695), .ZN(n20685) );
  OAI21_X1 U22827 ( .B1(n20686), .B2(n20680), .A(n20685), .ZN(U222) );
  AOI22_X1 U22828 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n20695), .ZN(n20687) );
  OAI21_X1 U22829 ( .B1(n20688), .B2(n20680), .A(n20687), .ZN(U221) );
  INV_X1 U22830 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20690) );
  AOI22_X1 U22831 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n20695), .ZN(n20689) );
  OAI21_X1 U22832 ( .B1(n20690), .B2(n20680), .A(n20689), .ZN(U220) );
  INV_X1 U22833 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20692) );
  AOI22_X1 U22834 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20695), .ZN(n20691) );
  OAI21_X1 U22835 ( .B1(n20692), .B2(n20680), .A(n20691), .ZN(U219) );
  INV_X1 U22836 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20694) );
  AOI22_X1 U22837 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n20695), .ZN(n20693) );
  OAI21_X1 U22838 ( .B1(n20694), .B2(n20680), .A(n20693), .ZN(U218) );
  INV_X1 U22839 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U22840 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n20682), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n20695), .ZN(n20696) );
  OAI21_X1 U22841 ( .B1(n20697), .B2(n20680), .A(n20696), .ZN(U217) );
  INV_X1 U22842 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20699) );
  OAI222_X1 U22843 ( .A1(U214), .A2(n20700), .B1(n20680), .B2(n20699), .C1(
        U212), .C2(n20698), .ZN(U216) );
  OAI22_X1 U22844 ( .A1(n22850), .A2(n20701), .B1(P1_W_R_N_REG_SCAN_IN), .B2(
        n22853), .ZN(n20702) );
  INV_X1 U22845 ( .A(n20702), .ZN(P1_U3483) );
  OAI21_X1 U22846 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n21435), .A(n21436), 
        .ZN(n20703) );
  INV_X1 U22847 ( .A(n22370), .ZN(n22321) );
  AOI211_X1 U22848 ( .C1(n20704), .C2(n20703), .A(n22321), .B(n21915), .ZN(
        n20705) );
  OAI21_X1 U22849 ( .B1(n20705), .B2(n21936), .A(n21927), .ZN(n20709) );
  AOI21_X1 U22850 ( .B1(n22370), .B2(n21871), .A(n20767), .ZN(n20706) );
  OAI21_X1 U22851 ( .B1(n20707), .B2(n21932), .A(n20706), .ZN(n20708) );
  MUX2_X1 U22852 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20709), .S(n20708), 
        .Z(P3_U3296) );
  INV_X1 U22853 ( .A(n20711), .ZN(n20713) );
  NOR2_X4 U22854 ( .A1(n20713), .A2(n21193), .ZN(n20750) );
  AOI22_X1 U22855 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20732), .ZN(n20715) );
  OAI21_X1 U22856 ( .B1(n20716), .B2(n20763), .A(n20715), .ZN(P3_U2768) );
  AOI22_X1 U22857 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20732), .ZN(n20717) );
  OAI21_X1 U22858 ( .B1(n20718), .B2(n20763), .A(n20717), .ZN(P3_U2769) );
  AOI22_X1 U22859 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20732), .ZN(n20719) );
  OAI21_X1 U22860 ( .B1(n20720), .B2(n20763), .A(n20719), .ZN(P3_U2770) );
  AOI22_X1 U22861 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20732), .ZN(n20721) );
  OAI21_X1 U22862 ( .B1(n20722), .B2(n20763), .A(n20721), .ZN(P3_U2771) );
  AOI22_X1 U22863 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20732), .ZN(n20723) );
  OAI21_X1 U22864 ( .B1(n21265), .B2(n20763), .A(n20723), .ZN(P3_U2772) );
  AOI22_X1 U22865 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20732), .ZN(n20724) );
  OAI21_X1 U22866 ( .B1(n21291), .B2(n20763), .A(n20724), .ZN(P3_U2773) );
  AOI22_X1 U22867 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20732), .ZN(n20725) );
  OAI21_X1 U22868 ( .B1(n21292), .B2(n20763), .A(n20725), .ZN(P3_U2774) );
  AOI22_X1 U22869 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20732), .ZN(n20726) );
  OAI21_X1 U22870 ( .B1(n20727), .B2(n20763), .A(n20726), .ZN(P3_U2775) );
  AOI22_X1 U22871 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20732), .ZN(n20728) );
  OAI21_X1 U22872 ( .B1(n20729), .B2(n20763), .A(n20728), .ZN(P3_U2776) );
  AOI22_X1 U22873 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20732), .ZN(n20730) );
  OAI21_X1 U22874 ( .B1(n20731), .B2(n20763), .A(n20730), .ZN(P3_U2777) );
  AOI22_X1 U22875 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20761), .ZN(n20733) );
  OAI21_X1 U22876 ( .B1(n21300), .B2(n20763), .A(n20733), .ZN(P3_U2778) );
  AOI22_X1 U22877 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20761), .ZN(n20734) );
  OAI21_X1 U22878 ( .B1(n20735), .B2(n20763), .A(n20734), .ZN(P3_U2779) );
  AOI22_X1 U22879 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20761), .ZN(n20736) );
  OAI21_X1 U22880 ( .B1(n20737), .B2(n20763), .A(n20736), .ZN(P3_U2780) );
  AOI22_X1 U22881 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20761), .ZN(n20738) );
  OAI21_X1 U22882 ( .B1(n21312), .B2(n20763), .A(n20738), .ZN(P3_U2781) );
  AOI22_X1 U22883 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20750), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20761), .ZN(n20739) );
  OAI21_X1 U22884 ( .B1(n20740), .B2(n20763), .A(n20739), .ZN(P3_U2782) );
  AOI22_X1 U22885 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20761), .ZN(n20741) );
  OAI21_X1 U22886 ( .B1(n21380), .B2(n20763), .A(n20741), .ZN(P3_U2783) );
  AOI22_X1 U22887 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20761), .ZN(n20742) );
  OAI21_X1 U22888 ( .B1(n21367), .B2(n20763), .A(n20742), .ZN(P3_U2784) );
  AOI22_X1 U22889 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20761), .ZN(n20743) );
  OAI21_X1 U22890 ( .B1(n21244), .B2(n20763), .A(n20743), .ZN(P3_U2785) );
  AOI22_X1 U22891 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20761), .ZN(n20744) );
  OAI21_X1 U22892 ( .B1(n21235), .B2(n20763), .A(n20744), .ZN(P3_U2786) );
  AOI22_X1 U22893 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20761), .ZN(n20745) );
  OAI21_X1 U22894 ( .B1(n21219), .B2(n20763), .A(n20745), .ZN(P3_U2787) );
  AOI22_X1 U22895 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20761), .ZN(n20746) );
  OAI21_X1 U22896 ( .B1(n20747), .B2(n20763), .A(n20746), .ZN(P3_U2788) );
  AOI22_X1 U22897 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20761), .ZN(n20748) );
  OAI21_X1 U22898 ( .B1(n20749), .B2(n20763), .A(n20748), .ZN(P3_U2789) );
  AOI22_X1 U22899 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20761), .ZN(n20751) );
  OAI21_X1 U22900 ( .B1(n21195), .B2(n20763), .A(n20751), .ZN(P3_U2790) );
  AOI22_X1 U22901 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20761), .ZN(n20752) );
  OAI21_X1 U22902 ( .B1(n21252), .B2(n20763), .A(n20752), .ZN(P3_U2791) );
  AOI22_X1 U22903 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20761), .ZN(n20753) );
  OAI21_X1 U22904 ( .B1(n21213), .B2(n20763), .A(n20753), .ZN(P3_U2792) );
  AOI22_X1 U22905 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20761), .ZN(n20754) );
  OAI21_X1 U22906 ( .B1(n20755), .B2(n20763), .A(n20754), .ZN(P3_U2793) );
  AOI22_X1 U22907 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20761), .ZN(n20756) );
  OAI21_X1 U22908 ( .B1(n21251), .B2(n20763), .A(n20756), .ZN(P3_U2794) );
  AOI22_X1 U22909 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20761), .ZN(n20757) );
  OAI21_X1 U22910 ( .B1(n20758), .B2(n20763), .A(n20757), .ZN(P3_U2795) );
  AOI22_X1 U22911 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20761), .ZN(n20759) );
  OAI21_X1 U22912 ( .B1(n21253), .B2(n20763), .A(n20759), .ZN(P3_U2796) );
  AOI22_X1 U22913 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20761), .ZN(n20760) );
  OAI21_X1 U22914 ( .B1(n21353), .B2(n20763), .A(n20760), .ZN(P3_U2797) );
  AOI22_X1 U22915 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20750), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20761), .ZN(n20762) );
  OAI21_X1 U22916 ( .B1(n21360), .B2(n20763), .A(n20762), .ZN(P3_U2798) );
  NOR2_X1 U22917 ( .A1(n21385), .A2(n21392), .ZN(n21413) );
  NOR2_X1 U22918 ( .A1(n20764), .A2(n21413), .ZN(n21390) );
  INV_X1 U22919 ( .A(n21390), .ZN(n21386) );
  NAND2_X1 U22920 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n21435), .ZN(n20765) );
  AOI211_X4 U22921 ( .C1(n22370), .C2(n22314), .A(n20770), .B(n20765), .ZN(
        n21141) );
  AND2_X1 U22922 ( .A1(n21917), .A2(n20766), .ZN(n21930) );
  NOR4_X2 U22923 ( .A1(n21866), .A2(n20767), .A3(n11264), .A4(n21930), .ZN(
        n20940) );
  AOI22_X1 U22924 ( .A1(n21141), .A2(n20768), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n20940), .ZN(n20775) );
  INV_X1 U22925 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20861) );
  NAND2_X1 U22926 ( .A1(n21155), .A2(n11264), .ZN(n20802) );
  INV_X1 U22927 ( .A(n20940), .ZN(n21187) );
  OAI21_X1 U22928 ( .B1(n20861), .B2(n20802), .A(n21168), .ZN(n20773) );
  INV_X1 U22929 ( .A(n11264), .ZN(n21920) );
  AOI21_X1 U22930 ( .B1(n21155), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n21920), .ZN(n20876) );
  OAI211_X1 U22931 ( .C1(n21436), .C2(n21435), .A(n22370), .B(n22314), .ZN(
        n20769) );
  INV_X1 U22932 ( .A(n20769), .ZN(n21914) );
  AOI211_X4 U22933 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n21435), .A(n21914), .B(
        n20770), .ZN(n21161) );
  OAI22_X1 U22934 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n21102), .B1(n21184), 
        .B2(n20771), .ZN(n20772) );
  AOI221_X1 U22935 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20773), .C1(
        n11315), .C2(n20876), .A(n20772), .ZN(n20774) );
  OAI211_X1 U22936 ( .C1(n21386), .C2(n21190), .A(n20775), .B(n20774), .ZN(
        P3_U2670) );
  NOR2_X1 U22937 ( .A1(n21920), .A2(n21155), .ZN(n20922) );
  INV_X1 U22938 ( .A(n20922), .ZN(n20983) );
  NOR3_X1 U22939 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20797) );
  AOI211_X1 U22940 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20776), .A(n20797), .B(
        n21183), .ZN(n20781) );
  NOR2_X1 U22941 ( .A1(n21413), .A2(n21891), .ZN(n21406) );
  NOR2_X1 U22942 ( .A1(n20777), .A2(n21406), .ZN(n21399) );
  AOI22_X1 U22943 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n21159), .B1(
        P3_REIP_REG_2__SCAN_IN), .B2(n20940), .ZN(n20779) );
  NAND2_X1 U22944 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .ZN(n20788) );
  OAI211_X1 U22945 ( .C1(P3_REIP_REG_2__SCAN_IN), .C2(P3_REIP_REG_1__SCAN_IN), 
        .A(n20941), .B(n20788), .ZN(n20778) );
  OAI211_X1 U22946 ( .C1(n21399), .C2(n21190), .A(n20779), .B(n20778), .ZN(
        n20780) );
  AOI211_X1 U22947 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n21161), .A(n20781), .B(
        n20780), .ZN(n20784) );
  NAND2_X1 U22948 ( .A1(n20861), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20978) );
  INV_X1 U22949 ( .A(n20978), .ZN(n20980) );
  OAI221_X1 U22950 ( .B1(n20980), .B2(n20785), .C1(n20978), .C2(n20782), .A(
        n21179), .ZN(n20783) );
  OAI211_X1 U22951 ( .C1(n20983), .C2(n20785), .A(n20784), .B(n20783), .ZN(
        P3_U2669) );
  OAI21_X1 U22952 ( .B1(n21385), .B2(n21408), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n21419) );
  NAND2_X1 U22953 ( .A1(n21419), .A2(n20786), .ZN(n21427) );
  NOR2_X1 U22954 ( .A1(n20793), .A2(n20788), .ZN(n20821) );
  NOR2_X1 U22955 ( .A1(n21102), .A2(n20821), .ZN(n20789) );
  INV_X1 U22956 ( .A(n20789), .ZN(n20787) );
  OAI22_X1 U22957 ( .A1(n21184), .A2(n20796), .B1(n20788), .B2(n20787), .ZN(
        n20795) );
  NOR2_X1 U22958 ( .A1(n20940), .A2(n20789), .ZN(n20817) );
  AOI21_X1 U22959 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20980), .A(
        n20860), .ZN(n20791) );
  XOR2_X1 U22960 ( .A(n20791), .B(n20790), .Z(n20792) );
  OAI22_X1 U22961 ( .A1(n20817), .A2(n20793), .B1(n21920), .B2(n20792), .ZN(
        n20794) );
  AOI211_X1 U22962 ( .C1(n20803), .C2(n21427), .A(n20795), .B(n20794), .ZN(
        n20799) );
  NAND2_X1 U22963 ( .A1(n20797), .A2(n20796), .ZN(n20801) );
  OAI211_X1 U22964 ( .C1(n20797), .C2(n20796), .A(n21141), .B(n20801), .ZN(
        n20798) );
  OAI211_X1 U22965 ( .C1(n21168), .C2(n20800), .A(n20799), .B(n20798), .ZN(
        P3_U2668) );
  NOR2_X1 U22966 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20801), .ZN(n20824) );
  AOI211_X1 U22967 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20801), .A(n20824), .B(
        n21183), .ZN(n20811) );
  AOI211_X1 U22968 ( .C1(n20818), .C2(n20861), .A(n20812), .B(n20802), .ZN(
        n20810) );
  INV_X1 U22969 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n20806) );
  OAI21_X1 U22970 ( .B1(n20804), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n20803), .ZN(n20805) );
  OAI211_X1 U22971 ( .C1(n21184), .C2(n20806), .A(n21822), .B(n20805), .ZN(
        n20809) );
  NAND3_X1 U22972 ( .A1(n20941), .A2(n20821), .A3(n20816), .ZN(n20807) );
  OAI21_X1 U22973 ( .B1(n21168), .B2(n20813), .A(n20807), .ZN(n20808) );
  NOR4_X1 U22974 ( .A1(n20811), .A2(n20810), .A3(n20809), .A4(n20808), .ZN(
        n20815) );
  OAI211_X1 U22975 ( .C1(n20922), .C2(n20813), .A(n20812), .B(n20876), .ZN(
        n20814) );
  OAI211_X1 U22976 ( .C1(n20817), .C2(n20816), .A(n20815), .B(n20814), .ZN(
        P3_U2667) );
  AOI21_X1 U22977 ( .B1(n20818), .B2(n20861), .A(n20860), .ZN(n20820) );
  XOR2_X1 U22978 ( .A(n20820), .B(n20819), .Z(n20831) );
  AOI22_X1 U22979 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_5__SCAN_IN), .ZN(n20830) );
  NAND2_X1 U22980 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n20821), .ZN(n20827) );
  NOR2_X1 U22981 ( .A1(n20822), .A2(n20827), .ZN(n20845) );
  OAI21_X1 U22982 ( .B1(n20845), .B2(n21102), .A(n21187), .ZN(n20853) );
  INV_X1 U22983 ( .A(n20845), .ZN(n20832) );
  NAND2_X1 U22984 ( .A1(n20941), .A2(n20832), .ZN(n20826) );
  NAND2_X1 U22985 ( .A1(n20824), .A2(n20823), .ZN(n20833) );
  OAI211_X1 U22986 ( .C1(n20824), .C2(n20823), .A(n21141), .B(n20833), .ZN(
        n20825) );
  OAI211_X1 U22987 ( .C1(n20827), .C2(n20826), .A(n21822), .B(n20825), .ZN(
        n20828) );
  AOI21_X1 U22988 ( .B1(P3_REIP_REG_5__SCAN_IN), .B2(n20853), .A(n20828), .ZN(
        n20829) );
  OAI211_X1 U22989 ( .C1(n21920), .C2(n20831), .A(n20830), .B(n20829), .ZN(
        P3_U2666) );
  NOR3_X1 U22990 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n21102), .A3(n20832), .ZN(
        n20854) );
  AOI211_X1 U22991 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n21159), .A(
        n21866), .B(n20854), .ZN(n20841) );
  NOR2_X1 U22992 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20833), .ZN(n20848) );
  AOI211_X1 U22993 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20833), .A(n20848), .B(
        n21183), .ZN(n20834) );
  AOI21_X1 U22994 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n21161), .A(n20834), .ZN(
        n20840) );
  AOI21_X1 U22995 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20983), .A(
        n20837), .ZN(n20835) );
  AOI22_X1 U22996 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20853), .B1(n20835), 
        .B2(n20876), .ZN(n20839) );
  NAND2_X1 U22997 ( .A1(n11159), .A2(n20980), .ZN(n20842) );
  NAND3_X1 U22998 ( .A1(n21179), .A2(n20837), .A3(n20842), .ZN(n20838) );
  NAND4_X1 U22999 ( .A1(n20841), .A2(n20840), .A3(n20839), .A4(n20838), .ZN(
        P3_U2665) );
  NAND2_X1 U23000 ( .A1(n21155), .A2(n20842), .ZN(n20844) );
  XOR2_X1 U23001 ( .A(n20844), .B(n20843), .Z(n20856) );
  NAND2_X1 U23002 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20845), .ZN(n20858) );
  NOR3_X1 U23003 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n21102), .A3(n20858), .ZN(
        n20846) );
  AOI211_X1 U23004 ( .C1(n21161), .C2(P3_EBX_REG_7__SCAN_IN), .A(n21866), .B(
        n20846), .ZN(n20850) );
  NAND2_X1 U23005 ( .A1(n20848), .A2(n20847), .ZN(n20857) );
  OAI211_X1 U23006 ( .C1(n20848), .C2(n20847), .A(n21141), .B(n20857), .ZN(
        n20849) );
  OAI211_X1 U23007 ( .C1(n21168), .C2(n20851), .A(n20850), .B(n20849), .ZN(
        n20852) );
  AOI221_X1 U23008 ( .B1(n20854), .B2(P3_REIP_REG_7__SCAN_IN), .C1(n20853), 
        .C2(P3_REIP_REG_7__SCAN_IN), .A(n20852), .ZN(n20855) );
  OAI21_X1 U23009 ( .B1(n20856), .B2(n21920), .A(n20855), .ZN(P3_U2664) );
  INV_X1 U23010 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20870) );
  NOR2_X1 U23011 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20857), .ZN(n20882) );
  OR2_X1 U23012 ( .A1(n21183), .A2(n20882), .ZN(n20872) );
  AOI21_X1 U23013 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n20857), .A(n20872), .ZN(
        n20868) );
  NOR2_X1 U23014 ( .A1(n21541), .A2(n20858), .ZN(n20859) );
  NAND2_X1 U23015 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n20859), .ZN(n20887) );
  AOI21_X1 U23016 ( .B1(n20941), .B2(n20887), .A(n20940), .ZN(n20896) );
  AOI21_X1 U23017 ( .B1(n20941), .B2(n20859), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n20866) );
  AOI21_X1 U23018 ( .B1(n20862), .B2(n20861), .A(n20860), .ZN(n20864) );
  XOR2_X1 U23019 ( .A(n20864), .B(n20863), .Z(n20865) );
  OAI22_X1 U23020 ( .A1(n20896), .A2(n20866), .B1(n21920), .B2(n20865), .ZN(
        n20867) );
  AOI211_X1 U23021 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n21161), .A(n20868), .B(
        n20867), .ZN(n20869) );
  OAI211_X1 U23022 ( .C1(n20870), .C2(n21168), .A(n20869), .B(n21822), .ZN(
        P3_U2663) );
  AOI21_X1 U23023 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n20983), .A(
        n20878), .ZN(n20877) );
  OAI22_X1 U23024 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20872), .B1(n20871), .B2(
        n21168), .ZN(n20875) );
  INV_X1 U23025 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20881) );
  AOI21_X1 U23026 ( .B1(n21141), .B2(n20882), .A(n21161), .ZN(n20873) );
  OAI22_X1 U23027 ( .A1(n20896), .A2(n20888), .B1(n20881), .B2(n20873), .ZN(
        n20874) );
  AOI211_X1 U23028 ( .C1(n20877), .C2(n20876), .A(n20875), .B(n20874), .ZN(
        n20880) );
  OAI211_X1 U23029 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20884), .A(
        n21179), .B(n20878), .ZN(n20879) );
  NAND4_X1 U23030 ( .A1(n20880), .A2(n21822), .A3(n20895), .A4(n20879), .ZN(
        P3_U2662) );
  NAND2_X1 U23031 ( .A1(n20882), .A2(n20881), .ZN(n20883) );
  AOI211_X1 U23032 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20883), .A(n20905), .B(
        n21183), .ZN(n20893) );
  OAI21_X1 U23033 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20884), .A(
        n21155), .ZN(n20885) );
  XNOR2_X1 U23034 ( .A(n20886), .B(n20885), .ZN(n20891) );
  NOR2_X1 U23035 ( .A1(n20888), .A2(n20887), .ZN(n20898) );
  NOR2_X1 U23036 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n21102), .ZN(n20889) );
  AOI22_X1 U23037 ( .A1(n21161), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n20898), 
        .B2(n20889), .ZN(n20890) );
  OAI211_X1 U23038 ( .C1(n21920), .C2(n20891), .A(n20890), .B(n21822), .ZN(
        n20892) );
  AOI211_X1 U23039 ( .C1(n21159), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20893), .B(n20892), .ZN(n20894) );
  OAI221_X1 U23040 ( .B1(n20897), .B2(n20896), .C1(n20897), .C2(n20895), .A(
        n20894), .ZN(P3_U2661) );
  INV_X1 U23041 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20911) );
  NAND2_X1 U23042 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n20898), .ZN(n20900) );
  NOR2_X1 U23043 ( .A1(n20899), .A2(n20900), .ZN(n20912) );
  OAI21_X1 U23044 ( .B1(n21102), .B2(n20912), .A(n21187), .ZN(n20977) );
  OAI21_X1 U23045 ( .B1(n21102), .B2(n20900), .A(n20899), .ZN(n20909) );
  OAI21_X1 U23046 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20901), .A(
        n21155), .ZN(n20903) );
  AOI21_X1 U23047 ( .B1(n20904), .B2(n20903), .A(n21920), .ZN(n20902) );
  OAI21_X1 U23048 ( .B1(n20904), .B2(n20903), .A(n20902), .ZN(n20907) );
  NAND2_X1 U23049 ( .A1(n20905), .A2(n20911), .ZN(n20917) );
  OAI211_X1 U23050 ( .C1(n20905), .C2(n20911), .A(n21141), .B(n20917), .ZN(
        n20906) );
  OAI211_X1 U23051 ( .C1(n21168), .C2(n11310), .A(n20907), .B(n20906), .ZN(
        n20908) );
  AOI21_X1 U23052 ( .B1(n20977), .B2(n20909), .A(n20908), .ZN(n20910) );
  OAI211_X1 U23053 ( .C1(n21184), .C2(n20911), .A(n20910), .B(n21822), .ZN(
        P3_U2660) );
  INV_X1 U23054 ( .A(n20977), .ZN(n21059) );
  NOR2_X1 U23055 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n21046), .ZN(n20932) );
  AOI211_X1 U23056 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n21159), .A(
        n21866), .B(n20932), .ZN(n20921) );
  OAI21_X1 U23057 ( .B1(n20913), .B2(n20978), .A(n21155), .ZN(n20915) );
  OAI21_X1 U23058 ( .B1(n20916), .B2(n20915), .A(n11264), .ZN(n20914) );
  AOI21_X1 U23059 ( .B1(n20916), .B2(n20915), .A(n20914), .ZN(n20919) );
  AOI211_X1 U23060 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20917), .A(n20927), .B(
        n21183), .ZN(n20918) );
  AOI211_X1 U23061 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n21161), .A(n20919), .B(
        n20918), .ZN(n20920) );
  OAI211_X1 U23062 ( .C1(n21059), .C2(n20925), .A(n20921), .B(n20920), .ZN(
        P3_U2659) );
  NOR2_X1 U23063 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21920), .ZN(
        n20924) );
  INV_X1 U23064 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20923) );
  AOI21_X1 U23065 ( .B1(n20924), .B2(n20923), .A(n20922), .ZN(n20936) );
  NOR3_X1 U23066 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n20925), .A3(n21046), 
        .ZN(n20926) );
  AOI211_X1 U23067 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n21159), .A(
        n21866), .B(n20926), .ZN(n20934) );
  INV_X1 U23068 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20930) );
  OAI211_X1 U23069 ( .C1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n20937), .A(
        n21179), .B(n20935), .ZN(n20929) );
  NAND2_X1 U23070 ( .A1(n20927), .A2(n20930), .ZN(n20944) );
  OAI211_X1 U23071 ( .C1(n20927), .C2(n20930), .A(n21141), .B(n20944), .ZN(
        n20928) );
  OAI211_X1 U23072 ( .C1(n20930), .C2(n21184), .A(n20929), .B(n20928), .ZN(
        n20931) );
  AOI221_X1 U23073 ( .B1(n20932), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n20977), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n20931), .ZN(n20933) );
  OAI211_X1 U23074 ( .C1(n20936), .C2(n20935), .A(n20934), .B(n20933), .ZN(
        P3_U2658) );
  OAI21_X1 U23075 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20937), .A(
        n21155), .ZN(n20938) );
  XOR2_X1 U23076 ( .A(n20939), .B(n20938), .Z(n20949) );
  AOI21_X1 U23077 ( .B1(n21161), .B2(P3_EBX_REG_14__SCAN_IN), .A(n21866), .ZN(
        n20948) );
  NAND2_X1 U23078 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_12__SCAN_IN), 
        .ZN(n20943) );
  NOR2_X1 U23079 ( .A1(n20942), .A2(n20943), .ZN(n20969) );
  NOR2_X1 U23080 ( .A1(n20941), .A2(n20940), .ZN(n21060) );
  OAI21_X1 U23081 ( .B1(n20969), .B2(n21060), .A(n21059), .ZN(n20957) );
  INV_X1 U23082 ( .A(n20957), .ZN(n20967) );
  AOI221_X1 U23083 ( .B1(n20943), .B2(n20942), .C1(n21046), .C2(n20942), .A(
        n20967), .ZN(n20946) );
  AOI211_X1 U23084 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20944), .A(n20959), .B(
        n21183), .ZN(n20945) );
  AOI211_X1 U23085 ( .C1(n21159), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20946), .B(n20945), .ZN(n20947) );
  OAI211_X1 U23086 ( .C1(n21920), .C2(n20949), .A(n20948), .B(n20947), .ZN(
        P3_U2657) );
  OAI21_X1 U23087 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20950), .A(
        n21155), .ZN(n20952) );
  OAI21_X1 U23088 ( .B1(n20953), .B2(n20952), .A(n11264), .ZN(n20951) );
  AOI21_X1 U23089 ( .B1(n20953), .B2(n20952), .A(n20951), .ZN(n20956) );
  INV_X1 U23090 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20958) );
  NAND3_X1 U23091 ( .A1(n20969), .A2(n21076), .A3(n20954), .ZN(n20966) );
  OAI211_X1 U23092 ( .C1(n21184), .C2(n20958), .A(n21822), .B(n20966), .ZN(
        n20955) );
  AOI211_X1 U23093 ( .C1(P3_REIP_REG_15__SCAN_IN), .C2(n20957), .A(n20956), 
        .B(n20955), .ZN(n20961) );
  NAND2_X1 U23094 ( .A1(n20959), .A2(n20958), .ZN(n20968) );
  OAI211_X1 U23095 ( .C1(n20959), .C2(n20958), .A(n21141), .B(n20968), .ZN(
        n20960) );
  OAI211_X1 U23096 ( .C1(n21168), .C2(n20962), .A(n20961), .B(n20960), .ZN(
        P3_U2656) );
  OAI21_X1 U23097 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20963), .A(
        n21155), .ZN(n20964) );
  XOR2_X1 U23098 ( .A(n20965), .B(n20964), .Z(n20975) );
  AOI22_X1 U23099 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n20974) );
  AOI21_X1 U23100 ( .B1(n20967), .B2(n20966), .A(n21837), .ZN(n20972) );
  AOI211_X1 U23101 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20968), .A(n20991), .B(
        n21183), .ZN(n20971) );
  NAND2_X1 U23102 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n20969), .ZN(n20976) );
  NOR3_X1 U23103 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20976), .A3(n21046), 
        .ZN(n20970) );
  NOR4_X1 U23104 ( .A1(n21866), .A2(n20972), .A3(n20971), .A4(n20970), .ZN(
        n20973) );
  OAI211_X1 U23105 ( .C1(n21920), .C2(n20975), .A(n20974), .B(n20973), .ZN(
        P3_U2655) );
  INV_X1 U23106 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n20994) );
  NOR2_X1 U23107 ( .A1(n21837), .A2(n20976), .ZN(n20986) );
  NAND2_X1 U23108 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n20986), .ZN(n21005) );
  INV_X1 U23109 ( .A(n21060), .ZN(n21185) );
  AOI21_X1 U23110 ( .B1(n21005), .B2(n21185), .A(n20977), .ZN(n21004) );
  INV_X1 U23111 ( .A(n21004), .ZN(n21009) );
  OAI21_X1 U23112 ( .B1(n20979), .B2(n20978), .A(n21155), .ZN(n20995) );
  OAI221_X1 U23113 ( .B1(n20984), .B2(n20981), .C1(n20984), .C2(n20980), .A(
        n11264), .ZN(n20982) );
  AOI22_X1 U23114 ( .A1(n20984), .A2(n20995), .B1(n20983), .B2(n20982), .ZN(
        n20989) );
  NAND3_X1 U23115 ( .A1(n20986), .A2(n21076), .A3(n20985), .ZN(n20987) );
  OAI211_X1 U23116 ( .C1(n21184), .C2(n20990), .A(n21822), .B(n20987), .ZN(
        n20988) );
  AOI211_X1 U23117 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n21009), .A(n20989), 
        .B(n20988), .ZN(n20993) );
  NAND2_X1 U23118 ( .A1(n20991), .A2(n20990), .ZN(n20999) );
  OAI211_X1 U23119 ( .C1(n20991), .C2(n20990), .A(n21141), .B(n20999), .ZN(
        n20992) );
  OAI211_X1 U23120 ( .C1(n21168), .C2(n20994), .A(n20993), .B(n20992), .ZN(
        P3_U2654) );
  NOR3_X1 U23121 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n21005), .A3(n21046), 
        .ZN(n21010) );
  AOI211_X1 U23122 ( .C1(n21161), .C2(P3_EBX_REG_18__SCAN_IN), .A(n21866), .B(
        n21010), .ZN(n21003) );
  INV_X1 U23123 ( .A(n20996), .ZN(n20998) );
  INV_X1 U23124 ( .A(n20995), .ZN(n20997) );
  AOI221_X1 U23125 ( .B1(n20998), .B2(n20997), .C1(n20996), .C2(n20995), .A(
        n21920), .ZN(n21001) );
  AOI211_X1 U23126 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20999), .A(n21015), .B(
        n21183), .ZN(n21000) );
  AOI211_X1 U23127 ( .C1(n21159), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n21001), .B(n21000), .ZN(n21002) );
  OAI211_X1 U23128 ( .C1(n21004), .C2(n21821), .A(n21003), .B(n21002), .ZN(
        P3_U2653) );
  NOR2_X1 U23129 ( .A1(n21821), .A2(n21005), .ZN(n21020) );
  NAND3_X1 U23130 ( .A1(n21020), .A2(n21076), .A3(n21006), .ZN(n21007) );
  OAI211_X1 U23131 ( .C1(n21184), .C2(n21014), .A(n21822), .B(n21007), .ZN(
        n21008) );
  AOI221_X1 U23132 ( .B1(n21010), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n21009), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n21008), .ZN(n21019) );
  OAI211_X1 U23133 ( .C1(n21013), .C2(n21012), .A(n11264), .B(n21026), .ZN(
        n21018) );
  NAND2_X1 U23134 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n21159), .ZN(
        n21017) );
  NAND2_X1 U23135 ( .A1(n21015), .A2(n21014), .ZN(n21022) );
  OAI211_X1 U23136 ( .C1(n21015), .C2(n21014), .A(n21141), .B(n21022), .ZN(
        n21016) );
  NAND4_X1 U23137 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        P3_U2652) );
  AOI22_X1 U23138 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n21031) );
  NAND2_X1 U23139 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n21020), .ZN(n21021) );
  NOR2_X1 U23140 ( .A1(n21021), .A2(n21046), .ZN(n21025) );
  NOR2_X1 U23141 ( .A1(n21801), .A2(n21021), .ZN(n21045) );
  OAI21_X1 U23142 ( .B1(n21045), .B2(n21060), .A(n21059), .ZN(n21024) );
  AOI211_X1 U23143 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n21022), .A(n21037), .B(
        n21183), .ZN(n21023) );
  AOI221_X1 U23144 ( .B1(n21025), .B2(n21801), .C1(n21024), .C2(
        P3_REIP_REG_20__SCAN_IN), .A(n21023), .ZN(n21030) );
  NAND2_X1 U23145 ( .A1(n21028), .A2(n21027), .ZN(n21034) );
  OAI211_X1 U23146 ( .C1(n21028), .C2(n21027), .A(n11264), .B(n21034), .ZN(
        n21029) );
  NAND3_X1 U23147 ( .A1(n21031), .A2(n21030), .A3(n21029), .ZN(P3_U2651) );
  NAND3_X1 U23148 ( .A1(n21045), .A2(n21076), .A3(n21032), .ZN(n21033) );
  OAI211_X1 U23149 ( .C1(n21045), .C2(n21060), .A(n21059), .B(n21033), .ZN(
        n21049) );
  NAND2_X1 U23150 ( .A1(n21033), .A2(n21032), .ZN(n21042) );
  NAND2_X1 U23151 ( .A1(n21155), .A2(n21034), .ZN(n21035) );
  NAND2_X1 U23152 ( .A1(n21036), .A2(n21035), .ZN(n21051) );
  OAI211_X1 U23153 ( .C1(n21036), .C2(n21035), .A(n11264), .B(n21051), .ZN(
        n21039) );
  NAND2_X1 U23154 ( .A1(n21037), .A2(n21044), .ZN(n21047) );
  OAI211_X1 U23155 ( .C1(n21037), .C2(n21044), .A(n21141), .B(n21047), .ZN(
        n21038) );
  OAI211_X1 U23156 ( .C1(n21168), .C2(n21040), .A(n21039), .B(n21038), .ZN(
        n21041) );
  AOI21_X1 U23157 ( .B1(n21049), .B2(n21042), .A(n21041), .ZN(n21043) );
  OAI21_X1 U23158 ( .B1(n21184), .B2(n21044), .A(n21043), .ZN(P3_U2650) );
  AOI22_X1 U23159 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n21056) );
  NAND2_X1 U23160 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n21045), .ZN(n21057) );
  NOR2_X1 U23161 ( .A1(n21057), .A2(n21046), .ZN(n21050) );
  NOR2_X1 U23162 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n21047), .ZN(n21067) );
  AOI211_X1 U23163 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n21047), .A(n21067), .B(
        n21183), .ZN(n21048) );
  AOI221_X1 U23164 ( .B1(n21050), .B2(n21058), .C1(n21049), .C2(
        P3_REIP_REG_22__SCAN_IN), .A(n21048), .ZN(n21055) );
  NAND2_X1 U23165 ( .A1(n21155), .A2(n21051), .ZN(n21052) );
  NAND2_X1 U23166 ( .A1(n21053), .A2(n21052), .ZN(n21063) );
  OAI211_X1 U23167 ( .C1(n21053), .C2(n21052), .A(n11264), .B(n21063), .ZN(
        n21054) );
  NAND3_X1 U23168 ( .A1(n21056), .A2(n21055), .A3(n21054), .ZN(P3_U2649) );
  NOR2_X1 U23169 ( .A1(n21058), .A2(n21057), .ZN(n21069) );
  AND2_X1 U23170 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n21069), .ZN(n21077) );
  OAI21_X1 U23171 ( .B1(n21077), .B2(n21060), .A(n21059), .ZN(n21088) );
  OAI22_X1 U23172 ( .A1(n21061), .A2(n21168), .B1(n21184), .B2(n21066), .ZN(
        n21062) );
  AOI21_X1 U23173 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(n21088), .A(n21062), 
        .ZN(n21073) );
  NAND2_X1 U23174 ( .A1(n21155), .A2(n21063), .ZN(n21065) );
  NAND2_X1 U23175 ( .A1(n21065), .A2(n21064), .ZN(n21080) );
  OAI211_X1 U23176 ( .C1(n21065), .C2(n21064), .A(n11264), .B(n21080), .ZN(
        n21072) );
  NAND2_X1 U23177 ( .A1(n21067), .A2(n21066), .ZN(n21074) );
  OAI211_X1 U23178 ( .C1(n21067), .C2(n21066), .A(n21141), .B(n21074), .ZN(
        n21071) );
  NAND3_X1 U23179 ( .A1(n21069), .A2(n21076), .A3(n21068), .ZN(n21070) );
  NAND4_X1 U23180 ( .A1(n21073), .A2(n21072), .A3(n21071), .A4(n21070), .ZN(
        P3_U2648) );
  NOR2_X1 U23181 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n21074), .ZN(n21094) );
  AOI21_X1 U23182 ( .B1(n21074), .B2(P3_EBX_REG_24__SCAN_IN), .A(n21183), .ZN(
        n21075) );
  AOI21_X1 U23183 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n21161), .A(n21075), .ZN(
        n21085) );
  NAND2_X1 U23184 ( .A1(n21077), .A2(n21076), .ZN(n21086) );
  NOR2_X1 U23185 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n21086), .ZN(n21089) );
  NOR2_X1 U23186 ( .A1(n21078), .A2(n21168), .ZN(n21079) );
  AOI211_X1 U23187 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n21088), .A(n21089), 
        .B(n21079), .ZN(n21084) );
  NAND2_X1 U23188 ( .A1(n21155), .A2(n21080), .ZN(n21081) );
  NAND2_X1 U23189 ( .A1(n21082), .A2(n21081), .ZN(n21090) );
  OAI211_X1 U23190 ( .C1(n21082), .C2(n21081), .A(n11264), .B(n21090), .ZN(
        n21083) );
  OAI211_X1 U23191 ( .C1(n21094), .C2(n21085), .A(n21084), .B(n21083), .ZN(
        P3_U2647) );
  NOR2_X1 U23192 ( .A1(n21089), .A2(n21088), .ZN(n21101) );
  AOI22_X1 U23193 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n21097) );
  NAND2_X1 U23194 ( .A1(n21155), .A2(n21090), .ZN(n21091) );
  NAND2_X1 U23195 ( .A1(n21092), .A2(n21091), .ZN(n21108) );
  OAI211_X1 U23196 ( .C1(n21092), .C2(n21091), .A(n11264), .B(n21108), .ZN(
        n21096) );
  NAND2_X1 U23197 ( .A1(n21094), .A2(n21093), .ZN(n21103) );
  OAI211_X1 U23198 ( .C1(n21094), .C2(n21093), .A(n21141), .B(n21103), .ZN(
        n21095) );
  AND3_X1 U23199 ( .A1(n21097), .A2(n21096), .A3(n21095), .ZN(n21098) );
  OAI221_X1 U23200 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n21116), .C1(n21099), 
        .C2(n21101), .A(n21098), .ZN(P3_U2646) );
  NAND2_X1 U23201 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n21100), .ZN(n21113) );
  NOR2_X1 U23202 ( .A1(n21100), .A2(n21099), .ZN(n21114) );
  OAI21_X1 U23203 ( .B1(n21114), .B2(n21102), .A(n21101), .ZN(n21138) );
  NOR2_X1 U23204 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n21103), .ZN(n21122) );
  AOI211_X1 U23205 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n21103), .A(n21122), .B(
        n21183), .ZN(n21107) );
  OAI22_X1 U23206 ( .A1(n21105), .A2(n21168), .B1(n21184), .B2(n21104), .ZN(
        n21106) );
  AOI211_X1 U23207 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n21138), .A(n21107), 
        .B(n21106), .ZN(n21112) );
  NAND2_X1 U23208 ( .A1(n21155), .A2(n21108), .ZN(n21110) );
  NAND2_X1 U23209 ( .A1(n21110), .A2(n21109), .ZN(n21118) );
  OAI211_X1 U23210 ( .C1(n21110), .C2(n21109), .A(n11264), .B(n21118), .ZN(
        n21111) );
  OAI211_X1 U23211 ( .C1(n21113), .C2(n21116), .A(n21112), .B(n21111), .ZN(
        P3_U2645) );
  AOI22_X1 U23212 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n21126) );
  INV_X1 U23213 ( .A(n21114), .ZN(n21115) );
  AOI22_X1 U23214 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n21138), .B1(n21156), 
        .B2(n21117), .ZN(n21125) );
  NAND2_X1 U23215 ( .A1(n21155), .A2(n21118), .ZN(n21119) );
  NAND2_X1 U23216 ( .A1(n21120), .A2(n21119), .ZN(n21130) );
  OAI211_X1 U23217 ( .C1(n21120), .C2(n21119), .A(n11264), .B(n21130), .ZN(
        n21124) );
  INV_X1 U23218 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n21121) );
  NAND2_X1 U23219 ( .A1(n21122), .A2(n21121), .ZN(n21127) );
  OAI211_X1 U23220 ( .C1(n21122), .C2(n21121), .A(n21141), .B(n21127), .ZN(
        n21123) );
  NAND4_X1 U23221 ( .A1(n21126), .A2(n21125), .A3(n21124), .A4(n21123), .ZN(
        P3_U2644) );
  AOI22_X1 U23222 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n21159), .B1(
        n21161), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n21137) );
  NOR2_X1 U23223 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n21127), .ZN(n21140) );
  AOI211_X1 U23224 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n21127), .A(n21140), .B(
        n21183), .ZN(n21128) );
  AOI21_X1 U23225 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n21138), .A(n21128), 
        .ZN(n21136) );
  INV_X1 U23226 ( .A(n21129), .ZN(n21132) );
  NAND2_X1 U23227 ( .A1(n21155), .A2(n21130), .ZN(n21131) );
  NAND2_X1 U23228 ( .A1(n21132), .A2(n21131), .ZN(n21147) );
  OAI211_X1 U23229 ( .C1(n21132), .C2(n21131), .A(n11264), .B(n21147), .ZN(
        n21135) );
  NAND2_X1 U23230 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n21133) );
  OAI211_X1 U23231 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n21156), .B(n21133), .ZN(n21134) );
  NAND4_X1 U23232 ( .A1(n21137), .A2(n21136), .A3(n21135), .A4(n21134), .ZN(
        P3_U2643) );
  NAND3_X1 U23233 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n21139) );
  AOI21_X1 U23234 ( .B1(n21139), .B2(n21185), .A(n21138), .ZN(n21174) );
  INV_X1 U23235 ( .A(n21140), .ZN(n21142) );
  NAND2_X1 U23236 ( .A1(n21140), .A2(n21144), .ZN(n21160) );
  NAND2_X1 U23237 ( .A1(n21141), .A2(n21160), .ZN(n21157) );
  AOI21_X1 U23238 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n21142), .A(n21157), .ZN(
        n21146) );
  NAND4_X1 U23239 ( .A1(n21156), .A2(P3_REIP_REG_28__SCAN_IN), .A3(
        P3_REIP_REG_27__SCAN_IN), .A4(n21153), .ZN(n21143) );
  OAI21_X1 U23240 ( .B1(n21144), .B2(n21184), .A(n21143), .ZN(n21145) );
  AOI211_X1 U23241 ( .C1(n21159), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n21146), .B(n21145), .ZN(n21152) );
  NAND2_X1 U23242 ( .A1(n21155), .A2(n21147), .ZN(n21149) );
  NAND2_X1 U23243 ( .A1(n21150), .A2(n21149), .ZN(n21154) );
  OAI211_X1 U23244 ( .C1(n21150), .C2(n21149), .A(n11264), .B(n21154), .ZN(
        n21151) );
  OAI211_X1 U23245 ( .C1(n21174), .C2(n21153), .A(n21152), .B(n21151), .ZN(
        P3_U2642) );
  NAND2_X1 U23246 ( .A1(n21155), .A2(n21154), .ZN(n21177) );
  XNOR2_X1 U23247 ( .A(n21178), .B(n21177), .ZN(n21164) );
  NAND4_X1 U23248 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n21156), .A3(
        P3_REIP_REG_29__SCAN_IN), .A4(P3_REIP_REG_27__SCAN_IN), .ZN(n21165) );
  NOR2_X1 U23249 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n21165), .ZN(n21176) );
  OAI22_X1 U23250 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n21157), .B1(n21174), 
        .B2(n21166), .ZN(n21158) );
  AOI211_X1 U23251 ( .C1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n21159), .A(
        n21176), .B(n21158), .ZN(n21163) );
  NOR2_X1 U23252 ( .A1(n21183), .A2(n21160), .ZN(n21173) );
  OAI21_X1 U23253 ( .B1(n21161), .B2(n21173), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n21162) );
  OAI211_X1 U23254 ( .C1(n21920), .C2(n21164), .A(n21163), .B(n21162), .ZN(
        P3_U2641) );
  INV_X1 U23255 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21172) );
  NOR3_X1 U23256 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n21166), .A3(n21165), 
        .ZN(n21171) );
  OAI22_X1 U23257 ( .A1(n21169), .A2(n21168), .B1(n21167), .B2(n21184), .ZN(
        n21170) );
  AOI211_X1 U23258 ( .C1(n21173), .C2(n21172), .A(n21171), .B(n21170), .ZN(
        n21182) );
  INV_X1 U23259 ( .A(n21174), .ZN(n21175) );
  OAI21_X1 U23260 ( .B1(n21176), .B2(n21175), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n21181) );
  NAND3_X1 U23261 ( .A1(n21179), .A2(n21178), .A3(n21177), .ZN(n21180) );
  NAND3_X1 U23262 ( .A1(n21182), .A2(n21181), .A3(n21180), .ZN(P3_U2640) );
  NAND2_X1 U23263 ( .A1(n21184), .A2(n21183), .ZN(n21186) );
  AOI22_X1 U23264 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n21186), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n21185), .ZN(n21189) );
  NAND3_X1 U23265 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n21187), .A3(
        n21402), .ZN(n21188) );
  OAI211_X1 U23266 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n21190), .A(
        n21189), .B(n21188), .ZN(P3_U2671) );
  NOR4_X1 U23267 ( .A1(n21219), .A2(n21235), .A3(n21367), .A4(n21195), .ZN(
        n21196) );
  NAND4_X1 U23268 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(n21196), .ZN(n21249) );
  NOR3_X1 U23269 ( .A1(n21294), .A2(n21369), .A3(n21249), .ZN(n21355) );
  NAND2_X1 U23270 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n21355), .ZN(n21362) );
  NAND2_X1 U23271 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21217), .ZN(n21208) );
  NOR2_X1 U23272 ( .A1(n21251), .A2(n21208), .ZN(n21202) );
  NAND2_X1 U23273 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n21202), .ZN(n21201) );
  NAND2_X1 U23274 ( .A1(n21201), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n21200) );
  NAND2_X1 U23275 ( .A1(n21379), .A2(n21197), .ZN(n21241) );
  AOI22_X1 U23276 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21377), .B1(n21376), .B2(
        n21198), .ZN(n21199) );
  OAI221_X1 U23277 ( .B1(n21201), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n21200), 
        .C2(n21313), .A(n21199), .ZN(P3_U2722) );
  INV_X1 U23278 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n21205) );
  INV_X1 U23279 ( .A(n21201), .ZN(n21349) );
  AOI21_X1 U23280 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n21370), .A(n21202), .ZN(
        n21204) );
  OAI222_X1 U23281 ( .A1(n21241), .A2(n21205), .B1(n21349), .B2(n21204), .C1(
        n21373), .C2(n21203), .ZN(P3_U2723) );
  NAND2_X1 U23282 ( .A1(n21370), .A2(n21208), .ZN(n21211) );
  AOI22_X1 U23283 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21377), .B1(n21376), .B2(
        n21206), .ZN(n21207) );
  OAI221_X1 U23284 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n21208), .C1(n21251), 
        .C2(n21211), .A(n21207), .ZN(P3_U2724) );
  INV_X1 U23285 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n21212) );
  NOR2_X1 U23286 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n21217), .ZN(n21210) );
  OAI222_X1 U23287 ( .A1(n21241), .A2(n21212), .B1(n21211), .B2(n21210), .C1(
        n21373), .C2(n21209), .ZN(P3_U2725) );
  INV_X1 U23288 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n21218) );
  OAI21_X1 U23289 ( .B1(n21213), .B2(n21313), .A(n21362), .ZN(n21214) );
  INV_X1 U23290 ( .A(n21214), .ZN(n21216) );
  OAI222_X1 U23291 ( .A1(n21241), .A2(n21218), .B1(n21217), .B2(n21216), .C1(
        n21373), .C2(n21215), .ZN(P3_U2726) );
  NAND2_X1 U23292 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n21220) );
  NOR2_X1 U23293 ( .A1(n21294), .A2(n21369), .ZN(n21368) );
  NAND2_X1 U23294 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n21368), .ZN(n21243) );
  NOR3_X1 U23295 ( .A1(n21219), .A2(n21235), .A3(n21246), .ZN(n21233) );
  INV_X1 U23296 ( .A(n21233), .ZN(n21230) );
  NOR2_X1 U23297 ( .A1(n21220), .A2(n21230), .ZN(n21225) );
  AOI21_X1 U23298 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n21370), .A(n21225), .ZN(
        n21221) );
  OAI222_X1 U23299 ( .A1(n21241), .A2(n21222), .B1(n21355), .B2(n21221), .C1(
        n21373), .C2(n21728), .ZN(P3_U2728) );
  AOI22_X1 U23300 ( .A1(n21233), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n21370), .ZN(n21224) );
  OAI222_X1 U23301 ( .A1(n21226), .A2(n21241), .B1(n21225), .B2(n21224), .C1(
        n21373), .C2(n21223), .ZN(P3_U2729) );
  NAND2_X1 U23302 ( .A1(n21230), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n21229) );
  AOI22_X1 U23303 ( .A1(n21377), .A2(BUF2_REG_5__SCAN_IN), .B1(n21376), .B2(
        n21227), .ZN(n21228) );
  OAI221_X1 U23304 ( .B1(n21230), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n21229), 
        .C2(n21313), .A(n21228), .ZN(P3_U2730) );
  AOI22_X1 U23305 ( .A1(n21236), .A2(P3_EAX_REG_3__SCAN_IN), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n21370), .ZN(n21232) );
  OAI222_X1 U23306 ( .A1(n21234), .A2(n21241), .B1(n21233), .B2(n21232), .C1(
        n21373), .C2(n21231), .ZN(P3_U2731) );
  NOR2_X1 U23307 ( .A1(n21235), .A2(n21246), .ZN(n21240) );
  AOI21_X1 U23308 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n21370), .A(n21236), .ZN(
        n21239) );
  INV_X1 U23309 ( .A(n21237), .ZN(n21238) );
  OAI222_X1 U23310 ( .A1(n21242), .A2(n21241), .B1(n21240), .B2(n21239), .C1(
        n21373), .C2(n21238), .ZN(P3_U2732) );
  OAI21_X1 U23311 ( .B1(n21313), .B2(n21244), .A(n21243), .ZN(n21245) );
  AOI22_X1 U23312 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21377), .B1(n21246), .B2(
        n21245), .ZN(n21247) );
  OAI21_X1 U23313 ( .B1(n21248), .B2(n21373), .A(n21247), .ZN(P3_U2733) );
  NAND4_X1 U23314 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_20__SCAN_IN), .ZN(n21293)
         );
  NAND4_X1 U23315 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n21250)
         );
  NOR4_X1 U23316 ( .A1(n21253), .A2(n21252), .A3(n21251), .A4(n21250), .ZN(
        n21356) );
  NOR2_X1 U23317 ( .A1(n21294), .A2(n21344), .ZN(n21286) );
  INV_X1 U23318 ( .A(n21286), .ZN(n21274) );
  NOR2_X1 U23319 ( .A1(n21293), .A2(n21274), .ZN(n21270) );
  INV_X1 U23320 ( .A(n21270), .ZN(n21260) );
  NAND2_X1 U23321 ( .A1(n21370), .A2(n21260), .ZN(n21268) );
  NOR2_X2 U23322 ( .A1(n21254), .A2(n21370), .ZN(n21343) );
  OAI22_X1 U23323 ( .A1(n21257), .A2(n21373), .B1(n21256), .B2(n21341), .ZN(
        n21258) );
  AOI21_X1 U23324 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n21343), .A(n21258), .ZN(
        n21259) );
  OAI221_X1 U23325 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21260), .C1(n21291), 
        .C2(n21268), .A(n21259), .ZN(P3_U2714) );
  NAND4_X1 U23326 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(n21286), .ZN(n21276) );
  INV_X1 U23327 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n21261) );
  OAI22_X1 U23328 ( .A1(n21262), .A2(n21373), .B1(n21261), .B2(n21341), .ZN(
        n21263) );
  AOI21_X1 U23329 ( .B1(BUF2_REG_4__SCAN_IN), .B2(n21343), .A(n21263), .ZN(
        n21264) );
  OAI221_X1 U23330 ( .B1(P3_EAX_REG_20__SCAN_IN), .B2(n21276), .C1(n21265), 
        .C2(n21268), .A(n21264), .ZN(P3_U2715) );
  AOI22_X1 U23331 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n21342), .B1(n21376), .B2(
        n21266), .ZN(n21273) );
  NAND2_X1 U23332 ( .A1(n21267), .A2(n21379), .ZN(n21381) );
  OAI21_X1 U23333 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n21381), .A(n21268), .ZN(
        n21269) );
  AOI22_X1 U23334 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n21343), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n21269), .ZN(n21272) );
  NAND3_X1 U23335 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n21270), .A3(n21292), 
        .ZN(n21271) );
  NAND3_X1 U23336 ( .A1(n21273), .A2(n21272), .A3(n21271), .ZN(P3_U2713) );
  AOI22_X1 U23337 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n21342), .ZN(n21278) );
  NAND2_X1 U23338 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .ZN(n21275) );
  NOR2_X1 U23339 ( .A1(n21275), .A2(n21274), .ZN(n21284) );
  OAI211_X1 U23340 ( .C1(n21284), .C2(P3_EAX_REG_19__SCAN_IN), .A(n21370), .B(
        n21276), .ZN(n21277) );
  OAI211_X1 U23341 ( .C1(n21279), .C2(n21373), .A(n21278), .B(n21277), .ZN(
        P3_U2716) );
  AOI22_X1 U23342 ( .A1(n21286), .A2(P3_EAX_REG_17__SCAN_IN), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n21370), .ZN(n21283) );
  AOI22_X1 U23343 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n21342), .B1(n21376), .B2(
        n21280), .ZN(n21282) );
  NAND2_X1 U23344 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n21343), .ZN(n21281) );
  OAI211_X1 U23345 ( .C1(n21284), .C2(n21283), .A(n21282), .B(n21281), .ZN(
        P3_U2717) );
  AOI22_X1 U23346 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n21342), .ZN(n21288) );
  NAND2_X1 U23347 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n21286), .ZN(n21285) );
  OAI211_X1 U23348 ( .C1(n21286), .C2(P3_EAX_REG_17__SCAN_IN), .A(n21370), .B(
        n21285), .ZN(n21287) );
  OAI211_X1 U23349 ( .C1(n21289), .C2(n21373), .A(n21288), .B(n21287), .ZN(
        P3_U2718) );
  AOI22_X1 U23350 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n21343), .B1(n21376), .B2(
        n21290), .ZN(n21297) );
  NAND2_X1 U23351 ( .A1(n21337), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n21336) );
  NOR2_X1 U23352 ( .A1(n21294), .A2(n21336), .ZN(n21331) );
  NAND2_X1 U23353 ( .A1(n21331), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n21330) );
  OAI211_X1 U23354 ( .C1(n21295), .C2(P3_EAX_REG_25__SCAN_IN), .A(n21370), .B(
        n21299), .ZN(n21296) );
  OAI211_X1 U23355 ( .C1(n21341), .C2(n21298), .A(n21297), .B(n21296), .ZN(
        P3_U2710) );
  AOI22_X1 U23356 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n21342), .ZN(n21303) );
  AOI211_X1 U23357 ( .C1(n21300), .C2(n21299), .A(n21326), .B(n21313), .ZN(
        n21301) );
  INV_X1 U23358 ( .A(n21301), .ZN(n21302) );
  OAI211_X1 U23359 ( .C1(n21304), .C2(n21373), .A(n21303), .B(n21302), .ZN(
        P3_U2709) );
  NAND2_X1 U23360 ( .A1(n21326), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n21325) );
  INV_X1 U23361 ( .A(n21325), .ZN(n21320) );
  NAND2_X1 U23362 ( .A1(n21320), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n21319) );
  NOR2_X2 U23363 ( .A1(n21319), .A2(n21312), .ZN(n21311) );
  NAND2_X1 U23364 ( .A1(n21311), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n21307) );
  OAI22_X1 U23365 ( .A1(n21313), .A2(n21311), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n21381), .ZN(n21305) );
  AOI22_X1 U23366 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n21342), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n21305), .ZN(n21306) );
  OAI21_X1 U23367 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n21307), .A(n21306), .ZN(
        P3_U2704) );
  AOI22_X1 U23368 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n21342), .ZN(n21309) );
  OAI211_X1 U23369 ( .C1(n21311), .C2(P3_EAX_REG_30__SCAN_IN), .A(n21370), .B(
        n21307), .ZN(n21308) );
  OAI211_X1 U23370 ( .C1(n21310), .C2(n21373), .A(n21309), .B(n21308), .ZN(
        P3_U2705) );
  INV_X1 U23371 ( .A(n21311), .ZN(n21315) );
  OAI21_X1 U23372 ( .B1(n21313), .B2(n21312), .A(n21319), .ZN(n21314) );
  AOI22_X1 U23373 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n21342), .B1(n21315), .B2(
        n21314), .ZN(n21318) );
  AOI22_X1 U23374 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n21343), .B1(n21376), .B2(
        n21316), .ZN(n21317) );
  NAND2_X1 U23375 ( .A1(n21318), .A2(n21317), .ZN(P3_U2706) );
  AOI22_X1 U23376 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n21342), .ZN(n21322) );
  OAI211_X1 U23377 ( .C1(n21320), .C2(P3_EAX_REG_28__SCAN_IN), .A(n21370), .B(
        n21319), .ZN(n21321) );
  OAI211_X1 U23378 ( .C1(n21323), .C2(n21373), .A(n21322), .B(n21321), .ZN(
        P3_U2707) );
  AOI22_X1 U23379 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n21343), .B1(n21376), .B2(
        n21324), .ZN(n21328) );
  OAI211_X1 U23380 ( .C1(n21326), .C2(P3_EAX_REG_27__SCAN_IN), .A(n21370), .B(
        n21325), .ZN(n21327) );
  OAI211_X1 U23381 ( .C1(n21341), .C2(n21329), .A(n21328), .B(n21327), .ZN(
        P3_U2708) );
  AOI22_X1 U23382 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n21342), .ZN(n21333) );
  OAI211_X1 U23383 ( .C1(n21331), .C2(P3_EAX_REG_24__SCAN_IN), .A(n21370), .B(
        n21330), .ZN(n21332) );
  OAI211_X1 U23384 ( .C1(n21334), .C2(n21373), .A(n21333), .B(n21332), .ZN(
        P3_U2711) );
  AOI22_X1 U23385 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n21343), .B1(n21376), .B2(
        n21335), .ZN(n21339) );
  OAI211_X1 U23386 ( .C1(n21337), .C2(P3_EAX_REG_23__SCAN_IN), .A(n21370), .B(
        n21336), .ZN(n21338) );
  OAI211_X1 U23387 ( .C1(n21341), .C2(n21340), .A(n21339), .B(n21338), .ZN(
        P3_U2712) );
  AOI22_X1 U23388 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n21343), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n21342), .ZN(n21347) );
  OAI211_X1 U23389 ( .C1(n21345), .C2(P3_EAX_REG_16__SCAN_IN), .A(n21370), .B(
        n21344), .ZN(n21346) );
  OAI211_X1 U23390 ( .C1(n21348), .C2(n21373), .A(n21347), .B(n21346), .ZN(
        P3_U2719) );
  NAND2_X1 U23391 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n21349), .ZN(n21354) );
  NAND2_X1 U23392 ( .A1(n21370), .A2(n21350), .ZN(n21359) );
  AOI22_X1 U23393 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n21377), .B1(n21376), .B2(
        n21351), .ZN(n21352) );
  OAI221_X1 U23394 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n21354), .C1(n21353), 
        .C2(n21359), .A(n21352), .ZN(P3_U2721) );
  NAND2_X1 U23395 ( .A1(n21356), .A2(n21355), .ZN(n21361) );
  AOI22_X1 U23396 ( .A1(n21376), .A2(n21357), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n21377), .ZN(n21358) );
  OAI221_X1 U23397 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n21361), .C1(n21360), 
        .C2(n21359), .A(n21358), .ZN(P3_U2720) );
  NAND2_X1 U23398 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n21377), .ZN(n21365) );
  OAI211_X1 U23399 ( .C1(n21363), .C2(P3_EAX_REG_8__SCAN_IN), .A(n21370), .B(
        n21362), .ZN(n21364) );
  OAI211_X1 U23400 ( .C1(n21366), .C2(n21373), .A(n21365), .B(n21364), .ZN(
        P3_U2727) );
  AOI22_X1 U23401 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n21377), .B1(n21368), .B2(
        n21367), .ZN(n21372) );
  NAND3_X1 U23402 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n21370), .A3(n21369), .ZN(
        n21371) );
  OAI211_X1 U23403 ( .C1(n21374), .C2(n21373), .A(n21372), .B(n21371), .ZN(
        P3_U2734) );
  AOI22_X1 U23404 ( .A1(n21377), .A2(BUF2_REG_0__SCAN_IN), .B1(n21376), .B2(
        n21375), .ZN(n21378) );
  OAI221_X1 U23405 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n21381), .C1(n21380), 
        .C2(n21379), .A(n21378), .ZN(P3_U2735) );
  NOR2_X1 U23406 ( .A1(n21382), .A2(n21778), .ZN(n21387) );
  AOI22_X1 U23407 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21859), .B1(
        n21387), .B2(n21385), .ZN(n21896) );
  AOI222_X1 U23408 ( .A1(n21472), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21896), 
        .B2(n21426), .C1(n21385), .C2(n21428), .ZN(n21383) );
  AOI22_X1 U23409 ( .A1(n21431), .A2(n21385), .B1(n21383), .B2(n21429), .ZN(
        P3_U3290) );
  NAND3_X1 U23410 ( .A1(n21409), .A2(n21384), .A3(n21410), .ZN(n21815) );
  AOI21_X1 U23411 ( .B1(n21385), .B2(n21859), .A(n21814), .ZN(n21397) );
  INV_X1 U23412 ( .A(n21397), .ZN(n21417) );
  OAI22_X1 U23413 ( .A1(n21387), .A2(n21386), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21417), .ZN(n21894) );
  AOI22_X1 U23414 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21388), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21481), .ZN(n21403) );
  NOR2_X1 U23415 ( .A1(n21389), .A2(n21472), .ZN(n21393) );
  AOI222_X1 U23416 ( .A1(n21894), .A2(n21426), .B1(n21390), .B2(n21428), .C1(
        n21403), .C2(n21393), .ZN(n21391) );
  AOI22_X1 U23417 ( .A1(n21431), .A2(n21392), .B1(n21391), .B2(n21429), .ZN(
        P3_U3289) );
  INV_X1 U23418 ( .A(n21393), .ZN(n21404) );
  AOI22_X1 U23419 ( .A1(n21396), .A2(n21395), .B1(n21394), .B2(n21410), .ZN(
        n21420) );
  OAI211_X1 U23420 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n21859), .A(
        n21415), .B(n21420), .ZN(n21400) );
  AOI222_X1 U23421 ( .A1(n21400), .A2(n21406), .B1(n21667), .B2(n21399), .C1(
        n21398), .C2(n21397), .ZN(n21890) );
  OAI222_X1 U23422 ( .A1(n21404), .A2(n21403), .B1(n21402), .B2(n21890), .C1(
        n21401), .C2(n21926), .ZN(n21405) );
  AOI22_X1 U23423 ( .A1(n21428), .A2(n21406), .B1(n21429), .B2(n21405), .ZN(
        n21407) );
  OAI21_X1 U23424 ( .B1(n21891), .B2(n21429), .A(n21407), .ZN(P3_U3288) );
  AND2_X1 U23425 ( .A1(n21408), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n21424) );
  NAND2_X1 U23426 ( .A1(n21410), .A2(n21409), .ZN(n21423) );
  NAND2_X1 U23427 ( .A1(n21888), .A2(n21891), .ZN(n21412) );
  OAI211_X1 U23428 ( .C1(n21413), .C2(n21412), .A(n21667), .B(n21411), .ZN(
        n21416) );
  OAI22_X1 U23429 ( .A1(n18317), .A2(n21416), .B1(n21415), .B2(n21414), .ZN(
        n21422) );
  OAI22_X1 U23430 ( .A1(n21420), .A2(n21419), .B1(n21418), .B2(n21417), .ZN(
        n21421) );
  AOI211_X1 U23431 ( .C1(n21424), .C2(n21423), .A(n21422), .B(n21421), .ZN(
        n21887) );
  INV_X1 U23432 ( .A(n21887), .ZN(n21425) );
  AOI22_X1 U23433 ( .A1(n21428), .A2(n21427), .B1(n21426), .B2(n21425), .ZN(
        n21430) );
  AOI22_X1 U23434 ( .A1(n21431), .A2(n21888), .B1(n21430), .B2(n21429), .ZN(
        P3_U3285) );
  NOR3_X1 U23435 ( .A1(n21433), .A2(n21432), .A3(n21882), .ZN(n21446) );
  XNOR2_X1 U23436 ( .A(n21435), .B(n21434), .ZN(n21437) );
  OAI21_X1 U23437 ( .B1(n21437), .B2(n21436), .A(n22370), .ZN(n21873) );
  NOR3_X1 U23438 ( .A1(n21438), .A2(n21881), .A3(n21873), .ZN(n21445) );
  INV_X1 U23439 ( .A(n21439), .ZN(n21441) );
  AOI211_X1 U23440 ( .C1(n21442), .C2(n21441), .A(n21877), .B(n21440), .ZN(
        n21443) );
  NAND3_X1 U23441 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21529) );
  NOR2_X1 U23442 ( .A1(n21448), .A2(n21529), .ZN(n21536) );
  AOI21_X1 U23443 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n21518) );
  INV_X1 U23444 ( .A(n21518), .ZN(n21497) );
  NAND2_X1 U23445 ( .A1(n21536), .A2(n21497), .ZN(n21540) );
  NOR2_X1 U23446 ( .A1(n21559), .A2(n21540), .ZN(n21607) );
  NAND2_X1 U23447 ( .A1(n21458), .A2(n21607), .ZN(n21642) );
  NOR2_X1 U23448 ( .A1(n21449), .A2(n21642), .ZN(n21455) );
  NAND2_X1 U23449 ( .A1(n21667), .A2(n21455), .ZN(n21627) );
  NAND3_X1 U23450 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n21536), .ZN(n21537) );
  NOR2_X1 U23451 ( .A1(n21559), .A2(n21537), .ZN(n21858) );
  NAND2_X1 U23452 ( .A1(n21458), .A2(n21858), .ZN(n21802) );
  OAI21_X1 U23453 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21849), .A(
        n21815), .ZN(n21493) );
  OAI22_X1 U23454 ( .A1(n21562), .A2(n21885), .B1(n21784), .B2(n21563), .ZN(
        n21582) );
  NAND2_X1 U23455 ( .A1(n21458), .A2(n21582), .ZN(n21631) );
  OAI21_X1 U23456 ( .B1(n21802), .B2(n21493), .A(n21631), .ZN(n21451) );
  NAND2_X1 U23457 ( .A1(n21451), .A2(n21459), .ZN(n21452) );
  AOI21_X1 U23458 ( .B1(n21627), .B2(n21452), .A(n21808), .ZN(n21794) );
  NAND2_X1 U23459 ( .A1(n21859), .A2(n21886), .ZN(n21847) );
  OAI21_X1 U23460 ( .B1(n21802), .B2(n21453), .A(n21849), .ZN(n21454) );
  OAI21_X1 U23461 ( .B1(n21455), .B2(n21886), .A(n21454), .ZN(n21780) );
  OAI22_X1 U23462 ( .A1(n21752), .A2(n21784), .B1(n21456), .B2(n21885), .ZN(
        n21457) );
  AOI211_X1 U23463 ( .C1(n21460), .C2(n21847), .A(n21780), .B(n21457), .ZN(
        n21636) );
  INV_X1 U23464 ( .A(n21858), .ZN(n21848) );
  NOR2_X1 U23465 ( .A1(n21472), .A2(n21848), .ZN(n21860) );
  AND2_X1 U23466 ( .A1(n21458), .A2(n21860), .ZN(n21606) );
  NAND2_X1 U23467 ( .A1(n21459), .A2(n21606), .ZN(n21777) );
  AOI221_X1 U23468 ( .B1(n21460), .B2(n21778), .C1(n21777), .C2(n21778), .A(
        n21808), .ZN(n21461) );
  AOI211_X1 U23469 ( .C1(n21636), .C2(n21461), .A(n21866), .B(n21634), .ZN(
        n21462) );
  AOI211_X1 U23470 ( .C1(n21464), .C2(n21794), .A(n21463), .B(n21462), .ZN(
        n21465) );
  OAI21_X1 U23471 ( .B1(n21466), .B2(n21790), .A(n21465), .ZN(P3_U2841) );
  NAND2_X1 U23472 ( .A1(n21841), .A2(n21783), .ZN(n21617) );
  AND2_X1 U23473 ( .A1(n21866), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n21468) );
  INV_X1 U23474 ( .A(n21687), .ZN(n21796) );
  AOI221_X1 U23475 ( .B1(n21859), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C1(
        n21796), .C2(n21472), .A(n21808), .ZN(n21467) );
  AOI211_X1 U23476 ( .C1(n21754), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n21468), .B(n21467), .ZN(n21469) );
  OAI221_X1 U23477 ( .B1(n21471), .B2(n21617), .C1(n21470), .C2(n21547), .A(
        n21469), .ZN(P3_U2862) );
  NAND3_X1 U23478 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n21687), .A3(
        n21472), .ZN(n21474) );
  OAI211_X1 U23479 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n21849), .A(
        n21481), .B(n21831), .ZN(n21473) );
  OAI211_X1 U23480 ( .C1(n21475), .C2(n21487), .A(n21474), .B(n21473), .ZN(
        n21477) );
  AOI22_X1 U23481 ( .A1(n21841), .A2(n21477), .B1(n21722), .B2(n21476), .ZN(
        n21479) );
  NAND2_X1 U23482 ( .A1(n21866), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n21478) );
  OAI211_X1 U23483 ( .C1(n21761), .C2(n21481), .A(n21479), .B(n21478), .ZN(
        P3_U2861) );
  NAND2_X1 U23484 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21480) );
  OAI21_X1 U23485 ( .B1(n21480), .B2(n21492), .A(n21497), .ZN(n21484) );
  NOR3_X1 U23486 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21481), .A3(
        n21493), .ZN(n21483) );
  NOR2_X1 U23487 ( .A1(n21861), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21803) );
  INV_X1 U23488 ( .A(n21803), .ZN(n21495) );
  AOI211_X1 U23489 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21495), .A(
        n21814), .B(n21492), .ZN(n21482) );
  AOI211_X1 U23490 ( .C1(n21667), .C2(n21484), .A(n21483), .B(n21482), .ZN(
        n21486) );
  AOI221_X1 U23491 ( .B1(n21487), .B2(n21486), .C1(n21485), .C2(n21486), .A(
        n21808), .ZN(n21488) );
  AOI211_X1 U23492 ( .C1(n21722), .C2(n21490), .A(n21489), .B(n21488), .ZN(
        n21491) );
  OAI21_X1 U23493 ( .B1(n21492), .B2(n21761), .A(n21491), .ZN(P3_U2860) );
  NAND2_X1 U23494 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21494) );
  OAI22_X1 U23495 ( .A1(n21518), .A2(n21886), .B1(n21494), .B2(n21493), .ZN(
        n21535) );
  NOR2_X1 U23496 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n21535), .ZN(
        n21500) );
  INV_X1 U23497 ( .A(n21494), .ZN(n21496) );
  AOI21_X1 U23498 ( .B1(n21496), .B2(n21495), .A(n21814), .ZN(n21517) );
  OAI21_X1 U23499 ( .B1(n21886), .B2(n21497), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21498) );
  OAI21_X1 U23500 ( .B1(n21517), .B2(n21498), .A(n21841), .ZN(n21505) );
  OAI22_X1 U23501 ( .A1(n21500), .A2(n21505), .B1(n21547), .B2(n21499), .ZN(
        n21501) );
  AOI21_X1 U23502 ( .B1(n21722), .B2(n21502), .A(n21501), .ZN(n21504) );
  NAND2_X1 U23503 ( .A1(n21866), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n21503) );
  OAI211_X1 U23504 ( .C1(n21761), .C2(n21507), .A(n21504), .B(n21503), .ZN(
        P3_U2859) );
  NOR3_X1 U23505 ( .A1(n21659), .A2(n21506), .A3(n21505), .ZN(n21512) );
  NAND2_X1 U23506 ( .A1(n21841), .A2(n21535), .ZN(n21528) );
  NOR3_X1 U23507 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21507), .A3(
        n21528), .ZN(n21511) );
  AOI22_X1 U23508 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21754), .B1(
        n21722), .B2(n21508), .ZN(n21509) );
  INV_X1 U23509 ( .A(n21509), .ZN(n21510) );
  NOR4_X1 U23510 ( .A1(n21513), .A2(n21512), .A3(n21511), .A4(n21510), .ZN(
        n21514) );
  OAI21_X1 U23511 ( .B1(n21547), .B2(n21515), .A(n21514), .ZN(P3_U2858) );
  NAND2_X1 U23512 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21516) );
  NOR2_X1 U23513 ( .A1(n21516), .A2(n21528), .ZN(n21521) );
  AOI211_X1 U23514 ( .C1(n21529), .C2(n21815), .A(n21517), .B(n21808), .ZN(
        n21520) );
  OAI21_X1 U23515 ( .B1(n21518), .B2(n21529), .A(n21667), .ZN(n21519) );
  AOI21_X1 U23516 ( .B1(n21520), .B2(n21519), .A(n21866), .ZN(n21527) );
  MUX2_X1 U23517 ( .A(n21521), .B(n21527), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n21522) );
  AOI21_X1 U23518 ( .B1(n21722), .B2(n21523), .A(n21522), .ZN(n21525) );
  OAI211_X1 U23519 ( .C1(n21547), .C2(n21526), .A(n21525), .B(n21524), .ZN(
        P3_U2857) );
  AOI22_X1 U23520 ( .A1(n21866), .A2(P3_REIP_REG_6__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21527), .ZN(n21533) );
  NOR3_X1 U23521 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n21529), .A3(
        n21528), .ZN(n21530) );
  AOI21_X1 U23522 ( .B1(n21531), .B2(n21722), .A(n21530), .ZN(n21532) );
  OAI211_X1 U23523 ( .C1(n21547), .C2(n21534), .A(n21533), .B(n21532), .ZN(
        P3_U2856) );
  NAND2_X1 U23524 ( .A1(n21536), .A2(n21535), .ZN(n21558) );
  AOI21_X1 U23525 ( .B1(n21537), .B2(n21815), .A(n11322), .ZN(n21538) );
  INV_X1 U23526 ( .A(n21538), .ZN(n21539) );
  AOI211_X1 U23527 ( .C1(n21667), .C2(n21540), .A(n21803), .B(n21539), .ZN(
        n21549) );
  AOI211_X1 U23528 ( .C1(n11322), .C2(n21558), .A(n21549), .B(n21808), .ZN(
        n21543) );
  OAI22_X1 U23529 ( .A1(n21822), .A2(n21541), .B1(n11322), .B2(n21761), .ZN(
        n21542) );
  AOI211_X1 U23530 ( .C1(n21544), .C2(n21722), .A(n21543), .B(n21542), .ZN(
        n21545) );
  OAI21_X1 U23531 ( .B1(n21547), .B2(n21546), .A(n21545), .ZN(P3_U2855) );
  NOR3_X1 U23532 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n11322), .A3(
        n21558), .ZN(n21551) );
  NOR3_X1 U23533 ( .A1(n21659), .A2(n21549), .A3(n21548), .ZN(n21550) );
  AOI211_X1 U23534 ( .C1(n21756), .C2(n21552), .A(n21551), .B(n21550), .ZN(
        n21557) );
  AOI22_X1 U23535 ( .A1(n21866), .A2(P3_REIP_REG_8__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n21754), .ZN(n21556) );
  AOI22_X1 U23536 ( .A1(n21865), .A2(n21554), .B1(n21722), .B2(n21553), .ZN(
        n21555) );
  OAI211_X1 U23537 ( .C1(n21557), .C2(n21808), .A(n21556), .B(n21555), .ZN(
        P3_U2854) );
  OAI21_X1 U23538 ( .B1(n21614), .B2(n21582), .A(n21841), .ZN(n21870) );
  AOI22_X1 U23539 ( .A1(n21866), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n21865), 
        .B2(n21560), .ZN(n21570) );
  AOI21_X1 U23540 ( .B1(n21561), .B2(n21858), .A(n21859), .ZN(n21580) );
  NAND2_X1 U23541 ( .A1(n21784), .A2(n21885), .ZN(n21811) );
  AOI21_X1 U23542 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21860), .A(
        n21861), .ZN(n21565) );
  NOR2_X1 U23543 ( .A1(n21607), .A2(n21886), .ZN(n21573) );
  AOI211_X1 U23544 ( .C1(n21783), .C2(n21562), .A(n21573), .B(n21808), .ZN(
        n21564) );
  NAND2_X1 U23545 ( .A1(n21756), .A2(n21563), .ZN(n21804) );
  NAND2_X1 U23546 ( .A1(n21564), .A2(n21804), .ZN(n21863) );
  AOI211_X1 U23547 ( .C1(n21567), .C2(n21811), .A(n21565), .B(n21863), .ZN(
        n21852) );
  OAI21_X1 U23548 ( .B1(n21567), .B2(n21566), .A(n21667), .ZN(n21574) );
  OAI211_X1 U23549 ( .C1(n21861), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21852), .B(n21574), .ZN(n21568) );
  OAI211_X1 U23550 ( .C1(n21580), .C2(n21568), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n21822), .ZN(n21569) );
  OAI211_X1 U23551 ( .C1(n21571), .C2(n21870), .A(n21570), .B(n21569), .ZN(
        P3_U2851) );
  AOI21_X1 U23552 ( .B1(n21572), .B2(n21860), .A(n21861), .ZN(n21591) );
  NOR2_X1 U23553 ( .A1(n21591), .A2(n21592), .ZN(n21584) );
  AOI21_X1 U23554 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n21859), .ZN(n21579) );
  INV_X1 U23555 ( .A(n21573), .ZN(n21575) );
  NAND2_X1 U23556 ( .A1(n21575), .A2(n21574), .ZN(n21589) );
  OAI22_X1 U23557 ( .A1(n21577), .A2(n21885), .B1(n21576), .B2(n21784), .ZN(
        n21578) );
  NOR4_X1 U23558 ( .A1(n21580), .A2(n21579), .A3(n21589), .A4(n21578), .ZN(
        n21842) );
  OAI21_X1 U23559 ( .B1(n21614), .B2(n21582), .A(n21581), .ZN(n21583) );
  AOI22_X1 U23560 ( .A1(n21584), .A2(n21842), .B1(n21592), .B2(n21583), .ZN(
        n21586) );
  AOI22_X1 U23561 ( .A1(n21841), .A2(n21586), .B1(n21865), .B2(n21585), .ZN(
        n21588) );
  OAI211_X1 U23562 ( .C1(n21761), .C2(n21592), .A(n21588), .B(n21587), .ZN(
        P3_U2850) );
  NAND2_X1 U23563 ( .A1(n21605), .A2(n21858), .ZN(n21590) );
  AOI21_X1 U23564 ( .B1(n21849), .B2(n21590), .A(n21589), .ZN(n21593) );
  AOI21_X1 U23565 ( .B1(n21667), .B2(n21592), .A(n21591), .ZN(n21840) );
  OAI211_X1 U23566 ( .C1(n21796), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n21593), .B(n21840), .ZN(n21594) );
  AOI22_X1 U23567 ( .A1(n21756), .A2(n21595), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n21594), .ZN(n21603) );
  NAND3_X1 U23568 ( .A1(n21605), .A2(n21614), .A3(n21596), .ZN(n21602) );
  OAI22_X1 U23569 ( .A1(n21598), .A2(n21790), .B1(n21617), .B2(n21597), .ZN(
        n21599) );
  AOI211_X1 U23570 ( .C1(n21754), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n21600), .B(n21599), .ZN(n21601) );
  OAI221_X1 U23571 ( .B1(n21808), .B2(n21603), .C1(n21808), .C2(n21602), .A(
        n21601), .ZN(P3_U2848) );
  NAND2_X1 U23572 ( .A1(n21604), .A2(n21756), .ZN(n21623) );
  INV_X1 U23573 ( .A(n21623), .ZN(n21615) );
  NAND3_X1 U23574 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21605), .A3(
        n21858), .ZN(n21610) );
  AOI21_X1 U23575 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21861), .A(
        n21606), .ZN(n21609) );
  AOI21_X1 U23576 ( .B1(n21612), .B2(n21607), .A(n21886), .ZN(n21608) );
  AOI211_X1 U23577 ( .C1(n21849), .C2(n21610), .A(n21609), .B(n21608), .ZN(
        n21611) );
  INV_X1 U23578 ( .A(n21611), .ZN(n21830) );
  AND2_X1 U23579 ( .A1(n21830), .A2(n21612), .ZN(n21613) );
  AOI22_X1 U23580 ( .A1(n21616), .A2(n21615), .B1(n21614), .B2(n21613), .ZN(
        n21626) );
  NOR3_X1 U23581 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21618), .A3(
        n21617), .ZN(n21620) );
  AOI211_X1 U23582 ( .C1(n21865), .C2(n21621), .A(n21620), .B(n21619), .ZN(
        n21625) );
  INV_X1 U23583 ( .A(n21622), .ZN(n21805) );
  OAI211_X1 U23584 ( .C1(n21805), .C2(n21885), .A(n21841), .B(n21623), .ZN(
        n21832) );
  OAI211_X1 U23585 ( .C1(n21830), .C2(n21832), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n21822), .ZN(n21624) );
  OAI211_X1 U23586 ( .C1(n21626), .C2(n21808), .A(n21625), .B(n21624), .ZN(
        P3_U2847) );
  OAI21_X1 U23587 ( .B1(n21861), .B2(n21777), .A(n21627), .ZN(n21628) );
  NOR2_X1 U23588 ( .A1(n21630), .A2(n21802), .ZN(n21632) );
  AOI22_X1 U23589 ( .A1(n21629), .A2(n21628), .B1(n21632), .B2(n21849), .ZN(
        n21679) );
  OAI21_X1 U23590 ( .B1(n21631), .B2(n21630), .A(n21679), .ZN(n21762) );
  INV_X1 U23591 ( .A(n21762), .ZN(n21769) );
  INV_X1 U23592 ( .A(n21632), .ZN(n21691) );
  NOR3_X1 U23593 ( .A1(n21803), .A2(n21641), .A3(n21691), .ZN(n21644) );
  AOI21_X1 U23594 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n21861), .A(
        n21644), .ZN(n21633) );
  AOI21_X1 U23595 ( .B1(n21634), .B2(n21847), .A(n21633), .ZN(n21635) );
  AOI22_X1 U23596 ( .A1(n21769), .A2(n21641), .B1(n21636), .B2(n21635), .ZN(
        n21638) );
  AOI22_X1 U23597 ( .A1(n21841), .A2(n21638), .B1(n21865), .B2(n21637), .ZN(
        n21640) );
  NAND2_X1 U23598 ( .A1(n21866), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n21639) );
  OAI211_X1 U23599 ( .C1(n21761), .C2(n21641), .A(n21640), .B(n21639), .ZN(
        P3_U2840) );
  OAI21_X1 U23600 ( .B1(n21679), .B2(n21655), .A(n21654), .ZN(n21648) );
  INV_X1 U23601 ( .A(n21642), .ZN(n21806) );
  NAND3_X1 U23602 ( .A1(n21643), .A2(n21806), .A3(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21668) );
  OAI21_X1 U23603 ( .B1(n21814), .B2(n21644), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21645) );
  AOI21_X1 U23604 ( .B1(n21667), .B2(n21668), .A(n21645), .ZN(n21760) );
  OAI221_X1 U23605 ( .B1(n21659), .B2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), 
        .C1(n21659), .C2(n21760), .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n21657) );
  AOI222_X1 U23606 ( .A1(n21648), .A2(n21657), .B1(n21783), .B2(n21647), .C1(
        n21756), .C2(n21646), .ZN(n21653) );
  OAI22_X1 U23607 ( .A1(n21654), .A2(n21761), .B1(n21790), .B2(n21649), .ZN(
        n21650) );
  INV_X1 U23608 ( .A(n21650), .ZN(n21652) );
  NAND2_X1 U23609 ( .A1(n21866), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n21651) );
  OAI211_X1 U23610 ( .C1(n21653), .C2(n21808), .A(n21652), .B(n21651), .ZN(
        P3_U2837) );
  NOR2_X1 U23611 ( .A1(n21655), .A2(n21654), .ZN(n21656) );
  AOI21_X1 U23612 ( .B1(n21656), .B2(n21762), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21665) );
  INV_X1 U23613 ( .A(n21657), .ZN(n21658) );
  NAND2_X1 U23614 ( .A1(n21756), .A2(n21681), .ZN(n21669) );
  OAI211_X1 U23615 ( .C1(n21659), .C2(n21658), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n21669), .ZN(n21660) );
  AOI22_X1 U23616 ( .A1(n21841), .A2(n21660), .B1(n21722), .B2(n21666), .ZN(
        n21664) );
  AOI22_X1 U23617 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n21754), .B1(
        n21865), .B2(n21661), .ZN(n21663) );
  OAI211_X1 U23618 ( .C1(n21665), .C2(n21664), .A(n21663), .B(n21662), .ZN(
        P3_U2836) );
  AOI22_X1 U23619 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21754), .B1(
        n21722), .B2(n21666), .ZN(n21672) );
  NOR2_X1 U23620 ( .A1(n21691), .A2(n21678), .ZN(n21702) );
  OAI21_X1 U23621 ( .B1(n21678), .B2(n21668), .A(n21667), .ZN(n21701) );
  AND2_X1 U23622 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21701), .ZN(
        n21685) );
  OAI211_X1 U23623 ( .C1(n21702), .C2(n21814), .A(n21685), .B(n21669), .ZN(
        n21670) );
  OAI21_X1 U23624 ( .B1(n21803), .B2(n21670), .A(n21841), .ZN(n21671) );
  NAND2_X1 U23625 ( .A1(n21689), .A2(n21762), .ZN(n21739) );
  AOI22_X1 U23626 ( .A1(n21672), .A2(n21671), .B1(n21739), .B2(n21738), .ZN(
        n21673) );
  AOI21_X1 U23627 ( .B1(n21865), .B2(n21674), .A(n21673), .ZN(n21676) );
  NAND2_X1 U23628 ( .A1(n21676), .A2(n21675), .ZN(P3_U2835) );
  NOR3_X1 U23629 ( .A1(n21679), .A2(n21678), .A3(n21677), .ZN(n21718) );
  AOI21_X1 U23630 ( .B1(n21734), .B2(n21756), .A(n21718), .ZN(n21680) );
  OAI21_X1 U23631 ( .B1(n21885), .B2(n21729), .A(n21680), .ZN(n21709) );
  NAND3_X1 U23632 ( .A1(n21692), .A2(n21841), .A3(n21709), .ZN(n21699) );
  NOR2_X1 U23633 ( .A1(n21681), .A2(n21703), .ZN(n21683) );
  NAND3_X1 U23634 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21702), .A3(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21684) );
  NAND2_X1 U23635 ( .A1(n21684), .A2(n21778), .ZN(n21700) );
  OAI211_X1 U23636 ( .C1(n21685), .C2(n21886), .A(n21841), .B(n21700), .ZN(
        n21686) );
  AOI211_X1 U23637 ( .C1(n21743), .C2(n21687), .A(n21705), .B(n21686), .ZN(
        n21694) );
  NAND2_X1 U23638 ( .A1(n21689), .A2(n21688), .ZN(n21690) );
  OAI21_X1 U23639 ( .B1(n21691), .B2(n21690), .A(n21849), .ZN(n21693) );
  AOI211_X1 U23640 ( .C1(n21694), .C2(n21693), .A(n21866), .B(n21692), .ZN(
        n21695) );
  AOI211_X1 U23641 ( .C1(n21865), .C2(n21697), .A(n21696), .B(n21695), .ZN(
        n21698) );
  NAND2_X1 U23642 ( .A1(n21699), .A2(n21698), .ZN(P3_U2833) );
  NAND2_X1 U23643 ( .A1(n21866), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n21711) );
  OAI211_X1 U23644 ( .C1(n21859), .C2(n21702), .A(n21701), .B(n21700), .ZN(
        n21733) );
  AOI211_X1 U23645 ( .C1(n21831), .C2(n21703), .A(n21733), .B(n21706), .ZN(
        n21715) );
  INV_X1 U23646 ( .A(n21715), .ZN(n21704) );
  OAI22_X1 U23647 ( .A1(n21808), .A2(n21707), .B1(n21761), .B2(n21706), .ZN(
        n21708) );
  OAI21_X1 U23648 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n21709), .A(
        n21708), .ZN(n21710) );
  OAI211_X1 U23649 ( .C1(n21712), .C2(n21790), .A(n21711), .B(n21710), .ZN(
        P3_U2832) );
  NOR2_X1 U23650 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21713), .ZN(
        n21719) );
  NAND2_X1 U23651 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n21831), .ZN(
        n21714) );
  OAI22_X1 U23652 ( .A1(n21716), .A2(n21784), .B1(n21715), .B2(n21714), .ZN(
        n21717) );
  AOI21_X1 U23653 ( .B1(n21719), .B2(n21718), .A(n21717), .ZN(n21726) );
  AOI21_X1 U23654 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21754), .A(
        n21720), .ZN(n21725) );
  AOI22_X1 U23655 ( .A1(n21865), .A2(n21723), .B1(n21722), .B2(n21721), .ZN(
        n21724) );
  OAI211_X1 U23656 ( .C1(n21726), .C2(n21808), .A(n21725), .B(n21724), .ZN(
        P3_U2831) );
  OAI21_X1 U23657 ( .B1(n21740), .B2(n21728), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n21732) );
  AOI21_X1 U23658 ( .B1(n21732), .B2(n21731), .A(n21730), .ZN(n21737) );
  AOI211_X1 U23659 ( .C1(n21738), .C2(n21847), .A(n21754), .B(n21733), .ZN(
        n21736) );
  OR2_X1 U23660 ( .A1(n21734), .A2(n21784), .ZN(n21735) );
  NAND3_X1 U23661 ( .A1(n21737), .A2(n21736), .A3(n21735), .ZN(n21746) );
  NAND2_X1 U23662 ( .A1(n21746), .A2(n21745), .ZN(n21751) );
  OR3_X1 U23663 ( .A1(n21748), .A2(n21790), .A3(n21747), .ZN(n21749) );
  OAI221_X1 U23664 ( .B1(n21866), .B2(n21751), .C1(n21822), .C2(n21750), .A(
        n21749), .ZN(P3_U2834) );
  NAND2_X1 U23665 ( .A1(n21753), .A2(n21752), .ZN(n21755) );
  AOI21_X1 U23666 ( .B1(n21756), .B2(n21755), .A(n21754), .ZN(n21757) );
  OAI21_X1 U23667 ( .B1(n21758), .B2(n21885), .A(n21757), .ZN(n21772) );
  INV_X1 U23668 ( .A(n21772), .ZN(n21759) );
  AOI21_X1 U23669 ( .B1(n21760), .B2(n21759), .A(n21866), .ZN(n21771) );
  INV_X1 U23670 ( .A(n21771), .ZN(n21767) );
  NAND3_X1 U23671 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21762), .A3(
        n21761), .ZN(n21765) );
  AOI22_X1 U23672 ( .A1(n21866), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n21865), 
        .B2(n21763), .ZN(n21764) );
  OAI221_X1 U23673 ( .B1(n21767), .B2(n21766), .C1(n21767), .C2(n21765), .A(
        n21764), .ZN(P3_U2839) );
  NOR4_X1 U23674 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21769), .A3(
        n21808), .A4(n21768), .ZN(n21770) );
  AOI21_X1 U23675 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n21866), .A(n21770), 
        .ZN(n21774) );
  OAI211_X1 U23676 ( .C1(n21831), .C2(n21772), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21771), .ZN(n21773) );
  OAI211_X1 U23677 ( .C1(n21775), .C2(n21790), .A(n21774), .B(n21773), .ZN(
        P3_U2838) );
  INV_X1 U23678 ( .A(n21776), .ZN(n21782) );
  AOI21_X1 U23679 ( .B1(n21778), .B2(n21777), .A(n21808), .ZN(n21779) );
  INV_X1 U23680 ( .A(n21779), .ZN(n21781) );
  AOI211_X1 U23681 ( .C1(n21783), .C2(n21782), .A(n21781), .B(n21780), .ZN(
        n21785) );
  AOI221_X1 U23682 ( .B1(n21786), .B2(n21785), .C1(n21784), .C2(n21785), .A(
        n21866), .ZN(n21798) );
  AOI22_X1 U23683 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21798), .B1(
        n21794), .B2(n21787), .ZN(n21789) );
  OAI211_X1 U23684 ( .C1(n21791), .C2(n21790), .A(n21789), .B(n21788), .ZN(
        P3_U2843) );
  INV_X1 U23685 ( .A(n21792), .ZN(n21795) );
  AOI22_X1 U23686 ( .A1(n21865), .A2(n21795), .B1(n21794), .B2(n21793), .ZN(
        n21800) );
  NOR3_X1 U23687 ( .A1(n21796), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n21915), .ZN(n21797) );
  OAI21_X1 U23688 ( .B1(n21798), .B2(n21797), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21799) );
  OAI211_X1 U23689 ( .C1(n21801), .C2(n21822), .A(n21800), .B(n21799), .ZN(
        P3_U2842) );
  NOR3_X1 U23690 ( .A1(n21803), .A2(n21802), .A3(n21833), .ZN(n21813) );
  NAND3_X1 U23691 ( .A1(n21805), .A2(n21807), .A3(n21804), .ZN(n21810) );
  AOI21_X1 U23692 ( .B1(n21807), .B2(n21806), .A(n21886), .ZN(n21809) );
  AOI211_X1 U23693 ( .C1(n21811), .C2(n21810), .A(n21809), .B(n21808), .ZN(
        n21812) );
  OAI21_X1 U23694 ( .B1(n21814), .B2(n21813), .A(n21812), .ZN(n21826) );
  OAI221_X1 U23695 ( .B1(n21826), .B2(n21816), .C1(n21826), .C2(n21815), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21823) );
  NOR2_X1 U23696 ( .A1(n21817), .A2(n21870), .ZN(n21834) );
  AOI22_X1 U23697 ( .A1(n21865), .A2(n21819), .B1(n21834), .B2(n21818), .ZN(
        n21820) );
  OAI221_X1 U23698 ( .B1(n21866), .B2(n21823), .C1(n21822), .C2(n21821), .A(
        n21820), .ZN(P3_U2844) );
  NOR2_X1 U23699 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21833), .ZN(
        n21824) );
  AOI22_X1 U23700 ( .A1(n21865), .A2(n21825), .B1(n21834), .B2(n21824), .ZN(
        n21829) );
  NAND3_X1 U23701 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21822), .A3(
        n21826), .ZN(n21827) );
  NAND3_X1 U23702 ( .A1(n21829), .A2(n21828), .A3(n21827), .ZN(P3_U2845) );
  OAI221_X1 U23703 ( .B1(n21832), .B2(n21831), .C1(n21832), .C2(n21830), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21838) );
  AOI22_X1 U23704 ( .A1(n21835), .A2(n21865), .B1(n21834), .B2(n21833), .ZN(
        n21836) );
  OAI221_X1 U23705 ( .B1(n21866), .B2(n21838), .C1(n21822), .C2(n21837), .A(
        n21836), .ZN(P3_U2846) );
  AOI22_X1 U23706 ( .A1(n21866), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n21865), 
        .B2(n21839), .ZN(n21845) );
  NAND3_X1 U23707 ( .A1(n21842), .A2(n21841), .A3(n21840), .ZN(n21843) );
  NAND3_X1 U23708 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21822), .A3(
        n21843), .ZN(n21844) );
  OAI211_X1 U23709 ( .C1(n21846), .C2(n21870), .A(n21845), .B(n21844), .ZN(
        P3_U2849) );
  NAND2_X1 U23710 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21850), .ZN(
        n21857) );
  AOI22_X1 U23711 ( .A1(n21849), .A2(n21848), .B1(n21869), .B2(n21847), .ZN(
        n21851) );
  AOI211_X1 U23712 ( .C1(n21852), .C2(n21851), .A(n21866), .B(n21850), .ZN(
        n21853) );
  AOI21_X1 U23713 ( .B1(n21854), .B2(n21865), .A(n21853), .ZN(n21856) );
  OAI211_X1 U23714 ( .C1(n21857), .C2(n21870), .A(n21856), .B(n21855), .ZN(
        P3_U2852) );
  OAI22_X1 U23715 ( .A1(n21861), .A2(n21860), .B1(n21859), .B2(n21858), .ZN(
        n21862) );
  OAI21_X1 U23716 ( .B1(n21863), .B2(n21862), .A(n21822), .ZN(n21868) );
  AOI22_X1 U23717 ( .A1(n21866), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21865), 
        .B2(n21864), .ZN(n21867) );
  OAI221_X1 U23718 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21870), .C1(
        n21869), .C2(n21868), .A(n21867), .ZN(P3_U2853) );
  NAND2_X1 U23719 ( .A1(n22321), .A2(n21871), .ZN(n21925) );
  INV_X1 U23720 ( .A(n21872), .ZN(n21919) );
  INV_X1 U23721 ( .A(n21873), .ZN(n21875) );
  NOR3_X1 U23722 ( .A1(n21875), .A2(n21874), .A3(n21881), .ZN(n21938) );
  AOI221_X1 U23723 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(n21938), .C1(
        P3_MORE_REG_SCAN_IN), .C2(n21938), .A(n21876), .ZN(n21912) );
  NAND2_X1 U23724 ( .A1(n21879), .A2(n21878), .ZN(n21880) );
  AOI22_X1 U23725 ( .A1(n21883), .A2(n21882), .B1(n21881), .B2(n21880), .ZN(
        n21884) );
  OAI221_X1 U23726 ( .B1(n11369), .B2(n21886), .C1(n11369), .C2(n21885), .A(
        n21884), .ZN(n21939) );
  INV_X1 U23727 ( .A(n21909), .ZN(n21889) );
  MUX2_X1 U23728 ( .A(n21888), .B(n21887), .S(n21889), .Z(n21907) );
  AOI22_X1 U23729 ( .A1(n21909), .A2(n21891), .B1(n21890), .B2(n21889), .ZN(
        n21902) );
  OR3_X1 U23730 ( .A1(n21896), .A2(n21895), .A3(n21892), .ZN(n21893) );
  AOI22_X1 U23731 ( .A1(n21896), .A2(n21895), .B1(n21894), .B2(n21893), .ZN(
        n21898) );
  OAI21_X1 U23732 ( .B1(n21909), .B2(n21898), .A(n21897), .ZN(n21901) );
  AND2_X1 U23733 ( .A1(n21902), .A2(n21901), .ZN(n21899) );
  OAI221_X1 U23734 ( .B1(n21902), .B2(n21901), .C1(n21900), .C2(n21899), .A(
        n21904), .ZN(n21906) );
  AOI21_X1 U23735 ( .B1(n21904), .B2(n21903), .A(n21902), .ZN(n21905) );
  AOI222_X1 U23736 ( .A1(n21907), .A2(n21906), .B1(n21907), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21906), .C2(n21905), .ZN(
        n21908) );
  AOI211_X1 U23737 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n21909), .A(
        n21939), .B(n21908), .ZN(n21911) );
  NAND3_X1 U23738 ( .A1(n21912), .A2(n21911), .A3(n21910), .ZN(n21931) );
  AOI211_X1 U23739 ( .C1(n21914), .C2(n21913), .A(n21937), .B(n21931), .ZN(
        n21921) );
  AOI21_X1 U23740 ( .B1(n22321), .B2(n21915), .A(n21921), .ZN(n21935) );
  NAND3_X1 U23741 ( .A1(n21917), .A2(n21935), .A3(n21916), .ZN(n21918) );
  NAND4_X1 U23742 ( .A1(n21920), .A2(n21925), .A3(n21919), .A4(n21918), .ZN(
        P3_U2997) );
  NOR2_X1 U23743 ( .A1(n21921), .A2(n21936), .ZN(n21924) );
  OAI21_X1 U23744 ( .B1(n21924), .B2(n21923), .A(n21922), .ZN(P3_U3282) );
  OAI211_X1 U23745 ( .C1(n21927), .C2(n21926), .A(n21936), .B(n21925), .ZN(
        n21928) );
  INV_X1 U23746 ( .A(n21928), .ZN(n21929) );
  AOI211_X1 U23747 ( .C1(n21932), .C2(n21931), .A(n21930), .B(n21929), .ZN(
        n21933) );
  OAI221_X1 U23748 ( .B1(n21936), .B2(n21935), .C1(n21936), .C2(n21934), .A(
        n21933), .ZN(P3_U2996) );
  NOR2_X1 U23749 ( .A1(n21938), .A2(n21937), .ZN(n21942) );
  MUX2_X1 U23750 ( .A(P3_MORE_REG_SCAN_IN), .B(n21939), .S(n21942), .Z(
        P3_U3295) );
  INV_X1 U23751 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21941) );
  OAI21_X1 U23752 ( .B1(n21942), .B2(n21941), .A(n21940), .ZN(P3_U2637) );
  AOI211_X1 U23753 ( .C1(n21945), .C2(n22325), .A(n21944), .B(n21943), .ZN(
        n21951) );
  OAI211_X1 U23754 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n21947), .A(n21946), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n21948) );
  AOI21_X1 U23755 ( .B1(n21948), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n22297), 
        .ZN(n21950) );
  NAND2_X1 U23756 ( .A1(n21951), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21949) );
  OAI21_X1 U23757 ( .B1(n21951), .B2(n21950), .A(n21949), .ZN(P1_U3485) );
  AOI22_X1 U23758 ( .A1(n21953), .A2(n22099), .B1(n22098), .B2(n21952), .ZN(
        n21964) );
  NAND2_X1 U23759 ( .A1(n22108), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21963) );
  NAND2_X1 U23760 ( .A1(n22005), .A2(n22012), .ZN(n21956) );
  INV_X1 U23761 ( .A(n21979), .ZN(n21994) );
  NOR3_X1 U23762 ( .A1(n21954), .A2(n21995), .A3(n21994), .ZN(n22050) );
  INV_X1 U23763 ( .A(n22050), .ZN(n21955) );
  NAND4_X1 U23764 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21958), .A3(
        n21957), .A4(n22060), .ZN(n21962) );
  OAI21_X1 U23765 ( .B1(n21960), .B2(n21959), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21961) );
  NAND4_X1 U23766 ( .A1(n21964), .A2(n21963), .A3(n21962), .A4(n21961), .ZN(
        P1_U3017) );
  NOR3_X1 U23767 ( .A1(n14517), .A2(n21969), .A3(n22049), .ZN(n21965) );
  AOI211_X1 U23768 ( .C1(n21969), .C2(n22045), .A(n21965), .B(n22015), .ZN(
        n21975) );
  NOR2_X1 U23769 ( .A1(n22049), .A2(n21978), .ZN(n21976) );
  NOR2_X1 U23770 ( .A1(n22067), .A2(n22111), .ZN(n21967) );
  AND2_X1 U23771 ( .A1(n22108), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n21966) );
  NOR3_X1 U23772 ( .A1(n21976), .A2(n21967), .A3(n21966), .ZN(n21973) );
  INV_X1 U23773 ( .A(n21968), .ZN(n21971) );
  NOR3_X1 U23774 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n21969), .A3(
        n21994), .ZN(n21970) );
  AOI21_X1 U23775 ( .B1(n22099), .B2(n21971), .A(n21970), .ZN(n21972) );
  OAI211_X1 U23776 ( .C1(n21975), .C2(n21974), .A(n21973), .B(n21972), .ZN(
        P1_U3029) );
  AOI211_X1 U23777 ( .C1(n21977), .C2(n22045), .A(n21976), .B(n22015), .ZN(
        n21991) );
  AOI22_X1 U23778 ( .A1(n22126), .A2(n22098), .B1(n22108), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n21985) );
  AOI22_X1 U23779 ( .A1(n21980), .A2(n21979), .B1(n22005), .B2(n21978), .ZN(
        n21993) );
  AOI211_X1 U23780 ( .C1(n21986), .C2(n21992), .A(n21993), .B(n21981), .ZN(
        n21982) );
  AOI21_X1 U23781 ( .B1(n21983), .B2(n22099), .A(n21982), .ZN(n21984) );
  OAI211_X1 U23782 ( .C1(n21991), .C2(n21986), .A(n21985), .B(n21984), .ZN(
        P1_U3027) );
  INV_X1 U23783 ( .A(n21987), .ZN(n21988) );
  AOI222_X1 U23784 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n22108), .B1(n22098), 
        .B2(n21989), .C1(n22099), .C2(n21988), .ZN(n21990) );
  OAI221_X1 U23785 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21993), .C1(
        n21992), .C2(n21991), .A(n21990), .ZN(P1_U3028) );
  NOR3_X1 U23786 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21995), .A3(
        n21994), .ZN(n22008) );
  AOI21_X1 U23787 ( .B1(n21995), .B2(n22045), .A(n22015), .ZN(n22011) );
  OAI21_X1 U23788 ( .B1(n22012), .B2(n22049), .A(n22011), .ZN(n22000) );
  NOR2_X1 U23789 ( .A1(n22008), .A2(n22000), .ZN(n22048) );
  AOI22_X1 U23790 ( .A1(n22156), .A2(n22098), .B1(n22108), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n21998) );
  AOI22_X1 U23791 ( .A1(n21996), .A2(n22099), .B1(n22060), .B2(n21999), .ZN(
        n21997) );
  OAI211_X1 U23792 ( .C1(n22048), .C2(n21999), .A(n21998), .B(n21997), .ZN(
        P1_U3025) );
  AOI22_X1 U23793 ( .A1(n22001), .A2(n22099), .B1(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n22000), .ZN(n22010) );
  INV_X1 U23794 ( .A(n22002), .ZN(n22003) );
  NAND3_X1 U23795 ( .A1(n22005), .A2(n22004), .A3(n22003), .ZN(n22006) );
  OAI21_X1 U23796 ( .B1(n22145), .B2(n22067), .A(n22006), .ZN(n22007) );
  AOI211_X1 U23797 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n22108), .A(n22008), .B(
        n22007), .ZN(n22009) );
  NAND2_X1 U23798 ( .A1(n22010), .A2(n22009), .ZN(P1_U3026) );
  NAND2_X1 U23799 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n22060), .ZN(
        n22023) );
  NAND3_X1 U23800 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n22012), .A3(
        n22011), .ZN(n22013) );
  OAI21_X1 U23801 ( .B1(n22015), .B2(n22014), .A(n22013), .ZN(n22029) );
  AOI222_X1 U23802 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22108), .B1(n22098), 
        .B2(n22017), .C1(n22099), .C2(n22016), .ZN(n22018) );
  OAI221_X1 U23803 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n22023), .C1(
        n22024), .C2(n22029), .A(n22018), .ZN(P1_U3024) );
  INV_X1 U23804 ( .A(n22019), .ZN(n22020) );
  AOI21_X1 U23805 ( .B1(n22021), .B2(n22098), .A(n22020), .ZN(n22028) );
  INV_X1 U23806 ( .A(n22022), .ZN(n22026) );
  AOI221_X1 U23807 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n22030), .C2(n22024), .A(
        n22023), .ZN(n22025) );
  AOI21_X1 U23808 ( .B1(n22026), .B2(n22099), .A(n22025), .ZN(n22027) );
  OAI211_X1 U23809 ( .C1(n22030), .C2(n22029), .A(n22028), .B(n22027), .ZN(
        P1_U3023) );
  NAND2_X1 U23810 ( .A1(n22033), .A2(n22060), .ZN(n22037) );
  INV_X1 U23811 ( .A(n22031), .ZN(n22032) );
  AOI21_X1 U23812 ( .B1(n22179), .B2(n22098), .A(n22032), .ZN(n22036) );
  OAI21_X1 U23813 ( .B1(n22033), .B2(n22071), .A(n22048), .ZN(n22040) );
  AOI22_X1 U23814 ( .A1(n22034), .A2(n22099), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n22040), .ZN(n22035) );
  OAI211_X1 U23815 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n22037), .A(
        n22036), .B(n22035), .ZN(P1_U3022) );
  AOI22_X1 U23816 ( .A1(n22189), .A2(n22098), .B1(n22108), .B2(
        P1_REIP_REG_10__SCAN_IN), .ZN(n22042) );
  AOI221_X1 U23817 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n22038), .C2(n14002), .A(
        n22037), .ZN(n22039) );
  AOI21_X1 U23818 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n22040), .A(
        n22039), .ZN(n22041) );
  OAI211_X1 U23819 ( .C1(n22084), .C2(n22043), .A(n22042), .B(n22041), .ZN(
        P1_U3021) );
  INV_X1 U23820 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n22218) );
  NOR2_X1 U23821 ( .A1(n22044), .A2(n22218), .ZN(n22056) );
  NOR2_X1 U23822 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n22046), .ZN(
        n22061) );
  NAND2_X1 U23823 ( .A1(n22046), .A2(n22045), .ZN(n22047) );
  OAI211_X1 U23824 ( .C1(n22051), .C2(n22049), .A(n22048), .B(n22047), .ZN(
        n22062) );
  AOI21_X1 U23825 ( .B1(n22050), .B2(n22061), .A(n22062), .ZN(n22054) );
  NAND3_X1 U23826 ( .A1(n22051), .A2(n22060), .A3(n22053), .ZN(n22052) );
  OAI21_X1 U23827 ( .B1(n22054), .B2(n22053), .A(n22052), .ZN(n22055) );
  AOI211_X1 U23828 ( .C1(n22213), .C2(n22098), .A(n22056), .B(n22055), .ZN(
        n22057) );
  OAI21_X1 U23829 ( .B1(n22058), .B2(n22084), .A(n22057), .ZN(P1_U3019) );
  AOI21_X1 U23830 ( .B1(n22202), .B2(n22098), .A(n22059), .ZN(n22064) );
  AOI22_X1 U23831 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n22062), .B1(
        n22061), .B2(n22060), .ZN(n22063) );
  OAI211_X1 U23832 ( .C1(n22065), .C2(n22084), .A(n22064), .B(n22063), .ZN(
        P1_U3020) );
  OAI22_X1 U23833 ( .A1(n22068), .A2(n22084), .B1(n22067), .B2(n22066), .ZN(
        n22069) );
  INV_X1 U23834 ( .A(n22069), .ZN(n22077) );
  NAND2_X1 U23835 ( .A1(n22108), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n22076) );
  OAI21_X1 U23836 ( .B1(n22073), .B2(n22071), .A(n22070), .ZN(n22081) );
  NAND2_X1 U23837 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n22081), .ZN(
        n22075) );
  INV_X1 U23838 ( .A(n22079), .ZN(n22090) );
  NAND3_X1 U23839 ( .A1(n22073), .A2(n22072), .A3(n22090), .ZN(n22074) );
  NAND4_X1 U23840 ( .A1(n22077), .A2(n22076), .A3(n22075), .A4(n22074), .ZN(
        P1_U3013) );
  OAI21_X1 U23841 ( .B1(n22079), .B2(n22078), .A(n14281), .ZN(n22080) );
  AOI22_X1 U23842 ( .A1(n22081), .A2(n22080), .B1(n22098), .B2(n22254), .ZN(
        n22083) );
  NAND2_X1 U23843 ( .A1(n22108), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n22082) );
  OAI211_X1 U23844 ( .C1(n22085), .C2(n22084), .A(n22083), .B(n22082), .ZN(
        P1_U3014) );
  AOI22_X1 U23845 ( .A1(n22087), .A2(n22099), .B1(n22098), .B2(n22086), .ZN(
        n22094) );
  NAND2_X1 U23846 ( .A1(n22108), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n22093) );
  OAI21_X1 U23847 ( .B1(n22089), .B2(n22088), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n22092) );
  NAND3_X1 U23848 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n14000), .A3(
        n22090), .ZN(n22091) );
  NAND4_X1 U23849 ( .A1(n22094), .A2(n22093), .A3(n22092), .A4(n22091), .ZN(
        P1_U3015) );
  INV_X1 U23850 ( .A(n22095), .ZN(n22100) );
  INV_X1 U23851 ( .A(n22096), .ZN(n22097) );
  AOI22_X1 U23852 ( .A1(n22100), .A2(n22099), .B1(n22098), .B2(n22097), .ZN(
        n22110) );
  AOI21_X1 U23853 ( .B1(n22103), .B2(n22102), .A(n22101), .ZN(n22107) );
  NOR3_X1 U23854 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n22105), .A3(
        n22104), .ZN(n22106) );
  AOI211_X1 U23855 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n22108), .A(n22107), 
        .B(n22106), .ZN(n22109) );
  NAND2_X1 U23856 ( .A1(n22110), .A2(n22109), .ZN(P1_U3009) );
  AOI21_X1 U23857 ( .B1(n22214), .B2(n14610), .A(n22190), .ZN(n22122) );
  INV_X1 U23858 ( .A(n22111), .ZN(n22112) );
  AOI22_X1 U23859 ( .A1(n22255), .A2(n22112), .B1(n22272), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n22121) );
  INV_X1 U23860 ( .A(n22113), .ZN(n22114) );
  AOI22_X1 U23861 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n22263), .B1(
        n22253), .B2(n22114), .ZN(n22116) );
  NAND3_X1 U23862 ( .A1(n22214), .A2(n22124), .A3(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n22115) );
  OAI211_X1 U23863 ( .C1(n14673), .C2(n22117), .A(n22116), .B(n22115), .ZN(
        n22118) );
  AOI21_X1 U23864 ( .B1(n22119), .B2(n22147), .A(n22118), .ZN(n22120) );
  OAI211_X1 U23865 ( .C1(n22122), .C2(n22124), .A(n22121), .B(n22120), .ZN(
        P1_U2838) );
  AOI21_X1 U23866 ( .B1(n22214), .B2(n22139), .A(n22190), .ZN(n22151) );
  NOR3_X1 U23867 ( .A1(n14610), .A2(n22124), .A3(n22123), .ZN(n22125) );
  AOI21_X1 U23868 ( .B1(n22125), .B2(n22214), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n22134) );
  AOI21_X1 U23869 ( .B1(n22263), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n22251), .ZN(n22128) );
  NAND2_X1 U23870 ( .A1(n22255), .A2(n22126), .ZN(n22127) );
  OAI211_X1 U23871 ( .C1(n22249), .C2(n22129), .A(n22128), .B(n22127), .ZN(
        n22130) );
  AOI21_X1 U23872 ( .B1(n22132), .B2(n22131), .A(n22130), .ZN(n22133) );
  OAI21_X1 U23873 ( .B1(n22151), .B2(n22134), .A(n22133), .ZN(n22135) );
  AOI21_X1 U23874 ( .B1(n22136), .B2(n22147), .A(n22135), .ZN(n22137) );
  OAI21_X1 U23875 ( .B1(n22138), .B2(n22267), .A(n22137), .ZN(P1_U2836) );
  NOR3_X1 U23876 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n22139), .A3(n22200), .ZN(
        n22140) );
  AOI211_X1 U23877 ( .C1(n22263), .C2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n22251), .B(n22140), .ZN(n22144) );
  INV_X1 U23878 ( .A(n22141), .ZN(n22142) );
  AOI22_X1 U23879 ( .A1(n22272), .A2(P1_EBX_REG_5__SCAN_IN), .B1(n22142), .B2(
        n22253), .ZN(n22143) );
  OAI211_X1 U23880 ( .C1(n22278), .C2(n22145), .A(n22144), .B(n22143), .ZN(
        n22146) );
  AOI21_X1 U23881 ( .B1(n22148), .B2(n22147), .A(n22146), .ZN(n22149) );
  OAI21_X1 U23882 ( .B1(n22151), .B2(n22150), .A(n22149), .ZN(P1_U2835) );
  AOI21_X1 U23883 ( .B1(n22214), .B2(n22163), .A(n22190), .ZN(n22174) );
  AOI21_X1 U23884 ( .B1(n22152), .B2(n22214), .A(P1_REIP_REG_6__SCAN_IN), .ZN(
        n22162) );
  OAI22_X1 U23885 ( .A1(n22249), .A2(n22154), .B1(n22153), .B2(n22246), .ZN(
        n22155) );
  AOI211_X1 U23886 ( .C1(n22255), .C2(n22156), .A(n22251), .B(n22155), .ZN(
        n22161) );
  INV_X1 U23887 ( .A(n22157), .ZN(n22158) );
  AOI22_X1 U23888 ( .A1(n22159), .A2(n22256), .B1(n22158), .B2(n22253), .ZN(
        n22160) );
  OAI211_X1 U23889 ( .C1(n22174), .C2(n22162), .A(n22161), .B(n22160), .ZN(
        P1_U2834) );
  NOR3_X1 U23890 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n22163), .A3(n22200), .ZN(
        n22164) );
  AOI211_X1 U23891 ( .C1(n22263), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n22251), .B(n22164), .ZN(n22168) );
  INV_X1 U23892 ( .A(n22165), .ZN(n22166) );
  AOI22_X1 U23893 ( .A1(n22272), .A2(P1_EBX_REG_7__SCAN_IN), .B1(n22166), .B2(
        n22253), .ZN(n22167) );
  OAI211_X1 U23894 ( .C1(n22278), .C2(n22169), .A(n22168), .B(n22167), .ZN(
        n22170) );
  AOI21_X1 U23895 ( .B1(n22171), .B2(n22256), .A(n22170), .ZN(n22172) );
  OAI21_X1 U23896 ( .B1(n22174), .B2(n22173), .A(n22172), .ZN(P1_U2833) );
  NOR3_X1 U23897 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n22175), .A3(n22200), .ZN(
        n22176) );
  AOI211_X1 U23898 ( .C1(n22263), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n22176), .B(n22251), .ZN(n22177) );
  OAI21_X1 U23899 ( .B1(n22249), .B2(n14252), .A(n22177), .ZN(n22178) );
  AOI21_X1 U23900 ( .B1(n22179), .B2(n22255), .A(n22178), .ZN(n22180) );
  OAI21_X1 U23901 ( .B1(n22181), .B2(n22268), .A(n22180), .ZN(n22182) );
  AOI21_X1 U23902 ( .B1(n22183), .B2(n22253), .A(n22182), .ZN(n22184) );
  OAI21_X1 U23903 ( .B1(n22186), .B2(n22185), .A(n22184), .ZN(P1_U2831) );
  AND2_X1 U23904 ( .A1(n22201), .A2(n22214), .ZN(n22187) );
  AOI22_X1 U23905 ( .A1(n22255), .A2(n22189), .B1(n22188), .B2(n22187), .ZN(
        n22199) );
  OAI21_X1 U23906 ( .B1(n22190), .B2(n22201), .A(n22273), .ZN(n22212) );
  OAI22_X1 U23907 ( .A1(n22212), .A2(n22192), .B1(n22191), .B2(n22249), .ZN(
        n22193) );
  AOI211_X1 U23908 ( .C1(n22263), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n22251), .B(n22193), .ZN(n22198) );
  OAI22_X1 U23909 ( .A1(n22195), .A2(n22268), .B1(n22194), .B2(n22267), .ZN(
        n22196) );
  INV_X1 U23910 ( .A(n22196), .ZN(n22197) );
  NAND3_X1 U23911 ( .A1(n22199), .A2(n22198), .A3(n22197), .ZN(P1_U2830) );
  NOR3_X1 U23912 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n22201), .A3(n22200), 
        .ZN(n22209) );
  INV_X1 U23913 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n22204) );
  AOI22_X1 U23914 ( .A1(n22202), .A2(n22255), .B1(n22272), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n22203) );
  OAI211_X1 U23915 ( .C1(n22246), .C2(n22204), .A(n22203), .B(n22264), .ZN(
        n22208) );
  OAI22_X1 U23916 ( .A1(n22206), .A2(n22267), .B1(n22268), .B2(n22205), .ZN(
        n22207) );
  NOR3_X1 U23917 ( .A1(n22209), .A2(n22208), .A3(n22207), .ZN(n22210) );
  OAI21_X1 U23918 ( .B1(n22212), .B2(n22211), .A(n22210), .ZN(P1_U2829) );
  AOI22_X1 U23919 ( .A1(n22213), .A2(n22255), .B1(n22272), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n22224) );
  NAND3_X1 U23920 ( .A1(n22218), .A2(n22215), .A3(n22214), .ZN(n22216) );
  OAI21_X1 U23921 ( .B1(n22218), .B2(n22217), .A(n22216), .ZN(n22219) );
  AOI211_X1 U23922 ( .C1(n22263), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n22251), .B(n22219), .ZN(n22223) );
  AOI22_X1 U23923 ( .A1(n22221), .A2(n22253), .B1(n22256), .B2(n22220), .ZN(
        n22222) );
  NAND3_X1 U23924 ( .A1(n22224), .A2(n22223), .A3(n22222), .ZN(P1_U2828) );
  NAND2_X1 U23925 ( .A1(n22273), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n22226) );
  AOI21_X1 U23926 ( .B1(n22226), .B2(n22225), .A(n22235), .ZN(n22227) );
  AOI211_X1 U23927 ( .C1(n22272), .C2(P1_EBX_REG_15__SCAN_IN), .A(n22251), .B(
        n22227), .ZN(n22233) );
  OAI22_X1 U23928 ( .A1(n22229), .A2(n22268), .B1(n22278), .B2(n22228), .ZN(
        n22230) );
  AOI21_X1 U23929 ( .B1(n22231), .B2(n22253), .A(n22230), .ZN(n22232) );
  OAI211_X1 U23930 ( .C1(n22234), .C2(n22246), .A(n22233), .B(n22232), .ZN(
        P1_U2825) );
  AOI21_X1 U23931 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(n22273), .A(n22235), 
        .ZN(n22245) );
  OAI22_X1 U23932 ( .A1(n22249), .A2(n22237), .B1(n22246), .B2(n22236), .ZN(
        n22238) );
  AOI211_X1 U23933 ( .C1(n22253), .C2(n22239), .A(n22251), .B(n22238), .ZN(
        n22244) );
  OAI22_X1 U23934 ( .A1(n22241), .A2(n22268), .B1(n22278), .B2(n22240), .ZN(
        n22242) );
  INV_X1 U23935 ( .A(n22242), .ZN(n22243) );
  OAI211_X1 U23936 ( .C1(n22259), .C2(n22245), .A(n22244), .B(n22243), .ZN(
        P1_U2824) );
  OAI22_X1 U23937 ( .A1(n22249), .A2(n22248), .B1(n22247), .B2(n22246), .ZN(
        n22250) );
  AOI211_X1 U23938 ( .C1(n22253), .C2(n22252), .A(n22251), .B(n22250), .ZN(
        n22262) );
  AOI22_X1 U23939 ( .A1(n22257), .A2(n22256), .B1(n22255), .B2(n22254), .ZN(
        n22261) );
  OAI21_X1 U23940 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n22259), .A(n22258), 
        .ZN(n22260) );
  NAND3_X1 U23941 ( .A1(n22262), .A2(n22261), .A3(n22260), .ZN(P1_U2823) );
  NAND2_X1 U23942 ( .A1(n22263), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n22265) );
  OAI211_X1 U23943 ( .C1(n22267), .C2(n22266), .A(n22265), .B(n22264), .ZN(
        n22271) );
  NOR2_X1 U23944 ( .A1(n22269), .A2(n22268), .ZN(n22270) );
  AOI211_X1 U23945 ( .C1(n22272), .C2(P1_EBX_REG_19__SCAN_IN), .A(n22271), .B(
        n22270), .ZN(n22277) );
  NAND2_X1 U23946 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n22275), .ZN(n22274) );
  OAI211_X1 U23947 ( .C1(P1_REIP_REG_19__SCAN_IN), .C2(n22275), .A(n22274), 
        .B(n22273), .ZN(n22276) );
  OAI211_X1 U23948 ( .C1(n22279), .C2(n22278), .A(n22277), .B(n22276), .ZN(
        P1_U2821) );
  OAI21_X1 U23949 ( .B1(n22281), .B2(n14721), .A(n22280), .ZN(P1_U2806) );
  AOI22_X1 U23950 ( .A1(n13179), .A2(n22298), .B1(n14517), .B2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n22282) );
  OAI21_X1 U23951 ( .B1(n22283), .B2(n22289), .A(n22282), .ZN(n22285) );
  AOI22_X1 U23952 ( .A1(n22286), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n22285), .B2(n22284), .ZN(n22287) );
  OAI21_X1 U23953 ( .B1(n22289), .B2(n22288), .A(n22287), .ZN(P1_U3474) );
  NAND2_X1 U23954 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n22605), .ZN(n22292) );
  OAI211_X1 U23955 ( .C1(n22293), .C2(n22292), .A(n22291), .B(n22290), .ZN(
        P1_U3163) );
  OAI21_X1 U23956 ( .B1(n22295), .B2(n13173), .A(n22294), .ZN(P1_U3466) );
  AOI21_X1 U23957 ( .B1(n22298), .B2(n22297), .A(n22296), .ZN(n22299) );
  OAI22_X1 U23958 ( .A1(n22301), .A2(n22300), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n22299), .ZN(n22302) );
  OAI21_X1 U23959 ( .B1(n22304), .B2(n22303), .A(n22302), .ZN(P1_U3161) );
  INV_X1 U23960 ( .A(n22305), .ZN(n22306) );
  OAI21_X1 U23961 ( .B1(n22308), .B2(n22590), .A(n22306), .ZN(P1_U2805) );
  OAI21_X1 U23962 ( .B1(n22308), .B2(n22307), .A(n22306), .ZN(P1_U3465) );
  INV_X1 U23963 ( .A(n22309), .ZN(n22310) );
  OAI21_X1 U23964 ( .B1(n22312), .B2(n19841), .A(n22310), .ZN(P2_U2818) );
  OAI21_X1 U23965 ( .B1(n22312), .B2(n22311), .A(n22310), .ZN(P2_U3592) );
  INV_X1 U23966 ( .A(n22313), .ZN(n22315) );
  OAI21_X1 U23967 ( .B1(n22317), .B2(n22314), .A(n22315), .ZN(P3_U2636) );
  OAI21_X1 U23968 ( .B1(n22317), .B2(n22316), .A(n22315), .ZN(P3_U3281) );
  INV_X1 U23969 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22318) );
  AOI21_X1 U23970 ( .B1(HOLD), .B2(n22319), .A(n22318), .ZN(n22322) );
  AOI21_X1 U23971 ( .B1(n22321), .B2(P3_STATE_REG_1__SCAN_IN), .A(n22320), 
        .ZN(n22383) );
  AOI21_X1 U23972 ( .B1(n22369), .B2(NA), .A(n22377), .ZN(n22381) );
  OAI22_X1 U23973 ( .A1(n22323), .A2(n22322), .B1(n22383), .B2(n22381), .ZN(
        P3_U3029) );
  OAI21_X1 U23974 ( .B1(NA), .B2(n22325), .A(n22324), .ZN(n22326) );
  OAI211_X1 U23975 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n22328), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n22326), .ZN(n22333) );
  INV_X1 U23976 ( .A(HOLD), .ZN(n22376) );
  NAND2_X1 U23977 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n22327), .ZN(n22337) );
  INV_X1 U23978 ( .A(n22337), .ZN(n22340) );
  NOR2_X1 U23979 ( .A1(n22328), .A2(n22337), .ZN(n22329) );
  MUX2_X1 U23980 ( .A(P1_STATE_REG_2__SCAN_IN), .B(n22329), .S(
        P1_STATE_REG_0__SCAN_IN), .Z(n22330) );
  AOI22_X1 U23981 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22340), .B1(n22330), 
        .B2(n22378), .ZN(n22332) );
  OAI211_X1 U23982 ( .C1(n22333), .C2(n22376), .A(n22332), .B(n22331), .ZN(
        P1_U3196) );
  OAI21_X1 U23983 ( .B1(n22335), .B2(n22376), .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n22341) );
  INV_X1 U23984 ( .A(n22341), .ZN(n22336) );
  NOR2_X1 U23985 ( .A1(n22334), .A2(n22376), .ZN(n22342) );
  AOI22_X1 U23986 ( .A1(n22336), .A2(P1_STATE_REG_0__SCAN_IN), .B1(n22342), 
        .B2(n22335), .ZN(n22339) );
  NAND3_X1 U23987 ( .A1(n22339), .A2(n22338), .A3(n22337), .ZN(P1_U3195) );
  NOR2_X1 U23988 ( .A1(n22340), .A2(n22343), .ZN(n22345) );
  AOI211_X1 U23989 ( .C1(NA), .C2(n22343), .A(n22342), .B(n22341), .ZN(n22344)
         );
  OAI22_X1 U23990 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n22345), .B1(n22853), 
        .B2(n22344), .ZN(P1_U3194) );
  NAND3_X1 U23991 ( .A1(n22347), .A2(HOLD), .A3(n22346), .ZN(n22353) );
  OAI21_X1 U23992 ( .B1(n22349), .B2(n22348), .A(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n22361) );
  OAI21_X1 U23993 ( .B1(n22350), .B2(n22378), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n22367) );
  AOI22_X1 U23994 ( .A1(n22355), .A2(n22351), .B1(n22361), .B2(n22367), .ZN(
        n22352) );
  NAND2_X1 U23995 ( .A1(n22353), .A2(n22352), .ZN(P2_U3209) );
  NOR2_X1 U23996 ( .A1(n22354), .A2(n22376), .ZN(n22364) );
  NOR3_X1 U23997 ( .A1(n22364), .A2(n22355), .A3(n22366), .ZN(n22357) );
  AOI211_X1 U23998 ( .C1(n22358), .C2(HOLD), .A(n22357), .B(n22356), .ZN(
        n22360) );
  NAND2_X1 U23999 ( .A1(n22359), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n22362) );
  NAND2_X1 U24000 ( .A1(n22360), .A2(n22362), .ZN(P2_U3210) );
  INV_X1 U24001 ( .A(n22361), .ZN(n22368) );
  OAI22_X1 U24002 ( .A1(NA), .A2(n22362), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22363) );
  OAI22_X1 U24003 ( .A1(n22364), .A2(n22363), .B1(HOLD), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n22365) );
  OAI22_X1 U24004 ( .A1(n22368), .A2(n22367), .B1(n22366), .B2(n22365), .ZN(
        P2_U3211) );
  OAI211_X1 U24005 ( .C1(n22376), .C2(n22377), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22374) );
  NOR2_X1 U24006 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n22385)
         );
  NOR3_X1 U24007 ( .A1(n22369), .A2(P3_STATE_REG_2__SCAN_IN), .A3(n22385), 
        .ZN(n22372) );
  NOR2_X1 U24008 ( .A1(n22370), .A2(n22369), .ZN(n22379) );
  AOI211_X1 U24009 ( .C1(n22372), .C2(n22375), .A(n22371), .B(n22379), .ZN(
        n22373) );
  OAI211_X1 U24010 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n22375), .A(n22374), 
        .B(n22373), .ZN(P3_U3030) );
  OAI22_X1 U24011 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n22377), .B2(n22376), .ZN(n22380)
         );
  OAI221_X1 U24012 ( .B1(n22380), .B2(n22379), .C1(n22380), .C2(n22378), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n22384) );
  INV_X1 U24013 ( .A(n22381), .ZN(n22382) );
  OAI22_X1 U24014 ( .A1(n22385), .A2(n22384), .B1(n22383), .B2(n22382), .ZN(
        P3_U3031) );
  NOR2_X1 U24015 ( .A1(n22478), .A2(n22386), .ZN(n22389) );
  AOI21_X1 U24016 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n22456), .A(n22389), 
        .ZN(n22387) );
  OAI21_X1 U24017 ( .B1(n22388), .B2(n22484), .A(n22387), .ZN(P1_U2937) );
  AOI21_X1 U24018 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n22456), .A(n22389), 
        .ZN(n22390) );
  OAI21_X1 U24019 ( .B1(n22391), .B2(n22484), .A(n22390), .ZN(P1_U2952) );
  NOR2_X1 U24020 ( .A1(n22478), .A2(n22392), .ZN(n22395) );
  AOI21_X1 U24021 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n22456), .A(n22395), 
        .ZN(n22393) );
  OAI21_X1 U24022 ( .B1(n22394), .B2(n22484), .A(n22393), .ZN(P1_U2938) );
  AOI21_X1 U24023 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n22456), .A(n22395), 
        .ZN(n22396) );
  OAI21_X1 U24024 ( .B1(n22397), .B2(n22484), .A(n22396), .ZN(P1_U2953) );
  NOR2_X1 U24025 ( .A1(n22478), .A2(n22398), .ZN(n22401) );
  AOI21_X1 U24026 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n22456), .A(n22401), 
        .ZN(n22399) );
  OAI21_X1 U24027 ( .B1(n22400), .B2(n22484), .A(n22399), .ZN(P1_U2939) );
  AOI21_X1 U24028 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n22456), .A(n22401), 
        .ZN(n22402) );
  OAI21_X1 U24029 ( .B1(n22403), .B2(n22484), .A(n22402), .ZN(P1_U2954) );
  NOR2_X1 U24030 ( .A1(n22478), .A2(n22404), .ZN(n22407) );
  AOI21_X1 U24031 ( .B1(P1_UWORD_REG_3__SCAN_IN), .B2(n22456), .A(n22407), 
        .ZN(n22405) );
  OAI21_X1 U24032 ( .B1(n22406), .B2(n22484), .A(n22405), .ZN(P1_U2940) );
  AOI21_X1 U24033 ( .B1(P1_LWORD_REG_3__SCAN_IN), .B2(n22456), .A(n22407), 
        .ZN(n22408) );
  OAI21_X1 U24034 ( .B1(n22409), .B2(n22484), .A(n22408), .ZN(P1_U2955) );
  INV_X1 U24035 ( .A(n22410), .ZN(n22411) );
  NOR2_X1 U24036 ( .A1(n22478), .A2(n22411), .ZN(n22415) );
  AOI21_X1 U24037 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n22456), .A(n22415), 
        .ZN(n22412) );
  OAI21_X1 U24038 ( .B1(n22413), .B2(n22484), .A(n22412), .ZN(P1_U2941) );
  AOI21_X1 U24039 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n22479), .A(n22415), 
        .ZN(n22416) );
  OAI21_X1 U24040 ( .B1(n22417), .B2(n22484), .A(n22416), .ZN(P1_U2956) );
  NOR2_X1 U24041 ( .A1(n22478), .A2(n22418), .ZN(n22421) );
  AOI21_X1 U24042 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n22479), .A(n22421), 
        .ZN(n22419) );
  OAI21_X1 U24043 ( .B1(n22420), .B2(n22484), .A(n22419), .ZN(P1_U2942) );
  AOI21_X1 U24044 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n22479), .A(n22421), 
        .ZN(n22422) );
  OAI21_X1 U24045 ( .B1(n13399), .B2(n22484), .A(n22422), .ZN(P1_U2957) );
  NOR2_X1 U24046 ( .A1(n22478), .A2(n22423), .ZN(n22426) );
  AOI21_X1 U24047 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n22479), .A(n22426), 
        .ZN(n22424) );
  OAI21_X1 U24048 ( .B1(n22425), .B2(n22484), .A(n22424), .ZN(P1_U2943) );
  AOI21_X1 U24049 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n22479), .A(n22426), 
        .ZN(n22427) );
  OAI21_X1 U24050 ( .B1(n15299), .B2(n22484), .A(n22427), .ZN(P1_U2958) );
  NOR2_X1 U24051 ( .A1(n22478), .A2(n22428), .ZN(n22431) );
  AOI21_X1 U24052 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n22479), .A(n22431), 
        .ZN(n22429) );
  OAI21_X1 U24053 ( .B1(n22430), .B2(n22484), .A(n22429), .ZN(P1_U2944) );
  AOI21_X1 U24054 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n22479), .A(n22431), 
        .ZN(n22432) );
  OAI21_X1 U24055 ( .B1(n13411), .B2(n22484), .A(n22432), .ZN(P1_U2959) );
  INV_X1 U24056 ( .A(n22433), .ZN(n22434) );
  NOR2_X1 U24057 ( .A1(n22478), .A2(n22434), .ZN(n22437) );
  AOI21_X1 U24058 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n22479), .A(n22437), 
        .ZN(n22435) );
  OAI21_X1 U24059 ( .B1(n22436), .B2(n22484), .A(n22435), .ZN(P1_U2945) );
  AOI21_X1 U24060 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n22479), .A(n22437), 
        .ZN(n22438) );
  OAI21_X1 U24061 ( .B1(n22439), .B2(n22484), .A(n22438), .ZN(P1_U2960) );
  INV_X1 U24062 ( .A(n22440), .ZN(n22441) );
  NOR2_X1 U24063 ( .A1(n22478), .A2(n22441), .ZN(n22444) );
  AOI21_X1 U24064 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n22456), .A(n22444), 
        .ZN(n22442) );
  OAI21_X1 U24065 ( .B1(n22443), .B2(n22484), .A(n22442), .ZN(P1_U2946) );
  AOI21_X1 U24066 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n22456), .A(n22444), 
        .ZN(n22445) );
  OAI21_X1 U24067 ( .B1(n22446), .B2(n22484), .A(n22445), .ZN(P1_U2961) );
  INV_X1 U24068 ( .A(n22447), .ZN(n22448) );
  NOR2_X1 U24069 ( .A1(n22478), .A2(n22448), .ZN(n22451) );
  AOI21_X1 U24070 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n22456), .A(n22451), 
        .ZN(n22449) );
  OAI21_X1 U24071 ( .B1(n22450), .B2(n22484), .A(n22449), .ZN(P1_U2947) );
  AOI21_X1 U24072 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n22456), .A(n22451), 
        .ZN(n22452) );
  OAI21_X1 U24073 ( .B1(n22453), .B2(n22484), .A(n22452), .ZN(P1_U2962) );
  INV_X1 U24074 ( .A(n22454), .ZN(n22455) );
  NOR2_X1 U24075 ( .A1(n22478), .A2(n22455), .ZN(n22459) );
  AOI21_X1 U24076 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n22456), .A(n22459), 
        .ZN(n22457) );
  OAI21_X1 U24077 ( .B1(n22458), .B2(n22484), .A(n22457), .ZN(P1_U2948) );
  AOI21_X1 U24078 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n22479), .A(n22459), 
        .ZN(n22460) );
  OAI21_X1 U24079 ( .B1(n22461), .B2(n22484), .A(n22460), .ZN(P1_U2963) );
  INV_X1 U24080 ( .A(n22462), .ZN(n22463) );
  NOR2_X1 U24081 ( .A1(n22478), .A2(n22463), .ZN(n22466) );
  AOI21_X1 U24082 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n22456), .A(n22466), 
        .ZN(n22464) );
  OAI21_X1 U24083 ( .B1(n22465), .B2(n22484), .A(n22464), .ZN(P1_U2949) );
  AOI21_X1 U24084 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n22479), .A(n22466), 
        .ZN(n22467) );
  OAI21_X1 U24085 ( .B1(n22468), .B2(n22484), .A(n22467), .ZN(P1_U2964) );
  INV_X1 U24086 ( .A(n22469), .ZN(n22470) );
  NOR2_X1 U24087 ( .A1(n22478), .A2(n22470), .ZN(n22473) );
  AOI21_X1 U24088 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n22456), .A(n22473), 
        .ZN(n22471) );
  OAI21_X1 U24089 ( .B1(n22472), .B2(n22484), .A(n22471), .ZN(P1_U2950) );
  AOI21_X1 U24090 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n22456), .A(n22473), 
        .ZN(n22474) );
  OAI21_X1 U24091 ( .B1(n22475), .B2(n22484), .A(n22474), .ZN(P1_U2965) );
  INV_X1 U24092 ( .A(n22476), .ZN(n22477) );
  NOR2_X1 U24093 ( .A1(n22478), .A2(n22477), .ZN(n22482) );
  AOI21_X1 U24094 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n22479), .A(n22482), 
        .ZN(n22480) );
  OAI21_X1 U24095 ( .B1(n22481), .B2(n22484), .A(n22480), .ZN(P1_U2951) );
  AOI21_X1 U24096 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n22456), .A(n22482), 
        .ZN(n22483) );
  OAI21_X1 U24097 ( .B1(n22485), .B2(n22484), .A(n22483), .ZN(P1_U2966) );
  NOR2_X1 U24098 ( .A1(n22487), .A2(n22486), .ZN(n22488) );
  NOR2_X1 U24099 ( .A1(n22844), .A2(n22607), .ZN(n22489) );
  NOR2_X1 U24100 ( .A1(n22607), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n22566) );
  AOI21_X1 U24101 ( .B1(n22490), .B2(n22489), .A(n22566), .ZN(n22498) );
  INV_X1 U24102 ( .A(n22498), .ZN(n22491) );
  NOR2_X1 U24103 ( .A1(n22515), .A2(n22593), .ZN(n22497) );
  NOR2_X1 U24104 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22492), .ZN(
        n22782) );
  AOI22_X1 U24105 ( .A1(n22844), .A2(n22598), .B1(n22782), .B2(n22608), .ZN(
        n22500) );
  INV_X1 U24106 ( .A(n22782), .ZN(n22495) );
  INV_X1 U24107 ( .A(n22507), .ZN(n22546) );
  NOR2_X1 U24108 ( .A1(n22493), .A2(n22605), .ZN(n22494) );
  AOI211_X1 U24109 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22495), .A(n22546), 
        .B(n22494), .ZN(n22496) );
  OAI21_X1 U24110 ( .B1(n22498), .B2(n22497), .A(n22496), .ZN(n22784) );
  AOI22_X1 U24111 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n22783), .B2(n22616), .ZN(n22499) );
  OAI211_X1 U24112 ( .C1(n22787), .C2(n22581), .A(n22500), .B(n22499), .ZN(
        P1_U3033) );
  NOR2_X1 U24113 ( .A1(n22796), .A2(n22607), .ZN(n22503) );
  AOI21_X1 U24114 ( .B1(n22503), .B2(n22502), .A(n22566), .ZN(n22509) );
  INV_X1 U24115 ( .A(n22509), .ZN(n22504) );
  NOR2_X1 U24116 ( .A1(n22515), .A2(n14636), .ZN(n22508) );
  NOR3_X1 U24117 ( .A1(n22584), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22519) );
  NAND2_X1 U24118 ( .A1(n22571), .A2(n22519), .ZN(n22505) );
  INV_X1 U24119 ( .A(n22505), .ZN(n22788) );
  AOI22_X1 U24120 ( .A1(n22796), .A2(n22616), .B1(n22608), .B2(n22788), .ZN(
        n22511) );
  NOR2_X1 U24121 ( .A1(n11710), .A2(n22605), .ZN(n22532) );
  AOI21_X1 U24122 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22505), .A(n22532), 
        .ZN(n22506) );
  OAI211_X1 U24123 ( .C1(n22509), .C2(n22508), .A(n22507), .B(n22506), .ZN(
        n22790) );
  AOI22_X1 U24124 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n22789), .B2(n22598), .ZN(n22510) );
  OAI211_X1 U24125 ( .C1(n22793), .C2(n22581), .A(n22511), .B(n22510), .ZN(
        P1_U3049) );
  INV_X1 U24126 ( .A(n22512), .ZN(n22514) );
  AOI21_X1 U24127 ( .B1(n22514), .B2(n22513), .A(n22607), .ZN(n22521) );
  INV_X1 U24128 ( .A(n22515), .ZN(n22517) );
  INV_X1 U24129 ( .A(n22519), .ZN(n22516) );
  NOR2_X1 U24130 ( .A1(n22571), .A2(n22516), .ZN(n22794) );
  AOI21_X1 U24131 ( .B1(n22517), .B2(n22603), .A(n22794), .ZN(n22522) );
  INV_X1 U24132 ( .A(n22522), .ZN(n22518) );
  AOI22_X1 U24133 ( .A1(n22795), .A2(n22616), .B1(n22794), .B2(n22608), .ZN(
        n22525) );
  OAI21_X1 U24134 ( .B1(n22563), .B2(n22519), .A(n22613), .ZN(n22520) );
  AOI21_X1 U24135 ( .B1(n22522), .B2(n22521), .A(n22520), .ZN(n22523) );
  AOI22_X1 U24136 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22797), .B1(
        n22796), .B2(n22598), .ZN(n22524) );
  OAI211_X1 U24137 ( .C1(n22800), .C2(n22581), .A(n22525), .B(n22524), .ZN(
        P1_U3057) );
  NOR2_X1 U24138 ( .A1(n22803), .A2(n22607), .ZN(n22527) );
  AOI21_X1 U24139 ( .B1(n22527), .B2(n22526), .A(n22566), .ZN(n22537) );
  INV_X1 U24140 ( .A(n22537), .ZN(n22529) );
  NOR2_X1 U24141 ( .A1(n22528), .A2(n14636), .ZN(n22536) );
  INV_X1 U24142 ( .A(n22530), .ZN(n22531) );
  NOR2_X1 U24143 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22531), .ZN(
        n22801) );
  AOI22_X1 U24144 ( .A1(n22803), .A2(n22616), .B1(n22801), .B2(n22608), .ZN(
        n22539) );
  INV_X1 U24145 ( .A(n22532), .ZN(n22533) );
  OAI211_X1 U24146 ( .C1(n13173), .C2(n22801), .A(n22533), .B(n22595), .ZN(
        n22534) );
  INV_X1 U24147 ( .A(n22534), .ZN(n22535) );
  OAI21_X1 U24148 ( .B1(n22537), .B2(n22536), .A(n22535), .ZN(n22804) );
  AOI22_X1 U24149 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n22802), .B2(n22598), .ZN(n22538) );
  OAI211_X1 U24150 ( .C1(n22807), .C2(n22581), .A(n22539), .B(n22538), .ZN(
        P1_U3081) );
  NOR2_X1 U24151 ( .A1(n22816), .A2(n22607), .ZN(n22541) );
  AOI21_X1 U24152 ( .B1(n22541), .B2(n22540), .A(n22566), .ZN(n22551) );
  INV_X1 U24153 ( .A(n22551), .ZN(n22545) );
  OR2_X1 U24154 ( .A1(n22542), .A2(n22586), .ZN(n22588) );
  INV_X1 U24155 ( .A(n22588), .ZN(n22543) );
  NOR3_X1 U24156 ( .A1(n22586), .A2(n22584), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n22562) );
  INV_X1 U24157 ( .A(n22562), .ZN(n22557) );
  NOR2_X1 U24158 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22557), .ZN(
        n22808) );
  AOI22_X1 U24159 ( .A1(n22816), .A2(n22616), .B1(n22808), .B2(n22608), .ZN(
        n22553) );
  INV_X1 U24160 ( .A(n22808), .ZN(n22548) );
  NAND2_X1 U24161 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n22588), .ZN(n22596) );
  INV_X1 U24162 ( .A(n22596), .ZN(n22547) );
  AOI211_X1 U24163 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n22548), .A(n22547), 
        .B(n22546), .ZN(n22549) );
  OAI21_X1 U24164 ( .B1(n22551), .B2(n22550), .A(n22549), .ZN(n22810) );
  AOI22_X1 U24165 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n22809), .B2(n22598), .ZN(n22552) );
  OAI211_X1 U24166 ( .C1(n22813), .C2(n22581), .A(n22553), .B(n22552), .ZN(
        P1_U3113) );
  NOR2_X1 U24167 ( .A1(n22571), .A2(n22557), .ZN(n22814) );
  AOI21_X1 U24168 ( .B1(n22556), .B2(n22603), .A(n22814), .ZN(n22558) );
  OAI22_X1 U24169 ( .A1(n22558), .A2(n22607), .B1(n22557), .B2(n22605), .ZN(
        n22815) );
  AOI22_X1 U24170 ( .A1(n22815), .A2(n22609), .B1(n22608), .B2(n22814), .ZN(
        n22565) );
  OAI211_X1 U24171 ( .C1(n11648), .C2(n22560), .A(n22559), .B(n22558), .ZN(
        n22561) );
  OAI211_X1 U24172 ( .C1(n22563), .C2(n22562), .A(n22613), .B(n22561), .ZN(
        n22817) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22598), .ZN(n22564) );
  OAI211_X1 U24174 ( .C1(n22601), .C2(n22820), .A(n22565), .B(n22564), .ZN(
        P1_U3121) );
  NAND3_X1 U24175 ( .A1(n22820), .A2(n22563), .A3(n22823), .ZN(n22568) );
  INV_X1 U24176 ( .A(n22566), .ZN(n22567) );
  NAND2_X1 U24177 ( .A1(n22568), .A2(n22567), .ZN(n22576) );
  AND2_X1 U24178 ( .A1(n22604), .A2(n14636), .ZN(n22574) );
  NAND2_X1 U24179 ( .A1(n22571), .A2(n22570), .ZN(n22822) );
  OAI22_X1 U24180 ( .A1(n22823), .A2(n22601), .B1(n22822), .B2(n22572), .ZN(
        n22573) );
  INV_X1 U24181 ( .A(n22573), .ZN(n22580) );
  INV_X1 U24182 ( .A(n22574), .ZN(n22575) );
  AOI22_X1 U24183 ( .A1(n22576), .A2(n22575), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22822), .ZN(n22577) );
  AOI22_X1 U24184 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22598), .ZN(n22579) );
  OAI211_X1 U24185 ( .C1(n22830), .C2(n22581), .A(n22580), .B(n22579), .ZN(
        P1_U3129) );
  NOR3_X1 U24186 ( .A1(n22586), .A2(n22585), .A3(n22584), .ZN(n22615) );
  INV_X1 U24187 ( .A(n22615), .ZN(n22606) );
  NOR2_X1 U24188 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n22606), .ZN(
        n22832) );
  NAND3_X1 U24189 ( .A1(n22604), .A2(n22593), .A3(n22563), .ZN(n22587) );
  OAI21_X1 U24190 ( .B1(n22589), .B2(n22588), .A(n22587), .ZN(n22831) );
  AOI22_X1 U24191 ( .A1(n22608), .A2(n22832), .B1(n22609), .B2(n22831), .ZN(
        n22600) );
  AOI21_X1 U24192 ( .B1(n22591), .B2(n22848), .A(n22590), .ZN(n22592) );
  AOI21_X1 U24193 ( .B1(n22593), .B2(n22604), .A(n22592), .ZN(n22594) );
  NOR2_X1 U24194 ( .A1(n22594), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n22597) );
  AOI22_X1 U24195 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n22834), .B2(n22598), .ZN(n22599) );
  OAI211_X1 U24196 ( .C1(n22601), .C2(n22848), .A(n22600), .B(n22599), .ZN(
        P1_U3145) );
  INV_X1 U24197 ( .A(n22602), .ZN(n22840) );
  AOI21_X1 U24198 ( .B1(n22604), .B2(n22603), .A(n22840), .ZN(n22610) );
  OAI22_X1 U24199 ( .A1(n22610), .A2(n22607), .B1(n22606), .B2(n22605), .ZN(
        n22842) );
  AOI22_X1 U24200 ( .A1(n22842), .A2(n22609), .B1(n22840), .B2(n22608), .ZN(
        n22618) );
  OAI21_X1 U24201 ( .B1(n22612), .B2(n22611), .A(n22610), .ZN(n22614) );
  OAI211_X1 U24202 ( .C1(n22563), .C2(n22615), .A(n22614), .B(n22613), .ZN(
        n22845) );
  AOI22_X1 U24203 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n22844), .B2(n22616), .ZN(n22617) );
  OAI211_X1 U24204 ( .C1(n22619), .C2(n22848), .A(n22618), .B(n22617), .ZN(
        P1_U3153) );
  AOI22_X1 U24205 ( .A1(n22844), .A2(n22637), .B1(n22782), .B2(n11263), .ZN(
        n22621) );
  AOI22_X1 U24206 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n22783), .B2(n22643), .ZN(n22620) );
  OAI211_X1 U24207 ( .C1(n22787), .C2(n22636), .A(n22621), .B(n22620), .ZN(
        P1_U3034) );
  AOI22_X1 U24208 ( .A1(n22796), .A2(n22643), .B1(n11263), .B2(n22788), .ZN(
        n22623) );
  AOI22_X1 U24209 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n22789), .B2(n22637), .ZN(n22622) );
  OAI211_X1 U24210 ( .C1(n22793), .C2(n22636), .A(n22623), .B(n22622), .ZN(
        P1_U3050) );
  AOI22_X1 U24211 ( .A1(n22795), .A2(n22643), .B1(n22794), .B2(n11263), .ZN(
        n22625) );
  AOI22_X1 U24212 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n22797), .B1(
        n22796), .B2(n22637), .ZN(n22624) );
  OAI211_X1 U24213 ( .C1(n22800), .C2(n22636), .A(n22625), .B(n22624), .ZN(
        P1_U3058) );
  AOI22_X1 U24214 ( .A1(n22803), .A2(n22643), .B1(n22801), .B2(n11263), .ZN(
        n22627) );
  AOI22_X1 U24215 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n22802), .B2(n22637), .ZN(n22626) );
  OAI211_X1 U24216 ( .C1(n22807), .C2(n22636), .A(n22627), .B(n22626), .ZN(
        P1_U3082) );
  AOI22_X1 U24217 ( .A1(n22816), .A2(n22643), .B1(n22808), .B2(n11263), .ZN(
        n22629) );
  AOI22_X1 U24218 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n22809), .B2(n22637), .ZN(n22628) );
  OAI211_X1 U24219 ( .C1(n22813), .C2(n22636), .A(n22629), .B(n22628), .ZN(
        P1_U3114) );
  AOI22_X1 U24220 ( .A1(n22815), .A2(n22642), .B1(n11263), .B2(n22814), .ZN(
        n22631) );
  AOI22_X1 U24221 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22637), .ZN(n22630) );
  OAI211_X1 U24222 ( .C1(n22640), .C2(n22820), .A(n22631), .B(n22630), .ZN(
        P1_U3122) );
  OAI22_X1 U24223 ( .A1(n22823), .A2(n22640), .B1(n22822), .B2(n22632), .ZN(
        n22633) );
  INV_X1 U24224 ( .A(n22633), .ZN(n22635) );
  AOI22_X1 U24225 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22637), .ZN(n22634) );
  OAI211_X1 U24226 ( .C1(n22830), .C2(n22636), .A(n22635), .B(n22634), .ZN(
        P1_U3130) );
  AOI22_X1 U24227 ( .A1(n11263), .A2(n22832), .B1(n22642), .B2(n22831), .ZN(
        n22639) );
  AOI22_X1 U24228 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n22834), .B2(n22637), .ZN(n22638) );
  OAI211_X1 U24229 ( .C1(n22640), .C2(n22848), .A(n22639), .B(n22638), .ZN(
        P1_U3146) );
  AOI22_X1 U24230 ( .A1(n22842), .A2(n22642), .B1(n22840), .B2(n11263), .ZN(
        n22645) );
  AOI22_X1 U24231 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n22844), .B2(n22643), .ZN(n22644) );
  OAI211_X1 U24232 ( .C1(n22646), .C2(n22848), .A(n22645), .B(n22644), .ZN(
        P1_U3154) );
  AOI22_X1 U24233 ( .A1(n22844), .A2(n22664), .B1(n22668), .B2(n22782), .ZN(
        n22648) );
  AOI22_X1 U24234 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n22783), .B2(n22670), .ZN(n22647) );
  OAI211_X1 U24235 ( .C1(n22787), .C2(n22663), .A(n22648), .B(n22647), .ZN(
        P1_U3035) );
  AOI22_X1 U24236 ( .A1(n22796), .A2(n22670), .B1(n22668), .B2(n22788), .ZN(
        n22650) );
  AOI22_X1 U24237 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n22664), .B2(n22789), .ZN(n22649) );
  OAI211_X1 U24238 ( .C1(n22793), .C2(n22663), .A(n22650), .B(n22649), .ZN(
        P1_U3051) );
  AOI22_X1 U24239 ( .A1(n22796), .A2(n22664), .B1(n22668), .B2(n22794), .ZN(
        n22652) );
  AOI22_X1 U24240 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n22797), .B1(
        n22795), .B2(n22670), .ZN(n22651) );
  OAI211_X1 U24241 ( .C1(n22800), .C2(n22663), .A(n22652), .B(n22651), .ZN(
        P1_U3059) );
  AOI22_X1 U24242 ( .A1(n22803), .A2(n22670), .B1(n22801), .B2(n22668), .ZN(
        n22654) );
  AOI22_X1 U24243 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n22664), .B2(n22802), .ZN(n22653) );
  OAI211_X1 U24244 ( .C1(n22807), .C2(n22663), .A(n22654), .B(n22653), .ZN(
        P1_U3083) );
  AOI22_X1 U24245 ( .A1(n22816), .A2(n22670), .B1(n22808), .B2(n22668), .ZN(
        n22656) );
  AOI22_X1 U24246 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n22664), .B2(n22809), .ZN(n22655) );
  OAI211_X1 U24247 ( .C1(n22813), .C2(n22663), .A(n22656), .B(n22655), .ZN(
        P1_U3115) );
  AOI22_X1 U24248 ( .A1(n22815), .A2(n22669), .B1(n22668), .B2(n22814), .ZN(
        n22658) );
  AOI22_X1 U24249 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22664), .ZN(n22657) );
  OAI211_X1 U24250 ( .C1(n22667), .C2(n22820), .A(n22658), .B(n22657), .ZN(
        P1_U3123) );
  OAI22_X1 U24251 ( .A1(n22823), .A2(n22667), .B1(n22822), .B2(n22659), .ZN(
        n22660) );
  INV_X1 U24252 ( .A(n22660), .ZN(n22662) );
  AOI22_X1 U24253 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22664), .ZN(n22661) );
  OAI211_X1 U24254 ( .C1(n22830), .C2(n22663), .A(n22662), .B(n22661), .ZN(
        P1_U3131) );
  AOI22_X1 U24255 ( .A1(n22668), .A2(n22832), .B1(n22669), .B2(n22831), .ZN(
        n22666) );
  AOI22_X1 U24256 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n22834), .B2(n22664), .ZN(n22665) );
  OAI211_X1 U24257 ( .C1(n22667), .C2(n22848), .A(n22666), .B(n22665), .ZN(
        P1_U3147) );
  AOI22_X1 U24258 ( .A1(n22842), .A2(n22669), .B1(n22840), .B2(n22668), .ZN(
        n22672) );
  AOI22_X1 U24259 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n22844), .B2(n22670), .ZN(n22671) );
  OAI211_X1 U24260 ( .C1(n22673), .C2(n22848), .A(n22672), .B(n22671), .ZN(
        P1_U3155) );
  AOI22_X1 U24261 ( .A1(n22844), .A2(n22691), .B1(n22782), .B2(n22695), .ZN(
        n22675) );
  AOI22_X1 U24262 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n22783), .B2(n22697), .ZN(n22674) );
  OAI211_X1 U24263 ( .C1(n22787), .C2(n22690), .A(n22675), .B(n22674), .ZN(
        P1_U3036) );
  AOI22_X1 U24264 ( .A1(n22796), .A2(n22697), .B1(n22695), .B2(n22788), .ZN(
        n22677) );
  AOI22_X1 U24265 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n22789), .B2(n22691), .ZN(n22676) );
  OAI211_X1 U24266 ( .C1(n22793), .C2(n22690), .A(n22677), .B(n22676), .ZN(
        P1_U3052) );
  AOI22_X1 U24267 ( .A1(n22796), .A2(n22691), .B1(n22794), .B2(n22695), .ZN(
        n22679) );
  AOI22_X1 U24268 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22797), .B1(
        n22795), .B2(n22697), .ZN(n22678) );
  OAI211_X1 U24269 ( .C1(n22800), .C2(n22690), .A(n22679), .B(n22678), .ZN(
        P1_U3060) );
  AOI22_X1 U24270 ( .A1(n22802), .A2(n22691), .B1(n22801), .B2(n22695), .ZN(
        n22681) );
  AOI22_X1 U24271 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n22803), .B2(n22697), .ZN(n22680) );
  OAI211_X1 U24272 ( .C1(n22807), .C2(n22690), .A(n22681), .B(n22680), .ZN(
        P1_U3084) );
  AOI22_X1 U24273 ( .A1(n22816), .A2(n22697), .B1(n22808), .B2(n22695), .ZN(
        n22683) );
  AOI22_X1 U24274 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n22809), .B2(n22691), .ZN(n22682) );
  OAI211_X1 U24275 ( .C1(n22813), .C2(n22690), .A(n22683), .B(n22682), .ZN(
        P1_U3116) );
  AOI22_X1 U24276 ( .A1(n22815), .A2(n22696), .B1(n22695), .B2(n22814), .ZN(
        n22685) );
  AOI22_X1 U24277 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22691), .ZN(n22684) );
  OAI211_X1 U24278 ( .C1(n22694), .C2(n22820), .A(n22685), .B(n22684), .ZN(
        P1_U3124) );
  OAI22_X1 U24279 ( .A1(n22823), .A2(n22694), .B1(n22822), .B2(n22686), .ZN(
        n22687) );
  INV_X1 U24280 ( .A(n22687), .ZN(n22689) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22691), .ZN(n22688) );
  OAI211_X1 U24282 ( .C1(n22830), .C2(n22690), .A(n22689), .B(n22688), .ZN(
        P1_U3132) );
  AOI22_X1 U24283 ( .A1(n22695), .A2(n22832), .B1(n22696), .B2(n22831), .ZN(
        n22693) );
  AOI22_X1 U24284 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n22834), .B2(n22691), .ZN(n22692) );
  OAI211_X1 U24285 ( .C1(n22694), .C2(n22848), .A(n22693), .B(n22692), .ZN(
        P1_U3148) );
  AOI22_X1 U24286 ( .A1(n22842), .A2(n22696), .B1(n22840), .B2(n22695), .ZN(
        n22699) );
  AOI22_X1 U24287 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n22844), .B2(n22697), .ZN(n22698) );
  OAI211_X1 U24288 ( .C1(n22700), .C2(n22848), .A(n22699), .B(n22698), .ZN(
        P1_U3156) );
  AOI22_X1 U24289 ( .A1(n22844), .A2(n22718), .B1(n22782), .B2(n22722), .ZN(
        n22702) );
  AOI22_X1 U24290 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n22783), .B2(n22724), .ZN(n22701) );
  OAI211_X1 U24291 ( .C1(n22787), .C2(n22717), .A(n22702), .B(n22701), .ZN(
        P1_U3037) );
  AOI22_X1 U24292 ( .A1(n22796), .A2(n22724), .B1(n22722), .B2(n22788), .ZN(
        n22704) );
  AOI22_X1 U24293 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n22789), .B2(n22718), .ZN(n22703) );
  OAI211_X1 U24294 ( .C1(n22793), .C2(n22717), .A(n22704), .B(n22703), .ZN(
        P1_U3053) );
  AOI22_X1 U24295 ( .A1(n22796), .A2(n22718), .B1(n22794), .B2(n22722), .ZN(
        n22706) );
  AOI22_X1 U24296 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22797), .B1(
        n22795), .B2(n22724), .ZN(n22705) );
  OAI211_X1 U24297 ( .C1(n22800), .C2(n22717), .A(n22706), .B(n22705), .ZN(
        P1_U3061) );
  AOI22_X1 U24298 ( .A1(n22803), .A2(n22724), .B1(n22801), .B2(n22722), .ZN(
        n22708) );
  AOI22_X1 U24299 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n22802), .B2(n22718), .ZN(n22707) );
  OAI211_X1 U24300 ( .C1(n22807), .C2(n22717), .A(n22708), .B(n22707), .ZN(
        P1_U3085) );
  AOI22_X1 U24301 ( .A1(n22816), .A2(n22724), .B1(n22808), .B2(n22722), .ZN(
        n22710) );
  AOI22_X1 U24302 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n22809), .B2(n22718), .ZN(n22709) );
  OAI211_X1 U24303 ( .C1(n22813), .C2(n22717), .A(n22710), .B(n22709), .ZN(
        P1_U3117) );
  AOI22_X1 U24304 ( .A1(n22815), .A2(n22723), .B1(n22722), .B2(n22814), .ZN(
        n22712) );
  AOI22_X1 U24305 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22718), .ZN(n22711) );
  OAI211_X1 U24306 ( .C1(n22721), .C2(n22820), .A(n22712), .B(n22711), .ZN(
        P1_U3125) );
  OAI22_X1 U24307 ( .A1(n22823), .A2(n22721), .B1(n22822), .B2(n22713), .ZN(
        n22714) );
  INV_X1 U24308 ( .A(n22714), .ZN(n22716) );
  AOI22_X1 U24309 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22718), .ZN(n22715) );
  OAI211_X1 U24310 ( .C1(n22830), .C2(n22717), .A(n22716), .B(n22715), .ZN(
        P1_U3133) );
  AOI22_X1 U24311 ( .A1(n22722), .A2(n22832), .B1(n22723), .B2(n22831), .ZN(
        n22720) );
  AOI22_X1 U24312 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n22834), .B2(n22718), .ZN(n22719) );
  OAI211_X1 U24313 ( .C1(n22721), .C2(n22848), .A(n22720), .B(n22719), .ZN(
        P1_U3149) );
  AOI22_X1 U24314 ( .A1(n22842), .A2(n22723), .B1(n22840), .B2(n22722), .ZN(
        n22726) );
  AOI22_X1 U24315 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22844), .B2(n22724), .ZN(n22725) );
  OAI211_X1 U24316 ( .C1(n22727), .C2(n22848), .A(n22726), .B(n22725), .ZN(
        P1_U3157) );
  AOI22_X1 U24317 ( .A1(n22844), .A2(n22745), .B1(n22782), .B2(n11122), .ZN(
        n22729) );
  AOI22_X1 U24318 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n22783), .B2(n22751), .ZN(n22728) );
  OAI211_X1 U24319 ( .C1(n22787), .C2(n22744), .A(n22729), .B(n22728), .ZN(
        P1_U3038) );
  AOI22_X1 U24320 ( .A1(n22796), .A2(n22751), .B1(n11122), .B2(n22788), .ZN(
        n22731) );
  AOI22_X1 U24321 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n22789), .B2(n22745), .ZN(n22730) );
  OAI211_X1 U24322 ( .C1(n22793), .C2(n22744), .A(n22731), .B(n22730), .ZN(
        P1_U3054) );
  AOI22_X1 U24323 ( .A1(n22796), .A2(n22745), .B1(n22794), .B2(n11122), .ZN(
        n22733) );
  AOI22_X1 U24324 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n22797), .B1(
        n22795), .B2(n22751), .ZN(n22732) );
  OAI211_X1 U24325 ( .C1(n22800), .C2(n22744), .A(n22733), .B(n22732), .ZN(
        P1_U3062) );
  AOI22_X1 U24326 ( .A1(n22802), .A2(n22745), .B1(n22801), .B2(n11122), .ZN(
        n22735) );
  AOI22_X1 U24327 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n22803), .B2(n22751), .ZN(n22734) );
  OAI211_X1 U24328 ( .C1(n22807), .C2(n22744), .A(n22735), .B(n22734), .ZN(
        P1_U3086) );
  AOI22_X1 U24329 ( .A1(n22816), .A2(n22751), .B1(n22808), .B2(n11122), .ZN(
        n22737) );
  AOI22_X1 U24330 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n22809), .B2(n22745), .ZN(n22736) );
  OAI211_X1 U24331 ( .C1(n22813), .C2(n22744), .A(n22737), .B(n22736), .ZN(
        P1_U3118) );
  AOI22_X1 U24332 ( .A1(n22815), .A2(n22750), .B1(n11122), .B2(n22814), .ZN(
        n22739) );
  AOI22_X1 U24333 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22745), .ZN(n22738) );
  OAI211_X1 U24334 ( .C1(n22748), .C2(n22820), .A(n22739), .B(n22738), .ZN(
        P1_U3126) );
  OAI22_X1 U24335 ( .A1(n22823), .A2(n22748), .B1(n22822), .B2(n22740), .ZN(
        n22741) );
  INV_X1 U24336 ( .A(n22741), .ZN(n22743) );
  AOI22_X1 U24337 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22745), .ZN(n22742) );
  OAI211_X1 U24338 ( .C1(n22830), .C2(n22744), .A(n22743), .B(n22742), .ZN(
        P1_U3134) );
  AOI22_X1 U24339 ( .A1(n11122), .A2(n22832), .B1(n22750), .B2(n22831), .ZN(
        n22747) );
  AOI22_X1 U24340 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n22834), .B2(n22745), .ZN(n22746) );
  OAI211_X1 U24341 ( .C1(n22748), .C2(n22848), .A(n22747), .B(n22746), .ZN(
        P1_U3150) );
  AOI22_X1 U24342 ( .A1(n22842), .A2(n22750), .B1(n22840), .B2(n11122), .ZN(
        n22753) );
  AOI22_X1 U24343 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n22844), .B2(n22751), .ZN(n22752) );
  OAI211_X1 U24344 ( .C1(n22754), .C2(n22848), .A(n22753), .B(n22752), .ZN(
        P1_U3158) );
  AOI22_X1 U24345 ( .A1(n22844), .A2(n22772), .B1(n22782), .B2(n11123), .ZN(
        n22756) );
  AOI22_X1 U24346 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n22783), .B2(n22778), .ZN(n22755) );
  OAI211_X1 U24347 ( .C1(n22787), .C2(n22771), .A(n22756), .B(n22755), .ZN(
        P1_U3039) );
  AOI22_X1 U24348 ( .A1(n22796), .A2(n22778), .B1(n11123), .B2(n22788), .ZN(
        n22758) );
  AOI22_X1 U24349 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n22789), .B2(n22772), .ZN(n22757) );
  OAI211_X1 U24350 ( .C1(n22793), .C2(n22771), .A(n22758), .B(n22757), .ZN(
        P1_U3055) );
  AOI22_X1 U24351 ( .A1(n22796), .A2(n22772), .B1(n22794), .B2(n11123), .ZN(
        n22760) );
  AOI22_X1 U24352 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n22797), .B1(
        n22795), .B2(n22778), .ZN(n22759) );
  OAI211_X1 U24353 ( .C1(n22800), .C2(n22771), .A(n22760), .B(n22759), .ZN(
        P1_U3063) );
  AOI22_X1 U24354 ( .A1(n22802), .A2(n22772), .B1(n22801), .B2(n11123), .ZN(
        n22762) );
  AOI22_X1 U24355 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n22803), .B2(n22778), .ZN(n22761) );
  OAI211_X1 U24356 ( .C1(n22807), .C2(n22771), .A(n22762), .B(n22761), .ZN(
        P1_U3087) );
  AOI22_X1 U24357 ( .A1(n22816), .A2(n22778), .B1(n22808), .B2(n11123), .ZN(
        n22764) );
  AOI22_X1 U24358 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n22809), .B2(n22772), .ZN(n22763) );
  OAI211_X1 U24359 ( .C1(n22813), .C2(n22771), .A(n22764), .B(n22763), .ZN(
        P1_U3119) );
  AOI22_X1 U24360 ( .A1(n22815), .A2(n22777), .B1(n11123), .B2(n22814), .ZN(
        n22766) );
  AOI22_X1 U24361 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22772), .ZN(n22765) );
  OAI211_X1 U24362 ( .C1(n22775), .C2(n22820), .A(n22766), .B(n22765), .ZN(
        P1_U3127) );
  OAI22_X1 U24363 ( .A1(n22823), .A2(n22775), .B1(n22822), .B2(n22767), .ZN(
        n22768) );
  INV_X1 U24364 ( .A(n22768), .ZN(n22770) );
  AOI22_X1 U24365 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22772), .ZN(n22769) );
  OAI211_X1 U24366 ( .C1(n22830), .C2(n22771), .A(n22770), .B(n22769), .ZN(
        P1_U3135) );
  AOI22_X1 U24367 ( .A1(n11123), .A2(n22832), .B1(n22777), .B2(n22831), .ZN(
        n22774) );
  AOI22_X1 U24368 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n22834), .B2(n22772), .ZN(n22773) );
  OAI211_X1 U24369 ( .C1(n22775), .C2(n22848), .A(n22774), .B(n22773), .ZN(
        P1_U3151) );
  AOI22_X1 U24370 ( .A1(n22842), .A2(n22777), .B1(n22840), .B2(n11123), .ZN(
        n22780) );
  AOI22_X1 U24371 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n22844), .B2(n22778), .ZN(n22779) );
  OAI211_X1 U24372 ( .C1(n22781), .C2(n22848), .A(n22780), .B(n22779), .ZN(
        P1_U3159) );
  AOI22_X1 U24373 ( .A1(n22844), .A2(n22833), .B1(n22782), .B2(n22839), .ZN(
        n22786) );
  AOI22_X1 U24374 ( .A1(n22784), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n22783), .B2(n22843), .ZN(n22785) );
  OAI211_X1 U24375 ( .C1(n22787), .C2(n22829), .A(n22786), .B(n22785), .ZN(
        P1_U3040) );
  AOI22_X1 U24376 ( .A1(n22796), .A2(n22843), .B1(n22839), .B2(n22788), .ZN(
        n22792) );
  AOI22_X1 U24377 ( .A1(n22790), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n22789), .B2(n22833), .ZN(n22791) );
  OAI211_X1 U24378 ( .C1(n22793), .C2(n22829), .A(n22792), .B(n22791), .ZN(
        P1_U3056) );
  AOI22_X1 U24379 ( .A1(n22795), .A2(n22843), .B1(n22794), .B2(n22839), .ZN(
        n22799) );
  AOI22_X1 U24380 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22797), .B1(
        n22796), .B2(n22833), .ZN(n22798) );
  OAI211_X1 U24381 ( .C1(n22800), .C2(n22829), .A(n22799), .B(n22798), .ZN(
        P1_U3064) );
  AOI22_X1 U24382 ( .A1(n22802), .A2(n22833), .B1(n22801), .B2(n22839), .ZN(
        n22806) );
  AOI22_X1 U24383 ( .A1(n22804), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n22803), .B2(n22843), .ZN(n22805) );
  OAI211_X1 U24384 ( .C1(n22807), .C2(n22829), .A(n22806), .B(n22805), .ZN(
        P1_U3088) );
  AOI22_X1 U24385 ( .A1(n22816), .A2(n22843), .B1(n22808), .B2(n22839), .ZN(
        n22812) );
  AOI22_X1 U24386 ( .A1(n22810), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n22809), .B2(n22833), .ZN(n22811) );
  OAI211_X1 U24387 ( .C1(n22813), .C2(n22829), .A(n22812), .B(n22811), .ZN(
        P1_U3120) );
  AOI22_X1 U24388 ( .A1(n22815), .A2(n22841), .B1(n22839), .B2(n22814), .ZN(
        n22819) );
  AOI22_X1 U24389 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n22817), .B1(
        n22816), .B2(n22833), .ZN(n22818) );
  OAI211_X1 U24390 ( .C1(n22838), .C2(n22820), .A(n22819), .B(n22818), .ZN(
        P1_U3128) );
  OAI22_X1 U24391 ( .A1(n22823), .A2(n22838), .B1(n22822), .B2(n22821), .ZN(
        n22824) );
  INV_X1 U24392 ( .A(n22824), .ZN(n22828) );
  AOI22_X1 U24393 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n22826), .B1(
        n22825), .B2(n22833), .ZN(n22827) );
  OAI211_X1 U24394 ( .C1(n22830), .C2(n22829), .A(n22828), .B(n22827), .ZN(
        P1_U3136) );
  AOI22_X1 U24395 ( .A1(n22839), .A2(n22832), .B1(n22841), .B2(n22831), .ZN(
        n22837) );
  AOI22_X1 U24396 ( .A1(n22835), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n22834), .B2(n22833), .ZN(n22836) );
  OAI211_X1 U24397 ( .C1(n22838), .C2(n22848), .A(n22837), .B(n22836), .ZN(
        P1_U3152) );
  AOI22_X1 U24398 ( .A1(n22842), .A2(n22841), .B1(n22840), .B2(n22839), .ZN(
        n22847) );
  AOI22_X1 U24399 ( .A1(n22845), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n22844), .B2(n22843), .ZN(n22846) );
  OAI211_X1 U24400 ( .C1(n22849), .C2(n22848), .A(n22847), .B(n22846), .ZN(
        P1_U3160) );
  AOI22_X1 U24401 ( .A1(n22853), .A2(n22852), .B1(n22851), .B2(n22850), .ZN(
        P1_U3486) );
  BUF_X1 U11239 ( .A(n15783), .Z(n11143) );
  CLKBUF_X1 U11259 ( .A(n13107), .Z(n13763) );
  CLKBUF_X1 U11262 ( .A(n13102), .Z(n11135) );
  CLKBUF_X1 U11263 ( .A(n12152), .Z(n12839) );
  NAND2_X1 U11270 ( .A1(n15263), .A2(n12406), .ZN(n12410) );
  CLKBUF_X1 U11274 ( .A(n11146), .Z(n14065) );
  NOR2_X2 U11283 ( .A1(n16671), .A2(n14022), .ZN(n16659) );
  CLKBUF_X1 U11292 ( .A(n12005), .Z(n20125) );
  CLKBUF_X1 U11307 ( .A(n16562), .Z(n11155) );
  CLKBUF_X1 U12024 ( .A(n17936), .Z(n17947) );
  CLKBUF_X1 U12467 ( .A(n15379), .Z(n19244) );
  CLKBUF_X1 U12488 ( .A(n18979), .Z(n18985) );
  XOR2_X1 U12589 ( .A(n14259), .B(n20607), .Z(n22065) );
  OR2_X1 U12590 ( .A1(n20294), .A2(n20293), .ZN(n22854) );
  CLKBUF_X1 U12885 ( .A(n18977), .Z(n21871) );
endmodule

