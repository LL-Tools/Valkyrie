

module b20_C_SARLock_k_128_6 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384;

  INV_X4 U4946 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X2 U4947 ( .A(n6959), .ZN(n6788) );
  CLKBUF_X1 U4948 ( .A(n5820), .Z(n4450) );
  AOI22_X1 U4949 ( .A1(n5820), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5819), .B2(
        n7099), .ZN(n5768) );
  OR2_X1 U4950 ( .A1(n5014), .A2(n5013), .ZN(n5016) );
  BUF_X2 U4952 ( .A(n6099), .Z(n6118) );
  NOR2_X1 U4953 ( .A1(n4544), .A2(n4807), .ZN(n4543) );
  CLKBUF_X2 U4954 ( .A(n6101), .Z(n4441) );
  CLKBUF_X1 U4955 ( .A(n8983), .Z(n4438) );
  NOR2_X1 U4956 ( .A1(n6604), .A2(n6603), .ZN(n8983) );
  AOI22_X1 U4957 ( .A1(n5981), .A2(keyinput1), .B1(n8211), .B2(keyinput89), 
        .ZN(n9514) );
  AOI22_X1 U4958 ( .A1(n9379), .A2(keyinput121), .B1(P1_ADDR_REG_14__SCAN_IN), 
        .B2(n9378), .ZN(n9377) );
  OAI221_X1 U4960 ( .B1(n5981), .B2(keyinput1), .C1(n8211), .C2(keyinput89), 
        .A(n9514), .ZN(n9515) );
  OAI221_X1 U4961 ( .B1(n9379), .B2(keyinput121), .C1(n9378), .C2(
        P1_ADDR_REG_14__SCAN_IN), .A(n9377), .ZN(n9380) );
  NOR2_X1 U4962 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5701) );
  INV_X2 U4963 ( .A(n6425), .ZN(n6579) );
  INV_X4 U4964 ( .A(n5065), .ZN(n5902) );
  NAND2_X1 U4965 ( .A1(n6536), .A2(n8865), .ZN(n8867) );
  INV_X2 U4966 ( .A(n6507), .ZN(n6581) );
  CLKBUF_X2 U4967 ( .A(n6101), .Z(n4442) );
  AOI21_X1 U4968 ( .B1(n9640), .B2(n10083), .A(n9639), .ZN(n4564) );
  AND2_X1 U4969 ( .A1(n5097), .A2(n4466), .ZN(n7608) );
  BUF_X1 U4970 ( .A(n5068), .Z(n6962) );
  NAND4_X1 U4971 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n7272)
         );
  OAI21_X1 U4972 ( .B1(n9538), .B2(n9158), .A(n9157), .ZN(n9225) );
  NAND2_X1 U4973 ( .A1(n5857), .A2(n8238), .ZN(n6983) );
  NAND2_X1 U4974 ( .A1(n4804), .A2(n4542), .ZN(n5122) );
  AND2_X1 U4975 ( .A1(n6927), .A2(n6926), .ZN(n8403) );
  NAND4_X2 U4976 ( .A1(n5565), .A2(n5564), .A3(n5563), .A4(n5562), .ZN(n8422)
         );
  INV_X1 U4977 ( .A(n7622), .ZN(n4444) );
  INV_X1 U4978 ( .A(n8535), .ZN(n8526) );
  OR2_X1 U4979 ( .A1(n9638), .A2(n4563), .ZN(n9681) );
  XNOR2_X1 U4980 ( .A(n5869), .B(n5868), .ZN(n5876) );
  AND2_X1 U4981 ( .A1(n5910), .A2(n9701), .ZN(n4439) );
  XNOR2_X1 U4982 ( .A(n5716), .B(n5715), .ZN(n5857) );
  CLKBUF_X2 U4983 ( .A(n6386), .Z(n4440) );
  NAND4_X1 U4984 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n6386)
         );
  XNOR2_X2 U4985 ( .A(n5016), .B(n5015), .ZN(n8242) );
  NAND2_X2 U4986 ( .A1(n5768), .A2(n5767), .ZN(n10014) );
  NAND2_X2 U4987 ( .A1(n4959), .A2(n4961), .ZN(n9538) );
  XNOR2_X2 U4988 ( .A(n5012), .B(n5011), .ZN(n8847) );
  NAND2_X4 U4990 ( .A1(n6845), .A2(n6844), .ZN(n6851) );
  NOR2_X2 U4991 ( .A1(n9782), .A2(n6433), .ZN(n7774) );
  NOR2_X2 U4992 ( .A1(n9783), .A2(n9784), .ZN(n9782) );
  OR2_X2 U4993 ( .A1(n7937), .A2(n6376), .ZN(n7018) );
  INV_X2 U4994 ( .A(n6376), .ZN(n5880) );
  NAND2_X1 U4995 ( .A1(n8273), .A2(n5909), .ZN(n6101) );
  OAI222_X1 U4996 ( .A1(n7385), .A2(P2_U3151), .B1(n8851), .B2(n6976), .C1(
        n6975), .C2(n8848), .ZN(P2_U3291) );
  OAI222_X1 U4997 ( .A1(n8277), .A2(n6974), .B1(n8275), .B2(n6976), .C1(n8274), 
        .C2(n9820), .ZN(P1_U3351) );
  OR2_X1 U4998 ( .A1(n6976), .A2(n5780), .ZN(n5767) );
  AND2_X2 U4999 ( .A1(n6374), .A2(n6593), .ZN(n6377) );
  AOI21_X2 U5000 ( .B1(n8580), .B2(n5551), .A(n5550), .ZN(n8589) );
  OR2_X4 U5001 ( .A1(n5876), .A2(n5875), .ZN(n6379) );
  NAND2_X1 U5002 ( .A1(n4896), .A2(n4894), .ZN(n8886) );
  NAND2_X2 U5003 ( .A1(n8649), .A2(n8650), .ZN(n8665) );
  XNOR2_X1 U5004 ( .A(n5450), .B(n5445), .ZN(n7824) );
  CLKBUF_X2 U5005 ( .A(n6851), .Z(n6919) );
  BUF_X1 U5006 ( .A(n9999), .Z(n4447) );
  NAND2_X1 U5007 ( .A1(n6849), .A2(n6848), .ZN(n6676) );
  CLKBUF_X2 U5008 ( .A(n5073), .Z(n6621) );
  INV_X2 U5009 ( .A(n6425), .ZN(n6564) );
  CLKBUF_X3 U5010 ( .A(n5206), .Z(n6356) );
  INV_X2 U5011 ( .A(n5072), .ZN(n5557) );
  INV_X2 U5012 ( .A(n6102), .ZN(n6084) );
  CLKBUF_X2 U5013 ( .A(n5577), .Z(n7642) );
  NAND2_X1 U5014 ( .A1(n5065), .A2(n8274), .ZN(n8277) );
  CLKBUF_X2 U5015 ( .A(n8274), .Z(P1_U3086) );
  INV_X1 U5016 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4683) );
  XNOR2_X1 U5017 ( .A(n9169), .B(n9168), .ZN(n9631) );
  OR2_X1 U5018 ( .A1(n9189), .A2(n9188), .ZN(n9634) );
  NAND2_X1 U5019 ( .A1(n9193), .A2(n4480), .ZN(n9190) );
  AOI21_X1 U5020 ( .B1(n6831), .B2(n6830), .A(n6829), .ZN(n6833) );
  NOR2_X1 U5021 ( .A1(n9233), .A2(n9232), .ZN(n9231) );
  AND2_X1 U5022 ( .A1(n6523), .A2(n6522), .ZN(n8864) );
  XNOR2_X1 U5023 ( .A(n5906), .B(n5905), .ZN(n9698) );
  OR2_X1 U5024 ( .A1(n8735), .A2(n8589), .ZN(n6807) );
  OAI21_X1 U5025 ( .B1(n10173), .B2(n4799), .A(n4798), .ZN(n10191) );
  INV_X1 U5026 ( .A(n4872), .ZN(n4871) );
  NAND2_X1 U5027 ( .A1(n7876), .A2(n6867), .ZN(n8175) );
  NAND2_X1 U5028 ( .A1(n5739), .A2(n5738), .ZN(n9146) );
  NAND2_X1 U5029 ( .A1(n5380), .A2(n5379), .ZN(n8703) );
  OAI21_X1 U5030 ( .B1(n5424), .B2(n5423), .A(n5435), .ZN(n7820) );
  OAI21_X1 U5031 ( .B1(n7305), .B2(n4883), .A(n4881), .ZN(n6430) );
  OR2_X1 U5032 ( .A1(n5579), .A2(n8560), .ZN(n5562) );
  OR2_X1 U5033 ( .A1(n5374), .A2(n5373), .ZN(n4773) );
  AOI21_X1 U5034 ( .B1(n7231), .B2(n7232), .A(n6854), .ZN(n7260) );
  AND2_X1 U5035 ( .A1(n5526), .A2(n8396), .ZN(n5546) );
  NAND2_X1 U5036 ( .A1(n5805), .A2(n5804), .ZN(n7990) );
  NAND2_X1 U5037 ( .A1(n4551), .A2(n5301), .ZN(n5316) );
  INV_X1 U5038 ( .A(n10014), .ZN(n7357) );
  AND2_X1 U5039 ( .A1(n5427), .A2(n5426), .ZN(n5439) );
  AND2_X1 U5040 ( .A1(n5784), .A2(n5783), .ZN(n10031) );
  NAND4_X2 U5041 ( .A1(n5058), .A2(n5057), .A3(n5056), .A4(n5055), .ZN(n8438)
         );
  OAI21_X1 U5042 ( .B1(n5599), .B2(n8218), .A(n7040), .ZN(n7009) );
  AND3_X1 U5043 ( .A1(n5040), .A2(n5039), .A3(n5038), .ZN(n6848) );
  NAND2_X2 U5044 ( .A1(n6383), .A2(n6385), .ZN(n4904) );
  INV_X2 U5045 ( .A(n5082), .ZN(n6627) );
  NAND4_X1 U5046 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n9005)
         );
  NAND2_X2 U5047 ( .A1(n6380), .A2(n6379), .ZN(n6383) );
  XNOR2_X1 U5048 ( .A(n5404), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8535) );
  INV_X1 U5049 ( .A(n6385), .ZN(n6507) );
  NAND2_X1 U5050 ( .A1(n5594), .A2(n5592), .ZN(n8287) );
  CLKBUF_X1 U5051 ( .A(n5205), .Z(n5579) );
  AND2_X1 U5052 ( .A1(n7018), .A2(n6378), .ZN(n6380) );
  NAND2_X1 U5053 ( .A1(n5019), .A2(n5020), .ZN(n5205) );
  OAI211_X1 U5054 ( .C1(n6375), .C2(n7017), .A(n6379), .B(n9972), .ZN(n6385)
         );
  NAND2_X4 U5055 ( .A1(n6379), .A2(n6377), .ZN(n6425) );
  CLKBUF_X1 U5056 ( .A(n5576), .Z(n7138) );
  NAND2_X1 U5057 ( .A1(n5842), .A2(n5877), .ZN(n7937) );
  NAND2_X1 U5058 ( .A1(n5848), .A2(n5847), .ZN(n6593) );
  NAND2_X1 U5059 ( .A1(n5736), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U5060 ( .A1(n5714), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U5061 ( .A1(n5721), .A2(n4463), .ZN(n8238) );
  OAI21_X1 U5062 ( .B1(n5867), .B2(n5866), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5869) );
  OR2_X1 U5063 ( .A1(n8223), .A2(n8229), .ZN(n5875) );
  XNOR2_X1 U5064 ( .A(n5844), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6374) );
  NAND2_X1 U5065 ( .A1(n5847), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  NAND2_X1 U5066 ( .A1(n4463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U5067 ( .A1(n5735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U5068 ( .A(n5103), .B(SI_3_), .ZN(n5101) );
  NAND2_X1 U5069 ( .A1(n5839), .A2(n4482), .ZN(n5847) );
  NAND2_X1 U5070 ( .A1(n5007), .A2(n5006), .ZN(n5570) );
  XNOR2_X1 U5071 ( .A(n5174), .B(SI_7_), .ZN(n5172) );
  INV_X2 U5072 ( .A(n8288), .ZN(n8851) );
  AND2_X1 U5073 ( .A1(n5202), .A2(n5201), .ZN(n5204) );
  INV_X2 U5074 ( .A(n9697), .ZN(n8275) );
  NOR2_X1 U5075 ( .A1(n5336), .A2(n5005), .ZN(n5006) );
  OR2_X1 U5076 ( .A1(n5138), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5157) );
  NOR2_X1 U5077 ( .A1(n4975), .A2(n5713), .ZN(n4974) );
  NOR2_X1 U5078 ( .A1(n4945), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4944) );
  AND3_X1 U5079 ( .A1(n4685), .A2(n4684), .A3(n4683), .ZN(n5002) );
  NAND2_X1 U5080 ( .A1(n7601), .A2(n4555), .ZN(n4801) );
  INV_X1 U5081 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4998) );
  NOR2_X2 U5082 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7142) );
  AND2_X1 U5083 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7601) );
  NOR2_X1 U5084 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7602) );
  OAI211_X1 U5085 ( .C1(n6910), .C2(n4908), .A(n4906), .B(1'b1), .ZN(n6914) );
  OAI21_X2 U5087 ( .B1(n8076), .B2(n4973), .A(n4459), .ZN(n9144) );
  OAI211_X1 U5088 ( .C1(n5780), .C2(n6970), .A(n5757), .B(n4989), .ZN(n9999)
         );
  XNOR2_X2 U5089 ( .A(n8563), .B(n8422), .ZN(n8264) );
  NOR3_X4 U5090 ( .A1(n8200), .A2(n4681), .A3(n9664), .ZN(n9583) );
  OR2_X4 U5091 ( .A1(n8146), .A2(n8197), .ZN(n8200) );
  INV_X1 U5092 ( .A(n4439), .ZN(n4448) );
  INV_X4 U5093 ( .A(n4439), .ZN(n4449) );
  INV_X2 U5094 ( .A(n7273), .ZN(n9992) );
  INV_X1 U5095 ( .A(n5754), .ZN(n5820) );
  CLKBUF_X1 U5096 ( .A(n5857), .Z(n4451) );
  NAND2_X4 U5097 ( .A1(n6983), .A2(n5065), .ZN(n5754) );
  NOR2_X2 U5098 ( .A1(n9213), .A2(n9640), .ZN(n4676) );
  INV_X1 U5099 ( .A(n4634), .ZN(n4633) );
  OAI21_X1 U5100 ( .B1(n4636), .B2(n6264), .A(n4635), .ZN(n4634) );
  OR2_X1 U5101 ( .A1(n6269), .A2(n6266), .ZN(n4635) );
  INV_X1 U5102 ( .A(n7272), .ZN(n7066) );
  NAND2_X1 U5103 ( .A1(n5299), .A2(n5298), .ZN(n4551) );
  INV_X1 U5104 ( .A(n5297), .ZN(n5298) );
  NAND2_X1 U5105 ( .A1(n4731), .A2(n6820), .ZN(n4730) );
  INV_X1 U5106 ( .A(n5371), .ZN(n4697) );
  NOR2_X1 U5107 ( .A1(n4621), .A2(n6246), .ZN(n4618) );
  INV_X1 U5108 ( .A(n4851), .ZN(n4849) );
  OR2_X1 U5109 ( .A1(n5215), .A2(n5214), .ZN(n5217) );
  AND2_X1 U5110 ( .A1(n7863), .A2(n5213), .ZN(n5214) );
  AND2_X1 U5111 ( .A1(n4556), .A2(n9925), .ZN(n6277) );
  NAND2_X1 U5112 ( .A1(n4557), .A2(n7362), .ZN(n4556) );
  INV_X1 U5113 ( .A(n8847), .ZN(n5019) );
  INV_X1 U5114 ( .A(n8242), .ZN(n5020) );
  INV_X1 U5115 ( .A(n10157), .ZN(n4579) );
  NOR2_X1 U5116 ( .A1(n10191), .A2(n8470), .ZN(n8471) );
  NOR2_X1 U5117 ( .A1(n10182), .A2(n8469), .ZN(n8470) );
  NOR2_X1 U5118 ( .A1(n10223), .A2(n8474), .ZN(n8475) );
  AND2_X1 U5119 ( .A1(n4720), .A2(n4719), .ZN(n4718) );
  NAND2_X1 U5120 ( .A1(n8803), .A2(n8598), .ZN(n4719) );
  OR2_X1 U5121 ( .A1(n5532), .A2(n4721), .ZN(n4720) );
  NAND2_X1 U5122 ( .A1(n5517), .A2(n5516), .ZN(n4721) );
  INV_X1 U5123 ( .A(n5516), .ZN(n4724) );
  AND2_X1 U5124 ( .A1(n5654), .A2(n8424), .ZN(n6787) );
  AND2_X1 U5125 ( .A1(n8665), .A2(n8652), .ZN(n4687) );
  OR2_X1 U5126 ( .A1(n5444), .A2(n8636), .ZN(n6780) );
  NAND2_X1 U5127 ( .A1(n4708), .A2(n7931), .ZN(n4707) );
  INV_X1 U5128 ( .A(n10301), .ZN(n4708) );
  AND2_X1 U5129 ( .A1(n5008), .A2(n4598), .ZN(n4597) );
  INV_X1 U5130 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4598) );
  OR2_X1 U5131 ( .A1(n9763), .A2(n8071), .ZN(n6307) );
  INV_X1 U5132 ( .A(n4760), .ZN(n4759) );
  OAI21_X1 U5133 ( .B1(n4762), .B2(n4761), .A(n5279), .ZN(n4760) );
  NOR2_X1 U5134 ( .A1(n5264), .A2(n4763), .ZN(n4762) );
  INV_X1 U5135 ( .A(n5243), .ZN(n4763) );
  XNOR2_X1 U5136 ( .A(n5241), .B(SI_10_), .ZN(n5240) );
  NAND2_X1 U5137 ( .A1(n4757), .A2(n4467), .ZN(n4752) );
  NAND2_X1 U5138 ( .A1(n5181), .A2(n5180), .ZN(n5196) );
  INV_X1 U5139 ( .A(n7787), .ZN(n4939) );
  INV_X1 U5140 ( .A(n7766), .ZN(n4940) );
  NAND2_X1 U5141 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  INV_X1 U5142 ( .A(n6880), .ZN(n4943) );
  NAND2_X1 U5143 ( .A1(n8526), .A2(n7823), .ZN(n6844) );
  NOR2_X1 U5144 ( .A1(n8730), .A2(n6626), .ZN(n6832) );
  INV_X1 U5145 ( .A(n5579), .ZN(n5551) );
  INV_X1 U5146 ( .A(n6356), .ZN(n5528) );
  INV_X1 U5147 ( .A(n5073), .ZN(n5137) );
  NAND2_X1 U5148 ( .A1(n5019), .A2(n8242), .ZN(n5073) );
  XNOR2_X1 U5149 ( .A(n8475), .B(n10233), .ZN(n10244) );
  INV_X1 U5150 ( .A(n4846), .ZN(n4842) );
  AND2_X1 U5151 ( .A1(n4845), .A2(n6746), .ZN(n4841) );
  AND2_X1 U5152 ( .A1(n5575), .A2(n5574), .ZN(n8635) );
  OR2_X1 U5153 ( .A1(n8641), .A2(n8622), .ZN(n6778) );
  OR2_X1 U5154 ( .A1(n8832), .A2(n8678), .ZN(n8649) );
  INV_X1 U5155 ( .A(n5107), .ZN(n6618) );
  INV_X1 U5156 ( .A(n8694), .ZN(n8720) );
  AOI21_X1 U5157 ( .B1(n7050), .B2(n7049), .A(n4982), .ZN(n7064) );
  NAND2_X1 U5158 ( .A1(n5880), .A2(n6593), .ZN(n7017) );
  XNOR2_X1 U5159 ( .A(n6384), .B(n6383), .ZN(n6392) );
  NAND2_X1 U5160 ( .A1(n4904), .A2(n7273), .ZN(n6381) );
  OAI21_X1 U5161 ( .B1(n6265), .B2(n4628), .A(n4626), .ZN(n6337) );
  AND2_X1 U5162 ( .A1(n4629), .A2(n4632), .ZN(n4628) );
  INV_X1 U5163 ( .A(n4627), .ZN(n4626) );
  AND4_X1 U5164 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n7565)
         );
  NAND2_X1 U5165 ( .A1(n8195), .A2(n4970), .ZN(n4973) );
  NAND2_X1 U5166 ( .A1(n8075), .A2(n8144), .ZN(n4970) );
  NAND2_X1 U5167 ( .A1(n7973), .A2(n7972), .ZN(n4965) );
  NAND2_X1 U5168 ( .A1(n6983), .A2(n5902), .ZN(n5780) );
  INV_X1 U5169 ( .A(n6983), .ZN(n5819) );
  OR2_X1 U5170 ( .A1(n7313), .A2(n7022), .ZN(n9612) );
  INV_X1 U5171 ( .A(n8921), .ZN(n9757) );
  NAND2_X1 U5172 ( .A1(n9693), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5851) );
  AOI21_X1 U5173 ( .B1(n4775), .B2(n4461), .A(n4764), .ZN(n5435) );
  NOR2_X1 U5174 ( .A1(n4765), .A2(n4771), .ZN(n4764) );
  XNOR2_X1 U5175 ( .A(n5167), .B(SI_6_), .ZN(n5165) );
  NAND2_X1 U5176 ( .A1(n5126), .A2(n5125), .ZN(n4554) );
  XNOR2_X1 U5177 ( .A(n5146), .B(SI_5_), .ZN(n5145) );
  OR2_X1 U5178 ( .A1(n5743), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5769) );
  NOR2_X1 U5179 ( .A1(n6853), .A2(n8438), .ZN(n6854) );
  AND2_X1 U5180 ( .A1(n6899), .A2(n6898), .ZN(n6900) );
  NOR2_X1 U5181 ( .A1(n6401), .A2(n6400), .ZN(n6402) );
  NAND2_X1 U5182 ( .A1(n8967), .A2(n6574), .ZN(n6613) );
  NOR2_X1 U5183 ( .A1(n6573), .A2(n6572), .ZN(n6574) );
  AND2_X1 U5184 ( .A1(n9215), .A2(n9164), .ZN(n9194) );
  NAND2_X1 U5185 ( .A1(n4565), .A2(n9200), .ZN(n9638) );
  OR2_X1 U5186 ( .A1(n9201), .A2(n9963), .ZN(n4565) );
  NAND2_X1 U5187 ( .A1(n4535), .A2(n6791), .ZN(n4534) );
  NAND2_X1 U5188 ( .A1(n9593), .A2(n7023), .ZN(n4648) );
  AOI21_X1 U5189 ( .B1(n6229), .B2(n6228), .A(n6227), .ZN(n6234) );
  MUX2_X1 U5190 ( .A(n6224), .B(n6223), .S(n7023), .Z(n6229) );
  NAND2_X1 U5191 ( .A1(n6810), .A2(n6809), .ZN(n4731) );
  NAND2_X1 U5192 ( .A1(n6806), .A2(n6805), .ZN(n4729) );
  OR2_X1 U5193 ( .A1(n4726), .A2(n6788), .ZN(n6803) );
  NOR2_X1 U5194 ( .A1(n10145), .A2(n4478), .ZN(n4787) );
  OAI21_X1 U5195 ( .B1(n4718), .B2(n6801), .A(n4457), .ZN(n4717) );
  OAI21_X1 U5196 ( .B1(n8717), .B2(n4697), .A(n5388), .ZN(n4696) );
  NOR2_X1 U5197 ( .A1(n4697), .A2(n4694), .ZN(n4693) );
  INV_X1 U5198 ( .A(n5349), .ZN(n4694) );
  NOR2_X1 U5199 ( .A1(n6422), .A2(n4885), .ZN(n4884) );
  INV_X1 U5200 ( .A(n6420), .ZN(n4885) );
  INV_X1 U5201 ( .A(n7306), .ZN(n4882) );
  NAND2_X1 U5202 ( .A1(n4645), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U5203 ( .A1(n4650), .A2(n4646), .ZN(n4645) );
  INV_X1 U5204 ( .A(n4618), .ZN(n4617) );
  AOI21_X1 U5205 ( .B1(n4618), .B2(n4622), .A(n4501), .ZN(n4616) );
  NOR2_X1 U5206 ( .A1(n4678), .A2(n8067), .ZN(n4677) );
  INV_X1 U5207 ( .A(n4679), .ZN(n4678) );
  INV_X1 U5208 ( .A(n5176), .ZN(n4755) );
  AOI21_X1 U5209 ( .B1(n4850), .B2(n4848), .A(n4847), .ZN(n6659) );
  NOR2_X1 U5210 ( .A1(n6813), .A2(n4849), .ZN(n4848) );
  OAI21_X1 U5211 ( .B1(n7202), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4613), .ZN(
        n7195) );
  NAND2_X1 U5212 ( .A1(n7202), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4613) );
  NAND2_X1 U5213 ( .A1(n7195), .A2(n7194), .ZN(n7193) );
  NAND2_X1 U5214 ( .A1(n7369), .A2(n7389), .ZN(n4605) );
  NAND2_X1 U5215 ( .A1(n7391), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4604) );
  NAND2_X1 U5216 ( .A1(n7727), .A2(n4615), .ZN(n7839) );
  OR2_X1 U5217 ( .A1(n7728), .A2(n7647), .ZN(n4615) );
  NAND2_X1 U5218 ( .A1(n10236), .A2(n4588), .ZN(n8489) );
  NAND2_X1 U5219 ( .A1(n8487), .A2(n10233), .ZN(n4588) );
  NOR2_X1 U5220 ( .A1(n4717), .A2(n4715), .ZN(n4714) );
  INV_X1 U5221 ( .A(n5498), .ZN(n4715) );
  INV_X1 U5222 ( .A(n4717), .ZN(n4712) );
  INV_X1 U5223 ( .A(n8631), .ZN(n4690) );
  INV_X1 U5224 ( .A(n8654), .ZN(n4691) );
  NAND2_X1 U5225 ( .A1(n4846), .A2(n6743), .ZN(n4845) );
  NAND2_X1 U5226 ( .A1(n5213), .A2(n4995), .ZN(n5218) );
  AND2_X1 U5227 ( .A1(n7796), .A2(n5217), .ZN(n5216) );
  NAND2_X1 U5228 ( .A1(n8433), .A2(n7802), .ZN(n6702) );
  NAND2_X1 U5229 ( .A1(n6862), .A2(n10286), .ZN(n6710) );
  NAND2_X1 U5230 ( .A1(n5051), .A2(n5041), .ZN(n6674) );
  OR2_X1 U5231 ( .A1(n8803), .A2(n8568), .ZN(n6799) );
  OR2_X1 U5232 ( .A1(n8339), .A2(n8719), .ZN(n6756) );
  OAI21_X1 U5233 ( .B1(n8107), .B2(n4514), .A(n5331), .ZN(n8158) );
  NOR3_X1 U5234 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U5235 ( .A1(n5009), .A2(n4948), .ZN(n4947) );
  NOR2_X1 U5236 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4948) );
  INV_X1 U5237 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5376) );
  OAI21_X1 U5238 ( .B1(n4629), .B2(n4633), .A(n4631), .ZN(n4627) );
  AOI21_X1 U5239 ( .B1(n6268), .B2(n4639), .A(n4641), .ZN(n4631) );
  OR2_X1 U5240 ( .A1(n5918), .A2(n7257), .ZN(n6262) );
  OR2_X1 U5241 ( .A1(n9655), .A2(n8899), .ZN(n9127) );
  INV_X1 U5242 ( .A(n9124), .ZN(n4831) );
  NOR2_X1 U5243 ( .A1(n9124), .A2(n4830), .ZN(n4834) );
  NOR2_X1 U5244 ( .A1(n6167), .A2(n6184), .ZN(n4830) );
  NAND2_X1 U5245 ( .A1(n9615), .A2(n4682), .ZN(n4681) );
  NOR2_X1 U5246 ( .A1(n9669), .A2(n9146), .ZN(n4682) );
  AND2_X1 U5247 ( .A1(n6232), .A2(n8187), .ZN(n6166) );
  AND2_X1 U5248 ( .A1(n6295), .A2(n6298), .ZN(n7707) );
  NAND2_X1 U5249 ( .A1(n6158), .A2(n6277), .ZN(n4625) );
  NAND2_X1 U5250 ( .A1(n4953), .A2(n4952), .ZN(n4951) );
  INV_X1 U5251 ( .A(n6386), .ZN(n4953) );
  NAND2_X1 U5252 ( .A1(n4727), .A2(n5520), .ZN(n5534) );
  NAND2_X1 U5253 ( .A1(n4737), .A2(n4735), .ZN(n5501) );
  AOI21_X1 U5254 ( .B1(n4739), .B2(n4741), .A(n4736), .ZN(n4735) );
  INV_X1 U5255 ( .A(n5485), .ZN(n4736) );
  NOR2_X1 U5256 ( .A1(n5395), .A2(n4769), .ZN(n4768) );
  INV_X1 U5257 ( .A(n5372), .ZN(n4769) );
  NAND2_X1 U5258 ( .A1(n4550), .A2(n4745), .ZN(n5352) );
  AOI21_X1 U5259 ( .B1(n4747), .B2(n4749), .A(n4517), .ZN(n4745) );
  NAND2_X1 U5260 ( .A1(n5316), .A2(n4747), .ZN(n4550) );
  NAND2_X1 U5261 ( .A1(n5263), .A2(n5249), .ZN(n5264) );
  NOR2_X1 U5262 ( .A1(n5244), .A2(n4840), .ZN(n4839) );
  INV_X1 U5263 ( .A(n5225), .ZN(n4840) );
  INV_X1 U5264 ( .A(n5240), .ZN(n5244) );
  AND2_X1 U5265 ( .A1(n5165), .A2(n5145), .ZN(n4734) );
  INV_X1 U5266 ( .A(n5148), .ZN(n4813) );
  OAI21_X1 U5267 ( .B1(n5902), .B2(P1_DATAO_REG_6__SCAN_IN), .A(n4732), .ZN(
        n5167) );
  NAND2_X1 U5268 ( .A1(n5902), .A2(n6997), .ZN(n4732) );
  AND2_X1 U5269 ( .A1(n8311), .A2(n6895), .ZN(n8314) );
  OR2_X1 U5270 ( .A1(n8361), .A2(n8358), .ZN(n6899) );
  INV_X1 U5271 ( .A(n6851), .ZN(n6921) );
  AND2_X1 U5272 ( .A1(n8179), .A2(n6869), .ZN(n6870) );
  NOR2_X1 U5273 ( .A1(n4910), .A2(n4907), .ZN(n4906) );
  NOR2_X1 U5274 ( .A1(n4912), .A2(n8637), .ZN(n4907) );
  INV_X1 U5275 ( .A(n8351), .ZN(n4910) );
  INV_X1 U5276 ( .A(n8433), .ZN(n6862) );
  AND2_X1 U5277 ( .A1(n5620), .A2(n7292), .ZN(n6944) );
  NOR2_X1 U5278 ( .A1(n8342), .A2(n4916), .ZN(n4915) );
  INV_X1 U5279 ( .A(n4918), .ZN(n4916) );
  INV_X1 U5280 ( .A(n8330), .ZN(n4921) );
  NAND2_X1 U5281 ( .A1(n4941), .A2(n4940), .ZN(n4937) );
  INV_X1 U5282 ( .A(n7765), .ZN(n4941) );
  INV_X1 U5283 ( .A(n8436), .ZN(n7761) );
  OR2_X1 U5284 ( .A1(n5026), .A2(n5013), .ZN(n5027) );
  INV_X1 U5285 ( .A(n5570), .ZN(n4595) );
  OR2_X1 U5286 ( .A1(n5072), .A2(n5200), .ZN(n5209) );
  NAND2_X1 U5287 ( .A1(n7390), .A2(n7389), .ZN(n10144) );
  NAND2_X1 U5288 ( .A1(n7388), .A2(n4789), .ZN(n4792) );
  XNOR2_X1 U5289 ( .A(n7369), .B(n4789), .ZN(n10130) );
  OR2_X1 U5290 ( .A1(n7373), .A2(n4789), .ZN(n4582) );
  OR2_X1 U5291 ( .A1(n10135), .A2(n10136), .ZN(n4580) );
  AND2_X1 U5292 ( .A1(n4580), .A2(n4510), .ZN(n10156) );
  NAND2_X1 U5293 ( .A1(n8448), .A2(n4599), .ZN(n7660) );
  OR2_X1 U5294 ( .A1(n8447), .A2(n7658), .ZN(n4599) );
  NAND2_X1 U5295 ( .A1(n4785), .A2(n4784), .ZN(n4783) );
  INV_X1 U5296 ( .A(n7634), .ZN(n4784) );
  XNOR2_X1 U5297 ( .A(n4469), .B(n7835), .ZN(n7736) );
  XNOR2_X1 U5298 ( .A(n7839), .B(n7835), .ZN(n7729) );
  NAND2_X1 U5299 ( .A1(n7729), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7841) );
  NOR2_X1 U5300 ( .A1(n4570), .A2(n8482), .ZN(n4569) );
  INV_X1 U5301 ( .A(n10170), .ZN(n4570) );
  NAND2_X1 U5302 ( .A1(n4574), .A2(n4573), .ZN(n4572) );
  INV_X1 U5303 ( .A(n4576), .ZN(n4574) );
  INV_X1 U5304 ( .A(n4528), .ZN(n4573) );
  NAND2_X1 U5305 ( .A1(n4800), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4799) );
  INV_X1 U5306 ( .A(n10192), .ZN(n4800) );
  NAND2_X1 U5307 ( .A1(n10186), .A2(n8484), .ZN(n10202) );
  NAND2_X1 U5308 ( .A1(n10202), .A2(n10203), .ZN(n10201) );
  NAND2_X1 U5309 ( .A1(n4778), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4777) );
  NAND2_X1 U5310 ( .A1(n10237), .A2(n10238), .ZN(n10236) );
  INV_X1 U5311 ( .A(n8515), .ZN(n4611) );
  AOI21_X1 U5312 ( .B1(n8515), .B2(n9447), .A(n4610), .ZN(n4607) );
  INV_X1 U5313 ( .A(n8524), .ZN(n4610) );
  NAND2_X1 U5314 ( .A1(n4716), .A2(n4718), .ZN(n8567) );
  NAND2_X1 U5315 ( .A1(n8597), .A2(n4722), .ZN(n4716) );
  INV_X1 U5316 ( .A(n6778), .ZN(n4865) );
  AOI21_X1 U5317 ( .B1(n8648), .B2(n5653), .A(n4986), .ZN(n8639) );
  NOR2_X1 U5318 ( .A1(n5652), .A2(n5651), .ZN(n4986) );
  AND2_X1 U5319 ( .A1(n6778), .A2(n6781), .ZN(n8638) );
  INV_X1 U5320 ( .A(n8704), .ZN(n5648) );
  AND4_X1 U5321 ( .A1(n5262), .A2(n5261), .A3(n5260), .A4(n5259), .ZN(n8134)
         );
  NAND2_X1 U5322 ( .A1(n4703), .A2(n4707), .ZN(n7928) );
  NAND2_X1 U5323 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  INV_X1 U5324 ( .A(n7942), .ZN(n4705) );
  OAI21_X1 U5325 ( .B1(n7679), .B2(n5156), .A(n5155), .ZN(n8247) );
  AND4_X1 U5326 ( .A1(n5162), .A2(n5161), .A3(n5160), .A4(n5159), .ZN(n7681)
         );
  XNOR2_X1 U5327 ( .A(n8438), .B(n10256), .ZN(n7576) );
  NAND2_X1 U5328 ( .A1(n5499), .A2(n5498), .ZN(n8597) );
  AND2_X1 U5329 ( .A1(n4858), .A2(n6792), .ZN(n4861) );
  NAND2_X1 U5330 ( .A1(n6791), .A2(n4859), .ZN(n4858) );
  NOR2_X1 U5331 ( .A1(n4540), .A2(n4864), .ZN(n4859) );
  INV_X1 U5332 ( .A(n4539), .ZN(n4862) );
  AND2_X1 U5333 ( .A1(n6631), .A2(n6630), .ZN(n8596) );
  AND2_X1 U5334 ( .A1(n6789), .A2(n6786), .ZN(n8623) );
  NAND2_X1 U5335 ( .A1(n8639), .A2(n8638), .ZN(n8754) );
  AND2_X1 U5336 ( .A1(n5415), .A2(n5414), .ZN(n8666) );
  NAND2_X1 U5337 ( .A1(n8666), .A2(n8665), .ZN(n8664) );
  NAND2_X1 U5338 ( .A1(n8160), .A2(n5349), .ZN(n8716) );
  AND4_X1 U5339 ( .A1(n5330), .A2(n5329), .A3(n5328), .A4(n5327), .ZN(n8161)
         );
  NAND2_X1 U5340 ( .A1(n4836), .A2(n6740), .ZN(n4835) );
  INV_X1 U5341 ( .A(n8042), .ZN(n4836) );
  NAND2_X1 U5342 ( .A1(n4706), .A2(n4700), .ZN(n4702) );
  NOR2_X1 U5343 ( .A1(n7942), .A2(n6874), .ZN(n4700) );
  OR2_X1 U5344 ( .A1(n5296), .A2(n4698), .ZN(n4701) );
  NOR2_X1 U5345 ( .A1(n5292), .A2(n4699), .ZN(n4698) );
  INV_X1 U5346 ( .A(n4707), .ZN(n4699) );
  AND2_X1 U5347 ( .A1(n6949), .A2(n6788), .ZN(n8694) );
  AND4_X1 U5348 ( .A1(n5311), .A2(n5310), .A3(n5309), .A4(n5308), .ZN(n8413)
         );
  INV_X1 U5349 ( .A(n8718), .ZN(n8695) );
  INV_X1 U5350 ( .A(n8635), .ZN(n8781) );
  NAND2_X1 U5351 ( .A1(n8035), .A2(n8026), .ZN(n5641) );
  NAND2_X1 U5352 ( .A1(n6721), .A2(n6720), .ZN(n8026) );
  AND2_X1 U5353 ( .A1(n5568), .A2(n4710), .ZN(n5014) );
  AND2_X1 U5354 ( .A1(n4709), .A2(n5008), .ZN(n4710) );
  NOR3_X1 U5355 ( .A1(n4947), .A2(P2_IR_REG_27__SCAN_IN), .A3(
        P2_IR_REG_28__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5356 ( .A1(n5589), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U5357 ( .A1(n5099), .A2(n4998), .ZN(n4945) );
  AND2_X1 U5358 ( .A1(n8930), .A2(n6535), .ZN(n8865) );
  AND2_X1 U5359 ( .A1(n6566), .A2(n6565), .ZN(n6592) );
  AND2_X1 U5360 ( .A1(n6453), .A2(n4876), .ZN(n4875) );
  AND2_X1 U5361 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  NAND2_X1 U5362 ( .A1(n4878), .A2(n4877), .ZN(n4876) );
  INV_X1 U5363 ( .A(n6430), .ZN(n6427) );
  OAI21_X1 U5364 ( .B1(n7066), .B2(n6385), .A(n6390), .ZN(n7049) );
  OAI22_X1 U5365 ( .A1(n6425), .A2(n9976), .B1(n9013), .B2(n6379), .ZN(n6389)
         );
  NAND2_X1 U5366 ( .A1(n6387), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6388) );
  INV_X1 U5367 ( .A(n6379), .ZN(n6387) );
  NOR2_X1 U5368 ( .A1(n6504), .A2(n6503), .ZN(n4899) );
  OR2_X1 U5369 ( .A1(n8878), .A2(n6505), .ZN(n4900) );
  NAND2_X1 U5370 ( .A1(n6527), .A2(n6528), .ZN(n4902) );
  INV_X1 U5371 ( .A(n8946), .ZN(n6528) );
  XNOR2_X1 U5372 ( .A(n6398), .B(n6383), .ZN(n6401) );
  NOR2_X1 U5373 ( .A1(n4869), .A2(n8916), .ZN(n4868) );
  NOR2_X1 U5374 ( .A1(n6487), .A2(n6488), .ZN(n4869) );
  AOI21_X1 U5375 ( .B1(n8929), .B2(n4892), .A(n4891), .ZN(n4890) );
  INV_X1 U5376 ( .A(n8930), .ZN(n4892) );
  INV_X1 U5377 ( .A(n6546), .ZN(n4891) );
  XOR2_X1 U5378 ( .A(n6556), .B(n6555), .Z(n8897) );
  NAND2_X1 U5379 ( .A1(n6470), .A2(n6472), .ZN(n6473) );
  INV_X1 U5380 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n4905) );
  INV_X1 U5381 ( .A(n4449), .ZN(n6004) );
  AND4_X1 U5382 ( .A1(n5943), .A2(n5942), .A3(n5941), .A4(n5940), .ZN(n8994)
         );
  AND4_X1 U5383 ( .A1(n5950), .A2(n5949), .A3(n5948), .A4(n5947), .ZN(n8971)
         );
  AND4_X1 U5384 ( .A1(n6034), .A2(n6033), .A3(n6032), .A4(n6031), .ZN(n7808)
         );
  OR2_X1 U5385 ( .A1(n4448), .A2(n6083), .ZN(n6086) );
  INV_X1 U5386 ( .A(n5919), .ZN(n6099) );
  NOR2_X1 U5387 ( .A1(n4658), .A2(n4657), .ZN(n4656) );
  INV_X1 U5388 ( .A(n9079), .ZN(n4657) );
  INV_X1 U5389 ( .A(n9077), .ZN(n4658) );
  INV_X1 U5390 ( .A(n4675), .ZN(n4671) );
  NOR2_X1 U5391 ( .A1(n9213), .A2(n4672), .ZN(n9113) );
  NAND2_X1 U5392 ( .A1(n4675), .A2(n4673), .ZN(n4672) );
  NOR2_X1 U5393 ( .A1(n6269), .A2(n9640), .ZN(n4673) );
  AND2_X1 U5394 ( .A1(n4676), .A2(n4674), .ZN(n9173) );
  NAND2_X1 U5395 ( .A1(n9215), .A2(n4485), .ZN(n9193) );
  AND2_X1 U5396 ( .A1(n6245), .A2(n9132), .ZN(n9216) );
  AOI21_X1 U5397 ( .B1(n9556), .B2(n4962), .A(n4515), .ZN(n4961) );
  NAND2_X1 U5398 ( .A1(n4966), .A2(n9150), .ZN(n9605) );
  NOR2_X1 U5399 ( .A1(n4969), .A2(n4968), .ZN(n4967) );
  NAND2_X1 U5400 ( .A1(n8070), .A2(n8075), .ZN(n4810) );
  NAND2_X1 U5401 ( .A1(n4810), .A2(n4808), .ZN(n8188) );
  NOR2_X1 U5402 ( .A1(n8195), .A2(n4809), .ZN(n4808) );
  INV_X1 U5403 ( .A(n6231), .ZN(n4809) );
  INV_X1 U5404 ( .A(n6166), .ZN(n8195) );
  NAND2_X1 U5405 ( .A1(n7966), .A2(n6307), .ZN(n8070) );
  AND2_X1 U5406 ( .A1(n6231), .A2(n6226), .ZN(n8075) );
  OR2_X1 U5407 ( .A1(n7898), .A2(n8989), .ZN(n4993) );
  NOR2_X2 U5408 ( .A1(n4993), .A2(n9763), .ZN(n8079) );
  NAND2_X1 U5409 ( .A1(n7708), .A2(n7707), .ZN(n4816) );
  NAND2_X1 U5410 ( .A1(n7532), .A2(n4560), .ZN(n7561) );
  AND2_X1 U5411 ( .A1(n6162), .A2(n6292), .ZN(n4560) );
  AND2_X1 U5412 ( .A1(n6210), .A2(n6292), .ZN(n7547) );
  NAND2_X1 U5413 ( .A1(n6161), .A2(n6290), .ZN(n7533) );
  NAND2_X1 U5414 ( .A1(n7533), .A2(n7547), .ZN(n7532) );
  OR2_X1 U5415 ( .A1(n6060), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U5416 ( .A1(n4827), .A2(n4825), .ZN(n7449) );
  NOR2_X1 U5417 ( .A1(n7476), .A2(n4826), .ZN(n4825) );
  INV_X1 U5418 ( .A(n5787), .ZN(n4826) );
  NAND2_X1 U5419 ( .A1(n7275), .A2(n6156), .ZN(n9945) );
  NAND2_X1 U5420 ( .A1(n5728), .A2(n5727), .ZN(n9649) );
  NAND2_X1 U5421 ( .A1(n5826), .A2(n5825), .ZN(n9664) );
  INV_X1 U5422 ( .A(n8197), .ZN(n9753) );
  NAND2_X1 U5423 ( .A1(n5862), .A2(n5718), .ZN(n4975) );
  NOR2_X1 U5424 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5718) );
  NAND2_X1 U5425 ( .A1(n5435), .A2(n5434), .ZN(n5450) );
  NAND2_X1 U5426 ( .A1(n4553), .A2(n5394), .ZN(n5418) );
  NAND2_X1 U5427 ( .A1(n4773), .A2(n4768), .ZN(n4553) );
  NAND2_X1 U5428 ( .A1(n4773), .A2(n5372), .ZN(n5396) );
  NAND2_X1 U5429 ( .A1(n4746), .A2(n5318), .ZN(n5334) );
  NAND2_X1 U5430 ( .A1(n5316), .A2(n5315), .ZN(n4746) );
  XNOR2_X1 U5431 ( .A(n5265), .B(n5264), .ZN(n7053) );
  NAND2_X1 U5432 ( .A1(n4838), .A2(n5243), .ZN(n5265) );
  XNOR2_X1 U5433 ( .A(n5245), .B(n5240), .ZN(n7031) );
  XNOR2_X1 U5434 ( .A(n5224), .B(n5223), .ZN(n7029) );
  OAI21_X1 U5435 ( .B1(n5173), .B2(n4467), .A(n4757), .ZN(n5224) );
  XNOR2_X1 U5436 ( .A(n5197), .B(n5196), .ZN(n7007) );
  AND2_X1 U5437 ( .A1(n4805), .A2(n5105), .ZN(n4804) );
  AND2_X1 U5438 ( .A1(n5766), .A2(n5769), .ZN(n7099) );
  NAND2_X1 U5439 ( .A1(n8368), .A2(n6882), .ZN(n8295) );
  NAND2_X1 U5440 ( .A1(n5474), .A2(n5473), .ZN(n8749) );
  INV_X1 U5441 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5442 ( .B1(n4938), .B2(n4940), .A(n6860), .ZN(n4936) );
  AND3_X1 U5443 ( .A1(n5460), .A2(n5459), .A3(n5458), .ZN(n8622) );
  AND3_X1 U5444 ( .A1(n5133), .A2(n5132), .A3(n5131), .ZN(n7611) );
  NAND2_X1 U5445 ( .A1(n5364), .A2(n5363), .ZN(n8711) );
  INV_X1 U5446 ( .A(n8423), .ZN(n8611) );
  NAND2_X1 U5447 ( .A1(n6855), .A2(n4444), .ZN(n4932) );
  NAND2_X1 U5448 ( .A1(n5455), .A2(n5454), .ZN(n8641) );
  AND3_X1 U5449 ( .A1(n5154), .A2(n5153), .A3(n5152), .ZN(n10276) );
  NAND2_X1 U5450 ( .A1(n4453), .A2(n5667), .ZN(n4548) );
  INV_X1 U5451 ( .A(n8161), .ZN(n8427) );
  OR2_X1 U5452 ( .A1(n5206), .A2(n5021), .ZN(n5022) );
  OR2_X1 U5453 ( .A1(n5205), .A2(n7503), .ZN(n5023) );
  OAI21_X1 U5454 ( .B1(n10244), .B2(n4794), .A(n4793), .ZN(n8521) );
  NAND2_X1 U5455 ( .A1(n4797), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4794) );
  INV_X1 U5456 ( .A(n8477), .ZN(n4797) );
  INV_X1 U5457 ( .A(n8476), .ZN(n4795) );
  AOI21_X1 U5458 ( .B1(n4594), .B2(n8528), .A(n4590), .ZN(n4589) );
  NAND2_X1 U5459 ( .A1(n4593), .A2(n4591), .ZN(n4590) );
  NOR2_X1 U5460 ( .A1(n8529), .A2(n8492), .ZN(n4594) );
  AOI21_X1 U5461 ( .B1(n10231), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n4592), .ZN(
        n4591) );
  OAI21_X1 U5462 ( .B1(n5587), .B2(n8635), .A(n5586), .ZN(n8559) );
  NOR2_X1 U5463 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  NOR2_X1 U5464 ( .A1(n6354), .A2(n8720), .ZN(n5584) );
  NAND2_X1 U5465 ( .A1(n5556), .A2(n5555), .ZN(n8563) );
  AOI21_X1 U5466 ( .B1(n8219), .B2(n6627), .A(n5508), .ZN(n8603) );
  NAND2_X1 U5467 ( .A1(n5649), .A2(n5648), .ZN(n8772) );
  NAND2_X1 U5468 ( .A1(n5270), .A2(n5269), .ZN(n8127) );
  AOI22_X1 U5469 ( .A1(n9698), .A2(n6627), .B1(n6618), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8793) );
  NOR2_X1 U5470 ( .A1(n8551), .A2(n6365), .ZN(n6373) );
  AND2_X1 U5471 ( .A1(n8550), .A2(n10272), .ZN(n6365) );
  NAND2_X1 U5472 ( .A1(n7820), .A2(n6627), .ZN(n4552) );
  INV_X1 U5473 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6971) );
  AND2_X1 U5474 ( .A1(n6614), .A2(n8968), .ZN(n6615) );
  NAND2_X1 U5475 ( .A1(n5742), .A2(n5741), .ZN(n8921) );
  NAND2_X1 U5476 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  AND2_X1 U5477 ( .A1(n8969), .A2(n8970), .ZN(n6559) );
  MUX2_X1 U5478 ( .A(n6274), .B(n6273), .S(n6376), .Z(n6333) );
  OAI21_X1 U5479 ( .B1(n6330), .B2(n7022), .A(n6600), .ZN(n6331) );
  NAND2_X1 U5480 ( .A1(n4665), .A2(n4664), .ZN(n9063) );
  NAND2_X1 U5481 ( .A1(n9862), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4664) );
  INV_X1 U5482 ( .A(n9863), .ZN(n4665) );
  NOR2_X1 U5483 ( .A1(n4996), .A2(n4964), .ZN(n4963) );
  INV_X1 U5484 ( .A(n7974), .ZN(n4964) );
  OAI21_X1 U5485 ( .B1(n9641), .B2(n10018), .A(n4564), .ZN(n4563) );
  MUX2_X1 U5486 ( .A(n6669), .B(n6668), .S(n6959), .Z(n6683) );
  OAI211_X1 U5487 ( .C1(n7417), .C2(n4643), .A(n4644), .B(n4642), .ZN(n6208)
         );
  NAND2_X1 U5488 ( .A1(n6189), .A2(n7023), .ZN(n4643) );
  NAND2_X1 U5489 ( .A1(n6065), .A2(n7023), .ZN(n4642) );
  NAND2_X1 U5490 ( .A1(n6196), .A2(n6266), .ZN(n4644) );
  NAND2_X1 U5491 ( .A1(n4536), .A2(n4533), .ZN(n6798) );
  NAND2_X1 U5492 ( .A1(n4534), .A2(n6794), .ZN(n4533) );
  AOI21_X1 U5493 ( .B1(n6230), .B2(n4647), .A(n6240), .ZN(n4646) );
  NOR2_X1 U5494 ( .A1(n4649), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U5495 ( .A1(n4730), .A2(n4483), .ZN(n6816) );
  NOR2_X1 U5496 ( .A1(n6814), .A2(n6813), .ZN(n6815) );
  NAND2_X1 U5497 ( .A1(n4730), .A2(n4484), .ZN(n6818) );
  INV_X1 U5498 ( .A(n4503), .ZN(n4847) );
  MUX2_X1 U5499 ( .A(n6263), .B(n6262), .S(n7023), .Z(n6264) );
  NAND2_X1 U5500 ( .A1(n4619), .A2(n4620), .ZN(n6252) );
  NAND2_X1 U5501 ( .A1(n4468), .A2(n9540), .ZN(n4619) );
  NOR2_X1 U5502 ( .A1(n7990), .A2(n8095), .ZN(n4679) );
  NAND2_X1 U5503 ( .A1(n5686), .A2(n5685), .ZN(n5688) );
  INV_X1 U5504 ( .A(n4748), .ZN(n4747) );
  OAI21_X1 U5505 ( .B1(n5315), .B2(n4749), .A(n5333), .ZN(n4748) );
  INV_X1 U5506 ( .A(n5318), .ZN(n4749) );
  NAND2_X1 U5507 ( .A1(n5276), .A2(n5263), .ZN(n4761) );
  NAND2_X1 U5508 ( .A1(n6657), .A2(n7514), .ZN(n6826) );
  XNOR2_X1 U5509 ( .A(n7202), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7191) );
  AND2_X1 U5510 ( .A1(n7163), .A2(n7160), .ZN(n7210) );
  NAND2_X1 U5511 ( .A1(n7148), .A2(n7193), .ZN(n7149) );
  OR2_X1 U5512 ( .A1(n10145), .A2(n4791), .ZN(n4790) );
  AOI21_X1 U5513 ( .B1(n7390), .B2(n4788), .A(n4787), .ZN(n4786) );
  NOR2_X1 U5514 ( .A1(n10145), .A2(n4789), .ZN(n4788) );
  AOI21_X1 U5515 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n7638), .A(n8455), .ZN(
        n7631) );
  NOR2_X1 U5516 ( .A1(n7631), .A2(n7700), .ZN(n7633) );
  NAND2_X1 U5517 ( .A1(n8464), .A2(n8463), .ZN(n8466) );
  NAND2_X1 U5518 ( .A1(n10183), .A2(n4614), .ZN(n8509) );
  OR2_X1 U5519 ( .A1(n10182), .A2(n8508), .ZN(n4614) );
  AND2_X1 U5520 ( .A1(n5650), .A2(n6766), .ZN(n8675) );
  INV_X1 U5521 ( .A(n4696), .ZN(n4695) );
  AND2_X1 U5522 ( .A1(n6761), .A2(n6744), .ZN(n6746) );
  NAND2_X1 U5523 ( .A1(n4471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U5524 ( .A1(n5378), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5402) );
  OR2_X1 U5525 ( .A1(n6450), .A2(n8087), .ZN(n6452) );
  AOI21_X1 U5526 ( .B1(n4882), .B2(n4884), .A(n4498), .ZN(n4881) );
  INV_X1 U5527 ( .A(n4884), .ZN(n4883) );
  OR2_X1 U5528 ( .A1(n6465), .A2(n6464), .ZN(n6466) );
  NAND2_X1 U5529 ( .A1(n4630), .A2(n6270), .ZN(n4629) );
  NAND2_X1 U5530 ( .A1(n4633), .A2(n4637), .ZN(n4630) );
  NAND2_X1 U5531 ( .A1(n4638), .A2(n6269), .ZN(n4637) );
  NAND2_X1 U5532 ( .A1(n6268), .A2(n4488), .ZN(n4632) );
  OAI21_X1 U5533 ( .B1(n4468), .B2(n4617), .A(n4616), .ZN(n6247) );
  NOR2_X1 U5534 ( .A1(n9885), .A2(n4667), .ZN(n9067) );
  AND2_X1 U5535 ( .A1(n9893), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4667) );
  INV_X1 U5536 ( .A(n9094), .ZN(n4655) );
  NOR2_X1 U5537 ( .A1(n5918), .A2(n9633), .ZN(n4675) );
  INV_X1 U5538 ( .A(n9135), .ZN(n4821) );
  AND2_X1 U5539 ( .A1(P1_REG3_REG_25__SCAN_IN), .A2(n5946), .ZN(n5936) );
  NAND2_X1 U5540 ( .A1(n4823), .A2(n9132), .ZN(n4822) );
  AND2_X1 U5541 ( .A1(n9130), .A2(n6251), .ZN(n9129) );
  NOR2_X1 U5542 ( .A1(n9567), .A2(n9122), .ZN(n4960) );
  INV_X1 U5543 ( .A(n9154), .ZN(n4962) );
  INV_X1 U5544 ( .A(n9616), .ZN(n4969) );
  INV_X1 U5545 ( .A(n9147), .ZN(n4968) );
  NAND2_X1 U5546 ( .A1(n8195), .A2(n4971), .ZN(n4972) );
  INV_X1 U5547 ( .A(n8144), .ZN(n4971) );
  NAND2_X1 U5548 ( .A1(n7568), .A2(n4481), .ZN(n7898) );
  NOR2_X1 U5549 ( .A1(n7344), .A2(n6160), .ZN(n6284) );
  NAND2_X1 U5550 ( .A1(n6195), .A2(n6082), .ZN(n6285) );
  AND2_X1 U5551 ( .A1(n4803), .A2(n7450), .ZN(n6290) );
  NAND2_X1 U5552 ( .A1(n6195), .A2(n4486), .ZN(n4803) );
  NAND2_X1 U5553 ( .A1(n4829), .A2(n4455), .ZN(n7451) );
  NAND2_X1 U5554 ( .A1(n7568), .A2(n4679), .ZN(n7810) );
  AND2_X1 U5555 ( .A1(n7539), .A2(n10058), .ZN(n7568) );
  OR2_X1 U5556 ( .A1(n7520), .A2(n7466), .ZN(n7454) );
  NOR2_X1 U5557 ( .A1(n9974), .A2(n4447), .ZN(n9955) );
  XNOR2_X1 U5558 ( .A(n5688), .B(n5689), .ZN(n5832) );
  NAND2_X1 U5559 ( .A1(n5503), .A2(n5502), .ZN(n5519) );
  INV_X1 U5560 ( .A(n5448), .ZN(n4744) );
  INV_X1 U5561 ( .A(n4766), .ZN(n4765) );
  OAI21_X1 U5562 ( .B1(n4768), .B2(n4767), .A(n5416), .ZN(n4766) );
  NAND2_X1 U5563 ( .A1(n5417), .A2(n5416), .ZN(n4772) );
  INV_X1 U5564 ( .A(n5373), .ZN(n4774) );
  INV_X1 U5565 ( .A(n5196), .ZN(n4751) );
  NOR2_X1 U5566 ( .A1(n5172), .A2(n4755), .ZN(n4750) );
  INV_X1 U5567 ( .A(n5101), .ZN(n4807) );
  INV_X1 U5568 ( .A(n5087), .ZN(n4806) );
  OAI21_X1 U5569 ( .B1(n5902), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5106), .ZN(
        n5123) );
  NAND2_X1 U5570 ( .A1(n5902), .A2(n6974), .ZN(n5106) );
  NAND2_X1 U5571 ( .A1(n7602), .A2(n5030), .ZN(n4802) );
  OAI21_X1 U5572 ( .B1(n6918), .B2(n4925), .A(n4922), .ZN(n6928) );
  AOI21_X1 U5573 ( .B1(n8395), .B2(n4924), .A(n4923), .ZN(n4922) );
  INV_X1 U5574 ( .A(n6917), .ZN(n4924) );
  INV_X1 U5575 ( .A(n8259), .ZN(n4923) );
  OR2_X1 U5576 ( .A1(n6885), .A2(n8161), .ZN(n6886) );
  AND2_X1 U5577 ( .A1(n4919), .A2(n8331), .ZN(n4918) );
  NAND2_X1 U5578 ( .A1(n8330), .A2(n4920), .ZN(n4919) );
  INV_X1 U5579 ( .A(n6886), .ZN(n4920) );
  OR2_X1 U5580 ( .A1(n6896), .A2(n8314), .ZN(n8358) );
  AOI21_X1 U5581 ( .B1(n8278), .B2(n8279), .A(n6904), .ZN(n6905) );
  XNOR2_X1 U5582 ( .A(n6851), .B(n6848), .ZN(n6850) );
  NAND2_X1 U5583 ( .A1(n6655), .A2(n7853), .ZN(n6664) );
  AND4_X1 U5584 ( .A1(n5193), .A2(n5192), .A3(n5191), .A4(n5190), .ZN(n6864)
         );
  NAND2_X1 U5585 ( .A1(n4587), .A2(n4586), .ZN(n4585) );
  NAND2_X1 U5586 ( .A1(n7642), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4586) );
  OR2_X1 U5587 ( .A1(n7642), .A2(n5017), .ZN(n4587) );
  NAND2_X1 U5588 ( .A1(n7210), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7213) );
  NAND2_X1 U5589 ( .A1(n4530), .A2(n4792), .ZN(n10146) );
  NAND2_X1 U5590 ( .A1(n4606), .A2(n4605), .ZN(n4603) );
  INV_X1 U5591 ( .A(n10141), .ZN(n4602) );
  NAND2_X1 U5592 ( .A1(n10141), .A2(n4604), .ZN(n4601) );
  OR2_X1 U5593 ( .A1(n5337), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5594 ( .A1(n7393), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U5595 ( .A1(n4581), .A2(n7381), .ZN(n8441) );
  NAND2_X1 U5596 ( .A1(n4578), .A2(n4577), .ZN(n4581) );
  AOI21_X1 U5597 ( .B1(n4510), .B2(n10136), .A(n7382), .ZN(n4577) );
  NAND2_X1 U5598 ( .A1(n10135), .A2(n4510), .ZN(n4578) );
  AOI21_X1 U5599 ( .B1(n8441), .B2(n8440), .A(n8439), .ZN(n8443) );
  NOR2_X1 U5600 ( .A1(n7692), .A2(n7872), .ZN(n7691) );
  NAND2_X1 U5601 ( .A1(n7689), .A2(n7661), .ZN(n7662) );
  NAND2_X1 U5602 ( .A1(n7735), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4782) );
  NOR2_X1 U5603 ( .A1(n7736), .A2(n5256), .ZN(n7827) );
  OR2_X1 U5604 ( .A1(n7831), .A2(n7830), .ZN(n8464) );
  NAND2_X1 U5605 ( .A1(n7841), .A2(n7842), .ZN(n8501) );
  XNOR2_X1 U5606 ( .A(n8466), .B(n8506), .ZN(n10173) );
  NAND2_X1 U5607 ( .A1(n10166), .A2(n8507), .ZN(n10184) );
  NAND2_X1 U5608 ( .A1(n10184), .A2(n10185), .ZN(n10183) );
  NAND2_X1 U5609 ( .A1(n4568), .A2(n4567), .ZN(n10187) );
  AOI21_X1 U5610 ( .B1(n4569), .B2(n4572), .A(n4525), .ZN(n4567) );
  NOR2_X1 U5611 ( .A1(n10173), .A2(n8467), .ZN(n10176) );
  XNOR2_X1 U5612 ( .A(n8509), .B(n10198), .ZN(n10200) );
  AND2_X1 U5613 ( .A1(n4777), .A2(n4475), .ZN(n10225) );
  NOR2_X1 U5614 ( .A1(n10225), .A2(n10224), .ZN(n10223) );
  NAND2_X1 U5615 ( .A1(n10201), .A2(n8485), .ZN(n10219) );
  NAND2_X1 U5616 ( .A1(n10219), .A2(n10220), .ZN(n10218) );
  NOR2_X1 U5617 ( .A1(n8497), .A2(P2_STATE_REG_SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5618 ( .A1(n10232), .A2(n8516), .ZN(n4593) );
  INV_X1 U5619 ( .A(n8489), .ZN(n8491) );
  AND2_X1 U5620 ( .A1(n4508), .A2(n4852), .ZN(n4851) );
  NAND2_X1 U5621 ( .A1(n8264), .A2(n4853), .ZN(n4852) );
  INV_X1 U5622 ( .A(n6807), .ZN(n4853) );
  OR2_X1 U5623 ( .A1(n8579), .A2(n6651), .ZN(n4850) );
  AND2_X1 U5624 ( .A1(n6656), .A2(n6804), .ZN(n6653) );
  NAND2_X1 U5625 ( .A1(n8579), .A2(n6807), .ZN(n5658) );
  NAND2_X1 U5626 ( .A1(n4713), .A2(n4711), .ZN(n6347) );
  NAND2_X1 U5627 ( .A1(n4712), .A2(n4456), .ZN(n4711) );
  NAND2_X1 U5628 ( .A1(n5499), .A2(n4714), .ZN(n4713) );
  NOR2_X1 U5629 ( .A1(n8589), .A2(n8718), .ZN(n5585) );
  AND2_X1 U5630 ( .A1(n5509), .A2(n8324), .ZN(n5526) );
  NOR2_X1 U5631 ( .A1(n5492), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5509) );
  OR2_X1 U5632 ( .A1(n5456), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5475) );
  OR2_X1 U5633 ( .A1(n5475), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5492) );
  AND3_X1 U5634 ( .A1(n5443), .A2(n5442), .A3(n5441), .ZN(n8636) );
  NAND2_X1 U5635 ( .A1(n4686), .A2(n4689), .ZN(n5462) );
  AOI21_X1 U5636 ( .B1(n4691), .B2(n8652), .A(n4690), .ZN(n4689) );
  NOR2_X1 U5637 ( .A1(n5408), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5427) );
  INV_X1 U5638 ( .A(n4855), .ZN(n4854) );
  OAI21_X1 U5639 ( .B1(n5648), .B2(n6748), .A(n8675), .ZN(n4855) );
  AND3_X1 U5640 ( .A1(n5433), .A2(n5432), .A3(n5431), .ZN(n8678) );
  NAND2_X1 U5641 ( .A1(n8715), .A2(n5371), .ZN(n8691) );
  NAND2_X1 U5642 ( .A1(n5365), .A2(n8344), .ZN(n5381) );
  NOR2_X1 U5643 ( .A1(n5325), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5342) );
  OR2_X1 U5644 ( .A1(n5306), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5325) );
  NOR2_X1 U5645 ( .A1(n5271), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5285) );
  OR2_X1 U5646 ( .A1(n5234), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5257) );
  OR2_X1 U5647 ( .A1(n5220), .A2(n5219), .ZN(n5221) );
  NAND2_X1 U5648 ( .A1(n5204), .A2(n9491), .ZN(n5234) );
  AOI21_X1 U5649 ( .B1(n8244), .B2(n5636), .A(n6707), .ZN(n7862) );
  INV_X1 U5650 ( .A(n6638), .ZN(n7863) );
  NOR2_X1 U5651 ( .A1(n5157), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5202) );
  INV_X1 U5652 ( .A(n7796), .ZN(n8246) );
  XNOR2_X1 U5653 ( .A(n7608), .B(n5632), .ZN(n7747) );
  INV_X1 U5654 ( .A(n6849), .ZN(n5051) );
  NAND2_X1 U5655 ( .A1(n7505), .A2(n5050), .ZN(n7509) );
  NAND2_X1 U5656 ( .A1(n6674), .A2(n6676), .ZN(n7505) );
  NAND2_X1 U5657 ( .A1(n5625), .A2(n8784), .ZN(n6671) );
  NAND2_X1 U5658 ( .A1(n4861), .A2(n4862), .ZN(n4856) );
  AOI21_X1 U5659 ( .B1(n8664), .B2(n8654), .A(n8655), .ZN(n4688) );
  AND4_X1 U5660 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n8719)
         );
  NAND2_X1 U5661 ( .A1(n8716), .A2(n8717), .ZN(n8715) );
  AOI21_X1 U5662 ( .B1(n5646), .B2(n4844), .A(n4843), .ZN(n4846) );
  INV_X1 U5663 ( .A(n6746), .ZN(n8717) );
  INV_X1 U5664 ( .A(n8158), .ZN(n5348) );
  NAND2_X1 U5665 ( .A1(n4837), .A2(n6734), .ZN(n8042) );
  NAND2_X1 U5666 ( .A1(n7994), .A2(n6735), .ZN(n4837) );
  AND2_X1 U5667 ( .A1(n6734), .A2(n6735), .ZN(n8000) );
  INV_X1 U5668 ( .A(n5009), .ZN(n4946) );
  INV_X1 U5669 ( .A(n4597), .ZN(n4596) );
  OR2_X1 U5670 ( .A1(n6076), .A2(n6058), .ZN(n6060) );
  AOI21_X1 U5671 ( .B1(n4898), .B2(n6505), .A(n4895), .ZN(n4894) );
  INV_X1 U5672 ( .A(n6510), .ZN(n4895) );
  NAND2_X1 U5673 ( .A1(n7776), .A2(n7775), .ZN(n4880) );
  NAND2_X1 U5674 ( .A1(n6534), .A2(n6533), .ZN(n8930) );
  XNOR2_X1 U5675 ( .A(n6406), .B(n6552), .ZN(n6408) );
  NAND2_X1 U5676 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U5677 ( .A1(n4904), .A2(n6403), .ZN(n6404) );
  NOR2_X1 U5678 ( .A1(n8936), .A2(n4899), .ZN(n4898) );
  OAI21_X1 U5679 ( .B1(n4875), .B2(n4873), .A(n4494), .ZN(n4872) );
  INV_X1 U5680 ( .A(n7984), .ZN(n4873) );
  NOR2_X1 U5681 ( .A1(n6115), .A2(n7248), .ZN(n6116) );
  NAND2_X1 U5682 ( .A1(n7305), .A2(n7306), .ZN(n7304) );
  OR2_X1 U5683 ( .A1(n6138), .A2(n6139), .ZN(n6334) );
  AND2_X1 U5684 ( .A1(n5957), .A2(n5956), .ZN(n8899) );
  AND2_X1 U5685 ( .A1(n5978), .A2(n5977), .ZN(n8938) );
  AND2_X1 U5686 ( .A1(n6120), .A2(n6119), .ZN(n6123) );
  NAND2_X1 U5687 ( .A1(n9042), .A2(n4489), .ZN(n9816) );
  NAND2_X1 U5688 ( .A1(n9816), .A2(n9817), .ZN(n9815) );
  AND2_X1 U5689 ( .A1(n9815), .A2(n4663), .ZN(n9832) );
  NAND2_X1 U5690 ( .A1(n7099), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4663) );
  NOR2_X1 U5691 ( .A1(n9721), .A2(n4660), .ZN(n9737) );
  NOR2_X1 U5692 ( .A1(n4662), .A2(n4661), .ZN(n4660) );
  NOR2_X1 U5693 ( .A1(n9737), .A2(n9738), .ZN(n9736) );
  NOR2_X1 U5694 ( .A1(n9736), .A2(n4659), .ZN(n7106) );
  AND2_X1 U5695 ( .A1(n9731), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U5696 ( .A1(n7106), .A2(n7105), .ZN(n7431) );
  NOR2_X1 U5697 ( .A1(n9707), .A2(n4666), .ZN(n9865) );
  AND2_X1 U5698 ( .A1(n9712), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4666) );
  AND2_X1 U5699 ( .A1(n9703), .A2(n7437), .ZN(n9857) );
  NOR2_X1 U5700 ( .A1(n9865), .A2(n9864), .ZN(n9863) );
  NOR2_X1 U5701 ( .A1(n9873), .A2(n4668), .ZN(n9887) );
  AND2_X1 U5702 ( .A1(n9881), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U5703 ( .A1(n9887), .A2(n9886), .ZN(n9885) );
  XNOR2_X1 U5704 ( .A(n9067), .B(n9066), .ZN(n9902) );
  OR2_X1 U5705 ( .A1(n9071), .A2(n9070), .ZN(n9078) );
  OR2_X1 U5706 ( .A1(n9070), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U5707 ( .A1(n4819), .A2(n4817), .ZN(n9180) );
  NAND2_X1 U5708 ( .A1(n4818), .A2(n9135), .ZN(n4817) );
  NAND2_X1 U5709 ( .A1(n9231), .A2(n4820), .ZN(n4819) );
  NOR2_X1 U5710 ( .A1(n4821), .A2(n9133), .ZN(n4820) );
  NAND2_X1 U5711 ( .A1(n6257), .A2(n9136), .ZN(n9188) );
  INV_X1 U5712 ( .A(n4824), .ZN(n9198) );
  AOI21_X1 U5713 ( .B1(n9231), .B2(n9132), .A(n4818), .ZN(n9196) );
  NOR2_X1 U5714 ( .A1(n9649), .A2(n9545), .ZN(n9226) );
  OR2_X1 U5715 ( .A1(n9664), .A2(n8995), .ZN(n9565) );
  NAND2_X1 U5716 ( .A1(n4833), .A2(n4452), .ZN(n9578) );
  NAND2_X1 U5717 ( .A1(n4831), .A2(n6184), .ZN(n4832) );
  NOR2_X1 U5718 ( .A1(n9578), .A2(n9579), .ZN(n9577) );
  NOR2_X1 U5719 ( .A1(n5984), .A2(n5912), .ZN(n5970) );
  AND2_X1 U5720 ( .A1(n6237), .A2(n6238), .ZN(n9594) );
  AND2_X1 U5721 ( .A1(n8190), .A2(n6233), .ZN(n9617) );
  OR2_X1 U5722 ( .A1(n9144), .A2(n9143), .ZN(n9148) );
  NAND2_X1 U5723 ( .A1(n6168), .A2(n6167), .ZN(n8190) );
  NOR2_X1 U5724 ( .A1(n8211), .A2(n6024), .ZN(n6014) );
  NAND2_X1 U5725 ( .A1(n7904), .A2(n6165), .ZN(n7965) );
  NAND2_X1 U5726 ( .A1(n4816), .A2(n4815), .ZN(n7893) );
  AND2_X1 U5727 ( .A1(n6163), .A2(n6295), .ZN(n4815) );
  NAND2_X1 U5728 ( .A1(n7893), .A2(n6219), .ZN(n7904) );
  AND2_X1 U5729 ( .A1(n6302), .A2(n6217), .ZN(n7891) );
  NOR2_X1 U5730 ( .A1(n6037), .A2(n7442), .ZN(n6030) );
  INV_X1 U5731 ( .A(n7566), .ZN(n4957) );
  NOR2_X1 U5732 ( .A1(n6053), .A2(n6043), .ZN(n6067) );
  NOR2_X1 U5733 ( .A1(n7454), .A2(n10048), .ZN(n7539) );
  OAI21_X1 U5734 ( .B1(n7515), .B2(n6194), .A(n6193), .ZN(n7417) );
  NAND2_X1 U5735 ( .A1(n4625), .A2(n6159), .ZN(n7344) );
  NAND2_X1 U5736 ( .A1(n4623), .A2(n4625), .ZN(n7347) );
  INV_X1 U5737 ( .A(n6159), .ZN(n4624) );
  NOR2_X1 U5738 ( .A1(n9939), .A2(n7407), .ZN(n7521) );
  OR2_X1 U5739 ( .A1(n6992), .A2(n5780), .ZN(n5772) );
  OAI21_X1 U5740 ( .B1(n9945), .B2(n6157), .A(n6280), .ZN(n9928) );
  NAND2_X1 U5741 ( .A1(n7276), .A2(n7323), .ZN(n7275) );
  AND2_X1 U5742 ( .A1(n9175), .A2(n9174), .ZN(n9628) );
  INV_X1 U5743 ( .A(n9217), .ZN(n9162) );
  NAND2_X1 U5744 ( .A1(n5732), .A2(n5731), .ZN(n9659) );
  NAND2_X1 U5745 ( .A1(n5824), .A2(n5823), .ZN(n9669) );
  INV_X1 U5746 ( .A(n7990), .ZN(n10070) );
  INV_X1 U5747 ( .A(n5850), .ZN(n7313) );
  XNOR2_X1 U5748 ( .A(n5901), .B(n5900), .ZN(n8272) );
  XNOR2_X1 U5749 ( .A(n5832), .B(SI_29_), .ZN(n6351) );
  XNOR2_X1 U5750 ( .A(n5682), .B(n5681), .ZN(n8234) );
  INV_X1 U5751 ( .A(n5847), .ZN(n5843) );
  AOI21_X1 U5752 ( .B1(n4740), .B2(n4742), .A(n5471), .ZN(n4739) );
  NAND2_X1 U5753 ( .A1(n5450), .A2(n4743), .ZN(n4738) );
  OAI21_X1 U5754 ( .B1(n5450), .B2(n5449), .A(n5448), .ZN(n5466) );
  OR2_X1 U5755 ( .A1(n5800), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U5756 ( .A1(n4758), .A2(n5263), .ZN(n5280) );
  OR2_X1 U5757 ( .A1(n5785), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5788) );
  AOI21_X1 U5758 ( .B1(n5165), .B2(n4813), .A(n4499), .ZN(n4812) );
  AND2_X1 U5759 ( .A1(n5777), .A2(n5781), .ZN(n9845) );
  XNOR2_X1 U5760 ( .A(n4669), .B(P1_IR_REG_1__SCAN_IN), .ZN(n7092) );
  NAND2_X1 U5761 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4669) );
  NAND2_X1 U5762 ( .A1(n4937), .A2(n4934), .ZN(n7786) );
  NOR2_X1 U5763 ( .A1(n7764), .A2(n4942), .ZN(n7788) );
  OR2_X1 U5764 ( .A1(n6928), .A2(n8258), .ZN(n6929) );
  AND2_X1 U5765 ( .A1(n5407), .A2(n5406), .ZN(n8768) );
  AND4_X1 U5766 ( .A1(n5387), .A2(n5386), .A3(n5385), .A4(n5384), .ZN(n8721)
         );
  NAND2_X1 U5767 ( .A1(n5199), .A2(n5198), .ZN(n10286) );
  AOI21_X1 U5768 ( .B1(n6921), .B2(n8784), .A(n6847), .ZN(n7225) );
  OR2_X1 U5769 ( .A1(n6876), .A2(n6875), .ZN(n6877) );
  NAND2_X1 U5770 ( .A1(n8130), .A2(n8129), .ZN(n8128) );
  NOR2_X1 U5771 ( .A1(n6911), .A2(n8424), .ZN(n4908) );
  XNOR2_X1 U5772 ( .A(n6915), .B(n8611), .ZN(n8323) );
  NAND2_X1 U5773 ( .A1(n8408), .A2(n6886), .ZN(n8332) );
  NAND2_X1 U5774 ( .A1(n4929), .A2(n4927), .ZN(n7605) );
  NAND2_X1 U5775 ( .A1(n4930), .A2(n4473), .ZN(n4929) );
  AND2_X1 U5776 ( .A1(n7259), .A2(n4473), .ZN(n4928) );
  NAND2_X1 U5777 ( .A1(n4917), .A2(n4918), .ZN(n8343) );
  OR2_X1 U5778 ( .A1(n8408), .A2(n4921), .ZN(n4917) );
  NAND2_X1 U5779 ( .A1(n6910), .A2(n4912), .ZN(n4911) );
  NAND2_X1 U5780 ( .A1(n8303), .A2(n8637), .ZN(n4909) );
  XNOR2_X1 U5781 ( .A(n6912), .B(n8599), .ZN(n8351) );
  INV_X1 U5782 ( .A(n4930), .ZN(n4926) );
  AOI21_X1 U5783 ( .B1(n7854), .B2(n7855), .A(n4500), .ZN(n7878) );
  NAND2_X1 U5784 ( .A1(n7878), .A2(n7877), .ZN(n7876) );
  NAND2_X1 U5785 ( .A1(n8128), .A2(n6880), .ZN(n8370) );
  AND2_X1 U5786 ( .A1(n6946), .A2(n6945), .ZN(n8390) );
  AOI21_X1 U5787 ( .B1(n4915), .B2(n4921), .A(n4513), .ZN(n4913) );
  INV_X1 U5788 ( .A(n4937), .ZN(n7764) );
  AND2_X1 U5789 ( .A1(n6883), .A2(n8413), .ZN(n6884) );
  INV_X1 U5790 ( .A(n8390), .ZN(n8415) );
  INV_X1 U5791 ( .A(n8636), .ZN(n8667) );
  INV_X1 U5792 ( .A(n8413), .ZN(n8428) );
  INV_X1 U5793 ( .A(n6864), .ZN(n5211) );
  NAND4_X1 U5794 ( .A1(n5210), .A2(n5209), .A3(n5208), .A4(n5207), .ZN(n8433)
         );
  INV_X1 U5795 ( .A(n7681), .ZN(n8434) );
  NAND4_X1 U5796 ( .A1(n5144), .A2(n5143), .A3(n5142), .A4(n5141), .ZN(n8435)
         );
  NAND3_X1 U5797 ( .A1(n5120), .A2(n5119), .A3(n4991), .ZN(n8436) );
  AND2_X1 U5798 ( .A1(n5118), .A2(n5117), .ZN(n4991) );
  OR2_X1 U5799 ( .A1(n7169), .A2(n6966), .ZN(n8492) );
  XNOR2_X1 U5800 ( .A(n4585), .B(n4584), .ZN(n10122) );
  AOI21_X1 U5801 ( .B1(n10123), .B2(n10122), .A(n4583), .ZN(n7187) );
  AND2_X1 U5802 ( .A1(n4585), .A2(n10118), .ZN(n4583) );
  XNOR2_X1 U5803 ( .A(n7130), .B(n4781), .ZN(n7186) );
  INV_X1 U5804 ( .A(n4603), .ZN(n10142) );
  NAND2_X1 U5805 ( .A1(n4580), .A2(n4582), .ZN(n10158) );
  AOI21_X1 U5806 ( .B1(n8453), .B2(n4465), .A(n8452), .ZN(n8455) );
  XNOR2_X1 U5807 ( .A(n7660), .B(n7700), .ZN(n7690) );
  NAND2_X1 U5808 ( .A1(n7690), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7689) );
  AOI21_X1 U5809 ( .B1(n7693), .B2(n7652), .A(n7651), .ZN(n7724) );
  NAND2_X1 U5810 ( .A1(n4571), .A2(n4569), .ZN(n10168) );
  AND2_X1 U5811 ( .A1(n4571), .A2(n4575), .ZN(n10169) );
  OR2_X1 U5812 ( .A1(n7833), .A2(n4572), .ZN(n4571) );
  INV_X1 U5813 ( .A(n4796), .ZN(n10243) );
  AOI21_X1 U5814 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8523), .A(n8521), .ZN(
        n8522) );
  NAND2_X1 U5815 ( .A1(n8523), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4612) );
  AND2_X1 U5816 ( .A1(n8545), .A2(n5561), .ZN(n8560) );
  OAI21_X1 U5817 ( .B1(n8573), .B2(n8635), .A(n8572), .ZN(n8734) );
  INV_X1 U5818 ( .A(n8571), .ZN(n8572) );
  NAND2_X1 U5819 ( .A1(n5491), .A2(n5490), .ZN(n8744) );
  NAND2_X1 U5820 ( .A1(n4863), .A2(n6786), .ZN(n8614) );
  NAND2_X1 U5821 ( .A1(n8754), .A2(n4864), .ZN(n4863) );
  OAI21_X1 U5822 ( .B1(n5649), .B2(n6748), .A(n4854), .ZN(n8765) );
  NAND2_X1 U5823 ( .A1(n5254), .A2(n5253), .ZN(n10307) );
  NAND2_X1 U5824 ( .A1(n5233), .A2(n5232), .ZN(n10301) );
  AND3_X2 U5825 ( .A1(n5071), .A2(n5070), .A3(n5069), .ZN(n10256) );
  AND2_X1 U5826 ( .A1(n8563), .A2(n10308), .ZN(n5588) );
  OAI21_X1 U5827 ( .B1(n8597), .B2(n5517), .A(n5516), .ZN(n8588) );
  NAND2_X1 U5828 ( .A1(n4860), .A2(n4861), .ZN(n8595) );
  OR2_X1 U5829 ( .A1(n4862), .A2(n8754), .ZN(n4860) );
  NAND2_X1 U5830 ( .A1(n8754), .A2(n6778), .ZN(n8624) );
  OR2_X1 U5831 ( .A1(n8776), .A2(n8775), .ZN(n8837) );
  NAND2_X1 U5832 ( .A1(n5340), .A2(n5339), .ZN(n8339) );
  NAND2_X1 U5833 ( .A1(n5645), .A2(n6632), .ZN(n8155) );
  NAND2_X1 U5834 ( .A1(n5324), .A2(n5323), .ZN(n8405) );
  NAND2_X1 U5835 ( .A1(n5305), .A2(n5304), .ZN(n8300) );
  NAND2_X1 U5836 ( .A1(n4702), .A2(n4701), .ZN(n8047) );
  NAND2_X1 U5837 ( .A1(n5284), .A2(n5283), .ZN(n8377) );
  INV_X1 U5838 ( .A(n5641), .ZN(n8027) );
  OR2_X1 U5839 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  INV_X1 U5840 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7005) );
  NOR2_X1 U5841 ( .A1(n5080), .A2(n4945), .ZN(n5128) );
  XNOR2_X1 U5842 ( .A(n5100), .B(n5099), .ZN(n7385) );
  NAND2_X1 U5843 ( .A1(n5829), .A2(n5828), .ZN(n9640) );
  NAND2_X1 U5844 ( .A1(n5817), .A2(n5816), .ZN(n9763) );
  AOI21_X1 U5845 ( .B1(n8903), .B2(n6488), .A(n6487), .ZN(n8915) );
  NAND2_X1 U5846 ( .A1(n5730), .A2(n5729), .ZN(n9655) );
  NAND2_X1 U5847 ( .A1(n4829), .A2(n5790), .ZN(n10048) );
  INV_X1 U5848 ( .A(n4899), .ZN(n4897) );
  INV_X1 U5849 ( .A(n4902), .ZN(n4901) );
  AOI21_X1 U5850 ( .B1(n4868), .B2(n6487), .A(n4493), .ZN(n4866) );
  NOR2_X2 U5851 ( .A1(n6604), .A2(n6590), .ZN(n8968) );
  NAND2_X1 U5852 ( .A1(n4888), .A2(n4886), .ZN(n8896) );
  AND2_X1 U5853 ( .A1(n8897), .A2(n4887), .ZN(n4886) );
  NAND2_X1 U5854 ( .A1(n4890), .A2(n4893), .ZN(n4887) );
  AND2_X1 U5855 ( .A1(n6601), .A2(n8023), .ZN(n9796) );
  AND4_X1 U5856 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n7709)
         );
  AND4_X1 U5857 ( .A1(n6057), .A2(n6056), .A3(n6055), .A4(n6054), .ZN(n7476)
         );
  AND4_X1 U5858 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n7475)
         );
  OR2_X1 U5859 ( .A1(n5919), .A2(n6109), .ZN(n6112) );
  OR2_X1 U5860 ( .A1(n6102), .A2(n9494), .ZN(n6103) );
  OR2_X1 U5861 ( .A1(n4441), .A2(n6094), .ZN(n6098) );
  NAND2_X1 U5862 ( .A1(n6084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5863 ( .A1(n9078), .A2(n4656), .ZN(n9095) );
  NAND2_X1 U5864 ( .A1(n9190), .A2(n4983), .ZN(n9169) );
  NAND2_X1 U5865 ( .A1(n5726), .A2(n5725), .ZN(n9643) );
  NOR2_X1 U5866 ( .A1(n9231), .A2(n9131), .ZN(n9210) );
  NAND2_X1 U5867 ( .A1(n9574), .A2(n9154), .ZN(n9557) );
  NAND2_X1 U5868 ( .A1(n4810), .A2(n6231), .ZN(n8140) );
  NAND2_X1 U5869 ( .A1(n5822), .A2(n5821), .ZN(n8197) );
  NAND2_X1 U5870 ( .A1(n4965), .A2(n7974), .ZN(n7976) );
  NAND2_X1 U5871 ( .A1(n5810), .A2(n5809), .ZN(n8989) );
  NAND2_X1 U5872 ( .A1(n4816), .A2(n6295), .ZN(n7806) );
  NAND2_X1 U5873 ( .A1(n5750), .A2(n5749), .ZN(n8067) );
  NAND2_X1 U5874 ( .A1(n7532), .A2(n6292), .ZN(n7559) );
  NAND2_X1 U5875 ( .A1(n7564), .A2(n7563), .ZN(n4958) );
  NAND2_X1 U5876 ( .A1(n4827), .A2(n5787), .ZN(n7466) );
  INV_X1 U5877 ( .A(n10031), .ZN(n7524) );
  INV_X1 U5878 ( .A(n9623), .ZN(n9957) );
  NAND2_X1 U5879 ( .A1(n9690), .A2(n6594), .ZN(n9949) );
  INV_X1 U5880 ( .A(n9970), .ZN(n9599) );
  NAND2_X1 U5881 ( .A1(n9121), .A2(n5861), .ZN(n9627) );
  INV_X1 U5882 ( .A(n5860), .ZN(n5861) );
  OAI21_X1 U5883 ( .B1(n4636), .B2(n10076), .A(n9624), .ZN(n5860) );
  NOR2_X1 U5884 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4651) );
  OAI21_X1 U5885 ( .B1(n5901), .B2(n5900), .A(n5899), .ZN(n5906) );
  OAI21_X1 U5886 ( .B1(n5418), .B2(n5417), .A(n5416), .ZN(n5424) );
  NAND2_X1 U5887 ( .A1(n4554), .A2(n5145), .ZN(n4814) );
  INV_X1 U5888 ( .A(n7092), .ZN(n9807) );
  NAND2_X1 U5889 ( .A1(n4546), .A2(n6839), .ZN(P2_U3296) );
  NAND2_X1 U5890 ( .A1(n4547), .A2(n6836), .ZN(n4546) );
  AND2_X1 U5891 ( .A1(n4589), .A2(n8496), .ZN(n8519) );
  OAI21_X1 U5892 ( .B1(n8552), .B2(n8777), .A(n6366), .ZN(n6367) );
  AOI21_X1 U5893 ( .B1(n4726), .B2(n6371), .A(n6370), .ZN(n6372) );
  NOR2_X1 U5894 ( .A1(n10309), .A2(n6369), .ZN(n6370) );
  OAI21_X1 U5895 ( .B1(n6970), .B2(n8851), .A(n4779), .ZN(P2_U3293) );
  NOR2_X1 U5896 ( .A1(n8848), .A2(n6971), .ZN(n4780) );
  NOR2_X1 U5897 ( .A1(n6614), .A2(n6591), .ZN(n6612) );
  NOR2_X1 U5898 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  INV_X1 U5899 ( .A(n9063), .ZN(n9061) );
  NAND2_X1 U5900 ( .A1(n4562), .A2(n4523), .ZN(P1_U3517) );
  NAND2_X1 U5901 ( .A1(n9681), .A2(n10092), .ZN(n4562) );
  INV_X1 U5902 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n4561) );
  INV_X1 U5903 ( .A(n6801), .ZN(n8576) );
  AND2_X1 U5904 ( .A1(n6807), .A2(n6808), .ZN(n6801) );
  NAND2_X1 U5905 ( .A1(n9134), .A2(n4822), .ZN(n4818) );
  NAND2_X2 U5906 ( .A1(n5068), .A2(n5902), .ZN(n5107) );
  NAND2_X1 U5907 ( .A1(n5747), .A2(n5746), .ZN(n6021) );
  AOI21_X1 U5908 ( .B1(n8592), .B2(n5551), .A(n5531), .ZN(n8568) );
  INV_X1 U5909 ( .A(n4688), .ZN(n8630) );
  NOR2_X1 U5910 ( .A1(n5570), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n5568) );
  AND2_X1 U5911 ( .A1(n4754), .A2(n5181), .ZN(n4757) );
  AND2_X1 U5912 ( .A1(n4832), .A2(n9123), .ZN(n4452) );
  INV_X1 U5913 ( .A(n7361), .ZN(n4557) );
  INV_X1 U5914 ( .A(n6769), .ZN(n5650) );
  AND2_X1 U5915 ( .A1(n8768), .A2(n8693), .ZN(n6769) );
  XOR2_X1 U5916 ( .A(n6665), .B(n8535), .Z(n4453) );
  INV_X1 U5917 ( .A(n6632), .ZN(n4844) );
  INV_X1 U5918 ( .A(n6786), .ZN(n4540) );
  NOR2_X1 U5919 ( .A1(n5570), .A2(n4491), .ZN(n5026) );
  NAND2_X1 U5920 ( .A1(n5724), .A2(n5723), .ZN(n6269) );
  INV_X1 U5921 ( .A(n6269), .ZN(n4636) );
  AND2_X1 U5922 ( .A1(n4901), .A2(n8864), .ZN(n4454) );
  NAND2_X1 U5923 ( .A1(n4900), .A2(n4897), .ZN(n8935) );
  AND2_X1 U5924 ( .A1(n4828), .A2(n5790), .ZN(n4455) );
  NAND2_X1 U5925 ( .A1(n4595), .A2(n4597), .ZN(n5566) );
  OAI21_X1 U5926 ( .B1(n8867), .B2(n4893), .A(n4890), .ZN(n8895) );
  AND2_X1 U5927 ( .A1(n6179), .A2(n9125), .ZN(n9567) );
  OR2_X1 U5928 ( .A1(n4723), .A2(n6801), .ZN(n4456) );
  INV_X1 U5929 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4652) );
  OR2_X1 U5930 ( .A1(n4725), .A2(n8589), .ZN(n4457) );
  NOR2_X1 U5931 ( .A1(n8371), .A2(n4943), .ZN(n4458) );
  AND2_X1 U5932 ( .A1(n4972), .A2(n8198), .ZN(n4459) );
  OR2_X1 U5933 ( .A1(n8200), .A2(n9146), .ZN(n4460) );
  AND3_X1 U5934 ( .A1(n4770), .A2(n4774), .A3(n5394), .ZN(n4461) );
  OR2_X1 U5935 ( .A1(n8076), .A2(n8075), .ZN(n4462) );
  INV_X1 U5936 ( .A(n6383), .ZN(n6577) );
  INV_X2 U5937 ( .A(n6577), .ZN(n6552) );
  INV_X1 U5938 ( .A(n4441), .ZN(n6108) );
  INV_X1 U5939 ( .A(n7389), .ZN(n4789) );
  INV_X1 U5940 ( .A(n10260), .ZN(n6846) );
  NAND3_X1 U5941 ( .A1(n4977), .A2(n4974), .A3(n4652), .ZN(n4463) );
  INV_X1 U5942 ( .A(n6748), .ZN(n6760) );
  AND2_X1 U5943 ( .A1(n8774), .A2(n8425), .ZN(n6748) );
  NOR2_X1 U5944 ( .A1(n5204), .A2(n5203), .ZN(n4464) );
  OR2_X1 U5945 ( .A1(n7392), .A2(n7655), .ZN(n4465) );
  OR2_X1 U5946 ( .A1(n5910), .A2(n5909), .ZN(n5919) );
  NAND2_X1 U5947 ( .A1(n5437), .A2(n5436), .ZN(n5444) );
  NAND2_X1 U5948 ( .A1(n5908), .A2(n5907), .ZN(n6138) );
  NAND2_X1 U5949 ( .A1(n9162), .A2(n9161), .ZN(n9215) );
  AND3_X1 U5950 ( .A1(n5096), .A2(n5095), .A3(n5094), .ZN(n4466) );
  NAND4_X2 U5951 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n6849)
         );
  INV_X1 U5952 ( .A(n6184), .ZN(n6233) );
  OR2_X1 U5953 ( .A1(n5196), .A2(n4755), .ZN(n4467) );
  INV_X1 U5954 ( .A(n4996), .ZN(n7975) );
  AND2_X1 U5955 ( .A1(n6307), .A2(n6276), .ZN(n4996) );
  AND2_X1 U5956 ( .A1(n9127), .A2(n6243), .ZN(n9540) );
  INV_X1 U5957 ( .A(n9540), .ZN(n4622) );
  AND2_X1 U5958 ( .A1(n6780), .A2(n6777), .ZN(n8655) );
  AND3_X1 U5959 ( .A1(n9567), .A2(n9122), .A3(n6241), .ZN(n4468) );
  AND2_X1 U5960 ( .A1(n4783), .A2(n4782), .ZN(n4469) );
  NOR2_X1 U5961 ( .A1(n8127), .A2(n8430), .ZN(n4470) );
  OR2_X1 U5962 ( .A1(n5566), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4471) );
  OR2_X1 U5963 ( .A1(n5630), .A2(n5629), .ZN(n4472) );
  NAND2_X1 U5964 ( .A1(n4909), .A2(n4911), .ZN(n8350) );
  NAND2_X1 U5965 ( .A1(n6629), .A2(n6628), .ZN(n6657) );
  NOR2_X1 U5966 ( .A1(n4541), .A2(n4540), .ZN(n4539) );
  NAND2_X1 U5967 ( .A1(n6856), .A2(n7608), .ZN(n4473) );
  XNOR2_X1 U5968 ( .A(n6910), .B(n6911), .ZN(n8303) );
  OAI21_X1 U5969 ( .B1(n4838), .B2(n4761), .A(n4759), .ZN(n5299) );
  NAND2_X1 U5970 ( .A1(n5355), .A2(n5354), .ZN(n5374) );
  NAND2_X1 U5971 ( .A1(n4814), .A2(n5148), .ZN(n5166) );
  AND2_X1 U5972 ( .A1(n4850), .A2(n4851), .ZN(n4474) );
  AND2_X1 U5973 ( .A1(n6710), .A2(n6702), .ZN(n6638) );
  INV_X1 U5974 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5066) );
  INV_X1 U5975 ( .A(n6755), .ZN(n4843) );
  NAND2_X1 U5976 ( .A1(n5577), .A2(n5576), .ZN(n5068) );
  OR2_X1 U5977 ( .A1(n10198), .A2(n8471), .ZN(n4475) );
  NAND2_X1 U5978 ( .A1(n8864), .A2(n6527), .ZN(n8945) );
  NAND2_X1 U5979 ( .A1(n9575), .A2(n9579), .ZN(n9574) );
  NAND2_X1 U5980 ( .A1(n9557), .A2(n9556), .ZN(n9555) );
  NAND2_X1 U5981 ( .A1(n4889), .A2(n8929), .ZN(n8928) );
  AND2_X1 U5982 ( .A1(n4796), .A2(n4795), .ZN(n4476) );
  NAND2_X1 U5983 ( .A1(n4566), .A2(n4998), .ZN(n5098) );
  OR3_X1 U5984 ( .A1(n5566), .A2(P2_IR_REG_22__SCAN_IN), .A3(n4946), .ZN(n4477) );
  OR2_X1 U5985 ( .A1(n4789), .A2(n4791), .ZN(n4478) );
  INV_X1 U5986 ( .A(n8095), .ZN(n10064) );
  NAND2_X1 U5987 ( .A1(n5799), .A2(n5798), .ZN(n8095) );
  NAND2_X1 U5988 ( .A1(n5178), .A2(n9390), .ZN(n5181) );
  OAI21_X1 U5989 ( .B1(n6264), .B2(n6269), .A(n4640), .ZN(n4639) );
  AND2_X1 U5990 ( .A1(n5271), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5991 ( .A1(n5644), .A2(n4835), .ZN(n8105) );
  AND2_X1 U5992 ( .A1(n9188), .A2(n9166), .ZN(n4480) );
  INV_X1 U5993 ( .A(n4676), .ZN(n9202) );
  AND2_X1 U5994 ( .A1(n8217), .A2(n4677), .ZN(n4481) );
  OR2_X1 U5995 ( .A1(n9649), .A2(n8971), .ZN(n9130) );
  INV_X1 U5996 ( .A(n7362), .ZN(n7118) );
  NAND2_X1 U5997 ( .A1(n6123), .A2(n6122), .ZN(n7362) );
  AND2_X1 U5998 ( .A1(n4988), .A2(n4905), .ZN(n4482) );
  AND2_X1 U5999 ( .A1(n4729), .A2(n6812), .ZN(n4483) );
  AND2_X1 U6000 ( .A1(n4729), .A2(n6348), .ZN(n4484) );
  AND2_X1 U6001 ( .A1(n9197), .A2(n9164), .ZN(n4485) );
  NAND2_X1 U6002 ( .A1(n6189), .A2(n6193), .ZN(n4486) );
  INV_X1 U6003 ( .A(n4621), .ZN(n4620) );
  OAI21_X1 U6004 ( .B1(n6242), .B2(n4622), .A(n6244), .ZN(n4621) );
  AND2_X1 U6005 ( .A1(n4900), .A2(n4898), .ZN(n4487) );
  AND2_X1 U6006 ( .A1(n4636), .A2(n4638), .ZN(n4488) );
  OR2_X1 U6007 ( .A1(n7098), .A2(n7097), .ZN(n4489) );
  NOR2_X1 U6008 ( .A1(n6787), .A2(n4865), .ZN(n4864) );
  OR2_X1 U6009 ( .A1(n6769), .A2(n6748), .ZN(n4490) );
  NAND2_X1 U6010 ( .A1(n6262), .A2(n6263), .ZN(n9168) );
  INV_X1 U6011 ( .A(n9168), .ZN(n4638) );
  INV_X1 U6012 ( .A(n9122), .ZN(n9579) );
  AND2_X1 U6013 ( .A1(n9565), .A2(n6146), .ZN(n9122) );
  INV_X1 U6014 ( .A(n6813), .ZN(n6656) );
  AND2_X1 U6015 ( .A1(n8552), .A2(n8421), .ZN(n6813) );
  INV_X1 U6016 ( .A(n6874), .ZN(n4704) );
  INV_X1 U6017 ( .A(n4723), .ZN(n4722) );
  OR2_X1 U6018 ( .A1(n5532), .A2(n4724), .ZN(n4723) );
  OR2_X1 U6019 ( .A1(n4947), .A2(n4596), .ZN(n4491) );
  OR2_X1 U6020 ( .A1(n4947), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4492) );
  NOR2_X1 U6021 ( .A1(n6493), .A2(n6492), .ZN(n4493) );
  NAND2_X1 U6022 ( .A1(n6460), .A2(n6459), .ZN(n4494) );
  OR2_X1 U6023 ( .A1(n5835), .A2(n5713), .ZN(n4495) );
  NAND2_X1 U6024 ( .A1(n5658), .A2(n8264), .ZN(n4496) );
  AND2_X1 U6025 ( .A1(n4738), .A2(n4740), .ZN(n4497) );
  INV_X1 U6026 ( .A(n4670), .ZN(n9174) );
  NOR3_X1 U6027 ( .A1(n9213), .A2(n9640), .A3(n4671), .ZN(n4670) );
  AND2_X1 U6028 ( .A1(n6424), .A2(n7472), .ZN(n4498) );
  AND2_X1 U6029 ( .A1(n5168), .A2(SI_6_), .ZN(n4499) );
  XNOR2_X1 U6030 ( .A(n5277), .B(SI_12_), .ZN(n5276) );
  INV_X1 U6031 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7000) );
  AND2_X1 U6032 ( .A1(n6863), .A2(n6862), .ZN(n4500) );
  INV_X1 U6033 ( .A(n4904), .ZN(n6514) );
  NAND2_X1 U6034 ( .A1(n6245), .A2(n9130), .ZN(n4501) );
  INV_X1 U6035 ( .A(n9134), .ZN(n9197) );
  AND2_X1 U6036 ( .A1(n6250), .A2(n9135), .ZN(n9134) );
  INV_X1 U6037 ( .A(n8438), .ZN(n6852) );
  OR2_X1 U6038 ( .A1(n10307), .A2(n8134), .ZN(n6721) );
  INV_X1 U6039 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U6040 ( .A1(n9216), .A2(n9130), .ZN(n4823) );
  AND2_X1 U6041 ( .A1(n9004), .A2(n6564), .ZN(n4502) );
  NAND2_X1 U6042 ( .A1(n7142), .A2(n5066), .ZN(n5080) );
  INV_X1 U6043 ( .A(n5080), .ZN(n4566) );
  AND2_X1 U6044 ( .A1(n6826), .A2(n6804), .ZN(n4503) );
  NAND2_X1 U6045 ( .A1(n4811), .A2(n4812), .ZN(n5173) );
  NOR2_X1 U6046 ( .A1(n6102), .A2(n9933), .ZN(n4504) );
  NOR2_X1 U6047 ( .A1(n8095), .A2(n7715), .ZN(n4505) );
  NAND2_X1 U6048 ( .A1(n8127), .A2(n8430), .ZN(n4506) );
  AND2_X1 U6049 ( .A1(n4605), .A2(n4604), .ZN(n4507) );
  NAND2_X1 U6050 ( .A1(n6812), .A2(n8422), .ZN(n4508) );
  OR2_X1 U6051 ( .A1(n5566), .A2(n4492), .ZN(n4509) );
  INV_X1 U6052 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9356) );
  INV_X1 U6053 ( .A(n6795), .ZN(n6630) );
  AND2_X1 U6054 ( .A1(n8809), .A2(n8611), .ZN(n6795) );
  INV_X1 U6055 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6972) );
  NAND2_X1 U6056 ( .A1(n4914), .A2(n4913), .ZN(n8310) );
  OAI22_X1 U6057 ( .A1(n5649), .A2(n4490), .B1(n4854), .B2(n6769), .ZN(n8648)
         );
  AND2_X1 U6058 ( .A1(n4579), .A2(n4582), .ZN(n4510) );
  NAND2_X1 U6059 ( .A1(n4965), .A2(n4963), .ZN(n8074) );
  AND4_X1 U6060 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n7931)
         );
  INV_X1 U6061 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n4661) );
  INV_X1 U6062 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4559) );
  INV_X1 U6063 ( .A(n6313), .ZN(n4649) );
  NAND2_X1 U6064 ( .A1(n6901), .A2(n6900), .ZN(n8278) );
  INV_X1 U6065 ( .A(n4741), .ZN(n4740) );
  OAI21_X1 U6066 ( .B1(n5445), .B2(n4742), .A(n5464), .ZN(n4741) );
  NAND2_X1 U6067 ( .A1(n4867), .A2(n4866), .ZN(n8956) );
  NAND2_X1 U6068 ( .A1(n4462), .A2(n8144), .ZN(n8196) );
  NAND2_X1 U6069 ( .A1(n9148), .A2(n9147), .ZN(n9610) );
  INV_X1 U6070 ( .A(n4870), .ZN(n8061) );
  XNOR2_X1 U6071 ( .A(n6920), .B(n8598), .ZN(n8395) );
  INV_X1 U6072 ( .A(n8395), .ZN(n4925) );
  NAND2_X1 U6073 ( .A1(n5734), .A2(n5733), .ZN(n9674) );
  NAND2_X1 U6074 ( .A1(n5545), .A2(n5544), .ZN(n8735) );
  INV_X1 U6075 ( .A(n8735), .ZN(n4725) );
  AND4_X1 U6076 ( .A1(n5370), .A2(n5369), .A3(n5368), .A4(n5367), .ZN(n8334)
         );
  AND2_X1 U6077 ( .A1(n9649), .A2(n9159), .ZN(n4511) );
  INV_X1 U6078 ( .A(n4680), .ZN(n9611) );
  NOR3_X1 U6079 ( .A1(n8200), .A2(n9146), .A3(n9674), .ZN(n4680) );
  NOR2_X1 U6080 ( .A1(n10176), .A2(n8468), .ZN(n4512) );
  INV_X1 U6081 ( .A(n8037), .ZN(n8429) );
  AND4_X1 U6082 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n8037)
         );
  AND2_X1 U6083 ( .A1(n6889), .A2(n8334), .ZN(n4513) );
  AND2_X1 U6084 ( .A1(n6546), .A2(n6545), .ZN(n8929) );
  INV_X1 U6085 ( .A(n8929), .ZN(n4893) );
  INV_X1 U6086 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n4684) );
  AND2_X1 U6087 ( .A1(n8405), .A2(n8427), .ZN(n4514) );
  INV_X1 U6088 ( .A(n4743), .ZN(n4742) );
  NOR2_X1 U6089 ( .A1(n5465), .A2(n4744), .ZN(n4743) );
  AND2_X1 U6090 ( .A1(n5481), .A2(n5480), .ZN(n8637) );
  NAND2_X1 U6091 ( .A1(n5831), .A2(n5830), .ZN(n9633) );
  INV_X1 U6092 ( .A(n9633), .ZN(n4674) );
  NOR2_X1 U6093 ( .A1(n9659), .A2(n9155), .ZN(n4515) );
  AND2_X1 U6094 ( .A1(n8772), .A2(n6760), .ZN(n4516) );
  AND2_X1 U6095 ( .A1(n5335), .A2(SI_15_), .ZN(n4517) );
  INV_X1 U6096 ( .A(n4771), .ZN(n4770) );
  NAND2_X1 U6097 ( .A1(n5423), .A2(n4772), .ZN(n4771) );
  INV_X1 U6098 ( .A(n4726), .ZN(n8552) );
  NAND2_X1 U6099 ( .A1(n6353), .A2(n6352), .ZN(n4726) );
  OR2_X1 U6100 ( .A1(n8200), .A2(n4681), .ZN(n4518) );
  NAND2_X1 U6101 ( .A1(n5525), .A2(n5524), .ZN(n8803) );
  AND2_X1 U6102 ( .A1(n7451), .A2(n7449), .ZN(n6195) );
  AND4_X1 U6103 ( .A1(n6049), .A2(n6048), .A3(n6047), .A4(n6046), .ZN(n7544)
         );
  INV_X1 U6104 ( .A(n7544), .ZN(n4828) );
  OR2_X1 U6105 ( .A1(n8300), .A2(n8428), .ZN(n4519) );
  INV_X1 U6106 ( .A(n5394), .ZN(n4767) );
  AND2_X1 U6107 ( .A1(n9078), .A2(n9077), .ZN(n4520) );
  INV_X1 U6109 ( .A(n10325), .ZN(n10323) );
  NAND2_X1 U6110 ( .A1(n7568), .A2(n10064), .ZN(n7567) );
  NAND2_X1 U6111 ( .A1(n7568), .A2(n4677), .ZN(n4521) );
  NOR2_X1 U6112 ( .A1(n7833), .A2(n4576), .ZN(n4522) );
  OR2_X1 U6113 ( .A1(n10092), .A2(n4561), .ZN(n4523) );
  NAND2_X1 U6114 ( .A1(n7304), .A2(n6420), .ZN(n7471) );
  NAND2_X1 U6115 ( .A1(n5222), .A2(n5221), .ZN(n7942) );
  NAND2_X1 U6116 ( .A1(n4958), .A2(n7566), .ZN(n7714) );
  INV_X1 U6117 ( .A(n7775), .ZN(n4877) );
  OR2_X1 U6118 ( .A1(n4942), .A2(n4939), .ZN(n4938) );
  INV_X1 U6119 ( .A(n4938), .ZN(n4934) );
  INV_X1 U6120 ( .A(n8482), .ZN(n4575) );
  AND2_X1 U6121 ( .A1(n4926), .A2(n7258), .ZN(n4524) );
  NOR2_X1 U6122 ( .A1(n8483), .A2(n8506), .ZN(n4525) );
  OR2_X1 U6123 ( .A1(n7417), .A2(n7414), .ZN(n4526) );
  OR2_X1 U6124 ( .A1(n4656), .A2(n4655), .ZN(n4527) );
  AND2_X1 U6125 ( .A1(n7836), .A2(n8504), .ZN(n4528) );
  AND2_X1 U6126 ( .A1(n4950), .A2(n4949), .ZN(n7325) );
  XOR2_X1 U6127 ( .A(n8526), .B(P2_REG1_REG_19__SCAN_IN), .Z(n4529) );
  AND2_X1 U6128 ( .A1(n10144), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4530) );
  AND2_X1 U6129 ( .A1(n4792), .A2(n10144), .ZN(n4531) );
  AND2_X1 U6130 ( .A1(n4603), .A2(n4602), .ZN(n4532) );
  INV_X1 U6131 ( .A(n9716), .ZN(n4662) );
  INV_X1 U6132 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4685) );
  XNOR2_X1 U6133 ( .A(n5032), .B(n5031), .ZN(n10118) );
  INV_X1 U6134 ( .A(n10118), .ZN(n4584) );
  AOI21_X1 U6135 ( .B1(n9142), .B2(n9947), .A(n9141), .ZN(n9630) );
  NAND2_X1 U6136 ( .A1(n7007), .A2(n5722), .ZN(n4827) );
  NAND2_X1 U6137 ( .A1(n6790), .A2(n6789), .ZN(n4535) );
  NAND2_X1 U6138 ( .A1(n4537), .A2(n6788), .ZN(n4536) );
  NAND2_X1 U6139 ( .A1(n4538), .A2(n6792), .ZN(n4537) );
  OAI21_X2 U6140 ( .B1(n6790), .B2(n6787), .A(n4539), .ZN(n4538) );
  INV_X1 U6141 ( .A(n6791), .ZN(n4541) );
  NAND2_X1 U6142 ( .A1(n5084), .A2(n5083), .ZN(n4545) );
  NAND2_X1 U6143 ( .A1(n4543), .A2(n5084), .ZN(n4542) );
  INV_X1 U6144 ( .A(n5083), .ZN(n4544) );
  NAND2_X1 U6145 ( .A1(n4545), .A2(n5087), .ZN(n5102) );
  OAI211_X1 U6146 ( .C1(n6835), .C2(n6844), .A(n4549), .B(n4548), .ZN(n4547)
         );
  NAND2_X1 U6147 ( .A1(n6835), .A2(n7500), .ZN(n4549) );
  NAND2_X2 U6148 ( .A1(n4552), .A2(n5425), .ZN(n8832) );
  NAND2_X1 U6149 ( .A1(n4734), .A2(n4554), .ZN(n4811) );
  XNOR2_X1 U6150 ( .A(n4554), .B(n5145), .ZN(n6992) );
  AND2_X4 U6151 ( .A1(n4802), .A2(n4801), .ZN(n5065) );
  INV_X1 U6152 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4555) );
  OAI21_X1 U6153 ( .B1(n5065), .B2(P2_DATAO_REG_3__SCAN_IN), .A(n4558), .ZN(
        n5103) );
  NAND2_X1 U6154 ( .A1(n5065), .A2(n4559), .ZN(n4558) );
  MUX2_X1 U6155 ( .A(n7744), .B(n7745), .S(n5065), .Z(n5398) );
  NAND2_X1 U6156 ( .A1(n4944), .A2(n4566), .ZN(n5149) );
  NAND2_X1 U6157 ( .A1(n7833), .A2(n4569), .ZN(n4568) );
  AND2_X1 U6158 ( .A1(n7834), .A2(n7835), .ZN(n4576) );
  NAND2_X1 U6159 ( .A1(n10130), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U6160 ( .A1(n4606), .A2(n4507), .ZN(n4600) );
  NAND2_X1 U6161 ( .A1(n4600), .A2(n4601), .ZN(n7654) );
  OAI21_X1 U6162 ( .B1(n4611), .B2(n10235), .A(n4607), .ZN(n4608) );
  NAND2_X1 U6163 ( .A1(n10235), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10234) );
  NAND2_X1 U6164 ( .A1(n4608), .A2(n4612), .ZN(n4609) );
  NAND2_X1 U6165 ( .A1(n10234), .A2(n8515), .ZN(n8525) );
  XNOR2_X1 U6166 ( .A(n4609), .B(n4529), .ZN(n8539) );
  NOR2_X1 U6167 ( .A1(n7404), .A2(n4624), .ZN(n4623) );
  NAND2_X1 U6168 ( .A1(n7347), .A2(n6192), .ZN(n7515) );
  NAND2_X1 U6169 ( .A1(n6269), .A2(n6266), .ZN(n4640) );
  INV_X1 U6170 ( .A(n4984), .ZN(n4641) );
  NAND2_X1 U6171 ( .A1(n6208), .A2(n7451), .ZN(n6209) );
  NAND4_X1 U6172 ( .A1(n6236), .A2(n9591), .A3(n6266), .A4(n6235), .ZN(n4650)
         );
  NAND3_X1 U6173 ( .A1(n4977), .A2(n4651), .A3(n4974), .ZN(n9693) );
  NAND2_X1 U6174 ( .A1(n4977), .A2(n4974), .ZN(n5720) );
  OR2_X1 U6175 ( .A1(n9071), .A2(n4654), .ZN(n4653) );
  NAND2_X1 U6176 ( .A1(n4653), .A2(n4527), .ZN(n9916) );
  MUX2_X1 U6177 ( .A(n9441), .B(P1_REG2_REG_1__SCAN_IN), .S(n7092), .Z(n9803)
         );
  NAND2_X1 U6178 ( .A1(n8666), .A2(n4687), .ZN(n4686) );
  NAND2_X1 U6179 ( .A1(n4692), .A2(n4695), .ZN(n5390) );
  NAND2_X1 U6180 ( .A1(n8160), .A2(n4693), .ZN(n4692) );
  INV_X1 U6181 ( .A(n5296), .ZN(n4706) );
  NAND3_X1 U6182 ( .A1(n4702), .A2(n4701), .A3(n4519), .ZN(n5313) );
  MUX2_X1 U6183 ( .A(n6788), .B(n6675), .S(n6674), .Z(n6680) );
  MUX2_X2 U6184 ( .A(n6785), .B(n6784), .S(n6959), .Z(n6790) );
  AOI21_X1 U6185 ( .B1(n6742), .B2(n6741), .A(n8104), .ZN(n6754) );
  OAI21_X1 U6186 ( .B1(n6670), .B2(n7853), .A(n6959), .ZN(n6673) );
  OAI211_X1 U6187 ( .C1(n6802), .C2(n8587), .A(n6801), .B(n6800), .ZN(n6810)
         );
  OAI21_X2 U6188 ( .B1(n6683), .B2(n6682), .A(n6681), .ZN(n6692) );
  INV_X1 U6189 ( .A(n6701), .ZN(n6719) );
  AOI21_X1 U6190 ( .B1(n6272), .B2(n6374), .A(n6271), .ZN(n6273) );
  NAND2_X2 U6191 ( .A1(n5910), .A2(n5909), .ZN(n6102) );
  OAI21_X1 U6192 ( .B1(n6333), .B2(n6593), .A(n6332), .ZN(n6345) );
  MUX2_X2 U6193 ( .A(n6700), .B(n6699), .S(n6959), .Z(n6701) );
  NAND2_X1 U6194 ( .A1(n6816), .A2(n6815), .ZN(n6817) );
  AOI21_X1 U6195 ( .B1(n6719), .B2(n6718), .A(n6717), .ZN(n6728) );
  OR2_X2 U6196 ( .A1(n5754), .A2(n5037), .ZN(n5751) );
  OR2_X2 U6197 ( .A1(n7334), .A2(n10014), .ZN(n7335) );
  NAND2_X1 U6198 ( .A1(n4977), .A2(n4976), .ZN(n5717) );
  NAND2_X1 U6199 ( .A1(n4726), .A2(n6354), .ZN(n6804) );
  NAND2_X1 U6200 ( .A1(n5534), .A2(n5533), .ZN(n5536) );
  NAND2_X1 U6201 ( .A1(n5519), .A2(n5518), .ZN(n4727) );
  NAND2_X1 U6202 ( .A1(n4728), .A2(n4729), .ZN(n6819) );
  INV_X1 U6203 ( .A(n4731), .ZN(n4728) );
  OAI21_X1 U6204 ( .B1(n5902), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4733), .ZN(
        n5146) );
  NAND2_X1 U6205 ( .A1(n5902), .A2(n5127), .ZN(n4733) );
  NAND2_X1 U6206 ( .A1(n5450), .A2(n4739), .ZN(n4737) );
  OAI21_X1 U6207 ( .B1(n5450), .B2(n4741), .A(n4739), .ZN(n5486) );
  NAND2_X1 U6208 ( .A1(n4751), .A2(n4750), .ZN(n4754) );
  NAND2_X1 U6209 ( .A1(n5173), .A2(n5172), .ZN(n4756) );
  NAND3_X1 U6210 ( .A1(n4753), .A2(n5223), .A3(n4752), .ZN(n5226) );
  NAND2_X1 U6211 ( .A1(n5173), .A2(n4757), .ZN(n4753) );
  NAND2_X1 U6212 ( .A1(n4756), .A2(n5176), .ZN(n5197) );
  NAND2_X1 U6213 ( .A1(n4838), .A2(n4762), .ZN(n4758) );
  INV_X1 U6214 ( .A(n5374), .ZN(n4775) );
  XNOR2_X1 U6215 ( .A(n7392), .B(n7396), .ZN(n7393) );
  AND2_X1 U6216 ( .A1(n4777), .A2(n4776), .ZN(n10209) );
  NAND2_X1 U6217 ( .A1(n10208), .A2(n10207), .ZN(n4776) );
  INV_X1 U6218 ( .A(n10208), .ZN(n4778) );
  OR2_X1 U6219 ( .A1(n7202), .A2(n7582), .ZN(n7157) );
  OR2_X1 U6220 ( .A1(n7202), .A2(n7141), .ZN(n7148) );
  AOI21_X1 U6221 ( .B1(n7202), .B2(P2_STATE_REG_SCAN_IN), .A(n4780), .ZN(n4779) );
  NAND2_X1 U6222 ( .A1(n5405), .A2(n7202), .ZN(n5069) );
  INV_X1 U6223 ( .A(n7202), .ZN(n4781) );
  XNOR2_X2 U6224 ( .A(n5067), .B(P2_IR_REG_2__SCAN_IN), .ZN(n7202) );
  INV_X1 U6225 ( .A(n4785), .ZN(n7635) );
  INV_X1 U6226 ( .A(n4783), .ZN(n7734) );
  OR2_X1 U6227 ( .A1(n7691), .A2(n7633), .ZN(n4785) );
  OAI21_X1 U6228 ( .B1(n7388), .B2(n4790), .A(n4786), .ZN(n10143) );
  INV_X1 U6229 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4791) );
  NAND2_X1 U6230 ( .A1(n8476), .A2(n4797), .ZN(n4793) );
  OR2_X1 U6231 ( .A1(n10244), .A2(n8478), .ZN(n4796) );
  NAND2_X1 U6232 ( .A1(n8468), .A2(n4800), .ZN(n4798) );
  NAND3_X1 U6233 ( .A1(n4802), .A2(P1_DATAO_REG_0__SCAN_IN), .A3(n4801), .ZN(
        n5033) );
  NAND2_X1 U6234 ( .A1(n5101), .A2(n4806), .ZN(n4805) );
  NAND2_X1 U6235 ( .A1(n5122), .A2(n5121), .ZN(n5126) );
  OAI21_X1 U6236 ( .B1(n9231), .B2(n4823), .A(n9132), .ZN(n4824) );
  NAND2_X1 U6237 ( .A1(n7029), .A2(n5722), .ZN(n4829) );
  NAND2_X1 U6238 ( .A1(n6168), .A2(n4834), .ZN(n4833) );
  NAND2_X1 U6239 ( .A1(n5226), .A2(n5225), .ZN(n5245) );
  NAND2_X1 U6240 ( .A1(n5226), .A2(n4839), .ZN(n4838) );
  OAI21_X1 U6241 ( .B1(n8105), .B2(n4842), .A(n4841), .ZN(n5647) );
  OAI21_X1 U6242 ( .B1(n5645), .B2(n6743), .A(n4846), .ZN(n8710) );
  NAND3_X1 U6243 ( .A1(n4857), .A2(n4856), .A3(n6630), .ZN(n5655) );
  NAND2_X1 U6244 ( .A1(n4861), .A2(n8754), .ZN(n4857) );
  NAND2_X1 U6245 ( .A1(n8903), .A2(n4868), .ZN(n4867) );
  OAI21_X1 U6246 ( .B1(n7774), .B2(n4879), .A(n4875), .ZN(n7983) );
  OAI21_X1 U6247 ( .B1(n7774), .B2(n4874), .A(n4871), .ZN(n4870) );
  NAND2_X1 U6248 ( .A1(n4878), .A2(n7984), .ZN(n4874) );
  OAI21_X1 U6249 ( .B1(n7774), .B2(n7776), .A(n7775), .ZN(n7953) );
  NAND2_X1 U6250 ( .A1(n6448), .A2(n4880), .ZN(n4879) );
  NAND2_X1 U6251 ( .A1(n8867), .A2(n4890), .ZN(n4888) );
  NAND2_X1 U6252 ( .A1(n8867), .A2(n8930), .ZN(n4889) );
  NAND2_X1 U6253 ( .A1(n8878), .A2(n4898), .ZN(n4896) );
  NAND2_X1 U6254 ( .A1(n4902), .A2(n8864), .ZN(n6536) );
  NAND2_X1 U6255 ( .A1(n4904), .A2(n4447), .ZN(n6396) );
  AOI22_X1 U6256 ( .A1(n4904), .A2(n7271), .B1(n7272), .B2(n6564), .ZN(n6391)
         );
  AOI22_X1 U6257 ( .A1(n10014), .A2(n4904), .B1(n9005), .B2(n6564), .ZN(n6410)
         );
  AOI22_X1 U6258 ( .A1(n7361), .A2(n4903), .B1(n7362), .B2(n6564), .ZN(n6414)
         );
  NAND2_X1 U6259 ( .A1(n10048), .A2(n4903), .ZN(n6435) );
  AOI21_X1 U6260 ( .B1(n7524), .B2(n4903), .A(n4502), .ZN(n6421) );
  NAND2_X1 U6261 ( .A1(n7961), .A2(n4903), .ZN(n6444) );
  NAND2_X1 U6262 ( .A1(n8095), .A2(n4903), .ZN(n6441) );
  NAND2_X1 U6263 ( .A1(n7990), .A2(n4903), .ZN(n6455) );
  NAND2_X1 U6264 ( .A1(n8067), .A2(n4903), .ZN(n6462) );
  NAND2_X1 U6265 ( .A1(n6021), .A2(n4903), .ZN(n6468) );
  NAND2_X1 U6266 ( .A1(n8989), .A2(n4903), .ZN(n6480) );
  NAND2_X1 U6267 ( .A1(n8921), .A2(n4903), .ZN(n6490) );
  NAND2_X1 U6268 ( .A1(n9146), .A2(n4903), .ZN(n6499) );
  NAND2_X1 U6269 ( .A1(n9669), .A2(n4903), .ZN(n6512) );
  NAND2_X1 U6270 ( .A1(n9659), .A2(n4903), .ZN(n6530) );
  NAND2_X1 U6271 ( .A1(n9655), .A2(n4903), .ZN(n6538) );
  NAND2_X1 U6272 ( .A1(n9649), .A2(n4903), .ZN(n6548) );
  NAND2_X1 U6273 ( .A1(n9643), .A2(n4903), .ZN(n6551) );
  NAND2_X1 U6274 ( .A1(n9640), .A2(n4903), .ZN(n6561) );
  NAND2_X1 U6275 ( .A1(n9633), .A2(n4903), .ZN(n6576) );
  NAND2_X1 U6276 ( .A1(n5839), .A2(n4988), .ZN(n5845) );
  NAND2_X1 U6277 ( .A1(n5020), .A2(n8847), .ZN(n5206) );
  NAND2_X1 U6278 ( .A1(n8847), .A2(n8242), .ZN(n5072) );
  INV_X1 U6279 ( .A(n6911), .ZN(n4912) );
  NAND2_X1 U6280 ( .A1(n8408), .A2(n4915), .ZN(n4914) );
  NAND2_X1 U6281 ( .A1(n6918), .A2(n6917), .ZN(n8394) );
  NAND2_X1 U6282 ( .A1(n7260), .A2(n7259), .ZN(n7258) );
  NAND2_X1 U6283 ( .A1(n7260), .A2(n4928), .ZN(n4927) );
  NAND2_X1 U6284 ( .A1(n7258), .A2(n4932), .ZN(n7484) );
  NAND2_X1 U6285 ( .A1(n4932), .A2(n4931), .ZN(n4930) );
  INV_X1 U6286 ( .A(n7485), .ZN(n4931) );
  NAND2_X1 U6287 ( .A1(n7765), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U6288 ( .A1(n4933), .A2(n4935), .ZN(n7854) );
  AND2_X1 U6289 ( .A1(n6858), .A2(n8435), .ZN(n4942) );
  NAND2_X1 U6290 ( .A1(n8128), .A2(n4458), .ZN(n8368) );
  NOR2_X2 U6291 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5756) );
  OAI21_X2 U6292 ( .B1(n9225), .B2(n4511), .A(n9160), .ZN(n9217) );
  NAND2_X1 U6293 ( .A1(n4951), .A2(n4949), .ZN(n7274) );
  NAND2_X1 U6294 ( .A1(n4440), .A2(n7273), .ZN(n4949) );
  NAND2_X1 U6295 ( .A1(n4951), .A2(n9961), .ZN(n4950) );
  INV_X1 U6296 ( .A(n7273), .ZN(n4952) );
  NAND2_X1 U6297 ( .A1(n4954), .A2(n7326), .ZN(n9953) );
  NAND2_X1 U6298 ( .A1(n7325), .A2(n7324), .ZN(n4954) );
  NAND2_X1 U6299 ( .A1(n4956), .A2(n4955), .ZN(n7815) );
  AOI21_X1 U6300 ( .B1(n7713), .B2(n4957), .A(n4505), .ZN(n4955) );
  NAND3_X1 U6301 ( .A1(n7564), .A2(n7563), .A3(n7713), .ZN(n4956) );
  NAND2_X1 U6302 ( .A1(n9575), .A2(n4960), .ZN(n4959) );
  NAND2_X1 U6303 ( .A1(n9148), .A2(n4967), .ZN(n4966) );
  NOR2_X1 U6304 ( .A1(n5713), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4976) );
  INV_X2 U6305 ( .A(n5835), .ZN(n4977) );
  AND2_X1 U6306 ( .A1(n9193), .A2(n9166), .ZN(n9189) );
  OAI21_X1 U6307 ( .B1(n5065), .B2(n5037), .A(n5036), .ZN(n5061) );
  NAND2_X1 U6308 ( .A1(n5065), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U6309 ( .A1(n8886), .A2(n8887), .ZN(n8885) );
  OR2_X1 U6310 ( .A1(n5072), .A2(n5042), .ZN(n5047) );
  NAND4_X1 U6311 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5625)
         );
  OAI21_X1 U6312 ( .B1(n6364), .B2(n8635), .A(n6363), .ZN(n8551) );
  AND2_X1 U6313 ( .A1(n6721), .A2(n6722), .ZN(n7929) );
  AND4_X4 U6314 ( .A1(n5079), .A2(n5078), .A3(n5077), .A4(n5076), .ZN(n7622)
         );
  OR2_X1 U6315 ( .A1(n6356), .A2(n5075), .ZN(n5076) );
  AOI21_X1 U6316 ( .B1(n8550), .B2(n7944), .A(n6362), .ZN(n6363) );
  OR2_X1 U6317 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  XNOR2_X1 U6318 ( .A(n9007), .B(n9999), .ZN(n7323) );
  AOI21_X2 U6319 ( .B1(n7242), .B2(n7244), .A(n7241), .ZN(n7305) );
  NAND2_X1 U6320 ( .A1(n5035), .A2(SI_0_), .ZN(n5060) );
  NOR2_X1 U6321 ( .A1(n6526), .A2(n6525), .ZN(n4978) );
  INV_X1 U6322 ( .A(n8839), .ZN(n6371) );
  AND2_X1 U6323 ( .A1(n5623), .A2(n5622), .ZN(n10311) );
  NOR2_X1 U6324 ( .A1(n8262), .A2(n8261), .ZN(n4979) );
  OR2_X1 U6325 ( .A1(n6983), .A2(n9807), .ZN(n4980) );
  OR2_X1 U6326 ( .A1(n10092), .A2(n5897), .ZN(n4981) );
  AND2_X1 U6327 ( .A1(n6391), .A2(n6577), .ZN(n4982) );
  OR2_X1 U6328 ( .A1(n4674), .A2(n9167), .ZN(n4983) );
  NAND2_X1 U6329 ( .A1(n6138), .A2(n6139), .ZN(n4984) );
  XNOR2_X1 U6330 ( .A(n5060), .B(n5061), .ZN(n5059) );
  AND2_X1 U6331 ( .A1(n6413), .A2(n6412), .ZN(n4985) );
  AND2_X1 U6332 ( .A1(n6118), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n4987) );
  AND3_X1 U6333 ( .A1(n5838), .A2(n5837), .A3(n5836), .ZN(n4988) );
  AND2_X1 U6334 ( .A1(n7473), .A2(n6423), .ZN(n6422) );
  OR2_X1 U6335 ( .A1(n6983), .A2(n7096), .ZN(n4989) );
  INV_X1 U6336 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5037) );
  NAND2_X1 U6337 ( .A1(n4496), .A2(n5660), .ZN(n8566) );
  INV_X1 U6338 ( .A(n8566), .ZN(n5664) );
  INV_X1 U6339 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5010) );
  INV_X1 U6340 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5034) );
  INV_X1 U6341 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  AND2_X1 U6342 ( .A1(n6037), .A2(n7442), .ZN(n4990) );
  NAND2_X1 U6343 ( .A1(n8896), .A2(n6559), .ZN(n8967) );
  INV_X1 U6344 ( .A(n10266), .ZN(n5632) );
  AND2_X1 U6345 ( .A1(n8087), .A2(n6449), .ZN(n4992) );
  NOR2_X1 U6346 ( .A1(n8360), .A2(n8361), .ZN(n4994) );
  NAND2_X1 U6347 ( .A1(n7865), .A2(n5212), .ZN(n4995) );
  INV_X1 U6348 ( .A(n6645), .ZN(n8157) );
  OR2_X1 U6349 ( .A1(n8744), .A2(n8599), .ZN(n4997) );
  INV_X1 U6350 ( .A(n6671), .ZN(n6670) );
  NAND2_X1 U6351 ( .A1(n6677), .A2(n6959), .ZN(n6678) );
  NAND2_X1 U6352 ( .A1(n6633), .A2(n6678), .ZN(n6679) );
  NOR2_X1 U6353 ( .A1(n6680), .A2(n6679), .ZN(n6682) );
  INV_X1 U6354 ( .A(n8035), .ZN(n6724) );
  NOR2_X1 U6355 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  AND2_X1 U6356 ( .A1(n8000), .A2(n6731), .ZN(n6732) );
  AND2_X1 U6357 ( .A1(n8044), .A2(n6736), .ZN(n6737) );
  NAND2_X1 U6358 ( .A1(n5650), .A2(n6749), .ZN(n6750) );
  NAND2_X1 U6359 ( .A1(n6751), .A2(n6959), .ZN(n6752) );
  NAND2_X1 U6360 ( .A1(n6753), .A2(n6752), .ZN(n6765) );
  MUX2_X1 U6361 ( .A(n6773), .B(n6772), .S(n6959), .Z(n6774) );
  NOR2_X1 U6362 ( .A1(n6793), .A2(n6788), .ZN(n6794) );
  OR2_X1 U6363 ( .A1(n8421), .A2(n6788), .ZN(n6805) );
  INV_X1 U6364 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5003) );
  NOR2_X1 U6365 ( .A1(n6819), .A2(n6820), .ZN(n6821) );
  NAND2_X1 U6366 ( .A1(n6817), .A2(n6788), .ZN(n6824) );
  INV_X1 U6367 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5008) );
  NOR2_X1 U6368 ( .A1(n8086), .A2(n7954), .ZN(n6447) );
  INV_X1 U6369 ( .A(n6471), .ZN(n6472) );
  NAND2_X1 U6370 ( .A1(n6824), .A2(n6823), .ZN(n6831) );
  INV_X1 U6371 ( .A(n8422), .ZN(n6348) );
  INV_X1 U6372 ( .A(n10007), .ZN(n6403) );
  INV_X1 U6373 ( .A(n6195), .ZN(n6065) );
  NAND2_X1 U6374 ( .A1(n6868), .A2(n7931), .ZN(n6869) );
  AOI21_X1 U6375 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n7391), .A(n10143), .ZN(
        n7392) );
  NOR2_X1 U6376 ( .A1(n10214), .A2(n8472), .ZN(n8474) );
  NOR2_X1 U6377 ( .A1(n8435), .A2(n10276), .ZN(n6687) );
  INV_X1 U6378 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5360) );
  OR2_X1 U6379 ( .A1(n6521), .A2(n6524), .ZN(n6522) );
  XNOR2_X1 U6380 ( .A(n6392), .B(n6393), .ZN(n7062) );
  NOR2_X1 U6381 ( .A1(n4504), .A2(n4987), .ZN(n6119) );
  INV_X1 U6382 ( .A(n9216), .ZN(n9161) );
  INV_X1 U6383 ( .A(n7887), .ZN(n6163) );
  INV_X1 U6384 ( .A(n5780), .ZN(n5722) );
  NAND2_X1 U6385 ( .A1(n6351), .A2(n5722), .ZN(n5834) );
  NAND2_X1 U6386 ( .A1(n5242), .A2(SI_10_), .ZN(n5243) );
  INV_X1 U6387 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5030) );
  INV_X1 U6388 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10127) );
  OR2_X1 U6389 ( .A1(n5381), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5408) );
  OR2_X1 U6390 ( .A1(n5257), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U6391 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5115) );
  AND2_X1 U6392 ( .A1(n6843), .A2(n6841), .ZN(n5669) );
  INV_X1 U6393 ( .A(n6739), .ZN(n5638) );
  NOR2_X1 U6394 ( .A1(n5337), .A2(n5336), .ZN(n5361) );
  AND2_X1 U6395 ( .A1(n5964), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5959) );
  INV_X1 U6396 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6058) );
  OR2_X1 U6397 ( .A1(n5992), .A2(n9298), .ZN(n5984) );
  NOR2_X1 U6398 ( .A1(n9379), .A2(n6008), .ZN(n6003) );
  OR2_X1 U6399 ( .A1(n9705), .A2(n9706), .ZN(n9703) );
  INV_X1 U6400 ( .A(n9173), .ZN(n9183) );
  AND2_X1 U6401 ( .A1(n5970), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5964) );
  OR2_X1 U6402 ( .A1(n6069), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U6403 ( .A1(n5834), .A2(n5833), .ZN(n5918) );
  NAND2_X1 U6404 ( .A1(n5247), .A2(n5246), .ZN(n5263) );
  NAND2_X1 U6405 ( .A1(n6881), .A2(n8037), .ZN(n6882) );
  NAND2_X1 U6406 ( .A1(n5439), .A2(n5438), .ZN(n5456) );
  INV_X1 U6407 ( .A(n8675), .ZN(n8687) );
  AND2_X1 U6408 ( .A1(n5342), .A2(n5341), .ZN(n5365) );
  INV_X1 U6409 ( .A(n10286), .ZN(n7802) );
  AND2_X1 U6410 ( .A1(n6944), .A2(n7010), .ZN(n6951) );
  NAND2_X1 U6411 ( .A1(n8956), .A2(n8958), .ZN(n6496) );
  INV_X1 U6412 ( .A(n6389), .ZN(n6390) );
  INV_X1 U6413 ( .A(n9664), .ZN(n8951) );
  INV_X1 U6414 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n7248) );
  INV_X1 U6415 ( .A(n9674), .ZN(n9615) );
  OR2_X1 U6416 ( .A1(n9968), .A2(n7281), .ZN(n9970) );
  INV_X1 U6417 ( .A(n7707), .ZN(n7814) );
  AND2_X1 U6418 ( .A1(n5225), .A2(n5186), .ZN(n5223) );
  INV_X1 U6419 ( .A(n6954), .ZN(n6955) );
  AOI21_X1 U6420 ( .B1(n8394), .B2(n8263), .A(n4979), .ZN(n8266) );
  AND2_X1 U6421 ( .A1(n6951), .A2(n6950), .ZN(n8410) );
  OAI22_X1 U6422 ( .A1(n7225), .A2(n7226), .B1(n6850), .B2(n6849), .ZN(n7231)
         );
  AND4_X1 U6423 ( .A1(n6625), .A2(n5583), .A3(n5582), .A4(n5581), .ZN(n6354)
         );
  NOR2_X1 U6424 ( .A1(n7206), .A2(n7207), .ZN(n7205) );
  AND2_X1 U6425 ( .A1(n6714), .A2(n6711), .ZN(n7867) );
  INV_X1 U6426 ( .A(n8714), .ZN(n8702) );
  NAND2_X1 U6427 ( .A1(n7010), .A2(n6932), .ZN(n8712) );
  INV_X1 U6428 ( .A(n8778), .ZN(n5678) );
  INV_X1 U6429 ( .A(n8777), .ZN(n8762) );
  NOR2_X1 U6430 ( .A1(n8559), .A2(n5588), .ZN(n5677) );
  INV_X1 U6431 ( .A(n8655), .ZN(n8652) );
  INV_X1 U6432 ( .A(n8227), .ZN(n7040) );
  XNOR2_X1 U6433 ( .A(n5595), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U6434 ( .A(n5229), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7700) );
  INV_X1 U6435 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6436 ( .A1(n6610), .A2(n6609), .ZN(n6611) );
  INV_X1 U6437 ( .A(n6331), .ZN(n6332) );
  AND4_X1 U6438 ( .A1(n5935), .A2(n5934), .A3(n5933), .A4(n5932), .ZN(n8993)
         );
  AND4_X1 U6439 ( .A1(n6029), .A2(n6028), .A3(n6027), .A4(n6026), .ZN(n7711)
         );
  INV_X1 U6440 ( .A(n9129), .ZN(n9232) );
  XNOR2_X1 U6441 ( .A(n5123), .B(SI_4_), .ZN(n5121) );
  NOR2_X1 U6442 ( .A1(n6956), .A2(n6955), .ZN(n6957) );
  INV_X1 U6443 ( .A(n8637), .ZN(n8424) );
  INV_X1 U6444 ( .A(n8721), .ZN(n8425) );
  INV_X1 U6445 ( .A(n7931), .ZN(n8432) );
  AND2_X1 U6446 ( .A1(n7300), .A2(n8712), .ZN(n8708) );
  INV_X1 U6447 ( .A(n6367), .ZN(n6368) );
  NAND2_X1 U6448 ( .A1(n5664), .A2(n5663), .ZN(n5665) );
  OR2_X1 U6449 ( .A1(n8770), .A2(n8769), .ZN(n8836) );
  OR2_X1 U6450 ( .A1(n10311), .A2(n10303), .ZN(n8841) );
  AND2_X1 U6451 ( .A1(n5603), .A2(n5602), .ZN(n8846) );
  INV_X1 U6452 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7011) );
  INV_X1 U6453 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6975) );
  AOI21_X1 U6454 ( .B1(n6613), .B2(n6612), .A(n6611), .ZN(n6617) );
  INV_X1 U6455 ( .A(n9649), .ZN(n9230) );
  INV_X1 U6456 ( .A(n8968), .ZN(n9791) );
  AND4_X1 U6457 ( .A1(n5928), .A2(n5927), .A3(n5926), .A4(n5925), .ZN(n9167)
         );
  AND2_X1 U6458 ( .A1(n7284), .A2(n9949), .ZN(n9968) );
  OR2_X1 U6459 ( .A1(n9968), .A2(n7270), .ZN(n9623) );
  OR2_X1 U6460 ( .A1(n7013), .A2(n7267), .ZN(n10109) );
  OR2_X1 U6461 ( .A1(n7013), .A2(n5896), .ZN(n10090) );
  INV_X1 U6462 ( .A(n5910), .ZN(n8273) );
  INV_X1 U6463 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6997) );
  INV_X1 U6464 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U6465 ( .A1(n5898), .A2(n4981), .ZN(P1_U3520) );
  INV_X1 U6466 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5624) );
  INV_X1 U6467 ( .A(n5149), .ZN(n5007) );
  NOR2_X1 U6468 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5001) );
  NOR2_X1 U6469 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5000) );
  NOR2_X1 U6470 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4999) );
  NAND4_X1 U6471 ( .A1(n5002), .A2(n5001), .A3(n5000), .A4(n4999), .ZN(n5336)
         );
  NOR2_X1 U6472 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5004) );
  NAND4_X1 U6473 ( .A1(n5004), .A2(n5360), .A3(n5376), .A4(n5003), .ZN(n5005)
         );
  INV_X1 U6474 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5015) );
  NAND2_X1 U6475 ( .A1(n5014), .A2(n5015), .ZN(n8293) );
  INV_X1 U6476 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5011) );
  INV_X1 U6477 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5013) );
  INV_X1 U6478 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5017) );
  OR2_X1 U6479 ( .A1(n5073), .A2(n5017), .ZN(n5025) );
  INV_X1 U6480 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6481 ( .A1(n5072), .A2(n5018), .ZN(n5024) );
  INV_X1 U6482 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7503) );
  INV_X1 U6483 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n5021) );
  XNOR2_X1 U6484 ( .A(n5027), .B(n5010), .ZN(n5577) );
  NAND2_X1 U6485 ( .A1(n4509), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5029) );
  INV_X1 U6486 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5028) );
  XNOR2_X1 U6487 ( .A(n5029), .B(n5028), .ZN(n5576) );
  INV_X1 U6488 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6979) );
  OR2_X1 U6489 ( .A1(n5107), .A2(n6979), .ZN(n5040) );
  INV_X1 U6490 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6491 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5031) );
  OR2_X1 U6492 ( .A1(n5068), .A2(n10118), .ZN(n5039) );
  NAND2_X1 U6493 ( .A1(n5068), .A2(n5065), .ZN(n5082) );
  OAI21_X1 U6494 ( .B1(n5065), .B2(n5034), .A(n5033), .ZN(n5035) );
  XNOR2_X1 U6495 ( .A(n5059), .B(SI_1_), .ZN(n6978) );
  OR2_X1 U6496 ( .A1(n5082), .A2(n6978), .ZN(n5038) );
  INV_X1 U6497 ( .A(n6848), .ZN(n5041) );
  INV_X1 U6498 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5042) );
  INV_X1 U6499 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5043) );
  OR2_X1 U6500 ( .A1(n5205), .A2(n5043), .ZN(n5046) );
  INV_X1 U6501 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7302) );
  OR2_X1 U6502 ( .A1(n5073), .A2(n7302), .ZN(n5045) );
  INV_X1 U6503 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7129) );
  OR2_X1 U6504 ( .A1(n5206), .A2(n7129), .ZN(n5044) );
  INV_X1 U6505 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n7178) );
  NAND2_X1 U6506 ( .A1(n5065), .A2(SI_0_), .ZN(n5049) );
  INV_X1 U6507 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5048) );
  XNOR2_X1 U6508 ( .A(n5049), .B(n5048), .ZN(n8852) );
  MUX2_X1 U6509 ( .A(n7178), .B(n8852), .S(n6962), .Z(n8784) );
  INV_X1 U6510 ( .A(n8784), .ZN(n7125) );
  NAND2_X1 U6511 ( .A1(n5625), .A2(n7125), .ZN(n5050) );
  NAND2_X1 U6512 ( .A1(n5051), .A2(n6848), .ZN(n5052) );
  NAND2_X1 U6513 ( .A1(n7509), .A2(n5052), .ZN(n7575) );
  NAND2_X1 U6514 ( .A1(n5137), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5058) );
  INV_X1 U6515 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5053) );
  OR2_X1 U6516 ( .A1(n5072), .A2(n5053), .ZN(n5057) );
  INV_X1 U6517 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6518 ( .A1(n5205), .A2(n5054), .ZN(n5056) );
  INV_X1 U6519 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7141) );
  OR2_X1 U6520 ( .A1(n5206), .A2(n7141), .ZN(n5055) );
  OR2_X1 U6521 ( .A1(n5107), .A2(n6971), .ZN(n5071) );
  NAND2_X1 U6522 ( .A1(n5059), .A2(SI_1_), .ZN(n5064) );
  INV_X1 U6523 ( .A(n5060), .ZN(n5062) );
  NAND2_X1 U6524 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  NAND2_X1 U6525 ( .A1(n5064), .A2(n5063), .ZN(n5084) );
  MUX2_X1 U6526 ( .A(n6969), .B(n6971), .S(n5065), .Z(n5085) );
  XNOR2_X2 U6527 ( .A(n5085), .B(SI_2_), .ZN(n5083) );
  XNOR2_X1 U6528 ( .A(n5084), .B(n5083), .ZN(n6970) );
  OR2_X1 U6529 ( .A1(n5082), .A2(n6970), .ZN(n5070) );
  OR2_X1 U6530 ( .A1(n7142), .A2(n5013), .ZN(n5067) );
  NAND2_X1 U6531 ( .A1(n7575), .A2(n7576), .ZN(n7550) );
  NAND2_X1 U6532 ( .A1(n6852), .A2(n10256), .ZN(n7551) );
  NAND2_X1 U6533 ( .A1(n5557), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5079) );
  INV_X1 U6534 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5074) );
  OR2_X1 U6535 ( .A1(n6621), .A2(n5074), .ZN(n5078) );
  OR2_X1 U6536 ( .A1(n5205), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5077) );
  INV_X1 U6537 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6538 ( .A1(n5080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U6539 ( .A(n5081), .B(n4998), .ZN(n7158) );
  OR2_X1 U6540 ( .A1(n5107), .A2(n4559), .ZN(n5089) );
  INV_X1 U6541 ( .A(n5085), .ZN(n5086) );
  NAND2_X1 U6542 ( .A1(n5086), .A2(SI_2_), .ZN(n5087) );
  XNOR2_X1 U6543 ( .A(n5102), .B(n5101), .ZN(n6973) );
  OR2_X1 U6544 ( .A1(n5082), .A2(n6973), .ZN(n5088) );
  OAI211_X1 U6545 ( .C1(n6962), .C2(n7158), .A(n5089), .B(n5088), .ZN(n10260)
         );
  NAND2_X1 U6546 ( .A1(n7622), .A2(n6846), .ZN(n5090) );
  AND2_X1 U6547 ( .A1(n7551), .A2(n5090), .ZN(n5091) );
  NAND2_X1 U6548 ( .A1(n7550), .A2(n5091), .ZN(n7618) );
  OR2_X1 U6549 ( .A1(n7622), .A2(n6846), .ZN(n7617) );
  INV_X1 U6550 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n7140) );
  OR2_X1 U6551 ( .A1(n6356), .A2(n7140), .ZN(n5097) );
  INV_X1 U6552 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5092) );
  OR2_X1 U6553 ( .A1(n5072), .A2(n5092), .ZN(n5096) );
  AND2_X1 U6554 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5093) );
  NOR2_X1 U6555 ( .A1(n5115), .A2(n5093), .ZN(n7486) );
  OR2_X1 U6556 ( .A1(n5205), .A2(n7486), .ZN(n5095) );
  NAND2_X1 U6557 ( .A1(n5137), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6558 ( .A1(n5098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5100) );
  INV_X1 U6559 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5099) );
  INV_X1 U6560 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6561 ( .A1(n5104), .A2(SI_3_), .ZN(n5105) );
  INV_X1 U6562 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6974) );
  XNOR2_X1 U6563 ( .A(n5122), .B(n5121), .ZN(n6976) );
  OR2_X1 U6564 ( .A1(n5082), .A2(n6976), .ZN(n5109) );
  OR2_X1 U6565 ( .A1(n5107), .A2(n6975), .ZN(n5108) );
  OAI211_X1 U6566 ( .C1(n6962), .C2(n7385), .A(n5109), .B(n5108), .ZN(n10266)
         );
  OR2_X1 U6567 ( .A1(n7608), .A2(n5632), .ZN(n5110) );
  AND2_X1 U6568 ( .A1(n7617), .A2(n5110), .ZN(n5111) );
  NAND2_X1 U6569 ( .A1(n7618), .A2(n5111), .ZN(n5113) );
  NAND2_X1 U6570 ( .A1(n7608), .A2(n5632), .ZN(n5112) );
  NAND2_X1 U6571 ( .A1(n5113), .A2(n5112), .ZN(n7752) );
  NAND2_X1 U6572 ( .A1(n5528), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5120) );
  OR2_X1 U6573 ( .A1(n6621), .A2(n4791), .ZN(n5119) );
  INV_X1 U6574 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5114) );
  OR2_X1 U6575 ( .A1(n5072), .A2(n5114), .ZN(n5118) );
  NAND2_X1 U6576 ( .A1(n5115), .A2(n10127), .ZN(n5138) );
  OR2_X1 U6577 ( .A1(n5115), .A2(n10127), .ZN(n5116) );
  AND2_X1 U6578 ( .A1(n5138), .A2(n5116), .ZN(n7607) );
  OR2_X1 U6579 ( .A1(n5205), .A2(n7607), .ZN(n5117) );
  INV_X1 U6580 ( .A(n5123), .ZN(n5124) );
  NAND2_X1 U6581 ( .A1(n5124), .A2(SI_4_), .ZN(n5125) );
  INV_X1 U6582 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5127) );
  OR2_X1 U6583 ( .A1(n5082), .A2(n6992), .ZN(n5133) );
  OR2_X1 U6584 ( .A1(n5107), .A2(n9356), .ZN(n5132) );
  OR2_X1 U6585 ( .A1(n5128), .A2(n5013), .ZN(n5130) );
  XNOR2_X1 U6586 ( .A(n5130), .B(n5129), .ZN(n7389) );
  OR2_X1 U6587 ( .A1(n6962), .A2(n7389), .ZN(n5131) );
  INV_X1 U6588 ( .A(n7611), .ZN(n10271) );
  NAND2_X1 U6589 ( .A1(n8436), .A2(n10271), .ZN(n5134) );
  NAND2_X1 U6590 ( .A1(n7752), .A2(n5134), .ZN(n5136) );
  NAND2_X1 U6591 ( .A1(n7761), .A2(n7611), .ZN(n5135) );
  NAND2_X1 U6592 ( .A1(n5136), .A2(n5135), .ZN(n7679) );
  NAND2_X1 U6593 ( .A1(n5137), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5144) );
  INV_X1 U6594 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7374) );
  OR2_X1 U6595 ( .A1(n6356), .A2(n7374), .ZN(n5143) );
  NAND2_X1 U6596 ( .A1(n5138), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5139) );
  AND2_X1 U6597 ( .A1(n5157), .A2(n5139), .ZN(n7685) );
  OR2_X1 U6598 ( .A1(n5205), .A2(n7685), .ZN(n5142) );
  INV_X1 U6599 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5140) );
  OR2_X1 U6600 ( .A1(n5072), .A2(n5140), .ZN(n5141) );
  INV_X1 U6601 ( .A(n5146), .ZN(n5147) );
  NAND2_X1 U6602 ( .A1(n5147), .A2(SI_5_), .ZN(n5148) );
  XNOR2_X1 U6603 ( .A(n5166), .B(n5165), .ZN(n6996) );
  OR2_X1 U6604 ( .A1(n5082), .A2(n6996), .ZN(n5154) );
  OR2_X1 U6605 ( .A1(n5107), .A2(n7000), .ZN(n5153) );
  NAND2_X1 U6606 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5150) );
  MUX2_X1 U6607 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5150), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5151) );
  OR2_X1 U6608 ( .A1(n5149), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5337) );
  NAND2_X1 U6609 ( .A1(n5151), .A2(n5337), .ZN(n7391) );
  OR2_X1 U6610 ( .A1(n6962), .A2(n7391), .ZN(n5152) );
  INV_X1 U6611 ( .A(n10276), .ZN(n7686) );
  NOR2_X1 U6612 ( .A1(n8435), .A2(n7686), .ZN(n5156) );
  NAND2_X1 U6613 ( .A1(n8435), .A2(n7686), .ZN(n5155) );
  NAND2_X1 U6614 ( .A1(n5557), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5162) );
  INV_X1 U6615 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7377) );
  OR2_X1 U6616 ( .A1(n6621), .A2(n7377), .ZN(n5161) );
  AND2_X1 U6617 ( .A1(n5157), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5158) );
  NOR2_X1 U6618 ( .A1(n5202), .A2(n5158), .ZN(n8252) );
  OR2_X1 U6619 ( .A1(n5579), .A2(n8252), .ZN(n5160) );
  INV_X1 U6620 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7656) );
  OR2_X1 U6621 ( .A1(n6356), .A2(n7656), .ZN(n5159) );
  NAND2_X1 U6622 ( .A1(n5337), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  INV_X1 U6623 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5163) );
  XNOR2_X1 U6624 ( .A(n5164), .B(n5163), .ZN(n7396) );
  INV_X1 U6625 ( .A(n5167), .ZN(n5168) );
  INV_X1 U6626 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n5169) );
  MUX2_X1 U6627 ( .A(n7005), .B(n5169), .S(n5902), .Z(n5174) );
  XNOR2_X1 U6628 ( .A(n5173), .B(n5172), .ZN(n7006) );
  OR2_X1 U6629 ( .A1(n7006), .A2(n5082), .ZN(n5171) );
  OR2_X1 U6630 ( .A1(n5107), .A2(n7005), .ZN(n5170) );
  OAI211_X1 U6631 ( .C1(n6962), .C2(n7396), .A(n5171), .B(n5170), .ZN(n8254)
         );
  NAND2_X1 U6632 ( .A1(n7681), .A2(n8254), .ZN(n6705) );
  INV_X1 U6633 ( .A(n8254), .ZN(n10281) );
  NAND2_X1 U6634 ( .A1(n8434), .A2(n10281), .ZN(n7800) );
  NAND2_X1 U6635 ( .A1(n6705), .A2(n7800), .ZN(n7796) );
  INV_X1 U6636 ( .A(n5174), .ZN(n5175) );
  NAND2_X1 U6637 ( .A1(n5175), .A2(SI_7_), .ZN(n5176) );
  INV_X1 U6638 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5177) );
  MUX2_X1 U6639 ( .A(n7011), .B(n5177), .S(n5902), .Z(n5178) );
  INV_X1 U6640 ( .A(SI_8_), .ZN(n9390) );
  INV_X1 U6641 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6642 ( .A1(n5179), .A2(SI_8_), .ZN(n5180) );
  INV_X1 U6643 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7033) );
  INV_X1 U6644 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5182) );
  MUX2_X1 U6645 ( .A(n7033), .B(n5182), .S(n5902), .Z(n5184) );
  INV_X1 U6646 ( .A(SI_9_), .ZN(n5183) );
  NAND2_X1 U6647 ( .A1(n5184), .A2(n5183), .ZN(n5225) );
  INV_X1 U6648 ( .A(n5184), .ZN(n5185) );
  NAND2_X1 U6649 ( .A1(n5185), .A2(SI_9_), .ZN(n5186) );
  NAND2_X1 U6650 ( .A1(n7029), .A2(n6627), .ZN(n5188) );
  INV_X2 U6651 ( .A(n6962), .ZN(n5405) );
  NOR2_X1 U6652 ( .A1(n5194), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5251) );
  OR2_X1 U6653 ( .A1(n5251), .A2(n5013), .ZN(n5229) );
  AOI22_X1 U6654 ( .A1(n6618), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5405), .B2(
        n7700), .ZN(n5187) );
  NAND2_X1 U6655 ( .A1(n5188), .A2(n5187), .ZN(n7884) );
  INV_X1 U6656 ( .A(n7884), .ZN(n10292) );
  NAND2_X1 U6657 ( .A1(n5557), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5193) );
  INV_X1 U6658 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7872) );
  OR2_X1 U6659 ( .A1(n6621), .A2(n7872), .ZN(n5192) );
  INV_X1 U6660 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n5201) );
  INV_X1 U6661 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n9491) );
  OR2_X1 U6662 ( .A1(n5204), .A2(n9491), .ZN(n5189) );
  AND2_X1 U6663 ( .A1(n5234), .A2(n5189), .ZN(n7882) );
  OR2_X1 U6664 ( .A1(n5205), .A2(n7882), .ZN(n5191) );
  INV_X1 U6665 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7643) );
  OR2_X1 U6666 ( .A1(n6356), .A2(n7643), .ZN(n5190) );
  NAND2_X1 U6667 ( .A1(n10292), .A2(n6864), .ZN(n5213) );
  NAND2_X1 U6668 ( .A1(n5194), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5195) );
  XNOR2_X1 U6669 ( .A(n5195), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8447) );
  AOI22_X1 U6670 ( .A1(n6618), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5405), .B2(
        n8447), .ZN(n5199) );
  NAND2_X1 U6671 ( .A1(n7007), .A2(n6627), .ZN(n5198) );
  NAND2_X1 U6672 ( .A1(n5137), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5210) );
  INV_X1 U6673 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5200) );
  NOR2_X1 U6674 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  OR2_X1 U6675 ( .A1(n5205), .A2(n4464), .ZN(n5208) );
  INV_X1 U6676 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7658) );
  OR2_X1 U6677 ( .A1(n5206), .A2(n7658), .ZN(n5207) );
  NAND2_X1 U6678 ( .A1(n10286), .A2(n8433), .ZN(n7865) );
  NAND2_X1 U6679 ( .A1(n5211), .A2(n7884), .ZN(n5212) );
  INV_X1 U6680 ( .A(n5218), .ZN(n5215) );
  NAND2_X1 U6681 ( .A1(n8247), .A2(n5216), .ZN(n5222) );
  INV_X1 U6682 ( .A(n5217), .ZN(n5220) );
  OR2_X1 U6683 ( .A1(n7681), .A2(n10281), .ZN(n7797) );
  AND2_X1 U6684 ( .A1(n7797), .A2(n5218), .ZN(n5219) );
  INV_X1 U6685 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7036) );
  INV_X1 U6686 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5227) );
  MUX2_X1 U6687 ( .A(n7036), .B(n5227), .S(n5902), .Z(n5241) );
  NAND2_X1 U6688 ( .A1(n7031), .A2(n6627), .ZN(n5233) );
  INV_X1 U6689 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6690 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U6691 ( .A1(n5230), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5231) );
  XNOR2_X1 U6692 ( .A(n5231), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7728) );
  AOI22_X1 U6693 ( .A1(n6618), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5405), .B2(
        n7728), .ZN(n5232) );
  NAND2_X1 U6694 ( .A1(n5557), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5239) );
  INV_X1 U6695 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7949) );
  OR2_X1 U6696 ( .A1(n6621), .A2(n7949), .ZN(n5238) );
  INV_X1 U6697 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7647) );
  OR2_X1 U6698 ( .A1(n6356), .A2(n7647), .ZN(n5237) );
  NAND2_X1 U6699 ( .A1(n5234), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5235) );
  AND2_X1 U6700 ( .A1(n5257), .A2(n5235), .ZN(n8123) );
  OR2_X1 U6701 ( .A1(n5579), .A2(n8123), .ZN(n5236) );
  AND2_X1 U6702 ( .A1(n10301), .A2(n8432), .ZN(n6874) );
  INV_X1 U6703 ( .A(n5241), .ZN(n5242) );
  INV_X1 U6704 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7054) );
  INV_X1 U6705 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9332) );
  MUX2_X1 U6706 ( .A(n7054), .B(n9332), .S(n5902), .Z(n5247) );
  INV_X1 U6707 ( .A(SI_11_), .ZN(n5246) );
  INV_X1 U6708 ( .A(n5247), .ZN(n5248) );
  NAND2_X1 U6709 ( .A1(n5248), .A2(SI_11_), .ZN(n5249) );
  NAND2_X1 U6710 ( .A1(n7053), .A2(n6627), .ZN(n5254) );
  NOR2_X1 U6711 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5250) );
  AND2_X1 U6712 ( .A1(n5251), .A2(n5250), .ZN(n5267) );
  OR2_X1 U6713 ( .A1(n5267), .A2(n5013), .ZN(n5252) );
  XNOR2_X1 U6714 ( .A(n5252), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7835) );
  AOI22_X1 U6715 ( .A1(n6618), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5405), .B2(
        n7835), .ZN(n5253) );
  NAND2_X1 U6716 ( .A1(n5557), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5262) );
  INV_X1 U6717 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5255) );
  OR2_X1 U6718 ( .A1(n6356), .A2(n5255), .ZN(n5261) );
  INV_X1 U6719 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5256) );
  OR2_X1 U6720 ( .A1(n6621), .A2(n5256), .ZN(n5260) );
  NAND2_X1 U6721 ( .A1(n5257), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5258) );
  AND2_X1 U6722 ( .A1(n5271), .A2(n5258), .ZN(n8183) );
  OR2_X1 U6723 ( .A1(n5579), .A2(n8183), .ZN(n5259) );
  INV_X1 U6724 ( .A(n8134), .ZN(n8431) );
  NOR2_X1 U6725 ( .A1(n10307), .A2(n8431), .ZN(n8031) );
  INV_X1 U6726 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9449) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5266) );
  MUX2_X1 U6728 ( .A(n9449), .B(n5266), .S(n5902), .Z(n5277) );
  XNOR2_X1 U6729 ( .A(n5280), .B(n5276), .ZN(n7072) );
  NAND2_X1 U6730 ( .A1(n7072), .A2(n6627), .ZN(n5270) );
  NAND2_X1 U6731 ( .A1(n5267), .A2(n4684), .ZN(n5281) );
  NAND2_X1 U6732 ( .A1(n5281), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5268) );
  XNOR2_X1 U6733 ( .A(n5268), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8504) );
  AOI22_X1 U6734 ( .A1(n6618), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5405), .B2(
        n8504), .ZN(n5269) );
  NAND2_X1 U6735 ( .A1(n5137), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5275) );
  INV_X1 U6736 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8101) );
  OR2_X1 U6737 ( .A1(n5072), .A2(n8101), .ZN(n5274) );
  NOR2_X1 U6738 ( .A1(n5285), .A2(n4479), .ZN(n8131) );
  OR2_X1 U6739 ( .A1(n5579), .A2(n8131), .ZN(n5273) );
  INV_X1 U6740 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8503) );
  OR2_X1 U6741 ( .A1(n6356), .A2(n8503), .ZN(n5272) );
  NAND4_X1 U6742 ( .A1(n5275), .A2(n5274), .A3(n5273), .A4(n5272), .ZN(n8430)
         );
  OR2_X1 U6743 ( .A1(n8031), .A2(n4470), .ZN(n7997) );
  INV_X1 U6744 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6745 ( .A1(n5278), .A2(SI_12_), .ZN(n5279) );
  MUX2_X1 U6746 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5902), .Z(n5300) );
  XNOR2_X1 U6747 ( .A(n5300), .B(SI_13_), .ZN(n5297) );
  XNOR2_X1 U6748 ( .A(n5299), .B(n5297), .ZN(n7222) );
  NAND2_X1 U6749 ( .A1(n7222), .A2(n6627), .ZN(n5284) );
  OR2_X1 U6750 ( .A1(n5281), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6751 ( .A1(n5282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5302) );
  XNOR2_X1 U6752 ( .A(n5302), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U6753 ( .A1(n6618), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5405), .B2(
        n10165), .ZN(n5283) );
  NAND2_X1 U6754 ( .A1(n5557), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5290) );
  INV_X1 U6755 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8467) );
  OR2_X1 U6756 ( .A1(n6621), .A2(n8467), .ZN(n5289) );
  INV_X1 U6757 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8011) );
  OR2_X1 U6758 ( .A1(n6356), .A2(n8011), .ZN(n5288) );
  INV_X1 U6759 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8372) );
  OR2_X1 U6760 ( .A1(n5285), .A2(n8372), .ZN(n5286) );
  NAND2_X1 U6761 ( .A1(n5285), .A2(n8372), .ZN(n5306) );
  AND2_X1 U6762 ( .A1(n5286), .A2(n5306), .ZN(n8375) );
  OR2_X1 U6763 ( .A1(n5579), .A2(n8375), .ZN(n5287) );
  OR2_X1 U6764 ( .A1(n8377), .A2(n8429), .ZN(n5295) );
  INV_X1 U6765 ( .A(n5295), .ZN(n5291) );
  OR2_X1 U6766 ( .A1(n7997), .A2(n5291), .ZN(n5292) );
  OR2_X1 U6767 ( .A1(n8377), .A2(n8037), .ZN(n6734) );
  NAND2_X1 U6768 ( .A1(n8377), .A2(n8037), .ZN(n6735) );
  NAND2_X1 U6769 ( .A1(n10307), .A2(n8431), .ZN(n8032) );
  AND2_X1 U6770 ( .A1(n4506), .A2(n8032), .ZN(n5293) );
  NOR2_X1 U6771 ( .A1(n4470), .A2(n5293), .ZN(n7998) );
  OR2_X1 U6772 ( .A1(n8000), .A2(n7998), .ZN(n5294) );
  AND2_X1 U6773 ( .A1(n5295), .A2(n5294), .ZN(n5296) );
  NAND2_X1 U6774 ( .A1(n5300), .A2(SI_13_), .ZN(n5301) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5902), .Z(n5317) );
  XNOR2_X1 U6776 ( .A(n5317), .B(SI_14_), .ZN(n5314) );
  XNOR2_X1 U6777 ( .A(n5316), .B(n5314), .ZN(n7238) );
  NAND2_X1 U6778 ( .A1(n7238), .A2(n6627), .ZN(n5305) );
  NAND2_X1 U6779 ( .A1(n5302), .A2(n4683), .ZN(n5303) );
  NAND2_X1 U6780 ( .A1(n5303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5320) );
  XNOR2_X1 U6781 ( .A(n5320), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U6782 ( .A1(n6618), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5405), .B2(
        n10182), .ZN(n5304) );
  NAND2_X1 U6783 ( .A1(n5557), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5311) );
  INV_X1 U6784 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8469) );
  OR2_X1 U6785 ( .A1(n6621), .A2(n8469), .ZN(n5310) );
  INV_X1 U6786 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8508) );
  OR2_X1 U6787 ( .A1(n6356), .A2(n8508), .ZN(n5309) );
  NAND2_X1 U6788 ( .A1(n5306), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5307) );
  AND2_X1 U6789 ( .A1(n5325), .A2(n5307), .ZN(n8298) );
  OR2_X1 U6790 ( .A1(n5579), .A2(n8298), .ZN(n5308) );
  NAND2_X1 U6791 ( .A1(n8300), .A2(n8428), .ZN(n5312) );
  NAND2_X1 U6792 ( .A1(n5313), .A2(n5312), .ZN(n8107) );
  INV_X1 U6793 ( .A(n5314), .ZN(n5315) );
  NAND2_X1 U6794 ( .A1(n5317), .A2(SI_14_), .ZN(n5318) );
  MUX2_X1 U6795 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n5902), .Z(n5335) );
  XNOR2_X1 U6796 ( .A(n5335), .B(SI_15_), .ZN(n5332) );
  XNOR2_X1 U6797 ( .A(n5334), .B(n5332), .ZN(n7340) );
  NAND2_X1 U6798 ( .A1(n7340), .A2(n6627), .ZN(n5324) );
  INV_X1 U6799 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6800 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  NAND2_X1 U6801 ( .A1(n5321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5322) );
  XNOR2_X1 U6802 ( .A(n5322), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U6803 ( .A1(n6618), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n10198), 
        .B2(n5405), .ZN(n5323) );
  NAND2_X1 U6804 ( .A1(n5557), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5330) );
  INV_X1 U6805 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8112) );
  OR2_X1 U6806 ( .A1(n6356), .A2(n8112), .ZN(n5329) );
  INV_X1 U6807 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n10207) );
  OR2_X1 U6808 ( .A1(n6621), .A2(n10207), .ZN(n5328) );
  AND2_X1 U6809 ( .A1(n5325), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5326) );
  NOR2_X1 U6810 ( .A1(n5342), .A2(n5326), .ZN(n8109) );
  OR2_X1 U6811 ( .A1(n5579), .A2(n8109), .ZN(n5327) );
  OR2_X1 U6812 ( .A1(n8405), .A2(n8427), .ZN(n5331) );
  INV_X1 U6813 ( .A(n5332), .ZN(n5333) );
  MUX2_X1 U6814 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n5902), .Z(n5353) );
  XNOR2_X1 U6815 ( .A(n5353), .B(SI_16_), .ZN(n5350) );
  XNOR2_X1 U6816 ( .A(n5352), .B(n5350), .ZN(n7495) );
  NAND2_X1 U6817 ( .A1(n7495), .A2(n6627), .ZN(n5340) );
  OR2_X1 U6818 ( .A1(n5361), .A2(n5013), .ZN(n5338) );
  XNOR2_X1 U6819 ( .A(n5338), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U6820 ( .A1(n6618), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5405), .B2(
        n10214), .ZN(n5339) );
  NAND2_X1 U6821 ( .A1(n5557), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5347) );
  INV_X1 U6822 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8472) );
  OR2_X1 U6823 ( .A1(n6621), .A2(n8472), .ZN(n5346) );
  INV_X1 U6824 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8512) );
  OR2_X1 U6825 ( .A1(n6356), .A2(n8512), .ZN(n5345) );
  INV_X1 U6826 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5341) );
  NOR2_X1 U6827 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  OR2_X1 U6828 ( .A1(n5365), .A2(n5343), .ZN(n8171) );
  INV_X1 U6829 ( .A(n8171), .ZN(n8337) );
  OR2_X1 U6830 ( .A1(n5579), .A2(n8337), .ZN(n5344) );
  NAND2_X1 U6831 ( .A1(n8339), .A2(n8719), .ZN(n6755) );
  NAND2_X1 U6832 ( .A1(n6756), .A2(n6755), .ZN(n6645) );
  NAND2_X1 U6833 ( .A1(n5348), .A2(n6645), .ZN(n8160) );
  INV_X1 U6834 ( .A(n8719), .ZN(n8426) );
  NAND2_X1 U6835 ( .A1(n8339), .A2(n8426), .ZN(n5349) );
  INV_X1 U6836 ( .A(n5350), .ZN(n5351) );
  NAND2_X1 U6837 ( .A1(n5352), .A2(n5351), .ZN(n5355) );
  NAND2_X1 U6838 ( .A1(n5353), .A2(SI_16_), .ZN(n5354) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7530) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7529) );
  MUX2_X1 U6841 ( .A(n7530), .B(n7529), .S(n5902), .Z(n5357) );
  INV_X1 U6842 ( .A(SI_17_), .ZN(n5356) );
  NAND2_X1 U6843 ( .A1(n5357), .A2(n5356), .ZN(n5372) );
  INV_X1 U6844 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6845 ( .A1(n5358), .A2(SI_17_), .ZN(n5359) );
  NAND2_X1 U6846 ( .A1(n5372), .A2(n5359), .ZN(n5373) );
  XNOR2_X1 U6847 ( .A(n5374), .B(n5373), .ZN(n7528) );
  NAND2_X1 U6848 ( .A1(n7528), .A2(n6627), .ZN(n5364) );
  NAND2_X1 U6849 ( .A1(n5361), .A2(n5360), .ZN(n5375) );
  NAND2_X1 U6850 ( .A1(n5375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5362) );
  XNOR2_X1 U6851 ( .A(n5362), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U6852 ( .A1(n6618), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5405), .B2(
        n10233), .ZN(n5363) );
  NAND2_X1 U6853 ( .A1(n5557), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5370) );
  INV_X1 U6854 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9447) );
  OR2_X1 U6855 ( .A1(n6356), .A2(n9447), .ZN(n5369) );
  INV_X1 U6856 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8478) );
  OR2_X1 U6857 ( .A1(n6621), .A2(n8478), .ZN(n5368) );
  INV_X1 U6858 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8344) );
  OR2_X1 U6859 ( .A1(n5365), .A2(n8344), .ZN(n5366) );
  AND2_X1 U6860 ( .A1(n5381), .A2(n5366), .ZN(n8713) );
  OR2_X1 U6861 ( .A1(n5579), .A2(n8713), .ZN(n5367) );
  OR2_X1 U6862 ( .A1(n8711), .A2(n8334), .ZN(n6761) );
  NAND2_X1 U6863 ( .A1(n8711), .A2(n8334), .ZN(n6744) );
  INV_X1 U6864 ( .A(n8334), .ZN(n8696) );
  NAND2_X1 U6865 ( .A1(n8711), .A2(n8696), .ZN(n5371) );
  INV_X1 U6866 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7630) );
  INV_X1 U6867 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9404) );
  MUX2_X1 U6868 ( .A(n7630), .B(n9404), .S(n5902), .Z(n5392) );
  XNOR2_X1 U6869 ( .A(n5392), .B(SI_18_), .ZN(n5391) );
  XNOR2_X1 U6870 ( .A(n5396), .B(n5391), .ZN(n7629) );
  NAND2_X1 U6871 ( .A1(n7629), .A2(n6627), .ZN(n5380) );
  INV_X1 U6872 ( .A(n5375), .ZN(n5377) );
  NAND2_X1 U6873 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  XNOR2_X1 U6874 ( .A(n5402), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8516) );
  AOI22_X1 U6875 ( .A1(n6618), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5405), .B2(
        n8516), .ZN(n5379) );
  NAND2_X1 U6876 ( .A1(n5137), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5387) );
  INV_X1 U6877 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9508) );
  OR2_X1 U6878 ( .A1(n5072), .A2(n9508), .ZN(n5386) );
  NAND2_X1 U6879 ( .A1(n5381), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5382) );
  AND2_X1 U6880 ( .A1(n5408), .A2(n5382), .ZN(n8699) );
  OR2_X1 U6881 ( .A1(n5579), .A2(n8699), .ZN(n5385) );
  INV_X1 U6882 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n5383) );
  OR2_X1 U6883 ( .A1(n6356), .A2(n5383), .ZN(n5384) );
  OR2_X1 U6884 ( .A1(n8703), .A2(n8425), .ZN(n5388) );
  NAND2_X1 U6885 ( .A1(n8703), .A2(n8425), .ZN(n5389) );
  NAND2_X1 U6886 ( .A1(n5390), .A2(n5389), .ZN(n8676) );
  INV_X1 U6887 ( .A(n5391), .ZN(n5395) );
  INV_X1 U6888 ( .A(n5392), .ZN(n5393) );
  NAND2_X1 U6889 ( .A1(n5393), .A2(SI_18_), .ZN(n5394) );
  INV_X1 U6890 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7745) );
  INV_X1 U6891 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7744) );
  INV_X1 U6892 ( .A(SI_19_), .ZN(n5397) );
  NAND2_X1 U6893 ( .A1(n5398), .A2(n5397), .ZN(n5416) );
  INV_X1 U6894 ( .A(n5398), .ZN(n5399) );
  NAND2_X1 U6895 ( .A1(n5399), .A2(SI_19_), .ZN(n5400) );
  NAND2_X1 U6896 ( .A1(n5416), .A2(n5400), .ZN(n5417) );
  XNOR2_X1 U6897 ( .A(n5418), .B(n5417), .ZN(n7743) );
  NAND2_X1 U6898 ( .A1(n7743), .A2(n6627), .ZN(n5407) );
  INV_X1 U6899 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6900 ( .A1(n5402), .A2(n5401), .ZN(n5403) );
  NAND2_X1 U6901 ( .A1(n5403), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5404) );
  AOI22_X1 U6902 ( .A1(n6618), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8535), .B2(
        n5405), .ZN(n5406) );
  AND2_X1 U6903 ( .A1(n5408), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5409) );
  OR2_X1 U6904 ( .A1(n5409), .A2(n5427), .ZN(n8682) );
  NAND2_X1 U6905 ( .A1(n5551), .A2(n8682), .ZN(n5413) );
  NAND2_X1 U6906 ( .A1(n5528), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5412) );
  INV_X1 U6907 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8684) );
  OR2_X1 U6908 ( .A1(n6621), .A2(n8684), .ZN(n5411) );
  NAND2_X1 U6909 ( .A1(n5557), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5410) );
  NAND4_X1 U6910 ( .A1(n5413), .A2(n5412), .A3(n5411), .A4(n5410), .ZN(n8693)
         );
  INV_X1 U6911 ( .A(n8768), .ZN(n8686) );
  INV_X1 U6912 ( .A(n8693), .ZN(n8364) );
  NAND2_X1 U6913 ( .A1(n8686), .A2(n8364), .ZN(n6766) );
  NAND2_X1 U6914 ( .A1(n8676), .A2(n8687), .ZN(n5415) );
  OR2_X1 U6915 ( .A1(n8768), .A2(n8364), .ZN(n5414) );
  INV_X1 U6916 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7821) );
  INV_X1 U6917 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7773) );
  MUX2_X1 U6918 ( .A(n7821), .B(n7773), .S(n5902), .Z(n5420) );
  INV_X1 U6919 ( .A(SI_20_), .ZN(n5419) );
  NAND2_X1 U6920 ( .A1(n5420), .A2(n5419), .ZN(n5434) );
  INV_X1 U6921 ( .A(n5420), .ZN(n5421) );
  NAND2_X1 U6922 ( .A1(n5421), .A2(SI_20_), .ZN(n5422) );
  AND2_X1 U6923 ( .A1(n5434), .A2(n5422), .ZN(n5423) );
  OR2_X1 U6924 ( .A1(n5107), .A2(n7821), .ZN(n5425) );
  INV_X1 U6925 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5426) );
  NOR2_X1 U6926 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  OR2_X1 U6927 ( .A1(n5439), .A2(n5428), .ZN(n8670) );
  NAND2_X1 U6928 ( .A1(n8670), .A2(n5551), .ZN(n5433) );
  NAND2_X1 U6929 ( .A1(n5137), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6930 ( .A1(n5557), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5429) );
  AND2_X1 U6931 ( .A1(n5430), .A2(n5429), .ZN(n5432) );
  NAND2_X1 U6932 ( .A1(n5528), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6933 ( .A1(n8832), .A2(n8678), .ZN(n8650) );
  INV_X1 U6934 ( .A(n8678), .ZN(n8657) );
  OR2_X1 U6935 ( .A1(n8832), .A2(n8657), .ZN(n8654) );
  INV_X1 U6936 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7851) );
  INV_X1 U6937 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7825) );
  MUX2_X1 U6938 ( .A(n7851), .B(n7825), .S(n5902), .Z(n5446) );
  XNOR2_X1 U6939 ( .A(n5446), .B(SI_21_), .ZN(n5445) );
  NAND2_X1 U6940 ( .A1(n7824), .A2(n6627), .ZN(n5437) );
  OR2_X1 U6941 ( .A1(n5107), .A2(n7851), .ZN(n5436) );
  INV_X1 U6942 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6943 ( .A1(n5439), .A2(n5438), .ZN(n5440) );
  NAND2_X1 U6944 ( .A1(n5456), .A2(n5440), .ZN(n8661) );
  NAND2_X1 U6945 ( .A1(n8661), .A2(n5551), .ZN(n5443) );
  AOI22_X1 U6946 ( .A1(n5528), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n5137), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U6947 ( .A1(n5557), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6948 ( .A1(n5444), .A2(n8636), .ZN(n6777) );
  OR2_X1 U6949 ( .A1(n5444), .A2(n8667), .ZN(n8631) );
  INV_X1 U6950 ( .A(n5445), .ZN(n5449) );
  INV_X1 U6951 ( .A(n5446), .ZN(n5447) );
  NAND2_X1 U6952 ( .A1(n5447), .A2(SI_21_), .ZN(n5448) );
  INV_X1 U6953 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7939) );
  INV_X1 U6954 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7938) );
  MUX2_X1 U6955 ( .A(n7939), .B(n7938), .S(n5902), .Z(n5451) );
  INV_X1 U6956 ( .A(SI_22_), .ZN(n9301) );
  NAND2_X1 U6957 ( .A1(n5451), .A2(n9301), .ZN(n5464) );
  INV_X1 U6958 ( .A(n5451), .ZN(n5452) );
  NAND2_X1 U6959 ( .A1(n5452), .A2(SI_22_), .ZN(n5453) );
  NAND2_X1 U6960 ( .A1(n5464), .A2(n5453), .ZN(n5465) );
  XNOR2_X1 U6961 ( .A(n5466), .B(n5465), .ZN(n7936) );
  NAND2_X1 U6962 ( .A1(n7936), .A2(n6627), .ZN(n5455) );
  OR2_X1 U6963 ( .A1(n5107), .A2(n7939), .ZN(n5454) );
  NAND2_X1 U6964 ( .A1(n5456), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U6965 ( .A1(n5475), .A2(n5457), .ZN(n8642) );
  NAND2_X1 U6966 ( .A1(n8642), .A2(n5551), .ZN(n5460) );
  AOI22_X1 U6967 ( .A1(n5528), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n5137), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U6968 ( .A1(n5557), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6969 ( .A1(n8641), .A2(n8622), .ZN(n6781) );
  INV_X1 U6970 ( .A(n8638), .ZN(n5461) );
  NAND2_X1 U6971 ( .A1(n5462), .A2(n5461), .ZN(n8633) );
  INV_X1 U6972 ( .A(n8622), .ZN(n8658) );
  OR2_X1 U6973 ( .A1(n8641), .A2(n8658), .ZN(n5463) );
  NAND2_X1 U6974 ( .A1(n8633), .A2(n5463), .ZN(n8619) );
  INV_X1 U6975 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8021) );
  INV_X1 U6976 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9354) );
  MUX2_X1 U6977 ( .A(n8021), .B(n9354), .S(n5902), .Z(n5468) );
  INV_X1 U6978 ( .A(SI_23_), .ZN(n5467) );
  NAND2_X1 U6979 ( .A1(n5468), .A2(n5467), .ZN(n5485) );
  INV_X1 U6980 ( .A(n5468), .ZN(n5469) );
  NAND2_X1 U6981 ( .A1(n5469), .A2(SI_23_), .ZN(n5470) );
  NAND2_X1 U6982 ( .A1(n5485), .A2(n5470), .ZN(n5471) );
  NAND2_X1 U6983 ( .A1(n4497), .A2(n5471), .ZN(n5472) );
  NAND2_X1 U6984 ( .A1(n5472), .A2(n5486), .ZN(n8022) );
  NAND2_X1 U6985 ( .A1(n8022), .A2(n6627), .ZN(n5474) );
  OR2_X1 U6986 ( .A1(n5107), .A2(n8021), .ZN(n5473) );
  NAND2_X1 U6987 ( .A1(n5475), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6988 ( .A1(n5492), .A2(n5476), .ZN(n8625) );
  NAND2_X1 U6989 ( .A1(n8625), .A2(n5551), .ZN(n5481) );
  INV_X1 U6990 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U6991 ( .A1(n5137), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U6992 ( .A1(n5557), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U6993 ( .C1(n6356), .C2(n8750), .A(n5478), .B(n5477), .ZN(n5479)
         );
  INV_X1 U6994 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6995 ( .A1(n8749), .A2(n8424), .ZN(n5482) );
  NAND2_X1 U6996 ( .A1(n8619), .A2(n5482), .ZN(n5484) );
  OR2_X1 U6997 ( .A1(n8749), .A2(n8424), .ZN(n5483) );
  NAND2_X1 U6998 ( .A1(n5484), .A2(n5483), .ZN(n8609) );
  INV_X1 U6999 ( .A(n8609), .ZN(n5497) );
  INV_X1 U7000 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8285) );
  INV_X1 U7001 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8153) );
  MUX2_X1 U7002 ( .A(n8285), .B(n8153), .S(n5902), .Z(n5487) );
  INV_X1 U7003 ( .A(SI_24_), .ZN(n9431) );
  NAND2_X1 U7004 ( .A1(n5487), .A2(n9431), .ZN(n5502) );
  INV_X1 U7005 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U7006 ( .A1(n5488), .A2(SI_24_), .ZN(n5489) );
  AND2_X1 U7007 ( .A1(n5502), .A2(n5489), .ZN(n5500) );
  XNOR2_X1 U7008 ( .A(n5501), .B(n5500), .ZN(n8152) );
  NAND2_X1 U7009 ( .A1(n8152), .A2(n6627), .ZN(n5491) );
  OR2_X1 U7010 ( .A1(n5107), .A2(n8285), .ZN(n5490) );
  AND2_X1 U7011 ( .A1(n5492), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5493) );
  OR2_X1 U7012 ( .A1(n5493), .A2(n5509), .ZN(n8613) );
  INV_X1 U7013 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U7014 ( .A1(n5137), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7015 ( .A1(n5557), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5494) );
  OAI211_X1 U7016 ( .C1(n6356), .C2(n9427), .A(n5495), .B(n5494), .ZN(n5496)
         );
  AOI21_X1 U7017 ( .B1(n8613), .B2(n5551), .A(n5496), .ZN(n8621) );
  INV_X1 U7018 ( .A(n8621), .ZN(n8599) );
  NAND2_X1 U7019 ( .A1(n5497), .A2(n4997), .ZN(n5499) );
  NAND2_X1 U7020 ( .A1(n8744), .A2(n8599), .ZN(n5498) );
  NAND2_X1 U7021 ( .A1(n5501), .A2(n5500), .ZN(n5503) );
  INV_X1 U7022 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8220) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8224) );
  MUX2_X1 U7024 ( .A(n8220), .B(n8224), .S(n5902), .Z(n5505) );
  INV_X1 U7025 ( .A(SI_25_), .ZN(n5504) );
  NAND2_X1 U7026 ( .A1(n5505), .A2(n5504), .ZN(n5520) );
  INV_X1 U7027 ( .A(n5505), .ZN(n5506) );
  NAND2_X1 U7028 ( .A1(n5506), .A2(SI_25_), .ZN(n5507) );
  AND2_X1 U7029 ( .A1(n5520), .A2(n5507), .ZN(n5518) );
  XNOR2_X1 U7030 ( .A(n5519), .B(n5518), .ZN(n8219) );
  NOR2_X1 U7031 ( .A1(n5107), .A2(n8220), .ZN(n5508) );
  INV_X1 U7032 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8324) );
  NOR2_X1 U7033 ( .A1(n5509), .A2(n8324), .ZN(n5510) );
  OR2_X1 U7034 ( .A1(n5526), .A2(n5510), .ZN(n8601) );
  NAND2_X1 U7035 ( .A1(n8601), .A2(n5551), .ZN(n5515) );
  INV_X1 U7036 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U7037 ( .A1(n5137), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5512) );
  NAND2_X1 U7038 ( .A1(n5557), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5511) );
  OAI211_X1 U7039 ( .C1(n8741), .C2(n6356), .A(n5512), .B(n5511), .ZN(n5513)
         );
  INV_X1 U7040 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7041 ( .A1(n5515), .A2(n5514), .ZN(n8423) );
  NOR2_X1 U7042 ( .A1(n8603), .A2(n8611), .ZN(n5517) );
  NAND2_X1 U7043 ( .A1(n8603), .A2(n8611), .ZN(n5516) );
  INV_X1 U7044 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8226) );
  INV_X1 U7045 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8230) );
  MUX2_X1 U7046 ( .A(n8226), .B(n8230), .S(n5902), .Z(n5521) );
  INV_X1 U7047 ( .A(SI_26_), .ZN(n9500) );
  NAND2_X1 U7048 ( .A1(n5521), .A2(n9500), .ZN(n5535) );
  INV_X1 U7049 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7050 ( .A1(n5522), .A2(SI_26_), .ZN(n5523) );
  AND2_X1 U7051 ( .A1(n5535), .A2(n5523), .ZN(n5533) );
  XNOR2_X1 U7052 ( .A(n5534), .B(n5533), .ZN(n8225) );
  NAND2_X1 U7053 ( .A1(n8225), .A2(n6627), .ZN(n5525) );
  OR2_X1 U7054 ( .A1(n5107), .A2(n8226), .ZN(n5524) );
  INV_X1 U7055 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8396) );
  NOR2_X1 U7056 ( .A1(n5526), .A2(n8396), .ZN(n5527) );
  OR2_X1 U7057 ( .A1(n5546), .A2(n5527), .ZN(n8592) );
  NAND2_X1 U7058 ( .A1(n5557), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7059 ( .A1(n5528), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5529) );
  OAI211_X1 U7060 ( .C1(n6621), .C2(n9306), .A(n5530), .B(n5529), .ZN(n5531)
         );
  INV_X1 U7061 ( .A(n8568), .ZN(n8598) );
  NOR2_X1 U7062 ( .A1(n8803), .A2(n8598), .ZN(n5532) );
  NAND2_X1 U7063 ( .A1(n5536), .A2(n5535), .ZN(n5541) );
  INV_X1 U7064 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5543) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5827) );
  MUX2_X1 U7066 ( .A(n5543), .B(n5827), .S(n5902), .Z(n5537) );
  INV_X1 U7067 ( .A(SI_27_), .ZN(n9507) );
  NAND2_X1 U7068 ( .A1(n5537), .A2(n9507), .ZN(n5552) );
  INV_X1 U7069 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U7070 ( .A1(n5538), .A2(SI_27_), .ZN(n5539) );
  AND2_X1 U7071 ( .A1(n5552), .A2(n5539), .ZN(n5540) );
  NAND2_X1 U7072 ( .A1(n5541), .A2(n5540), .ZN(n5553) );
  OR2_X1 U7073 ( .A1(n5541), .A2(n5540), .ZN(n5542) );
  NAND2_X1 U7074 ( .A1(n5553), .A2(n5542), .ZN(n8231) );
  NAND2_X1 U7075 ( .A1(n8231), .A2(n6627), .ZN(n5545) );
  OR2_X1 U7076 ( .A1(n5107), .A2(n5543), .ZN(n5544) );
  INV_X1 U7077 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9503) );
  OR2_X1 U7078 ( .A1(n5546), .A2(n9503), .ZN(n5547) );
  NAND2_X1 U7079 ( .A1(n9503), .A2(n5546), .ZN(n5560) );
  NAND2_X1 U7080 ( .A1(n5547), .A2(n5560), .ZN(n8580) );
  INV_X1 U7081 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8736) );
  NAND2_X1 U7082 ( .A1(n5137), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U7083 ( .A1(n5557), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5548) );
  OAI211_X1 U7084 ( .C1(n8736), .C2(n6356), .A(n5549), .B(n5548), .ZN(n5550)
         );
  NAND2_X1 U7085 ( .A1(n8735), .A2(n8589), .ZN(n6808) );
  INV_X1 U7086 ( .A(n8589), .ZN(n7493) );
  NAND2_X1 U7087 ( .A1(n5553), .A2(n5552), .ZN(n5682) );
  INV_X1 U7088 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5554) );
  INV_X1 U7089 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8237) );
  MUX2_X1 U7090 ( .A(n5554), .B(n8237), .S(n5902), .Z(n5684) );
  XNOR2_X1 U7091 ( .A(n5684), .B(SI_28_), .ZN(n5681) );
  NAND2_X1 U7092 ( .A1(n8234), .A2(n6627), .ZN(n5556) );
  OR2_X1 U7093 ( .A1(n5107), .A2(n5554), .ZN(n5555) );
  NAND2_X1 U7094 ( .A1(n5557), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5565) );
  INV_X1 U7095 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9490) );
  OR2_X1 U7096 ( .A1(n6356), .A2(n9490), .ZN(n5564) );
  INV_X1 U7097 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8561) );
  OR2_X1 U7098 ( .A1(n6621), .A2(n8561), .ZN(n5563) );
  INV_X1 U7099 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5559) );
  INV_X1 U7100 ( .A(n5560), .ZN(n5558) );
  NAND2_X1 U7101 ( .A1(n5559), .A2(n5558), .ZN(n8545) );
  NAND2_X1 U7102 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(n5560), .ZN(n5561) );
  XNOR2_X1 U7103 ( .A(n6347), .B(n8264), .ZN(n5587) );
  NAND2_X1 U7104 ( .A1(n5566), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5567) );
  XNOR2_X1 U7105 ( .A(n5567), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6838) );
  NAND2_X1 U7106 ( .A1(n8535), .A2(n6838), .ZN(n5575) );
  INV_X1 U7107 ( .A(n5568), .ZN(n5572) );
  NAND2_X1 U7108 ( .A1(n5572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5569) );
  XNOR2_X1 U7109 ( .A(n5569), .B(P2_IR_REG_21__SCAN_IN), .ZN(n7499) );
  NAND2_X1 U7110 ( .A1(n5570), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5571) );
  MUX2_X1 U7111 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5571), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n5573) );
  NAND2_X1 U7112 ( .A1(n5573), .A2(n5572), .ZN(n7823) );
  INV_X1 U7113 ( .A(n7823), .ZN(n5667) );
  NAND2_X1 U7114 ( .A1(n7499), .A2(n5667), .ZN(n5574) );
  OR2_X1 U7115 ( .A1(n7138), .A2(n7642), .ZN(n5578) );
  NAND2_X1 U7116 ( .A1(n6962), .A2(n5578), .ZN(n6949) );
  INV_X1 U7117 ( .A(n6949), .ZN(n8569) );
  NAND2_X2 U7118 ( .A1(n6838), .A2(n7499), .ZN(n6959) );
  NAND2_X1 U7119 ( .A1(n8569), .A2(n6788), .ZN(n8718) );
  OR2_X1 U7120 ( .A1(n5579), .A2(n8545), .ZN(n6625) );
  INV_X1 U7121 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5580) );
  OR2_X1 U7122 ( .A1(n6621), .A2(n5580), .ZN(n5583) );
  INV_X1 U7123 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6369) );
  OR2_X1 U7124 ( .A1(n5072), .A2(n6369), .ZN(n5582) );
  INV_X1 U7125 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9371) );
  OR2_X1 U7126 ( .A1(n6356), .A2(n9371), .ZN(n5581) );
  OR2_X1 U7127 ( .A1(n6838), .A2(n7499), .ZN(n10291) );
  INV_X1 U7128 ( .A(n10291), .ZN(n10308) );
  INV_X1 U7129 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U7130 ( .A1(n5616), .A2(n5615), .ZN(n5589) );
  INV_X1 U7131 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5590) );
  NAND2_X1 U7132 ( .A1(n5591), .A2(n5590), .ZN(n5594) );
  INV_X1 U7133 ( .A(P2_B_REG_SCAN_IN), .ZN(n5593) );
  XNOR2_X1 U7134 ( .A(n8287), .B(n5593), .ZN(n5599) );
  NAND2_X1 U7135 ( .A1(n5594), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7136 ( .A1(n4477), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5596) );
  MUX2_X1 U7137 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5596), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5598) );
  INV_X1 U7138 ( .A(n5026), .ZN(n5597) );
  NAND2_X1 U7139 ( .A1(n5598), .A2(n5597), .ZN(n8227) );
  INV_X1 U7140 ( .A(n7009), .ZN(n5601) );
  INV_X1 U7141 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7142 ( .A1(n5601), .A2(n5600), .ZN(n6843) );
  NAND2_X1 U7143 ( .A1(n8227), .A2(n8287), .ZN(n6841) );
  OR2_X1 U7144 ( .A1(n7009), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5603) );
  OR2_X1 U7145 ( .A1(n8218), .A2(n7040), .ZN(n5602) );
  NAND2_X1 U7146 ( .A1(n5669), .A2(n8846), .ZN(n5674) );
  NOR4_X1 U7147 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5612) );
  INV_X1 U7148 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n9411) );
  INV_X1 U7149 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9518) );
  INV_X1 U7150 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n9414) );
  INV_X1 U7151 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n9327) );
  NAND4_X1 U7152 ( .A1(n9411), .A2(n9518), .A3(n9414), .A4(n9327), .ZN(n5609)
         );
  NOR4_X1 U7153 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5607) );
  NOR4_X1 U7154 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5606) );
  NOR4_X1 U7155 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5605) );
  NOR4_X1 U7156 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5604) );
  NAND4_X1 U7157 ( .A1(n5607), .A2(n5606), .A3(n5605), .A4(n5604), .ZN(n5608)
         );
  NOR4_X1 U7158 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n5609), .A4(n5608), .ZN(n5611) );
  NOR4_X1 U7159 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5610) );
  AND3_X1 U7160 ( .A1(n5612), .A2(n5611), .A3(n5610), .ZN(n5613) );
  OR2_X1 U7161 ( .A1(n7009), .A2(n5613), .ZN(n5673) );
  INV_X1 U7162 ( .A(n5673), .ZN(n5619) );
  OR2_X1 U7163 ( .A1(n5674), .A2(n5619), .ZN(n6937) );
  NOR2_X1 U7164 ( .A1(n8227), .A2(n8287), .ZN(n5614) );
  NAND2_X1 U7165 ( .A1(n8218), .A2(n5614), .ZN(n7169) );
  XNOR2_X1 U7166 ( .A(n5616), .B(n5615), .ZN(n6960) );
  AND2_X1 U7167 ( .A1(n6960), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6965) );
  NAND2_X1 U7168 ( .A1(n7169), .A2(n6965), .ZN(n8845) );
  NOR2_X1 U7169 ( .A1(n6937), .A2(n8845), .ZN(n6931) );
  OR2_X1 U7170 ( .A1(n6844), .A2(n6959), .ZN(n6948) );
  INV_X1 U7171 ( .A(n7499), .ZN(n7853) );
  AND3_X1 U7172 ( .A1(n6838), .A2(n7853), .A3(n5667), .ZN(n5617) );
  NAND2_X1 U7173 ( .A1(n8535), .A2(n5617), .ZN(n6940) );
  NAND2_X1 U7174 ( .A1(n6948), .A2(n6940), .ZN(n5618) );
  NAND2_X1 U7175 ( .A1(n6931), .A2(n5618), .ZN(n5623) );
  NOR2_X1 U7176 ( .A1(n8846), .A2(n5619), .ZN(n5620) );
  INV_X1 U7177 ( .A(n5669), .ZN(n7292) );
  INV_X1 U7178 ( .A(n8845), .ZN(n7010) );
  AND2_X1 U7179 ( .A1(n8535), .A2(n7823), .ZN(n7500) );
  OR2_X1 U7180 ( .A1(n7500), .A2(n10291), .ZN(n8608) );
  AND2_X1 U7181 ( .A1(n10291), .A2(n6959), .ZN(n5621) );
  NAND2_X1 U7182 ( .A1(n6940), .A2(n5621), .ZN(n6923) );
  NAND2_X1 U7183 ( .A1(n8608), .A2(n6923), .ZN(n6936) );
  NAND2_X1 U7184 ( .A1(n6951), .A2(n6936), .ZN(n5622) );
  INV_X2 U7185 ( .A(n10311), .ZN(n10309) );
  MUX2_X1 U7186 ( .A(n5624), .B(n5677), .S(n10309), .Z(n5666) );
  NOR2_X1 U7187 ( .A1(n5625), .A2(n8784), .ZN(n6847) );
  INV_X1 U7188 ( .A(n6847), .ZN(n7502) );
  OR2_X1 U7189 ( .A1(n7505), .A2(n7502), .ZN(n5626) );
  NAND2_X1 U7190 ( .A1(n5626), .A2(n6674), .ZN(n7573) );
  INV_X1 U7191 ( .A(n7576), .ZN(n6633) );
  NAND2_X1 U7192 ( .A1(n7573), .A2(n6633), .ZN(n5628) );
  INV_X1 U7193 ( .A(n10256), .ZN(n5627) );
  NAND2_X1 U7194 ( .A1(n6852), .A2(n5627), .ZN(n6667) );
  NAND2_X1 U7195 ( .A1(n5628), .A2(n6667), .ZN(n7555) );
  XNOR2_X1 U7196 ( .A(n4444), .B(n10260), .ZN(n7554) );
  NAND2_X1 U7197 ( .A1(n7555), .A2(n7554), .ZN(n7616) );
  NAND2_X1 U7198 ( .A1(n7622), .A2(n10260), .ZN(n7615) );
  NAND2_X1 U7199 ( .A1(n7608), .A2(n10266), .ZN(n7749) );
  NAND2_X1 U7200 ( .A1(n7761), .A2(n10271), .ZN(n6690) );
  AND2_X1 U7201 ( .A1(n7749), .A2(n6690), .ZN(n5630) );
  NAND2_X1 U7202 ( .A1(n8436), .A2(n7611), .ZN(n6693) );
  INV_X1 U7203 ( .A(n6693), .ZN(n5629) );
  AND2_X1 U7204 ( .A1(n7615), .A2(n4472), .ZN(n5631) );
  NAND2_X1 U7205 ( .A1(n7616), .A2(n5631), .ZN(n7675) );
  NAND2_X1 U7206 ( .A1(n7747), .A2(n6693), .ZN(n5633) );
  NAND2_X1 U7207 ( .A1(n4472), .A2(n5633), .ZN(n7674) );
  INV_X1 U7208 ( .A(n7674), .ZN(n5634) );
  INV_X1 U7209 ( .A(n6687), .ZN(n6697) );
  NAND2_X1 U7210 ( .A1(n8435), .A2(n10276), .ZN(n6695) );
  NAND2_X1 U7211 ( .A1(n6697), .A2(n6695), .ZN(n7678) );
  NOR2_X1 U7212 ( .A1(n5634), .A2(n7678), .ZN(n5635) );
  AOI21_X1 U7213 ( .B1(n7675), .B2(n5635), .A(n6687), .ZN(n8245) );
  NAND2_X1 U7214 ( .A1(n8245), .A2(n8246), .ZN(n8244) );
  NAND2_X1 U7215 ( .A1(n6702), .A2(n7800), .ZN(n6712) );
  INV_X1 U7216 ( .A(n6712), .ZN(n5636) );
  INV_X1 U7217 ( .A(n6710), .ZN(n6707) );
  OR2_X1 U7218 ( .A1(n6864), .A2(n7884), .ZN(n6714) );
  NAND2_X1 U7219 ( .A1(n6864), .A2(n7884), .ZN(n6711) );
  NAND2_X1 U7220 ( .A1(n7862), .A2(n7867), .ZN(n7861) );
  NAND2_X1 U7221 ( .A1(n7861), .A2(n6714), .ZN(n7922) );
  OR2_X1 U7222 ( .A1(n10301), .A2(n7931), .ZN(n6871) );
  NAND2_X1 U7223 ( .A1(n6721), .A2(n6871), .ZN(n8025) );
  INV_X1 U7224 ( .A(n8430), .ZN(n7932) );
  OR2_X1 U7225 ( .A1(n8127), .A2(n7932), .ZN(n6730) );
  INV_X1 U7226 ( .A(n6730), .ZN(n5640) );
  OR2_X1 U7227 ( .A1(n8025), .A2(n5640), .ZN(n7993) );
  INV_X1 U7228 ( .A(n6734), .ZN(n5642) );
  OR2_X1 U7229 ( .A1(n7993), .A2(n5642), .ZN(n8041) );
  OR2_X1 U7230 ( .A1(n8300), .A2(n8413), .ZN(n6740) );
  INV_X1 U7231 ( .A(n6740), .ZN(n5643) );
  OR2_X1 U7232 ( .A1(n8041), .A2(n5643), .ZN(n5637) );
  NOR2_X1 U7233 ( .A1(n7922), .A2(n5637), .ZN(n5639) );
  NAND2_X1 U7234 ( .A1(n8300), .A2(n8413), .ZN(n6739) );
  NOR2_X1 U7235 ( .A1(n5639), .A2(n5638), .ZN(n5644) );
  NAND2_X1 U7236 ( .A1(n10307), .A2(n8134), .ZN(n6722) );
  NAND2_X1 U7237 ( .A1(n10301), .A2(n7931), .ZN(n7924) );
  NAND2_X1 U7238 ( .A1(n6722), .A2(n7924), .ZN(n6720) );
  XNOR2_X1 U7239 ( .A(n8127), .B(n8430), .ZN(n8035) );
  NAND2_X1 U7240 ( .A1(n5641), .A2(n6730), .ZN(n7994) );
  INV_X1 U7241 ( .A(n8105), .ZN(n5645) );
  NAND2_X1 U7242 ( .A1(n8405), .A2(n8161), .ZN(n6632) );
  OR2_X1 U7243 ( .A1(n8405), .A2(n8161), .ZN(n8154) );
  NAND2_X1 U7244 ( .A1(n6756), .A2(n8154), .ZN(n6743) );
  INV_X1 U7245 ( .A(n6743), .ZN(n5646) );
  NAND2_X1 U7246 ( .A1(n5647), .A2(n6744), .ZN(n8705) );
  INV_X1 U7247 ( .A(n8705), .ZN(n5649) );
  INV_X1 U7248 ( .A(n8703), .ZN(n8774) );
  NAND2_X1 U7249 ( .A1(n8703), .A2(n8721), .ZN(n6751) );
  NAND2_X1 U7250 ( .A1(n6760), .A2(n6751), .ZN(n8704) );
  AND2_X1 U7251 ( .A1(n8649), .A2(n6780), .ZN(n5653) );
  INV_X1 U7252 ( .A(n6780), .ZN(n5652) );
  NAND2_X1 U7253 ( .A1(n6777), .A2(n8650), .ZN(n6772) );
  INV_X1 U7254 ( .A(n6772), .ZN(n5651) );
  INV_X1 U7255 ( .A(n8749), .ZN(n5654) );
  NAND2_X1 U7256 ( .A1(n8749), .A2(n8637), .ZN(n6786) );
  NAND2_X1 U7257 ( .A1(n8744), .A2(n8621), .ZN(n6791) );
  OR2_X1 U7258 ( .A1(n8744), .A2(n8621), .ZN(n6792) );
  INV_X1 U7259 ( .A(n8603), .ZN(n8809) );
  AND2_X1 U7260 ( .A1(n8603), .A2(n8423), .ZN(n6796) );
  INV_X1 U7261 ( .A(n6796), .ZN(n6631) );
  NAND2_X1 U7262 ( .A1(n5655), .A2(n6631), .ZN(n8585) );
  INV_X1 U7263 ( .A(n8585), .ZN(n5656) );
  NAND2_X1 U7264 ( .A1(n5656), .A2(n6799), .ZN(n8575) );
  NAND2_X1 U7265 ( .A1(n8803), .A2(n8568), .ZN(n8574) );
  AND2_X1 U7266 ( .A1(n6801), .A2(n8574), .ZN(n5657) );
  NAND2_X1 U7267 ( .A1(n8575), .A2(n5657), .ZN(n8579) );
  INV_X1 U7268 ( .A(n5658), .ZN(n5659) );
  INV_X1 U7269 ( .A(n8264), .ZN(n6651) );
  NAND2_X1 U7270 ( .A1(n5659), .A2(n6651), .ZN(n5660) );
  OR2_X1 U7271 ( .A1(n6844), .A2(n7853), .ZN(n5662) );
  INV_X1 U7272 ( .A(n6838), .ZN(n7941) );
  OR2_X1 U7273 ( .A1(n8535), .A2(n7941), .ZN(n5661) );
  NAND2_X1 U7274 ( .A1(n5662), .A2(n5661), .ZN(n5668) );
  AND2_X1 U7275 ( .A1(n5668), .A2(n6948), .ZN(n7944) );
  NAND2_X1 U7276 ( .A1(n7500), .A2(n7941), .ZN(n10297) );
  INV_X1 U7277 ( .A(n10297), .ZN(n10272) );
  OR2_X1 U7278 ( .A1(n7944), .A2(n10272), .ZN(n10287) );
  INV_X1 U7279 ( .A(n10287), .ZN(n10303) );
  INV_X1 U7280 ( .A(n8841), .ZN(n5663) );
  NAND2_X1 U7281 ( .A1(n5666), .A2(n5665), .ZN(P2_U3455) );
  AOI21_X1 U7282 ( .B1(n5668), .B2(n5667), .A(n6788), .ZN(n5670) );
  NAND2_X1 U7283 ( .A1(n5669), .A2(n5670), .ZN(n7293) );
  NOR2_X1 U7284 ( .A1(n10297), .A2(n7499), .ZN(n6932) );
  INV_X1 U7285 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U7286 ( .A1(n8846), .A2(n5671), .ZN(n7294) );
  OAI21_X1 U7287 ( .B1(n7293), .B2(n6932), .A(n7294), .ZN(n5676) );
  AND2_X1 U7288 ( .A1(n6844), .A2(n6788), .ZN(n6934) );
  NOR2_X1 U7289 ( .A1(n8845), .A2(n6934), .ZN(n5672) );
  AND2_X1 U7290 ( .A1(n5673), .A2(n5672), .ZN(n7295) );
  AND2_X1 U7291 ( .A1(n5674), .A2(n7295), .ZN(n5675) );
  AND2_X2 U7292 ( .A1(n5676), .A2(n5675), .ZN(n10325) );
  MUX2_X1 U7293 ( .A(n9490), .B(n5677), .S(n10325), .Z(n5680) );
  NAND2_X1 U7294 ( .A1(n10325), .A2(n10287), .ZN(n8778) );
  NAND2_X1 U7295 ( .A1(n5664), .A2(n5678), .ZN(n5679) );
  NAND2_X1 U7296 ( .A1(n5680), .A2(n5679), .ZN(P2_U3487) );
  NAND2_X1 U7297 ( .A1(n5682), .A2(n5681), .ZN(n5686) );
  INV_X1 U7298 ( .A(SI_28_), .ZN(n5683) );
  NAND2_X1 U7299 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  INV_X1 U7300 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8241) );
  INV_X1 U7301 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9700) );
  MUX2_X1 U7302 ( .A(n8241), .B(n9700), .S(n5902), .Z(n5689) );
  INV_X1 U7303 ( .A(n5832), .ZN(n5687) );
  NAND2_X1 U7304 ( .A1(n5687), .A2(SI_29_), .ZN(n5693) );
  INV_X1 U7305 ( .A(n5688), .ZN(n5691) );
  INV_X1 U7306 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7307 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7308 ( .A1(n5693), .A2(n5692), .ZN(n5901) );
  INV_X1 U7309 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8849) );
  INV_X1 U7310 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8276) );
  MUX2_X1 U7311 ( .A(n8849), .B(n8276), .S(n5902), .Z(n5694) );
  INV_X1 U7312 ( .A(SI_30_), .ZN(n9413) );
  NAND2_X1 U7313 ( .A1(n5694), .A2(n9413), .ZN(n5899) );
  INV_X1 U7314 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7315 ( .A1(n5695), .A2(SI_30_), .ZN(n5696) );
  NAND2_X1 U7316 ( .A1(n5899), .A2(n5696), .ZN(n5900) );
  NOR2_X1 U7317 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5700) );
  NOR2_X2 U7319 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5698) );
  NOR2_X2 U7320 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5697) );
  AND4_X2 U7321 ( .A1(n5700), .A2(n5699), .A3(n5698), .A4(n5697), .ZN(n5708)
         );
  NAND2_X1 U7322 ( .A1(n5756), .A2(n5701), .ZN(n5743) );
  INV_X1 U7323 ( .A(n5743), .ZN(n5707) );
  INV_X1 U7325 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5704) );
  INV_X1 U7326 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5703) );
  INV_X1 U7327 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5702) );
  AND4_X2 U7328 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n5706)
         );
  NAND3_X2 U7329 ( .A1(n5708), .A2(n5707), .A3(n5706), .ZN(n5835) );
  NOR2_X1 U7330 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5712) );
  NOR2_X1 U7331 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5711) );
  NOR2_X1 U7332 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5710) );
  NOR2_X1 U7333 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5709) );
  NAND4_X1 U7334 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n5713)
         );
  INV_X1 U7335 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U7336 ( .A1(n5717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  INV_X1 U7337 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U7338 ( .A1(n5872), .A2(n5871), .ZN(n5714) );
  INV_X1 U7339 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7340 ( .A1(n5720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5719) );
  MUX2_X1 U7341 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5719), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5721) );
  NAND2_X1 U7342 ( .A1(n8272), .A2(n5722), .ZN(n5724) );
  OR2_X1 U7343 ( .A1(n5754), .A2(n8276), .ZN(n5723) );
  NAND2_X1 U7344 ( .A1(n8225), .A2(n5722), .ZN(n5726) );
  OR2_X1 U7345 ( .A1(n5754), .A2(n8230), .ZN(n5725) );
  INV_X1 U7346 ( .A(n9643), .ZN(n9214) );
  NAND2_X1 U7347 ( .A1(n8219), .A2(n5722), .ZN(n5728) );
  OR2_X1 U7348 ( .A1(n5754), .A2(n8224), .ZN(n5727) );
  NAND2_X1 U7349 ( .A1(n8152), .A2(n5722), .ZN(n5730) );
  OR2_X1 U7350 ( .A1(n5754), .A2(n8153), .ZN(n5729) );
  NAND2_X1 U7351 ( .A1(n8022), .A2(n5722), .ZN(n5732) );
  OR2_X1 U7352 ( .A1(n5754), .A2(n9354), .ZN(n5731) );
  INV_X1 U7353 ( .A(n9659), .ZN(n9564) );
  NAND2_X1 U7354 ( .A1(n7820), .A2(n5722), .ZN(n5734) );
  OR2_X1 U7355 ( .A1(n5754), .A2(n7773), .ZN(n5733) );
  NAND2_X1 U7356 ( .A1(n7743), .A2(n5722), .ZN(n5739) );
  NAND2_X1 U7357 ( .A1(n5835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5740) );
  INV_X1 U7358 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7359 ( .A1(n5740), .A2(n5837), .ZN(n5735) );
  INV_X1 U7360 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7361 ( .A1(n5818), .A2(n5838), .ZN(n5736) );
  XNOR2_X2 U7362 ( .A(n5737), .B(P1_IR_REG_19__SCAN_IN), .ZN(n6376) );
  AOI22_X1 U7363 ( .A1(n4450), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6376), .B2(
        n4443), .ZN(n5738) );
  NAND2_X1 U7364 ( .A1(n7528), .A2(n5722), .ZN(n5742) );
  XNOR2_X1 U7365 ( .A(n5740), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9100) );
  AOI22_X1 U7366 ( .A1(n4450), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n4443), .B2(
        n9100), .ZN(n5741) );
  NAND2_X1 U7367 ( .A1(n7238), .A2(n5722), .ZN(n5747) );
  NOR2_X1 U7368 ( .A1(n5769), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5773) );
  NOR2_X1 U7369 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5744) );
  NAND2_X1 U7370 ( .A1(n5773), .A2(n5744), .ZN(n5785) );
  NOR2_X1 U7371 ( .A1(n5788), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5791) );
  NOR2_X1 U7372 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5745) );
  NAND2_X1 U7373 ( .A1(n5791), .A2(n5745), .ZN(n5800) );
  OR2_X1 U7374 ( .A1(n5802), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7375 ( .A1(n5814), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5806) );
  XNOR2_X1 U7376 ( .A(n5806), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U7377 ( .A1(n9893), .A2(n4443), .B1(n4450), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5746) );
  INV_X1 U7378 ( .A(n6021), .ZN(n8217) );
  NAND2_X1 U7379 ( .A1(n7222), .A2(n5722), .ZN(n5750) );
  NAND2_X1 U7380 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U7381 ( .A(n5748), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9881) );
  AOI22_X1 U7382 ( .A1(n9881), .A2(n4443), .B1(n4450), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5749) );
  OAI211_X2 U7383 ( .C1(n5780), .C2(n6978), .A(n5751), .B(n4980), .ZN(n7273)
         );
  INV_X1 U7384 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9013) );
  INV_X1 U7385 ( .A(SI_0_), .ZN(n5752) );
  NOR2_X1 U7386 ( .A1(n5065), .A2(n5752), .ZN(n5753) );
  XNOR2_X1 U7387 ( .A(n5753), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n6967) );
  MUX2_X1 U7388 ( .A(n9013), .B(n6967), .S(n6983), .Z(n9976) );
  NAND2_X1 U7389 ( .A1(n9992), .A2(n9976), .ZN(n9974) );
  OR2_X1 U7390 ( .A1(n5754), .A2(n6969), .ZN(n5757) );
  OR2_X1 U7391 ( .A1(n5756), .A2(n5755), .ZN(n5759) );
  INV_X1 U7392 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5758) );
  XNOR2_X1 U7393 ( .A(n5759), .B(n5758), .ZN(n7096) );
  OR2_X1 U7394 ( .A1(n6973), .A2(n5780), .ZN(n5764) );
  NAND2_X1 U7395 ( .A1(n5759), .A2(n5758), .ZN(n5760) );
  NAND2_X1 U7396 ( .A1(n5760), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5761) );
  XNOR2_X1 U7397 ( .A(n5761), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U7398 ( .A1(n4443), .A2(n9038), .ZN(n5763) );
  OR2_X1 U7399 ( .A1(n5754), .A2(n6972), .ZN(n5762) );
  AND3_X2 U7400 ( .A1(n5764), .A2(n5763), .A3(n5762), .ZN(n10007) );
  NAND2_X1 U7401 ( .A1(n9955), .A2(n10007), .ZN(n7334) );
  NAND2_X1 U7402 ( .A1(n5743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5765) );
  MUX2_X1 U7403 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5765), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5766) );
  NAND2_X1 U7404 ( .A1(n5769), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5770) );
  XNOR2_X1 U7405 ( .A(n5770), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U7406 ( .A1(n4450), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n4443), .B2(
        n9835), .ZN(n5771) );
  NAND2_X1 U7407 ( .A1(n5772), .A2(n5771), .ZN(n7361) );
  OR2_X2 U7408 ( .A1(n7335), .A2(n7361), .ZN(n9939) );
  OR2_X1 U7409 ( .A1(n6996), .A2(n5780), .ZN(n5779) );
  OR2_X1 U7410 ( .A1(n5773), .A2(n5755), .ZN(n5776) );
  INV_X1 U7411 ( .A(n5776), .ZN(n5774) );
  NAND2_X1 U7412 ( .A1(n5774), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5777) );
  INV_X1 U7413 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7414 ( .A1(n5776), .A2(n5775), .ZN(n5781) );
  AOI22_X1 U7415 ( .A1(n4450), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n4443), .B2(
        n9845), .ZN(n5778) );
  NAND2_X1 U7416 ( .A1(n5779), .A2(n5778), .ZN(n7407) );
  OR2_X1 U7417 ( .A1(n7006), .A2(n5780), .ZN(n5784) );
  NAND2_X1 U7418 ( .A1(n5781), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5782) );
  XNOR2_X1 U7419 ( .A(n5782), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9716) );
  AOI22_X1 U7420 ( .A1(n4450), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n4443), .B2(
        n9716), .ZN(n5783) );
  NAND2_X1 U7421 ( .A1(n7521), .A2(n10031), .ZN(n7520) );
  NAND2_X1 U7422 ( .A1(n5785), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5786) );
  XNOR2_X1 U7423 ( .A(n5786), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9731) );
  AOI22_X1 U7424 ( .A1(n4450), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n4443), .B2(
        n9731), .ZN(n5787) );
  NAND2_X1 U7425 ( .A1(n5788), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5789) );
  XNOR2_X1 U7426 ( .A(n5789), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7434) );
  AOI22_X1 U7427 ( .A1(n4450), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n4443), .B2(
        n7434), .ZN(n5790) );
  NAND2_X1 U7428 ( .A1(n7031), .A2(n5722), .ZN(n5793) );
  OR2_X1 U7429 ( .A1(n5791), .A2(n5755), .ZN(n5795) );
  XNOR2_X1 U7430 ( .A(n5795), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U7431 ( .A1(n4450), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n4443), .B2(
        n9712), .ZN(n5792) );
  NAND2_X1 U7432 ( .A1(n5793), .A2(n5792), .ZN(n7961) );
  INV_X1 U7433 ( .A(n7961), .ZN(n10058) );
  NAND2_X1 U7434 ( .A1(n7053), .A2(n5722), .ZN(n5799) );
  INV_X1 U7435 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7436 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7437 ( .A1(n5796), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5797) );
  XNOR2_X1 U7438 ( .A(n5797), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U7439 ( .A1(n4443), .A2(n9862), .B1(n4450), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n5798) );
  NAND2_X1 U7440 ( .A1(n7072), .A2(n5722), .ZN(n5805) );
  NAND2_X1 U7441 ( .A1(n5800), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5801) );
  MUX2_X1 U7442 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5801), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5803) );
  AND2_X1 U7443 ( .A1(n5803), .A2(n5802), .ZN(n9062) );
  AOI22_X1 U7444 ( .A1(n4450), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9062), .B2(
        n4443), .ZN(n5804) );
  NAND2_X1 U7445 ( .A1(n7340), .A2(n5722), .ZN(n5810) );
  INV_X1 U7446 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7447 ( .A1(n5806), .A2(n5812), .ZN(n5807) );
  NAND2_X1 U7448 ( .A1(n5807), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5808) );
  XNOR2_X1 U7449 ( .A(n5808), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9905) );
  AOI22_X1 U7450 ( .A1(n9905), .A2(n4443), .B1(n4450), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7451 ( .A1(n7495), .A2(n5722), .ZN(n5817) );
  INV_X1 U7452 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7453 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  OAI21_X1 U7454 ( .B1(n5814), .B2(n5813), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5815) );
  XNOR2_X1 U7455 ( .A(n5815), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9084) );
  AOI22_X1 U7456 ( .A1(n9084), .A2(n4443), .B1(n4450), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5816) );
  NAND2_X1 U7457 ( .A1(n9757), .A2(n8079), .ZN(n8146) );
  NAND2_X1 U7458 ( .A1(n7629), .A2(n5722), .ZN(n5822) );
  XNOR2_X1 U7459 ( .A(n5818), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U7460 ( .A1(n4450), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n4443), .B2(
        n9920), .ZN(n5821) );
  NAND2_X1 U7461 ( .A1(n7824), .A2(n5722), .ZN(n5824) );
  OR2_X1 U7462 ( .A1(n5754), .A2(n7825), .ZN(n5823) );
  NAND2_X1 U7463 ( .A1(n7936), .A2(n5722), .ZN(n5826) );
  OR2_X1 U7464 ( .A1(n5754), .A2(n7938), .ZN(n5825) );
  NAND2_X1 U7465 ( .A1(n9564), .A2(n9583), .ZN(n9559) );
  OR2_X2 U7466 ( .A1(n9655), .A2(n9559), .ZN(n9545) );
  NAND2_X1 U7467 ( .A1(n9214), .A2(n9226), .ZN(n9213) );
  NAND2_X1 U7468 ( .A1(n8231), .A2(n5722), .ZN(n5829) );
  OR2_X1 U7469 ( .A1(n5754), .A2(n5827), .ZN(n5828) );
  NAND2_X1 U7470 ( .A1(n8234), .A2(n5722), .ZN(n5831) );
  OR2_X1 U7471 ( .A1(n5754), .A2(n8237), .ZN(n5830) );
  OR2_X1 U7472 ( .A1(n5754), .A2(n9700), .ZN(n5833) );
  INV_X1 U7473 ( .A(n9113), .ZN(n5849) );
  INV_X1 U7474 ( .A(n5835), .ZN(n5839) );
  INV_X1 U7475 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5836) );
  INV_X1 U7476 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7477 ( .A1(n5843), .A2(n5840), .ZN(n5867) );
  NAND2_X1 U7478 ( .A1(n5867), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5841) );
  INV_X1 U7479 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5865) );
  OR2_X1 U7480 ( .A1(n5841), .A2(n5865), .ZN(n5842) );
  NAND2_X1 U7481 ( .A1(n5841), .A2(n5865), .ZN(n5877) );
  INV_X1 U7482 ( .A(n6374), .ZN(n7826) );
  AND2_X1 U7483 ( .A1(n7937), .A2(n7826), .ZN(n5850) );
  NAND2_X1 U7484 ( .A1(n5845), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  MUX2_X1 U7485 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5846), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5848) );
  INV_X1 U7486 ( .A(n6593), .ZN(n7022) );
  INV_X1 U7487 ( .A(n9612), .ZN(n9975) );
  OAI211_X1 U7488 ( .C1(n4636), .C2(n4670), .A(n5849), .B(n9975), .ZN(n9121)
         );
  NAND2_X1 U7489 ( .A1(n5850), .A2(n7017), .ZN(n10076) );
  XNOR2_X2 U7490 ( .A(n5851), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5910) );
  XNOR2_X2 U7491 ( .A(n5852), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5909) );
  INV_X1 U7492 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7493 ( .A1(n4442), .A2(n5853), .ZN(n5856) );
  INV_X1 U7494 ( .A(n5909), .ZN(n9701) );
  INV_X1 U7495 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9115) );
  OR2_X1 U7496 ( .A1(n4449), .A2(n9115), .ZN(n5855) );
  INV_X1 U7497 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9438) );
  OR2_X1 U7498 ( .A1(n5919), .A2(n9438), .ZN(n5854) );
  AND3_X1 U7499 ( .A1(n5856), .A2(n5855), .A3(n5854), .ZN(n6139) );
  INV_X1 U7500 ( .A(n7937), .ZN(n6375) );
  AND2_X1 U7501 ( .A1(n6375), .A2(n6374), .ZN(n6981) );
  NAND2_X1 U7502 ( .A1(n6981), .A2(n8238), .ZN(n8972) );
  INV_X1 U7503 ( .A(P1_B_REG_SCAN_IN), .ZN(n5858) );
  NOR2_X1 U7504 ( .A1(n4451), .A2(n5858), .ZN(n5859) );
  OR2_X1 U7505 ( .A1(n8972), .A2(n5859), .ZN(n9138) );
  OR2_X1 U7506 ( .A1(n6139), .A2(n9138), .ZN(n9624) );
  NAND2_X1 U7507 ( .A1(n4495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5863) );
  XNOR2_X1 U7508 ( .A(n5863), .B(n5862), .ZN(n8223) );
  NAND2_X1 U7509 ( .A1(n8223), .A2(P1_B_REG_SCAN_IN), .ZN(n5870) );
  INV_X1 U7510 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7511 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  INV_X1 U7512 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5868) );
  MUX2_X1 U7513 ( .A(P1_B_REG_SCAN_IN), .B(n5870), .S(n5876), .Z(n5874) );
  XNOR2_X1 U7514 ( .A(n5872), .B(n5871), .ZN(n8229) );
  INV_X1 U7515 ( .A(n8229), .ZN(n5873) );
  NAND2_X1 U7516 ( .A1(n5874), .A2(n5873), .ZN(n9689) );
  NAND2_X1 U7517 ( .A1(n8229), .A2(n8223), .ZN(n9691) );
  OAI21_X1 U7518 ( .B1(n9689), .B2(P1_D_REG_1__SCAN_IN), .A(n9691), .ZN(n5894)
         );
  NAND2_X1 U7519 ( .A1(n5877), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7520 ( .A(n5878), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6329) );
  INV_X1 U7521 ( .A(n6329), .ZN(n6982) );
  NAND3_X1 U7522 ( .A1(n6379), .A2(P1_STATE_REG_SCAN_IN), .A3(n6982), .ZN(
        n6980) );
  NAND2_X1 U7523 ( .A1(n6981), .A2(n7017), .ZN(n6598) );
  INV_X1 U7524 ( .A(n6598), .ZN(n5879) );
  NOR2_X1 U7525 ( .A1(n6980), .A2(n5879), .ZN(n7268) );
  NOR2_X1 U7526 ( .A1(n9612), .A2(n5880), .ZN(n6594) );
  INV_X1 U7527 ( .A(n6594), .ZN(n5893) );
  NOR4_X1 U7528 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n5884) );
  NOR4_X1 U7529 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5883) );
  NOR4_X1 U7530 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n5882) );
  NOR4_X1 U7531 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5881) );
  AND4_X1 U7532 ( .A1(n5884), .A2(n5883), .A3(n5882), .A4(n5881), .ZN(n5890)
         );
  NOR2_X1 U7533 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .ZN(
        n5888) );
  NOR4_X1 U7534 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5887) );
  NOR4_X1 U7535 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5886) );
  NOR4_X1 U7536 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5885) );
  AND4_X1 U7537 ( .A1(n5888), .A2(n5887), .A3(n5886), .A4(n5885), .ZN(n5889)
         );
  NAND2_X1 U7538 ( .A1(n5890), .A2(n5889), .ZN(n6585) );
  INV_X1 U7539 ( .A(n6585), .ZN(n5891) );
  OR2_X1 U7540 ( .A1(n9689), .A2(n5891), .ZN(n5892) );
  NAND4_X1 U7541 ( .A1(n5894), .A2(n7268), .A3(n5893), .A4(n5892), .ZN(n7013)
         );
  OR2_X1 U7542 ( .A1(n9689), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7543 ( .A1(n5876), .A2(n8229), .ZN(n9692) );
  NAND2_X1 U7544 ( .A1(n5895), .A2(n9692), .ZN(n7267) );
  INV_X1 U7545 ( .A(n7267), .ZN(n5896) );
  INV_X2 U7546 ( .A(n10090), .ZN(n10092) );
  NAND2_X1 U7547 ( .A1(n9627), .A2(n10092), .ZN(n5898) );
  INV_X1 U7548 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5897) );
  INV_X1 U7549 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5903) );
  INV_X1 U7550 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9694) );
  MUX2_X1 U7551 ( .A(n5903), .B(n9694), .S(n5902), .Z(n5904) );
  XNOR2_X1 U7552 ( .A(n5904), .B(SI_31_), .ZN(n5905) );
  NAND2_X1 U7553 ( .A1(n9698), .A2(n5722), .ZN(n5908) );
  OR2_X1 U7554 ( .A1(n5754), .A2(n9694), .ZN(n5907) );
  NAND2_X1 U7555 ( .A1(n6108), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5917) );
  INV_X1 U7556 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9307) );
  OR2_X1 U7557 ( .A1(n5919), .A2(n9307), .ZN(n5916) );
  INV_X1 U7558 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U7559 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n6115) );
  NAND2_X1 U7560 ( .A1(n6116), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6076) );
  INV_X1 U7561 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6051) );
  INV_X1 U7562 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U7563 ( .A1(n6067), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6069) );
  INV_X1 U7564 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6035) );
  INV_X1 U7565 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7442) );
  NAND2_X1 U7566 ( .A1(n6030), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7567 ( .A1(n6014), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6008) );
  AND2_X1 U7568 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n5911) );
  NAND2_X1 U7569 ( .A1(n6003), .A2(n5911), .ZN(n5992) );
  INV_X1 U7570 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U7571 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5912) );
  NAND2_X1 U7572 ( .A1(n5959), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5951) );
  INV_X1 U7573 ( .A(n5951), .ZN(n5946) );
  NAND2_X1 U7574 ( .A1(n5936), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5938) );
  INV_X1 U7575 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9318) );
  NOR2_X1 U7576 ( .A1(n5938), .A2(n9318), .ZN(n5922) );
  NAND2_X1 U7577 ( .A1(n5922), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9171) );
  OR2_X1 U7578 ( .A1(n6102), .A2(n9171), .ZN(n5915) );
  INV_X1 U7579 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7580 ( .A1(n4449), .A2(n5913), .ZN(n5914) );
  AND4_X1 U7581 ( .A1(n5917), .A2(n5916), .A3(n5915), .A4(n5914), .ZN(n7257)
         );
  NAND2_X1 U7582 ( .A1(n5918), .A2(n7257), .ZN(n6263) );
  INV_X1 U7583 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9329) );
  NAND2_X1 U7584 ( .A1(n6118), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7585 ( .A1(n6004), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5920) );
  OAI211_X1 U7586 ( .C1(n4441), .C2(n9329), .A(n5921), .B(n5920), .ZN(n8992)
         );
  INV_X1 U7587 ( .A(n8992), .ZN(n9139) );
  OR2_X1 U7588 ( .A1(n6269), .A2(n9139), .ZN(n6324) );
  NAND2_X1 U7589 ( .A1(n6118), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5928) );
  INV_X1 U7590 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9376) );
  OR2_X1 U7591 ( .A1(n4442), .A2(n9376), .ZN(n5927) );
  INV_X1 U7592 ( .A(n5922), .ZN(n5931) );
  INV_X1 U7593 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7594 ( .A1(n5931), .A2(n5923), .ZN(n5924) );
  NAND2_X1 U7595 ( .A1(n9171), .A2(n5924), .ZN(n9184) );
  OR2_X1 U7596 ( .A1(n6102), .A2(n9184), .ZN(n5926) );
  INV_X1 U7597 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9185) );
  OR2_X1 U7598 ( .A1(n4449), .A2(n9185), .ZN(n5925) );
  OR2_X1 U7599 ( .A1(n9633), .A2(n9167), .ZN(n6257) );
  NAND2_X1 U7600 ( .A1(n9633), .A2(n9167), .ZN(n9136) );
  NAND2_X1 U7601 ( .A1(n6118), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5935) );
  INV_X1 U7602 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7603 ( .A1(n4441), .A2(n5929), .ZN(n5934) );
  NAND2_X1 U7604 ( .A1(n5938), .A2(n9318), .ZN(n5930) );
  NAND2_X1 U7605 ( .A1(n5931), .A2(n5930), .ZN(n9204) );
  OR2_X1 U7606 ( .A1(n6102), .A2(n9204), .ZN(n5933) );
  INV_X1 U7607 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9205) );
  OR2_X1 U7608 ( .A1(n4449), .A2(n9205), .ZN(n5932) );
  OR2_X1 U7609 ( .A1(n9640), .A2(n8993), .ZN(n6250) );
  NAND2_X1 U7610 ( .A1(n9640), .A2(n8993), .ZN(n9135) );
  NAND2_X1 U7611 ( .A1(n6108), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5943) );
  INV_X1 U7612 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9331) );
  OR2_X1 U7613 ( .A1(n5919), .A2(n9331), .ZN(n5942) );
  INV_X1 U7614 ( .A(n5936), .ZN(n5945) );
  INV_X1 U7615 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U7616 ( .A1(n5945), .A2(n9442), .ZN(n5937) );
  NAND2_X1 U7617 ( .A1(n5938), .A2(n5937), .ZN(n9219) );
  OR2_X1 U7618 ( .A1(n6102), .A2(n9219), .ZN(n5941) );
  INV_X1 U7619 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7620 ( .A1(n4449), .A2(n5939), .ZN(n5940) );
  OR2_X1 U7621 ( .A1(n9643), .A2(n8994), .ZN(n6245) );
  NAND2_X1 U7622 ( .A1(n9643), .A2(n8994), .ZN(n9132) );
  NAND2_X1 U7623 ( .A1(n6118), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5950) );
  INV_X1 U7624 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7625 ( .A1(n4442), .A2(n5944), .ZN(n5949) );
  OAI21_X1 U7626 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n5946), .A(n5945), .ZN(
        n9227) );
  OR2_X1 U7627 ( .A1(n6102), .A2(n9227), .ZN(n5948) );
  INV_X1 U7628 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9428) );
  OR2_X1 U7629 ( .A1(n4449), .A2(n9428), .ZN(n5947) );
  NAND2_X1 U7630 ( .A1(n9649), .A2(n8971), .ZN(n6251) );
  OR2_X1 U7631 ( .A1(n5959), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5952) );
  AND2_X1 U7632 ( .A1(n5952), .A2(n5951), .ZN(n9547) );
  NAND2_X1 U7633 ( .A1(n9547), .A2(n6084), .ZN(n5957) );
  INV_X1 U7634 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9360) );
  NAND2_X1 U7635 ( .A1(n6004), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7636 ( .A1(n6108), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5953) );
  OAI211_X1 U7637 ( .C1(n5919), .C2(n9360), .A(n5954), .B(n5953), .ZN(n5955)
         );
  INV_X1 U7638 ( .A(n5955), .ZN(n5956) );
  NAND2_X1 U7639 ( .A1(n9655), .A2(n8899), .ZN(n6243) );
  NOR2_X1 U7640 ( .A1(n5964), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5958) );
  OR2_X1 U7641 ( .A1(n5959), .A2(n5958), .ZN(n8871) );
  INV_X1 U7642 ( .A(n8871), .ZN(n9562) );
  INV_X1 U7643 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U7644 ( .A1(n6108), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5961) );
  INV_X1 U7645 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9430) );
  OR2_X1 U7646 ( .A1(n5919), .A2(n9430), .ZN(n5960) );
  OAI211_X1 U7647 ( .C1(n9493), .C2(n4449), .A(n5961), .B(n5960), .ZN(n5962)
         );
  AOI21_X1 U7648 ( .B1(n9562), .B2(n6084), .A(n5962), .ZN(n8947) );
  OR2_X1 U7649 ( .A1(n9659), .A2(n8947), .ZN(n6179) );
  NAND2_X1 U7650 ( .A1(n9659), .A2(n8947), .ZN(n9125) );
  NOR2_X1 U7651 ( .A1(n5970), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5963) );
  OR2_X1 U7652 ( .A1(n5964), .A2(n5963), .ZN(n9582) );
  INV_X1 U7653 ( .A(n9582), .ZN(n5969) );
  INV_X1 U7654 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5967) );
  NAND2_X1 U7655 ( .A1(n6118), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7656 ( .A1(n6004), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5965) );
  OAI211_X1 U7657 ( .C1(n5967), .C2(n4441), .A(n5966), .B(n5965), .ZN(n5968)
         );
  AOI21_X1 U7658 ( .B1(n5969), .B2(n6084), .A(n5968), .ZN(n8995) );
  NAND2_X1 U7659 ( .A1(n9664), .A2(n8995), .ZN(n6146) );
  INV_X1 U7660 ( .A(n5970), .ZN(n5972) );
  INV_X1 U7661 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8939) );
  INV_X1 U7662 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8890) );
  OAI21_X1 U7663 ( .B1(n5984), .B2(n8939), .A(n8890), .ZN(n5971) );
  NAND2_X1 U7664 ( .A1(n5972), .A2(n5971), .ZN(n9602) );
  OR2_X1 U7665 ( .A1(n9602), .A2(n6102), .ZN(n5978) );
  INV_X1 U7666 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U7667 ( .A1(n6118), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7668 ( .A1(n6004), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5973) );
  OAI211_X1 U7669 ( .C1(n5975), .C2(n4442), .A(n5974), .B(n5973), .ZN(n5976)
         );
  INV_X1 U7670 ( .A(n5976), .ZN(n5977) );
  OR2_X1 U7671 ( .A1(n9669), .A2(n8938), .ZN(n6237) );
  NAND2_X1 U7672 ( .A1(n9669), .A2(n8938), .ZN(n6238) );
  XNOR2_X1 U7673 ( .A(n5984), .B(P1_REG3_REG_20__SCAN_IN), .ZN(n9613) );
  INV_X1 U7674 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7675 ( .A1(n6118), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5980) );
  NAND2_X1 U7676 ( .A1(n6004), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5979) );
  OAI211_X1 U7677 ( .C1(n5981), .C2(n4441), .A(n5980), .B(n5979), .ZN(n5982)
         );
  AOI21_X1 U7678 ( .B1(n9613), .B2(n6084), .A(n5982), .ZN(n8889) );
  OR2_X1 U7679 ( .A1(n9674), .A2(n8889), .ZN(n9591) );
  NAND2_X1 U7680 ( .A1(n9674), .A2(n8889), .ZN(n9593) );
  NAND2_X1 U7681 ( .A1(n9591), .A2(n9593), .ZN(n9616) );
  NAND2_X1 U7682 ( .A1(n5992), .A2(n9298), .ZN(n5983) );
  AND2_X1 U7683 ( .A1(n5984), .A2(n5983), .ZN(n8879) );
  NAND2_X1 U7684 ( .A1(n8879), .A2(n6084), .ZN(n5990) );
  INV_X1 U7685 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7686 ( .A1(n6004), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7687 ( .A1(n6118), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5985) );
  OAI211_X1 U7688 ( .C1(n4442), .C2(n5987), .A(n5986), .B(n5985), .ZN(n5988)
         );
  INV_X1 U7689 ( .A(n5988), .ZN(n5989) );
  AND2_X1 U7690 ( .A1(n5990), .A2(n5989), .ZN(n8937) );
  OR2_X1 U7691 ( .A1(n9146), .A2(n8937), .ZN(n6235) );
  AND2_X1 U7692 ( .A1(n9146), .A2(n8937), .ZN(n6184) );
  NAND2_X1 U7693 ( .A1(n6235), .A2(n6233), .ZN(n8199) );
  NAND2_X1 U7694 ( .A1(n6003), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5991) );
  INV_X1 U7695 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8960) );
  NAND2_X1 U7696 ( .A1(n5991), .A2(n8960), .ZN(n5993) );
  NAND2_X1 U7697 ( .A1(n5993), .A2(n5992), .ZN(n8961) );
  OR2_X1 U7698 ( .A1(n8961), .A2(n6102), .ZN(n5998) );
  INV_X1 U7699 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U7700 ( .A1(n6118), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7701 ( .A1(n6004), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5994) );
  OAI211_X1 U7702 ( .C1(n9101), .C2(n4441), .A(n5995), .B(n5994), .ZN(n5996)
         );
  INV_X1 U7703 ( .A(n5996), .ZN(n5997) );
  AND2_X1 U7704 ( .A1(n5998), .A2(n5997), .ZN(n6495) );
  OR2_X1 U7705 ( .A1(n8197), .A2(n6495), .ZN(n6232) );
  NAND2_X1 U7706 ( .A1(n8197), .A2(n6495), .ZN(n8187) );
  INV_X1 U7707 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7708 ( .A(n6003), .B(n5999), .ZN(n8917) );
  INV_X1 U7709 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9081) );
  NAND2_X1 U7710 ( .A1(n6118), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6001) );
  OR2_X1 U7711 ( .A1(n4449), .A2(n9399), .ZN(n6000) );
  OAI211_X1 U7712 ( .C1(n9081), .C2(n4442), .A(n6001), .B(n6000), .ZN(n6002)
         );
  AOI21_X1 U7713 ( .B1(n8917), .B2(n6084), .A(n6002), .ZN(n8143) );
  OR2_X1 U7714 ( .A1(n8921), .A2(n8143), .ZN(n6231) );
  NAND2_X1 U7715 ( .A1(n8921), .A2(n8143), .ZN(n6226) );
  AOI21_X1 U7716 ( .B1(n9379), .B2(n6008), .A(n6003), .ZN(n8909) );
  INV_X1 U7717 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U7718 ( .A1(n6118), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U7719 ( .A1(n6004), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6005) );
  OAI211_X1 U7720 ( .C1(n9053), .C2(n4441), .A(n6006), .B(n6005), .ZN(n6007)
         );
  AOI21_X1 U7721 ( .B1(n8909), .B2(n6084), .A(n6007), .ZN(n8071) );
  NAND2_X1 U7722 ( .A1(n9763), .A2(n8071), .ZN(n6276) );
  INV_X1 U7723 ( .A(n8989), .ZN(n9769) );
  OAI21_X1 U7724 ( .B1(n6014), .B2(P1_REG3_REG_15__SCAN_IN), .A(n6008), .ZN(
        n8986) );
  INV_X1 U7725 ( .A(n8986), .ZN(n6012) );
  INV_X1 U7726 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U7727 ( .A1(n6118), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7728 ( .A1(n6108), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6009) );
  OAI211_X1 U7729 ( .C1(n4449), .C2(n7912), .A(n6010), .B(n6009), .ZN(n6011)
         );
  AOI21_X1 U7730 ( .B1(n6012), .B2(n6084), .A(n6011), .ZN(n7968) );
  INV_X1 U7731 ( .A(n7968), .ZN(n8999) );
  AND2_X1 U7732 ( .A1(n9769), .A2(n8999), .ZN(n6303) );
  INV_X1 U7733 ( .A(n6303), .ZN(n6221) );
  NAND2_X1 U7734 ( .A1(n8989), .A2(n7968), .ZN(n7964) );
  NAND2_X1 U7735 ( .A1(n6221), .A2(n7964), .ZN(n7972) );
  NAND2_X1 U7736 ( .A1(n6118), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6020) );
  INV_X1 U7737 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7738 ( .A1(n4449), .A2(n6013), .ZN(n6019) );
  NAND2_X1 U7739 ( .A1(n6024), .A2(n8211), .ZN(n6016) );
  INV_X1 U7740 ( .A(n6014), .ZN(n6015) );
  NAND2_X1 U7741 ( .A1(n6016), .A2(n6015), .ZN(n7899) );
  OR2_X1 U7742 ( .A1(n6102), .A2(n7899), .ZN(n6018) );
  INV_X1 U7743 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9050) );
  OR2_X1 U7744 ( .A1(n4442), .A2(n9050), .ZN(n6017) );
  AND4_X1 U7745 ( .A1(n6020), .A2(n6019), .A3(n6018), .A4(n6017), .ZN(n7908)
         );
  OR2_X1 U7746 ( .A1(n6021), .A2(n7908), .ZN(n6302) );
  NAND2_X1 U7747 ( .A1(n6021), .A2(n7908), .ZN(n6217) );
  NAND2_X1 U7748 ( .A1(n6108), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6029) );
  INV_X1 U7749 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7750 ( .A1(n5919), .A2(n6022), .ZN(n6028) );
  OR2_X1 U7751 ( .A1(n6030), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7752 ( .A1(n6024), .A2(n6023), .ZN(n8065) );
  OR2_X1 U7753 ( .A1(n6102), .A2(n8065), .ZN(n6027) );
  INV_X1 U7754 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6025) );
  OR2_X1 U7755 ( .A1(n4449), .A2(n6025), .ZN(n6026) );
  OR2_X1 U7756 ( .A1(n8067), .A2(n7711), .ZN(n6301) );
  NAND2_X1 U7757 ( .A1(n8067), .A2(n7711), .ZN(n7892) );
  NAND2_X1 U7758 ( .A1(n6301), .A2(n7892), .ZN(n7887) );
  NAND2_X1 U7759 ( .A1(n6118), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6034) );
  INV_X1 U7760 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7716) );
  OR2_X1 U7761 ( .A1(n4449), .A2(n7716), .ZN(n6033) );
  OR2_X1 U7762 ( .A1(n4990), .A2(n6030), .ZN(n7988) );
  OR2_X1 U7763 ( .A1(n6102), .A2(n7988), .ZN(n6032) );
  INV_X1 U7764 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7439) );
  OR2_X1 U7765 ( .A1(n4441), .A2(n7439), .ZN(n6031) );
  OR2_X1 U7766 ( .A1(n7990), .A2(n7808), .ZN(n6295) );
  NAND2_X1 U7767 ( .A1(n7990), .A2(n7808), .ZN(n6298) );
  NAND2_X1 U7768 ( .A1(n6118), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6042) );
  INV_X1 U7769 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7438) );
  OR2_X1 U7770 ( .A1(n4442), .A2(n7438), .ZN(n6041) );
  NAND2_X1 U7771 ( .A1(n6069), .A2(n6035), .ZN(n6036) );
  NAND2_X1 U7772 ( .A1(n6037), .A2(n6036), .ZN(n8093) );
  OR2_X1 U7773 ( .A1(n6102), .A2(n8093), .ZN(n6040) );
  INV_X1 U7774 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7775 ( .A1(n4449), .A2(n6038), .ZN(n6039) );
  OR2_X1 U7776 ( .A1(n8095), .A2(n7709), .ZN(n6294) );
  NAND2_X1 U7777 ( .A1(n8095), .A2(n7709), .ZN(n6293) );
  NAND2_X1 U7778 ( .A1(n6294), .A2(n6293), .ZN(n7713) );
  NAND2_X1 U7779 ( .A1(n6118), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6049) );
  INV_X1 U7780 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7087) );
  OR2_X1 U7781 ( .A1(n4441), .A2(n7087), .ZN(n6048) );
  INV_X1 U7782 ( .A(n6067), .ZN(n6045) );
  NAND2_X1 U7783 ( .A1(n6053), .A2(n6043), .ZN(n6044) );
  NAND2_X1 U7784 ( .A1(n6045), .A2(n6044), .ZN(n7782) );
  OR2_X1 U7785 ( .A1(n6102), .A2(n7782), .ZN(n6047) );
  INV_X1 U7786 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7460) );
  OR2_X1 U7787 ( .A1(n4449), .A2(n7460), .ZN(n6046) );
  NAND2_X1 U7788 ( .A1(n6118), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6057) );
  INV_X1 U7789 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7423) );
  OR2_X1 U7790 ( .A1(n4449), .A2(n7423), .ZN(n6056) );
  INV_X1 U7791 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6050) );
  OR2_X1 U7792 ( .A1(n4442), .A2(n6050), .ZN(n6055) );
  NAND2_X1 U7793 ( .A1(n6060), .A2(n6051), .ZN(n6052) );
  NAND2_X1 U7794 ( .A1(n6053), .A2(n6052), .ZN(n9795) );
  OR2_X1 U7795 ( .A1(n6102), .A2(n9795), .ZN(n6054) );
  AND2_X1 U7796 ( .A1(n7466), .A2(n7476), .ZN(n7414) );
  INV_X1 U7797 ( .A(n7414), .ZN(n6189) );
  NAND2_X1 U7798 ( .A1(n6108), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7799 ( .A1(n6118), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U7800 ( .A1(n6076), .A2(n6058), .ZN(n6059) );
  NAND2_X1 U7801 ( .A1(n6060), .A2(n6059), .ZN(n7522) );
  OR2_X1 U7802 ( .A1(n6102), .A2(n7522), .ZN(n6062) );
  OR2_X1 U7803 ( .A1(n4449), .A2(n4661), .ZN(n6061) );
  NAND4_X1 U7804 ( .A1(n6064), .A2(n6063), .A3(n6062), .A4(n6061), .ZN(n9004)
         );
  INV_X1 U7805 ( .A(n9004), .ZN(n7411) );
  NAND2_X1 U7806 ( .A1(n7524), .A2(n7411), .ZN(n6193) );
  NAND2_X1 U7807 ( .A1(n10048), .A2(n7544), .ZN(n7450) );
  NAND2_X1 U7808 ( .A1(n6118), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6073) );
  INV_X1 U7809 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6066) );
  OR2_X1 U7810 ( .A1(n4441), .A2(n6066), .ZN(n6072) );
  OR2_X1 U7811 ( .A1(n6067), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7812 ( .A1(n6069), .A2(n6068), .ZN(n7959) );
  OR2_X1 U7813 ( .A1(n6102), .A2(n7959), .ZN(n6071) );
  INV_X1 U7814 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7537) );
  OR2_X1 U7815 ( .A1(n4449), .A2(n7537), .ZN(n6070) );
  OR2_X1 U7816 ( .A1(n7961), .A2(n7565), .ZN(n6210) );
  NAND2_X1 U7817 ( .A1(n7961), .A2(n7565), .ZN(n6292) );
  AND2_X1 U7818 ( .A1(n10031), .A2(n9004), .ZN(n6194) );
  NAND2_X1 U7819 ( .A1(n6108), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6080) );
  INV_X1 U7820 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6074) );
  OR2_X1 U7821 ( .A1(n5919), .A2(n6074), .ZN(n6079) );
  OR2_X1 U7822 ( .A1(n6116), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U7823 ( .A1(n6076), .A2(n6075), .ZN(n7349) );
  OR2_X1 U7824 ( .A1(n6102), .A2(n7349), .ZN(n6078) );
  INV_X1 U7825 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7350) );
  OR2_X1 U7826 ( .A1(n4449), .A2(n7350), .ZN(n6077) );
  OR2_X1 U7827 ( .A1(n7407), .A2(n7475), .ZN(n6192) );
  INV_X1 U7828 ( .A(n6192), .ZN(n6081) );
  NOR2_X1 U7829 ( .A1(n6194), .A2(n6081), .ZN(n6082) );
  NAND2_X1 U7830 ( .A1(n6099), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6088) );
  INV_X1 U7831 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6986) );
  OR2_X1 U7832 ( .A1(n4442), .A2(n6986), .ZN(n6087) );
  INV_X1 U7833 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6083) );
  NOR2_X1 U7834 ( .A1(n7272), .A2(n9976), .ZN(n6153) );
  INV_X1 U7835 ( .A(n6153), .ZN(n9962) );
  NAND2_X1 U7836 ( .A1(n7272), .A2(n9976), .ZN(n6278) );
  NAND2_X1 U7837 ( .A1(n9962), .A2(n6278), .ZN(n7315) );
  NOR2_X1 U7838 ( .A1(n7315), .A2(n6374), .ZN(n6107) );
  NAND2_X1 U7839 ( .A1(n6118), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6092) );
  OR2_X1 U7840 ( .A1(n4442), .A2(n10095), .ZN(n6091) );
  INV_X1 U7841 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7097) );
  OR2_X1 U7842 ( .A1(n4449), .A2(n7097), .ZN(n6090) );
  OR2_X1 U7843 ( .A1(n6102), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6089) );
  NAND4_X2 U7844 ( .A1(n6092), .A2(n6091), .A3(n6090), .A4(n6089), .ZN(n9006)
         );
  NOR2_X1 U7845 ( .A1(n9006), .A2(n10007), .ZN(n6157) );
  INV_X1 U7846 ( .A(n6157), .ZN(n6093) );
  NAND2_X1 U7847 ( .A1(n9006), .A2(n10007), .ZN(n6280) );
  NAND2_X1 U7848 ( .A1(n6093), .A2(n6280), .ZN(n9954) );
  INV_X1 U7849 ( .A(n9954), .ZN(n9944) );
  INV_X1 U7850 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6094) );
  INV_X1 U7851 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9441) );
  OR2_X1 U7852 ( .A1(n4448), .A2(n9441), .ZN(n6097) );
  NAND2_X1 U7853 ( .A1(n6099), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7854 ( .A1(n6084), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7855 ( .A1(n6099), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6106) );
  INV_X1 U7856 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7095) );
  OR2_X1 U7857 ( .A1(n4449), .A2(n7095), .ZN(n6105) );
  INV_X1 U7858 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6100) );
  OR2_X1 U7859 ( .A1(n4441), .A2(n6100), .ZN(n6104) );
  INV_X1 U7860 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9494) );
  NAND4_X2 U7861 ( .A1(n6106), .A2(n6105), .A3(n6104), .A4(n6103), .ZN(n9007)
         );
  AND4_X1 U7862 ( .A1(n6107), .A2(n9944), .A3(n7274), .A4(n7323), .ZN(n6124)
         );
  NAND2_X1 U7863 ( .A1(n6108), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6113) );
  INV_X1 U7864 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7865 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n6115), .ZN(n7336) );
  OR2_X1 U7866 ( .A1(n6102), .A2(n7336), .ZN(n6111) );
  INV_X1 U7867 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7333) );
  OR2_X1 U7868 ( .A1(n4449), .A2(n7333), .ZN(n6110) );
  OR2_X1 U7869 ( .A1(n7357), .A2(n9005), .ZN(n9926) );
  NAND2_X1 U7870 ( .A1(n7357), .A2(n9005), .ZN(n9925) );
  AND2_X1 U7871 ( .A1(n9926), .A2(n9925), .ZN(n7330) );
  NAND2_X1 U7872 ( .A1(n7407), .A2(n7475), .ZN(n6191) );
  INV_X1 U7873 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6114) );
  OR2_X1 U7874 ( .A1(n4449), .A2(n6114), .ZN(n6120) );
  AND2_X1 U7875 ( .A1(n6115), .A2(n7248), .ZN(n6117) );
  OR2_X1 U7876 ( .A1(n6117), .A2(n6116), .ZN(n9933) );
  INV_X1 U7877 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6121) );
  OR2_X1 U7878 ( .A1(n4442), .A2(n6121), .ZN(n6122) );
  XNOR2_X1 U7879 ( .A(n7361), .B(n7362), .ZN(n9929) );
  NAND4_X1 U7880 ( .A1(n6124), .A2(n7330), .A3(n6191), .A4(n9929), .ZN(n6125)
         );
  NOR2_X1 U7881 ( .A1(n6285), .A2(n6125), .ZN(n6126) );
  NAND3_X1 U7882 ( .A1(n6290), .A2(n7547), .A3(n6126), .ZN(n6127) );
  NOR2_X1 U7883 ( .A1(n7713), .A2(n6127), .ZN(n6128) );
  NAND4_X1 U7884 ( .A1(n7891), .A2(n6163), .A3(n7707), .A4(n6128), .ZN(n6129)
         );
  NOR2_X1 U7885 ( .A1(n7972), .A2(n6129), .ZN(n6130) );
  NAND4_X1 U7886 ( .A1(n6166), .A2(n8075), .A3(n4996), .A4(n6130), .ZN(n6131)
         );
  NOR3_X1 U7887 ( .A1(n9616), .A2(n8199), .A3(n6131), .ZN(n6132) );
  NAND4_X1 U7888 ( .A1(n9567), .A2(n9122), .A3(n9594), .A4(n6132), .ZN(n6133)
         );
  NOR2_X1 U7889 ( .A1(n4622), .A2(n6133), .ZN(n6134) );
  NAND4_X1 U7890 ( .A1(n9134), .A2(n9216), .A3(n9129), .A4(n6134), .ZN(n6135)
         );
  NOR2_X1 U7891 ( .A1(n9188), .A2(n6135), .ZN(n6136) );
  NAND2_X1 U7892 ( .A1(n6269), .A2(n9139), .ZN(n6140) );
  AND4_X1 U7893 ( .A1(n4638), .A2(n6324), .A3(n6136), .A4(n6140), .ZN(n6137)
         );
  AND3_X1 U7894 ( .A1(n6334), .A2(n6137), .A3(n4984), .ZN(n6271) );
  INV_X1 U7895 ( .A(n6271), .ZN(n6178) );
  INV_X1 U7896 ( .A(n6139), .ZN(n6993) );
  NOR2_X1 U7897 ( .A1(n6269), .A2(n6993), .ZN(n6173) );
  AND2_X1 U7898 ( .A1(n6140), .A2(n6263), .ZN(n6323) );
  NAND2_X1 U7899 ( .A1(n6262), .A2(n6257), .ZN(n6322) );
  NAND2_X1 U7900 ( .A1(n9136), .A2(n9135), .ZN(n6258) );
  AND2_X1 U7901 ( .A1(n6250), .A2(n6245), .ZN(n6254) );
  INV_X1 U7902 ( .A(n6254), .ZN(n6317) );
  NAND2_X1 U7903 ( .A1(n6179), .A2(n9565), .ZN(n6141) );
  NAND2_X1 U7904 ( .A1(n6141), .A2(n9125), .ZN(n6182) );
  INV_X1 U7905 ( .A(n6182), .ZN(n6142) );
  NAND2_X1 U7906 ( .A1(n6142), .A2(n6243), .ZN(n6143) );
  AND3_X1 U7907 ( .A1(n9130), .A2(n9127), .A3(n6143), .ZN(n6151) );
  INV_X1 U7908 ( .A(n9593), .ZN(n6144) );
  NAND2_X1 U7909 ( .A1(n6237), .A2(n6144), .ZN(n6145) );
  AND2_X1 U7910 ( .A1(n6145), .A2(n6238), .ZN(n9123) );
  NAND2_X1 U7911 ( .A1(n9125), .A2(n6146), .ZN(n6180) );
  INV_X1 U7912 ( .A(n6180), .ZN(n6147) );
  NAND3_X1 U7913 ( .A1(n6243), .A2(n9123), .A3(n6147), .ZN(n6148) );
  INV_X1 U7914 ( .A(n6251), .ZN(n6246) );
  AOI21_X1 U7915 ( .B1(n6151), .B2(n6148), .A(n6246), .ZN(n6149) );
  NOR2_X1 U7916 ( .A1(n6317), .A2(n6149), .ZN(n6150) );
  OR2_X1 U7917 ( .A1(n6258), .A2(n6150), .ZN(n6320) );
  INV_X1 U7918 ( .A(n6151), .ZN(n6152) );
  NAND2_X1 U7919 ( .A1(n6237), .A2(n9591), .ZN(n9124) );
  OR2_X1 U7920 ( .A1(n6152), .A2(n9124), .ZN(n6314) );
  INV_X1 U7921 ( .A(n6302), .ZN(n7905) );
  NOR2_X1 U7922 ( .A1(n7972), .A2(n7905), .ZN(n6165) );
  NAND2_X1 U7923 ( .A1(n7274), .A2(n6153), .ZN(n6155) );
  OR2_X1 U7924 ( .A1(n4440), .A2(n9992), .ZN(n6154) );
  NAND2_X1 U7925 ( .A1(n6155), .A2(n6154), .ZN(n7276) );
  INV_X1 U7926 ( .A(n4447), .ZN(n7287) );
  OR2_X1 U7927 ( .A1(n9007), .A2(n7287), .ZN(n6156) );
  NAND2_X1 U7928 ( .A1(n9928), .A2(n9926), .ZN(n6158) );
  NAND2_X1 U7929 ( .A1(n7361), .A2(n7118), .ZN(n6159) );
  INV_X1 U7930 ( .A(n6191), .ZN(n6160) );
  OR2_X1 U7931 ( .A1(n6284), .A2(n6285), .ZN(n6161) );
  INV_X1 U7932 ( .A(n7713), .ZN(n6162) );
  NAND2_X1 U7933 ( .A1(n7561), .A2(n6294), .ZN(n7708) );
  INV_X1 U7934 ( .A(n7891), .ZN(n7916) );
  INV_X1 U7935 ( .A(n7892), .ZN(n6164) );
  NOR2_X1 U7936 ( .A1(n7916), .A2(n6164), .ZN(n6219) );
  NAND3_X1 U7937 ( .A1(n7965), .A2(n4996), .A3(n7964), .ZN(n7966) );
  NAND2_X1 U7938 ( .A1(n8188), .A2(n8187), .ZN(n6168) );
  INV_X1 U7939 ( .A(n8199), .ZN(n6167) );
  OAI21_X1 U7940 ( .B1(n6314), .B2(n9617), .A(n9132), .ZN(n6169) );
  AND2_X1 U7941 ( .A1(n6254), .A2(n6169), .ZN(n6170) );
  NOR2_X1 U7942 ( .A1(n6320), .A2(n6170), .ZN(n6171) );
  OR2_X1 U7943 ( .A1(n6322), .A2(n6171), .ZN(n6172) );
  OAI211_X1 U7944 ( .C1(n6138), .C2(n6173), .A(n6323), .B(n6172), .ZN(n6176)
         );
  INV_X1 U7945 ( .A(n6324), .ZN(n6174) );
  NAND2_X1 U7946 ( .A1(n6174), .A2(n6138), .ZN(n6175) );
  NAND4_X1 U7947 ( .A1(n6176), .A2(n6981), .A3(n4984), .A4(n6175), .ZN(n6177)
         );
  NAND2_X1 U7948 ( .A1(n6178), .A2(n6177), .ZN(n6274) );
  NAND2_X1 U7949 ( .A1(n6180), .A2(n6179), .ZN(n6181) );
  NAND2_X1 U7950 ( .A1(n7937), .A2(n6376), .ZN(n7023) );
  MUX2_X1 U7951 ( .A(n6182), .B(n6181), .S(n7023), .Z(n6242) );
  NAND2_X1 U7952 ( .A1(n6238), .A2(n9593), .ZN(n6183) );
  MUX2_X1 U7953 ( .A(n6183), .B(n9124), .S(n7023), .Z(n6240) );
  AND2_X1 U7954 ( .A1(n6235), .A2(n6232), .ZN(n6275) );
  NAND2_X1 U7955 ( .A1(n8187), .A2(n6226), .ZN(n6185) );
  AOI21_X1 U7956 ( .B1(n6275), .B2(n6185), .A(n6184), .ZN(n6313) );
  NAND2_X1 U7957 ( .A1(n7344), .A2(n6192), .ZN(n6186) );
  INV_X1 U7958 ( .A(n6194), .ZN(n6187) );
  AND2_X1 U7959 ( .A1(n6187), .A2(n6193), .ZN(n7410) );
  NAND3_X1 U7960 ( .A1(n6186), .A2(n7410), .A3(n6191), .ZN(n6188) );
  NAND3_X1 U7961 ( .A1(n6188), .A2(n7449), .A3(n6187), .ZN(n6190) );
  NAND3_X1 U7962 ( .A1(n6190), .A2(n7450), .A3(n6189), .ZN(n6196) );
  NAND2_X1 U7963 ( .A1(n6192), .A2(n6191), .ZN(n7404) );
  INV_X1 U7964 ( .A(n6210), .ZN(n6289) );
  AOI21_X1 U7965 ( .B1(n6208), .B2(n7450), .A(n6289), .ZN(n6216) );
  NAND4_X1 U7966 ( .A1(n6298), .A2(n6292), .A3(n6293), .A4(n7023), .ZN(n6215)
         );
  INV_X1 U7967 ( .A(n7709), .ZN(n7715) );
  NOR2_X1 U7968 ( .A1(n7715), .A2(n7023), .ZN(n6200) );
  INV_X1 U7969 ( .A(n7808), .ZN(n9002) );
  NOR2_X1 U7970 ( .A1(n9002), .A2(n7023), .ZN(n6197) );
  AOI21_X1 U7971 ( .B1(n8095), .B2(n6200), .A(n6197), .ZN(n6206) );
  NAND2_X1 U7972 ( .A1(n7715), .A2(n7023), .ZN(n6199) );
  INV_X1 U7973 ( .A(n7023), .ZN(n6266) );
  OAI22_X1 U7974 ( .A1(n8095), .A2(n6199), .B1(n7808), .B2(n6266), .ZN(n6198)
         );
  NAND2_X1 U7975 ( .A1(n10070), .A2(n6198), .ZN(n6205) );
  NOR2_X1 U7976 ( .A1(n6199), .A2(n7808), .ZN(n6203) );
  NAND2_X1 U7977 ( .A1(n6200), .A2(n7808), .ZN(n6201) );
  NAND2_X1 U7978 ( .A1(n8095), .A2(n6201), .ZN(n6202) );
  OAI21_X1 U7979 ( .B1(n8095), .B2(n6203), .A(n6202), .ZN(n6204) );
  OAI211_X1 U7980 ( .C1(n10070), .C2(n6206), .A(n6205), .B(n6204), .ZN(n6207)
         );
  NOR2_X1 U7981 ( .A1(n7887), .A2(n6207), .ZN(n6214) );
  NAND2_X1 U7982 ( .A1(n6209), .A2(n6292), .ZN(n6212) );
  AND4_X1 U7983 ( .A1(n6295), .A2(n6266), .A3(n6294), .A4(n6210), .ZN(n6211)
         );
  NAND2_X1 U7984 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  OAI211_X1 U7985 ( .C1(n6216), .C2(n6215), .A(n6214), .B(n6213), .ZN(n6220)
         );
  NAND3_X1 U7986 ( .A1(n6220), .A2(n7891), .A3(n6301), .ZN(n6218) );
  AND2_X1 U7987 ( .A1(n7964), .A2(n6217), .ZN(n6305) );
  AOI21_X1 U7988 ( .B1(n6218), .B2(n6305), .A(n6303), .ZN(n6224) );
  NAND2_X1 U7989 ( .A1(n6220), .A2(n6219), .ZN(n6222) );
  NAND3_X1 U7990 ( .A1(n6222), .A2(n6221), .A3(n6302), .ZN(n6223) );
  NOR2_X1 U7991 ( .A1(n7964), .A2(n6266), .ZN(n6225) );
  NOR2_X1 U7992 ( .A1(n7975), .A2(n6225), .ZN(n6228) );
  AOI21_X1 U7993 ( .B1(n6226), .B2(n6276), .A(n7023), .ZN(n6227) );
  NAND4_X1 U7994 ( .A1(n6234), .A2(n6275), .A3(n6307), .A4(n6231), .ZN(n6230)
         );
  NAND2_X1 U7995 ( .A1(n6232), .A2(n6231), .ZN(n6306) );
  OAI211_X1 U7996 ( .C1(n6234), .C2(n6306), .A(n6233), .B(n8187), .ZN(n6236)
         );
  MUX2_X1 U7997 ( .A(n6238), .B(n6237), .S(n6266), .Z(n6239) );
  MUX2_X1 U7998 ( .A(n9127), .B(n6243), .S(n7023), .Z(n6244) );
  NAND3_X1 U7999 ( .A1(n6247), .A2(n9132), .A3(n9135), .ZN(n6248) );
  NAND3_X1 U8000 ( .A1(n6257), .A2(n6250), .A3(n6248), .ZN(n6249) );
  NAND2_X1 U8001 ( .A1(n6249), .A2(n9136), .ZN(n6261) );
  INV_X1 U8002 ( .A(n6250), .ZN(n6256) );
  NAND2_X1 U8003 ( .A1(n6252), .A2(n6251), .ZN(n6253) );
  NAND3_X1 U8004 ( .A1(n6254), .A2(n9130), .A3(n6253), .ZN(n6255) );
  OAI21_X1 U8005 ( .B1(n6256), .B2(n9132), .A(n6255), .ZN(n6259) );
  OAI21_X1 U8006 ( .B1(n6259), .B2(n6258), .A(n6257), .ZN(n6260) );
  MUX2_X1 U8007 ( .A(n6261), .B(n6260), .S(n6266), .Z(n6265) );
  NAND2_X1 U8008 ( .A1(n6993), .A2(n8992), .ZN(n6267) );
  AND2_X1 U8009 ( .A1(n6334), .A2(n6267), .ZN(n6268) );
  AND2_X1 U8010 ( .A1(n6138), .A2(n8992), .ZN(n6270) );
  NAND2_X1 U8011 ( .A1(n6337), .A2(n6375), .ZN(n6272) );
  INV_X1 U8012 ( .A(n6275), .ZN(n6312) );
  INV_X1 U8013 ( .A(n6276), .ZN(n6310) );
  INV_X1 U8014 ( .A(n6277), .ZN(n6283) );
  AOI21_X1 U8015 ( .B1(n4440), .B2(n9992), .A(n7826), .ZN(n6281) );
  NAND2_X1 U8016 ( .A1(n9007), .A2(n7287), .ZN(n6279) );
  NAND4_X1 U8017 ( .A1(n6281), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n6282)
         );
  NOR2_X1 U8018 ( .A1(n6283), .A2(n6282), .ZN(n6288) );
  INV_X1 U8019 ( .A(n6284), .ZN(n6287) );
  INV_X1 U8020 ( .A(n6285), .ZN(n6286) );
  OAI21_X1 U8021 ( .B1(n6288), .B2(n6287), .A(n6286), .ZN(n6291) );
  AOI21_X1 U8022 ( .B1(n6291), .B2(n6290), .A(n6289), .ZN(n6297) );
  NAND2_X1 U8023 ( .A1(n6293), .A2(n6292), .ZN(n6296) );
  OAI211_X1 U8024 ( .C1(n6297), .C2(n6296), .A(n6295), .B(n6294), .ZN(n6299)
         );
  NAND3_X1 U8025 ( .A1(n6299), .A2(n7892), .A3(n6298), .ZN(n6300) );
  NAND3_X1 U8026 ( .A1(n6302), .A2(n6301), .A3(n6300), .ZN(n6304) );
  AOI21_X1 U8027 ( .B1(n6305), .B2(n6304), .A(n6303), .ZN(n6309) );
  INV_X1 U8028 ( .A(n6306), .ZN(n6308) );
  OAI211_X1 U8029 ( .C1(n6310), .C2(n6309), .A(n6308), .B(n6307), .ZN(n6311)
         );
  NOR2_X1 U8030 ( .A1(n6312), .A2(n6311), .ZN(n6316) );
  INV_X1 U8031 ( .A(n6314), .ZN(n6315) );
  OAI21_X1 U8032 ( .B1(n6316), .B2(n4649), .A(n6315), .ZN(n6318) );
  AOI21_X1 U8033 ( .B1(n6318), .B2(n9132), .A(n6317), .ZN(n6319) );
  NOR2_X1 U8034 ( .A1(n6320), .A2(n6319), .ZN(n6321) );
  NOR2_X1 U8035 ( .A1(n6322), .A2(n6321), .ZN(n6326) );
  INV_X1 U8036 ( .A(n6323), .ZN(n6325) );
  OAI211_X1 U8037 ( .C1(n6326), .C2(n6325), .A(n6324), .B(n4984), .ZN(n6327)
         );
  NAND2_X1 U8038 ( .A1(n6327), .A2(n6334), .ZN(n6328) );
  XNOR2_X1 U8039 ( .A(n6328), .B(n5880), .ZN(n6330) );
  AND2_X1 U8040 ( .A1(n6329), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6600) );
  OR2_X1 U8041 ( .A1(n4984), .A2(n7023), .ZN(n6336) );
  AND2_X1 U8042 ( .A1(n6600), .A2(n7937), .ZN(n6338) );
  AND2_X1 U8043 ( .A1(n7022), .A2(n6374), .ZN(n7014) );
  OAI211_X1 U8044 ( .C1(n6334), .C2(n5880), .A(n6338), .B(n7014), .ZN(n6335)
         );
  AOI21_X1 U8045 ( .B1(n6337), .B2(n6336), .A(n6335), .ZN(n6343) );
  INV_X1 U8046 ( .A(n6981), .ZN(n6588) );
  NOR2_X1 U8047 ( .A1(n6588), .A2(n7017), .ZN(n7020) );
  INV_X1 U8048 ( .A(n8238), .ZN(n9009) );
  INV_X1 U8049 ( .A(n4451), .ZN(n7074) );
  AND2_X1 U8050 ( .A1(n9009), .A2(n7074), .ZN(n9012) );
  NAND2_X1 U8051 ( .A1(n7020), .A2(n9012), .ZN(n6340) );
  INV_X1 U8052 ( .A(n6338), .ZN(n6339) );
  OAI211_X1 U8053 ( .C1(n6340), .C2(n6980), .A(P1_B_REG_SCAN_IN), .B(n6339), 
        .ZN(n6341) );
  INV_X1 U8054 ( .A(n6341), .ZN(n6342) );
  NAND2_X1 U8055 ( .A1(n6345), .A2(n6344), .ZN(P1_U3242) );
  INV_X1 U8056 ( .A(n8563), .ZN(n6812) );
  NAND2_X1 U8057 ( .A1(n8563), .A2(n8422), .ZN(n6346) );
  NAND2_X1 U8058 ( .A1(n6347), .A2(n6346), .ZN(n6350) );
  NAND2_X1 U8059 ( .A1(n6812), .A2(n6348), .ZN(n6349) );
  NAND2_X1 U8060 ( .A1(n6350), .A2(n6349), .ZN(n6355) );
  NAND2_X1 U8061 ( .A1(n6351), .A2(n6627), .ZN(n6353) );
  OR2_X1 U8062 ( .A1(n5107), .A2(n8241), .ZN(n6352) );
  INV_X1 U8063 ( .A(n6354), .ZN(n8421) );
  XNOR2_X1 U8064 ( .A(n6355), .B(n6653), .ZN(n6364) );
  XNOR2_X1 U8065 ( .A(n4474), .B(n6653), .ZN(n8550) );
  AND2_X1 U8066 ( .A1(n8422), .A2(n6788), .ZN(n6811) );
  INV_X1 U8067 ( .A(n6811), .ZN(n8570) );
  INV_X1 U8068 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9335) );
  OR2_X1 U8069 ( .A1(n6356), .A2(n9335), .ZN(n6360) );
  INV_X1 U8070 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8549) );
  OR2_X1 U8071 ( .A1(n6621), .A2(n8549), .ZN(n6359) );
  INV_X1 U8072 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6357) );
  OR2_X1 U8073 ( .A1(n5072), .A2(n6357), .ZN(n6358) );
  AND4_X1 U8074 ( .A1(n6625), .A2(n6360), .A3(n6359), .A4(n6358), .ZN(n7514)
         );
  NAND2_X1 U8075 ( .A1(n6962), .A2(P2_B_REG_SCAN_IN), .ZN(n6361) );
  NAND2_X1 U8076 ( .A1(n8694), .A2(n6361), .ZN(n8542) );
  OAI22_X1 U8077 ( .A1(n8570), .A2(n6949), .B1(n7514), .B2(n8542), .ZN(n6362)
         );
  NAND2_X1 U8078 ( .A1(n10325), .A2(n10308), .ZN(n8777) );
  NAND2_X1 U8079 ( .A1(n10323), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6366) );
  OAI21_X1 U8080 ( .B1(n6373), .B2(n10323), .A(n6368), .ZN(P2_U3488) );
  OR2_X1 U8081 ( .A1(n10311), .A2(n10291), .ZN(n8839) );
  OAI21_X1 U8082 ( .B1(n6373), .B2(n10311), .A(n6372), .ZN(P2_U3456) );
  NAND2_X1 U8083 ( .A1(n4440), .A2(n6564), .ZN(n6382) );
  NAND2_X1 U8084 ( .A1(n6377), .A2(n6376), .ZN(n9972) );
  INV_X1 U8085 ( .A(n6377), .ZN(n6378) );
  NAND2_X1 U8086 ( .A1(n6382), .A2(n6381), .ZN(n6384) );
  AOI22_X1 U8087 ( .A1(n4440), .A2(n6507), .B1(n6564), .B2(n7273), .ZN(n6393)
         );
  INV_X1 U8088 ( .A(n9976), .ZN(n7271) );
  NAND2_X1 U8089 ( .A1(n6391), .A2(n6388), .ZN(n7050) );
  NAND2_X1 U8090 ( .A1(n7062), .A2(n7064), .ZN(n7063) );
  INV_X1 U8091 ( .A(n6392), .ZN(n6394) );
  NAND2_X1 U8092 ( .A1(n7063), .A2(n6395), .ZN(n7043) );
  NAND2_X1 U8093 ( .A1(n9007), .A2(n6564), .ZN(n6397) );
  NAND2_X1 U8094 ( .A1(n6397), .A2(n6396), .ZN(n6398) );
  AOI22_X1 U8095 ( .A1(n9007), .A2(n6507), .B1(n6564), .B2(n4447), .ZN(n6399)
         );
  XNOR2_X1 U8096 ( .A(n6401), .B(n6399), .ZN(n7044) );
  INV_X1 U8097 ( .A(n6399), .ZN(n6400) );
  AOI21_X2 U8098 ( .B1(n7043), .B2(n7044), .A(n6402), .ZN(n7057) );
  NAND2_X1 U8099 ( .A1(n9006), .A2(n6579), .ZN(n6405) );
  INV_X1 U8100 ( .A(n9006), .ZN(n7327) );
  OAI22_X1 U8101 ( .A1(n7327), .A2(n6581), .B1(n10007), .B2(n6425), .ZN(n6407)
         );
  XNOR2_X1 U8102 ( .A(n6408), .B(n6407), .ZN(n7056) );
  OAI21_X1 U8103 ( .B1(n7057), .B2(n7056), .A(n6409), .ZN(n7115) );
  XNOR2_X1 U8104 ( .A(n6410), .B(n6552), .ZN(n6411) );
  INV_X1 U8105 ( .A(n9005), .ZN(n7358) );
  OAI22_X1 U8106 ( .A1(n7358), .A2(n6581), .B1(n7357), .B2(n6425), .ZN(n6412)
         );
  XOR2_X1 U8107 ( .A(n6411), .B(n6412), .Z(n7117) );
  NOR2_X1 U8108 ( .A1(n7115), .A2(n7117), .ZN(n7116) );
  INV_X1 U8109 ( .A(n6411), .ZN(n6413) );
  NOR2_X1 U8110 ( .A1(n7116), .A2(n4985), .ZN(n6416) );
  XNOR2_X1 U8111 ( .A(n6414), .B(n6383), .ZN(n6415) );
  NAND2_X1 U8112 ( .A1(n6416), .A2(n6415), .ZN(n7242) );
  OAI22_X1 U8113 ( .A1(n4557), .A2(n6425), .B1(n7118), .B2(n6581), .ZN(n7244)
         );
  NOR2_X1 U8114 ( .A1(n6416), .A2(n6415), .ZN(n7241) );
  INV_X1 U8115 ( .A(n7407), .ZN(n10028) );
  OAI22_X1 U8116 ( .A1(n10028), .A2(n6425), .B1(n7475), .B2(n6581), .ZN(n6418)
         );
  OAI22_X1 U8117 ( .A1(n10028), .A2(n6514), .B1(n7475), .B2(n6425), .ZN(n6417)
         );
  XNOR2_X1 U8118 ( .A(n6417), .B(n6383), .ZN(n6419) );
  XOR2_X1 U8119 ( .A(n6418), .B(n6419), .Z(n7306) );
  OR2_X1 U8120 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  XNOR2_X1 U8121 ( .A(n6421), .B(n6552), .ZN(n7473) );
  AOI22_X1 U8122 ( .A1(n7524), .A2(n6564), .B1(n6507), .B2(n9004), .ZN(n6423)
         );
  INV_X1 U8123 ( .A(n7473), .ZN(n6424) );
  INV_X1 U8124 ( .A(n6423), .ZN(n7472) );
  INV_X1 U8125 ( .A(n7466), .ZN(n10040) );
  OAI22_X1 U8126 ( .A1(n10040), .A2(n6514), .B1(n7476), .B2(n6425), .ZN(n6426)
         );
  XOR2_X1 U8127 ( .A(n6383), .B(n6426), .Z(n6428) );
  NAND2_X1 U8128 ( .A1(n6427), .A2(n6428), .ZN(n6432) );
  INV_X1 U8129 ( .A(n6428), .ZN(n6429) );
  NAND2_X1 U8130 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  NAND2_X1 U8131 ( .A1(n6432), .A2(n6431), .ZN(n9783) );
  OAI22_X1 U8132 ( .A1(n10040), .A2(n6425), .B1(n7476), .B2(n6581), .ZN(n9784)
         );
  INV_X1 U8133 ( .A(n6432), .ZN(n6433) );
  OR2_X1 U8134 ( .A1(n7544), .A2(n6425), .ZN(n6434) );
  NAND2_X1 U8135 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  XNOR2_X1 U8136 ( .A(n6436), .B(n6577), .ZN(n6439) );
  NOR2_X1 U8137 ( .A1(n7544), .A2(n6581), .ZN(n6437) );
  AOI21_X1 U8138 ( .B1(n10048), .B2(n6579), .A(n6437), .ZN(n6438) );
  NOR2_X1 U8139 ( .A1(n6439), .A2(n6438), .ZN(n7776) );
  NAND2_X1 U8140 ( .A1(n6439), .A2(n6438), .ZN(n7775) );
  OR2_X1 U8141 ( .A1(n7709), .A2(n6425), .ZN(n6440) );
  NAND2_X1 U8142 ( .A1(n6441), .A2(n6440), .ZN(n6442) );
  XNOR2_X1 U8143 ( .A(n6442), .B(n6552), .ZN(n8087) );
  OAI22_X1 U8144 ( .A1(n10064), .A2(n6425), .B1(n7709), .B2(n6581), .ZN(n6449)
         );
  OR2_X1 U8145 ( .A1(n7565), .A2(n6425), .ZN(n6443) );
  NAND2_X1 U8146 ( .A1(n6444), .A2(n6443), .ZN(n6445) );
  XNOR2_X1 U8147 ( .A(n6445), .B(n6577), .ZN(n8086) );
  NOR2_X1 U8148 ( .A1(n7565), .A2(n6581), .ZN(n6446) );
  AOI21_X1 U8149 ( .B1(n7961), .B2(n6564), .A(n6446), .ZN(n7954) );
  NOR2_X1 U8150 ( .A1(n4992), .A2(n6447), .ZN(n6448) );
  INV_X1 U8151 ( .A(n6449), .ZN(n8088) );
  AOI21_X1 U8152 ( .B1(n8086), .B2(n7954), .A(n8088), .ZN(n6450) );
  NAND3_X1 U8153 ( .A1(n8088), .A2(n8086), .A3(n7954), .ZN(n6451) );
  OAI22_X1 U8154 ( .A1(n10070), .A2(n6425), .B1(n7808), .B2(n6581), .ZN(n6458)
         );
  NAND2_X1 U8155 ( .A1(n9002), .A2(n6579), .ZN(n6454) );
  NAND2_X1 U8156 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  XNOR2_X1 U8157 ( .A(n6456), .B(n6383), .ZN(n6457) );
  XOR2_X1 U8158 ( .A(n6458), .B(n6457), .Z(n7984) );
  INV_X1 U8159 ( .A(n6457), .ZN(n6460) );
  INV_X1 U8160 ( .A(n6458), .ZN(n6459) );
  INV_X1 U8161 ( .A(n7711), .ZN(n9001) );
  NAND2_X1 U8162 ( .A1(n9001), .A2(n6579), .ZN(n6461) );
  NAND2_X1 U8163 ( .A1(n6462), .A2(n6461), .ZN(n6463) );
  XNOR2_X1 U8164 ( .A(n6463), .B(n6552), .ZN(n6465) );
  INV_X1 U8165 ( .A(n8067), .ZN(n10077) );
  OAI22_X1 U8166 ( .A1(n10077), .A2(n6425), .B1(n7711), .B2(n6581), .ZN(n6464)
         );
  XNOR2_X1 U8167 ( .A(n6465), .B(n6464), .ZN(n8062) );
  OAI21_X1 U8168 ( .B1(n8061), .B2(n8062), .A(n6466), .ZN(n6470) );
  OR2_X1 U8169 ( .A1(n7908), .A2(n6425), .ZN(n6467) );
  NAND2_X1 U8170 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  XNOR2_X1 U8171 ( .A(n6469), .B(n6552), .ZN(n6471) );
  XNOR2_X1 U8172 ( .A(n6470), .B(n6471), .ZN(n8208) );
  INV_X1 U8173 ( .A(n7908), .ZN(n9000) );
  AOI22_X1 U8174 ( .A1(n6021), .A2(n6579), .B1(n6507), .B2(n9000), .ZN(n8209)
         );
  NAND2_X1 U8175 ( .A1(n8208), .A2(n8209), .ZN(n8207) );
  NAND2_X1 U8176 ( .A1(n8207), .A2(n6473), .ZN(n8903) );
  INV_X1 U8177 ( .A(n9763), .ZN(n7978) );
  OAI22_X1 U8178 ( .A1(n7978), .A2(n6514), .B1(n8071), .B2(n6425), .ZN(n6474)
         );
  XNOR2_X1 U8179 ( .A(n6474), .B(n6552), .ZN(n8906) );
  NAND2_X1 U8180 ( .A1(n9763), .A2(n6579), .ZN(n6476) );
  OR2_X1 U8181 ( .A1(n8071), .A2(n6581), .ZN(n6475) );
  NAND2_X1 U8182 ( .A1(n6476), .A2(n6475), .ZN(n6482) );
  NAND2_X1 U8183 ( .A1(n8989), .A2(n6579), .ZN(n6478) );
  OR2_X1 U8184 ( .A1(n7968), .A2(n6581), .ZN(n6477) );
  NAND2_X1 U8185 ( .A1(n6478), .A2(n6477), .ZN(n8981) );
  OR2_X1 U8186 ( .A1(n7968), .A2(n6425), .ZN(n6479) );
  NAND2_X1 U8187 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  XNOR2_X1 U8188 ( .A(n6481), .B(n6383), .ZN(n6485) );
  AOI22_X1 U8189 ( .A1(n8906), .A2(n6482), .B1(n8981), .B2(n6485), .ZN(n6488)
         );
  INV_X1 U8190 ( .A(n6485), .ZN(n8904) );
  INV_X1 U8191 ( .A(n8981), .ZN(n6483) );
  INV_X1 U8192 ( .A(n6482), .ZN(n8905) );
  AOI21_X1 U8193 ( .B1(n8904), .B2(n6483), .A(n8905), .ZN(n6486) );
  NAND2_X1 U8194 ( .A1(n8905), .A2(n6483), .ZN(n6484) );
  OAI22_X1 U8195 ( .A1(n8906), .A2(n6486), .B1(n6485), .B2(n6484), .ZN(n6487)
         );
  OR2_X1 U8196 ( .A1(n8143), .A2(n6425), .ZN(n6489) );
  NAND2_X1 U8197 ( .A1(n6490), .A2(n6489), .ZN(n6491) );
  XNOR2_X1 U8198 ( .A(n6491), .B(n6383), .ZN(n6493) );
  OAI22_X1 U8199 ( .A1(n9757), .A2(n6425), .B1(n8143), .B2(n6581), .ZN(n6492)
         );
  XNOR2_X1 U8200 ( .A(n6493), .B(n6492), .ZN(n8916) );
  OAI22_X1 U8201 ( .A1(n9753), .A2(n6514), .B1(n6495), .B2(n6425), .ZN(n6494)
         );
  XOR2_X1 U8202 ( .A(n6552), .B(n6494), .Z(n8958) );
  INV_X1 U8203 ( .A(n6495), .ZN(n8996) );
  AOI22_X1 U8204 ( .A1(n8197), .A2(n6579), .B1(n6507), .B2(n8996), .ZN(n8957)
         );
  OAI21_X1 U8205 ( .B1(n8956), .B2(n8958), .A(n8957), .ZN(n6497) );
  NAND2_X1 U8206 ( .A1(n6497), .A2(n6496), .ZN(n8878) );
  INV_X1 U8207 ( .A(n8937), .ZN(n9145) );
  NAND2_X1 U8208 ( .A1(n9145), .A2(n6579), .ZN(n6498) );
  NAND2_X1 U8209 ( .A1(n6499), .A2(n6498), .ZN(n6500) );
  XNOR2_X1 U8210 ( .A(n6500), .B(n6552), .ZN(n8876) );
  NAND2_X1 U8211 ( .A1(n9146), .A2(n6579), .ZN(n6502) );
  NAND2_X1 U8212 ( .A1(n9145), .A2(n6507), .ZN(n6501) );
  NAND2_X1 U8213 ( .A1(n6502), .A2(n6501), .ZN(n8875) );
  NOR2_X1 U8214 ( .A1(n8876), .A2(n8875), .ZN(n6505) );
  INV_X1 U8215 ( .A(n8876), .ZN(n6504) );
  INV_X1 U8216 ( .A(n8875), .ZN(n6503) );
  OAI22_X1 U8217 ( .A1(n9615), .A2(n6514), .B1(n8889), .B2(n6425), .ZN(n6506)
         );
  XOR2_X1 U8218 ( .A(n6383), .B(n6506), .Z(n6509) );
  INV_X1 U8219 ( .A(n8889), .ZN(n9149) );
  AOI22_X1 U8220 ( .A1(n9674), .A2(n6579), .B1(n6507), .B2(n9149), .ZN(n6508)
         );
  NAND2_X1 U8221 ( .A1(n6509), .A2(n6508), .ZN(n6510) );
  OAI21_X1 U8222 ( .B1(n6509), .B2(n6508), .A(n6510), .ZN(n8936) );
  INV_X1 U8223 ( .A(n9669), .ZN(n8894) );
  OAI22_X1 U8224 ( .A1(n8894), .A2(n6425), .B1(n8938), .B2(n6581), .ZN(n6518)
         );
  INV_X1 U8225 ( .A(n8938), .ZN(n9151) );
  NAND2_X1 U8226 ( .A1(n9151), .A2(n6579), .ZN(n6511) );
  NAND2_X1 U8227 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  XNOR2_X1 U8228 ( .A(n6513), .B(n6383), .ZN(n6517) );
  XOR2_X1 U8229 ( .A(n6518), .B(n6517), .Z(n8887) );
  OAI22_X1 U8230 ( .A1(n8951), .A2(n6514), .B1(n8995), .B2(n6425), .ZN(n6515)
         );
  XOR2_X1 U8231 ( .A(n6552), .B(n6515), .Z(n6526) );
  AND2_X1 U8232 ( .A1(n8887), .A2(n6526), .ZN(n6516) );
  NAND2_X1 U8233 ( .A1(n8886), .A2(n6516), .ZN(n6523) );
  INV_X1 U8234 ( .A(n6526), .ZN(n6521) );
  INV_X1 U8235 ( .A(n6517), .ZN(n6520) );
  INV_X1 U8236 ( .A(n6518), .ZN(n6519) );
  NAND2_X1 U8237 ( .A1(n6520), .A2(n6519), .ZN(n6524) );
  INV_X1 U8238 ( .A(n6524), .ZN(n6525) );
  NAND2_X1 U8239 ( .A1(n8885), .A2(n4978), .ZN(n6527) );
  OAI22_X1 U8240 ( .A1(n8951), .A2(n6425), .B1(n8995), .B2(n6581), .ZN(n8946)
         );
  OR2_X1 U8241 ( .A1(n8947), .A2(n6425), .ZN(n6529) );
  NAND2_X1 U8242 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  XNOR2_X1 U8243 ( .A(n6531), .B(n6577), .ZN(n6534) );
  NOR2_X1 U8244 ( .A1(n8947), .A2(n6581), .ZN(n6532) );
  AOI21_X1 U8245 ( .B1(n9659), .B2(n6579), .A(n6532), .ZN(n6533) );
  OR2_X1 U8246 ( .A1(n6534), .A2(n6533), .ZN(n6535) );
  INV_X1 U8247 ( .A(n8899), .ZN(n9156) );
  NAND2_X1 U8248 ( .A1(n9156), .A2(n6579), .ZN(n6537) );
  NAND2_X1 U8249 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  XNOR2_X1 U8250 ( .A(n6539), .B(n6577), .ZN(n6541) );
  NOR2_X1 U8251 ( .A1(n8899), .A2(n6581), .ZN(n6540) );
  AOI21_X1 U8252 ( .B1(n9655), .B2(n6579), .A(n6540), .ZN(n6542) );
  NAND2_X1 U8253 ( .A1(n6541), .A2(n6542), .ZN(n6546) );
  INV_X1 U8254 ( .A(n6541), .ZN(n6544) );
  INV_X1 U8255 ( .A(n6542), .ZN(n6543) );
  NAND2_X1 U8256 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  OAI22_X1 U8257 ( .A1(n9230), .A2(n6425), .B1(n8971), .B2(n6581), .ZN(n6556)
         );
  OR2_X1 U8258 ( .A1(n8971), .A2(n6425), .ZN(n6547) );
  NAND2_X1 U8259 ( .A1(n6548), .A2(n6547), .ZN(n6549) );
  XNOR2_X1 U8260 ( .A(n6549), .B(n6383), .ZN(n6555) );
  OR2_X1 U8261 ( .A1(n8994), .A2(n6425), .ZN(n6550) );
  NAND2_X1 U8262 ( .A1(n6551), .A2(n6550), .ZN(n6553) );
  XNOR2_X1 U8263 ( .A(n6553), .B(n6552), .ZN(n6569) );
  NOR2_X1 U8264 ( .A1(n8994), .A2(n6581), .ZN(n6554) );
  AOI21_X1 U8265 ( .B1(n9643), .B2(n6579), .A(n6554), .ZN(n6570) );
  XNOR2_X1 U8266 ( .A(n6569), .B(n6570), .ZN(n8969) );
  INV_X1 U8267 ( .A(n6555), .ZN(n6558) );
  INV_X1 U8268 ( .A(n6556), .ZN(n6557) );
  NAND2_X1 U8269 ( .A1(n6558), .A2(n6557), .ZN(n8970) );
  OR2_X1 U8270 ( .A1(n8993), .A2(n6425), .ZN(n6560) );
  NAND2_X1 U8271 ( .A1(n6561), .A2(n6560), .ZN(n6562) );
  XNOR2_X1 U8272 ( .A(n6562), .B(n6577), .ZN(n6566) );
  INV_X1 U8273 ( .A(n6566), .ZN(n6568) );
  NOR2_X1 U8274 ( .A1(n8993), .A2(n6581), .ZN(n6563) );
  AOI21_X1 U8275 ( .B1(n9640), .B2(n6564), .A(n6563), .ZN(n6565) );
  INV_X1 U8276 ( .A(n6565), .ZN(n6567) );
  AOI21_X1 U8277 ( .B1(n6568), .B2(n6567), .A(n6592), .ZN(n8854) );
  INV_X1 U8278 ( .A(n8854), .ZN(n6573) );
  INV_X1 U8279 ( .A(n6569), .ZN(n6571) );
  OR2_X1 U8280 ( .A1(n6571), .A2(n6570), .ZN(n8855) );
  INV_X1 U8281 ( .A(n8855), .ZN(n6572) );
  OR2_X1 U8282 ( .A1(n9167), .A2(n6425), .ZN(n6575) );
  NAND2_X1 U8283 ( .A1(n6576), .A2(n6575), .ZN(n6578) );
  XNOR2_X1 U8284 ( .A(n6578), .B(n6577), .ZN(n6583) );
  NAND2_X1 U8285 ( .A1(n9633), .A2(n6579), .ZN(n6580) );
  OAI21_X1 U8286 ( .B1(n9167), .B2(n6581), .A(n6580), .ZN(n6582) );
  XNOR2_X1 U8287 ( .A(n6583), .B(n6582), .ZN(n6614) );
  INV_X1 U8288 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U8289 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  OR2_X1 U8290 ( .A1(n9689), .A2(n6586), .ZN(n6587) );
  NAND2_X1 U8291 ( .A1(n6587), .A2(n9691), .ZN(n7266) );
  OR2_X1 U8292 ( .A1(n7267), .A2(n7266), .ZN(n6604) );
  INV_X1 U8293 ( .A(n6980), .ZN(n9690) );
  NAND2_X1 U8294 ( .A1(n6588), .A2(n10076), .ZN(n6596) );
  INV_X1 U8295 ( .A(n6596), .ZN(n6589) );
  NAND2_X1 U8296 ( .A1(n9690), .A2(n6589), .ZN(n6590) );
  OR2_X1 U8297 ( .A1(n6592), .A2(n9791), .ZN(n6591) );
  NAND3_X1 U8298 ( .A1(n6614), .A2(n8968), .A3(n6592), .ZN(n6610) );
  NOR2_X1 U8299 ( .A1(n7313), .A2(n6593), .ZN(n7280) );
  NAND2_X1 U8300 ( .A1(n9690), .A2(n7280), .ZN(n6595) );
  OAI21_X2 U8301 ( .B1(n6604), .B2(n6595), .A(n9949), .ZN(n8988) );
  INV_X1 U8302 ( .A(n7020), .ZN(n7314) );
  NAND2_X1 U8303 ( .A1(n7022), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7771) );
  NAND3_X1 U8304 ( .A1(n7314), .A2(n6596), .A3(n7771), .ZN(n6597) );
  NAND2_X1 U8305 ( .A1(n6604), .A2(n6597), .ZN(n7045) );
  NAND3_X1 U8306 ( .A1(n7045), .A2(n6379), .A3(n6598), .ZN(n6599) );
  NAND2_X1 U8307 ( .A1(n6599), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6601) );
  INV_X1 U8308 ( .A(n6600), .ZN(n8023) );
  INV_X1 U8309 ( .A(n7017), .ZN(n6602) );
  NAND2_X1 U8310 ( .A1(n9690), .A2(n6602), .ZN(n6603) );
  OR2_X1 U8311 ( .A1(n7257), .A2(n8972), .ZN(n6606) );
  NAND2_X1 U8312 ( .A1(n6981), .A2(n9009), .ZN(n9140) );
  OR2_X1 U8313 ( .A1(n8993), .A2(n9140), .ZN(n6605) );
  NAND2_X1 U8314 ( .A1(n6606), .A2(n6605), .ZN(n9181) );
  INV_X1 U8315 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n8274) );
  AOI22_X1 U8316 ( .A1(n4438), .A2(n9181), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6607) );
  OAI21_X1 U8317 ( .B1(n9796), .B2(n9184), .A(n6607), .ZN(n6608) );
  AOI21_X1 U8318 ( .B1(n9633), .B2(n8988), .A(n6608), .ZN(n6609) );
  INV_X1 U8319 ( .A(n6613), .ZN(n8857) );
  NAND2_X1 U8320 ( .A1(n8857), .A2(n6615), .ZN(n6616) );
  NAND2_X1 U8321 ( .A1(n6617), .A2(n6616), .ZN(P1_U3220) );
  INV_X1 U8322 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6619) );
  OR2_X1 U8323 ( .A1(n6356), .A2(n6619), .ZN(n6624) );
  INV_X1 U8324 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6620) );
  OR2_X1 U8325 ( .A1(n6621), .A2(n6620), .ZN(n6623) );
  INV_X1 U8326 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9406) );
  OR2_X1 U8327 ( .A1(n5072), .A2(n9406), .ZN(n6622) );
  NAND4_X1 U8328 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n8544)
         );
  NOR2_X1 U8329 ( .A1(n8793), .A2(n8544), .ZN(n6829) );
  INV_X1 U8330 ( .A(n8793), .ZN(n8730) );
  INV_X1 U8331 ( .A(n8544), .ZN(n6626) );
  NAND2_X1 U8332 ( .A1(n8272), .A2(n6627), .ZN(n6629) );
  OR2_X1 U8333 ( .A1(n5107), .A2(n8849), .ZN(n6628) );
  NOR2_X1 U8334 ( .A1(n6657), .A2(n7514), .ZN(n6814) );
  INV_X1 U8335 ( .A(n6814), .ZN(n6827) );
  NAND2_X1 U8336 ( .A1(n6799), .A2(n8574), .ZN(n8587) );
  INV_X1 U8337 ( .A(n8587), .ZN(n8586) );
  NAND2_X1 U8338 ( .A1(n6792), .A2(n6791), .ZN(n8615) );
  INV_X1 U8339 ( .A(n6787), .ZN(n6789) );
  NAND2_X1 U8340 ( .A1(n8154), .A2(n6632), .ZN(n8104) );
  INV_X1 U8341 ( .A(n8104), .ZN(n8106) );
  AND2_X1 U8342 ( .A1(n6740), .A2(n6739), .ZN(n8044) );
  INV_X1 U8343 ( .A(n8044), .ZN(n8046) );
  AND2_X1 U8344 ( .A1(n6633), .A2(n7554), .ZN(n6635) );
  AND2_X1 U8345 ( .A1(n6671), .A2(n7502), .ZN(n8783) );
  INV_X1 U8346 ( .A(n7505), .ZN(n6634) );
  NAND4_X1 U8347 ( .A1(n6635), .A2(n8783), .A3(n6634), .A4(n7747), .ZN(n6637)
         );
  INV_X1 U8348 ( .A(n7678), .ZN(n7676) );
  XNOR2_X1 U8349 ( .A(n8436), .B(n10271), .ZN(n7753) );
  NAND2_X1 U8350 ( .A1(n7676), .A2(n7753), .ZN(n6636) );
  NOR2_X1 U8351 ( .A1(n6637), .A2(n6636), .ZN(n6639) );
  NAND4_X1 U8352 ( .A1(n6639), .A2(n8246), .A3(n7867), .A4(n6638), .ZN(n6640)
         );
  NAND2_X1 U8353 ( .A1(n6871), .A2(n7924), .ZN(n7943) );
  NOR2_X1 U8354 ( .A1(n6640), .A2(n7943), .ZN(n6641) );
  NAND4_X1 U8355 ( .A1(n8000), .A2(n7929), .A3(n6641), .A4(n8035), .ZN(n6642)
         );
  NOR2_X1 U8356 ( .A1(n8046), .A2(n6642), .ZN(n6643) );
  NAND2_X1 U8357 ( .A1(n8106), .A2(n6643), .ZN(n6644) );
  OR3_X1 U8358 ( .A1(n8717), .A2(n6645), .A3(n6644), .ZN(n6646) );
  NOR4_X1 U8359 ( .A1(n8665), .A2(n8687), .A3(n8704), .A4(n6646), .ZN(n6647)
         );
  NAND4_X1 U8360 ( .A1(n8623), .A2(n8638), .A3(n8655), .A4(n6647), .ZN(n6648)
         );
  NOR2_X1 U8361 ( .A1(n8615), .A2(n6648), .ZN(n6649) );
  NAND4_X1 U8362 ( .A1(n6801), .A2(n8586), .A3(n8596), .A4(n6649), .ZN(n6650)
         );
  NOR2_X1 U8363 ( .A1(n6651), .A2(n6650), .ZN(n6652) );
  NAND4_X1 U8364 ( .A1(n6827), .A2(n6653), .A3(n6652), .A4(n6826), .ZN(n6654)
         );
  NOR3_X1 U8365 ( .A1(n6829), .A2(n6832), .A3(n6654), .ZN(n6655) );
  AOI21_X1 U8366 ( .B1(n8793), .B2(n6657), .A(n6832), .ZN(n6658) );
  NAND2_X1 U8367 ( .A1(n6659), .A2(n6658), .ZN(n6662) );
  AOI21_X1 U8368 ( .B1(n8544), .B2(n6827), .A(n8793), .ZN(n6660) );
  NOR2_X1 U8369 ( .A1(n6660), .A2(n7853), .ZN(n6661) );
  NAND2_X1 U8370 ( .A1(n6662), .A2(n6661), .ZN(n6663) );
  NAND2_X1 U8371 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  NAND2_X1 U8372 ( .A1(n4444), .A2(n6846), .ZN(n6689) );
  NAND2_X1 U8373 ( .A1(n8438), .A2(n10256), .ZN(n6666) );
  NAND2_X1 U8374 ( .A1(n6689), .A2(n6666), .ZN(n6669) );
  NAND2_X1 U8375 ( .A1(n7615), .A2(n6667), .ZN(n6668) );
  NAND3_X1 U8376 ( .A1(n6676), .A2(n6838), .A3(n6671), .ZN(n6672) );
  AOI22_X1 U8377 ( .A1(n6673), .A2(n6672), .B1(n6847), .B2(n7853), .ZN(n6675)
         );
  INV_X1 U8378 ( .A(n6676), .ZN(n6677) );
  INV_X1 U8379 ( .A(n7608), .ZN(n8437) );
  NAND2_X1 U8380 ( .A1(n8437), .A2(n5632), .ZN(n6684) );
  MUX2_X1 U8381 ( .A(n7749), .B(n6684), .S(n6959), .Z(n6681) );
  INV_X1 U8382 ( .A(n7615), .ZN(n6685) );
  OAI211_X1 U8383 ( .C1(n6692), .C2(n6685), .A(n6693), .B(n6684), .ZN(n6686)
         );
  NAND2_X1 U8384 ( .A1(n6686), .A2(n6690), .ZN(n6688) );
  AOI21_X1 U8385 ( .B1(n6688), .B2(n6695), .A(n6687), .ZN(n6700) );
  INV_X1 U8386 ( .A(n6689), .ZN(n6691) );
  OAI211_X1 U8387 ( .C1(n6692), .C2(n6691), .A(n6690), .B(n7749), .ZN(n6694)
         );
  NAND2_X1 U8388 ( .A1(n6694), .A2(n6693), .ZN(n6698) );
  INV_X1 U8389 ( .A(n6695), .ZN(n6696) );
  AOI21_X1 U8390 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(n6699) );
  NAND2_X1 U8391 ( .A1(n6714), .A2(n6702), .ZN(n6704) );
  NAND2_X1 U8392 ( .A1(n6711), .A2(n6710), .ZN(n6703) );
  MUX2_X1 U8393 ( .A(n6704), .B(n6703), .S(n6959), .Z(n6709) );
  NOR2_X1 U8394 ( .A1(n6709), .A2(n7796), .ZN(n6718) );
  INV_X1 U8395 ( .A(n6705), .ZN(n6706) );
  NOR2_X1 U8396 ( .A1(n6707), .A2(n6706), .ZN(n6708) );
  OAI211_X1 U8397 ( .C1(n6709), .C2(n6708), .A(n7924), .B(n6711), .ZN(n6716)
         );
  NAND3_X1 U8398 ( .A1(n6712), .A2(n6711), .A3(n6710), .ZN(n6713) );
  NAND3_X1 U8399 ( .A1(n6871), .A2(n6714), .A3(n6713), .ZN(n6715) );
  MUX2_X1 U8400 ( .A(n6716), .B(n6715), .S(n6959), .Z(n6717) );
  MUX2_X1 U8401 ( .A(n8025), .B(n6720), .S(n6959), .Z(n6727) );
  MUX2_X1 U8402 ( .A(n6722), .B(n6721), .S(n6959), .Z(n6723) );
  INV_X1 U8403 ( .A(n6723), .ZN(n6725) );
  OAI21_X1 U8404 ( .B1(n6728), .B2(n6727), .A(n6726), .ZN(n6733) );
  NAND2_X1 U8405 ( .A1(n8127), .A2(n7932), .ZN(n6729) );
  MUX2_X1 U8406 ( .A(n6730), .B(n6729), .S(n6959), .Z(n6731) );
  NAND2_X1 U8407 ( .A1(n6733), .A2(n6732), .ZN(n6738) );
  MUX2_X1 U8408 ( .A(n6735), .B(n6734), .S(n6959), .Z(n6736) );
  NAND2_X1 U8409 ( .A1(n6738), .A2(n6737), .ZN(n6742) );
  MUX2_X1 U8410 ( .A(n6740), .B(n6739), .S(n6959), .Z(n6741) );
  OAI211_X1 U8411 ( .C1(n6754), .C2(n6743), .A(n6788), .B(n6755), .ZN(n6747)
         );
  AOI21_X1 U8412 ( .B1(n6751), .B2(n6744), .A(n6959), .ZN(n6745) );
  AOI21_X1 U8413 ( .B1(n6747), .B2(n6746), .A(n6745), .ZN(n6763) );
  NOR2_X1 U8414 ( .A1(n6748), .A2(n6959), .ZN(n6749) );
  OR2_X2 U8415 ( .A1(n6763), .A2(n6750), .ZN(n6753) );
  INV_X1 U8416 ( .A(n6754), .ZN(n6759) );
  NOR2_X1 U8417 ( .A1(n4843), .A2(n4844), .ZN(n6758) );
  INV_X1 U8418 ( .A(n6756), .ZN(n6757) );
  AOI211_X1 U8419 ( .C1(n6759), .C2(n6758), .A(n6788), .B(n6757), .ZN(n6762)
         );
  OAI211_X1 U8420 ( .C1(n6763), .C2(n6762), .A(n6761), .B(n6760), .ZN(n6764)
         );
  NAND3_X1 U8421 ( .A1(n6765), .A2(n6766), .A3(n6764), .ZN(n6776) );
  INV_X1 U8422 ( .A(n8650), .ZN(n6768) );
  INV_X1 U8423 ( .A(n6766), .ZN(n6767) );
  NOR2_X1 U8424 ( .A1(n6768), .A2(n6767), .ZN(n6771) );
  NOR2_X1 U8425 ( .A1(n8665), .A2(n6769), .ZN(n6770) );
  MUX2_X1 U8426 ( .A(n6771), .B(n6770), .S(n6959), .Z(n6775) );
  NAND2_X1 U8427 ( .A1(n6780), .A2(n8649), .ZN(n6773) );
  AOI21_X2 U8428 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n6783) );
  NAND2_X1 U8429 ( .A1(n8638), .A2(n6777), .ZN(n6779) );
  OAI21_X1 U8430 ( .B1(n6783), .B2(n6779), .A(n6778), .ZN(n6785) );
  NAND2_X1 U8431 ( .A1(n8638), .A2(n6780), .ZN(n6782) );
  OAI211_X1 U8432 ( .C1(n6783), .C2(n6782), .A(n6786), .B(n6781), .ZN(n6784)
         );
  INV_X1 U8433 ( .A(n6792), .ZN(n6793) );
  MUX2_X1 U8434 ( .A(n6796), .B(n6795), .S(n6959), .Z(n6797) );
  AOI21_X1 U8435 ( .B1(n6798), .B2(n8596), .A(n6797), .ZN(n6802) );
  MUX2_X1 U8436 ( .A(n6799), .B(n8574), .S(n6959), .Z(n6800) );
  NAND2_X1 U8437 ( .A1(n6804), .A2(n6803), .ZN(n6806) );
  MUX2_X1 U8438 ( .A(n6808), .B(n6807), .S(n6959), .Z(n6809) );
  AOI21_X1 U8439 ( .B1(n8563), .B2(n6959), .A(n6811), .ZN(n6820) );
  AOI21_X1 U8440 ( .B1(n6818), .B2(n4503), .A(n6788), .ZN(n6822) );
  NOR2_X1 U8441 ( .A1(n6822), .A2(n6821), .ZN(n6823) );
  INV_X1 U8442 ( .A(n6831), .ZN(n6825) );
  NAND2_X1 U8443 ( .A1(n6825), .A2(n6959), .ZN(n6834) );
  INV_X1 U8444 ( .A(n6826), .ZN(n6828) );
  OAI21_X1 U8445 ( .B1(n6828), .B2(n6959), .A(n6827), .ZN(n6830) );
  AOI21_X2 U8446 ( .B1(n6834), .B2(n6833), .A(n6832), .ZN(n6835) );
  INV_X1 U8447 ( .A(n6960), .ZN(n7168) );
  NAND2_X1 U8448 ( .A1(n7168), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8019) );
  INV_X1 U8449 ( .A(n8019), .ZN(n6836) );
  NOR2_X1 U8450 ( .A1(n8845), .A2(n6948), .ZN(n6942) );
  INV_X1 U8451 ( .A(n7138), .ZN(n7133) );
  NAND3_X1 U8452 ( .A1(n6942), .A2(n7133), .A3(n7642), .ZN(n6837) );
  OAI211_X1 U8453 ( .C1(n6838), .C2(n8019), .A(n6837), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6839) );
  XNOR2_X1 U8454 ( .A(n7499), .B(n7823), .ZN(n6840) );
  AND2_X1 U8455 ( .A1(n6841), .A2(n6840), .ZN(n6842) );
  NAND2_X1 U8456 ( .A1(n6843), .A2(n6842), .ZN(n6845) );
  XNOR2_X1 U8457 ( .A(n10276), .B(n6919), .ZN(n6858) );
  XNOR2_X1 U8458 ( .A(n6846), .B(n6851), .ZN(n6855) );
  XNOR2_X1 U8459 ( .A(n6849), .B(n6850), .ZN(n7226) );
  XNOR2_X1 U8460 ( .A(n10256), .B(n6851), .ZN(n6853) );
  XNOR2_X1 U8461 ( .A(n6852), .B(n6853), .ZN(n7232) );
  XNOR2_X1 U8462 ( .A(n6855), .B(n7622), .ZN(n7259) );
  XNOR2_X1 U8463 ( .A(n10266), .B(n6851), .ZN(n6856) );
  XNOR2_X1 U8464 ( .A(n7608), .B(n6856), .ZN(n7485) );
  XNOR2_X1 U8465 ( .A(n7611), .B(n6851), .ZN(n6857) );
  XNOR2_X1 U8466 ( .A(n6857), .B(n8436), .ZN(n7606) );
  OAI22_X1 U8467 ( .A1(n7605), .A2(n7606), .B1(n6857), .B2(n8436), .ZN(n7765)
         );
  XNOR2_X1 U8468 ( .A(n6858), .B(n8435), .ZN(n7766) );
  XNOR2_X1 U8469 ( .A(n10281), .B(n6851), .ZN(n6859) );
  XNOR2_X1 U8470 ( .A(n6859), .B(n7681), .ZN(n7787) );
  OR2_X1 U8471 ( .A1(n6859), .A2(n8434), .ZN(n6860) );
  XNOR2_X1 U8472 ( .A(n7802), .B(n6851), .ZN(n6861) );
  XNOR2_X1 U8473 ( .A(n6861), .B(n6862), .ZN(n7855) );
  INV_X1 U8474 ( .A(n6861), .ZN(n6863) );
  XNOR2_X1 U8475 ( .A(n7884), .B(n6851), .ZN(n6865) );
  XNOR2_X1 U8476 ( .A(n6865), .B(n5211), .ZN(n7877) );
  INV_X1 U8477 ( .A(n6865), .ZN(n6866) );
  NAND2_X1 U8478 ( .A1(n6866), .A2(n5211), .ZN(n6867) );
  XNOR2_X1 U8479 ( .A(n7929), .B(n6919), .ZN(n8179) );
  XOR2_X1 U8480 ( .A(n6919), .B(n10301), .Z(n8176) );
  INV_X1 U8481 ( .A(n8176), .ZN(n6868) );
  NAND2_X1 U8482 ( .A1(n8175), .A2(n6870), .ZN(n6878) );
  INV_X1 U8483 ( .A(n6871), .ZN(n7923) );
  NOR2_X1 U8484 ( .A1(n8134), .A2(n6919), .ZN(n6872) );
  INV_X1 U8485 ( .A(n7929), .ZN(n7926) );
  AOI211_X1 U8486 ( .C1(n7923), .C2(n6919), .A(n6872), .B(n7926), .ZN(n6876)
         );
  NOR2_X1 U8487 ( .A1(n8134), .A2(n6921), .ZN(n6873) );
  AOI211_X1 U8488 ( .C1(n6921), .C2(n6874), .A(n6873), .B(n7929), .ZN(n6875)
         );
  NAND2_X1 U8489 ( .A1(n6878), .A2(n6877), .ZN(n8130) );
  XNOR2_X1 U8490 ( .A(n8127), .B(n6851), .ZN(n6879) );
  XNOR2_X1 U8491 ( .A(n6879), .B(n8430), .ZN(n8129) );
  OR2_X1 U8492 ( .A1(n6879), .A2(n7932), .ZN(n6880) );
  XNOR2_X1 U8493 ( .A(n8377), .B(n6851), .ZN(n6881) );
  XNOR2_X1 U8494 ( .A(n6881), .B(n8037), .ZN(n8371) );
  XNOR2_X1 U8495 ( .A(n8300), .B(n6919), .ZN(n6883) );
  XNOR2_X1 U8496 ( .A(n6883), .B(n8428), .ZN(n8294) );
  AOI21_X1 U8497 ( .B1(n8295), .B2(n8294), .A(n6884), .ZN(n8406) );
  XNOR2_X1 U8498 ( .A(n8405), .B(n6851), .ZN(n6885) );
  XNOR2_X1 U8499 ( .A(n6885), .B(n8427), .ZN(n8409) );
  NAND2_X1 U8500 ( .A1(n8406), .A2(n8409), .ZN(n8408) );
  XNOR2_X1 U8501 ( .A(n8339), .B(n6919), .ZN(n6887) );
  NAND2_X1 U8502 ( .A1(n6887), .A2(n8719), .ZN(n8330) );
  INV_X1 U8503 ( .A(n6887), .ZN(n6888) );
  NAND2_X1 U8504 ( .A1(n6888), .A2(n8426), .ZN(n8331) );
  XNOR2_X1 U8505 ( .A(n8711), .B(n6919), .ZN(n6889) );
  XNOR2_X1 U8506 ( .A(n6889), .B(n8334), .ZN(n8342) );
  XNOR2_X1 U8507 ( .A(n8703), .B(n6919), .ZN(n6893) );
  XNOR2_X1 U8508 ( .A(n6893), .B(n8425), .ZN(n8386) );
  XNOR2_X1 U8509 ( .A(n8768), .B(n6919), .ZN(n6894) );
  NAND2_X1 U8510 ( .A1(n6894), .A2(n8693), .ZN(n6892) );
  AND2_X1 U8511 ( .A1(n8386), .A2(n6892), .ZN(n8357) );
  XNOR2_X1 U8512 ( .A(n8832), .B(n6919), .ZN(n6897) );
  XNOR2_X1 U8513 ( .A(n6897), .B(n8678), .ZN(n8361) );
  INV_X1 U8514 ( .A(n8361), .ZN(n6890) );
  AND2_X1 U8515 ( .A1(n8357), .A2(n6890), .ZN(n6891) );
  NAND2_X1 U8516 ( .A1(n8310), .A2(n6891), .ZN(n6901) );
  INV_X1 U8517 ( .A(n6892), .ZN(n6896) );
  NAND2_X1 U8518 ( .A1(n6893), .A2(n8721), .ZN(n8311) );
  XNOR2_X1 U8519 ( .A(n6894), .B(n8693), .ZN(n8312) );
  INV_X1 U8520 ( .A(n8312), .ZN(n6895) );
  NAND2_X1 U8521 ( .A1(n6897), .A2(n8678), .ZN(n6898) );
  XOR2_X1 U8522 ( .A(n6919), .B(n5444), .Z(n6903) );
  INV_X1 U8523 ( .A(n6903), .ZN(n6902) );
  XNOR2_X1 U8524 ( .A(n6902), .B(n8667), .ZN(n8279) );
  NOR2_X1 U8525 ( .A1(n6903), .A2(n8667), .ZN(n6904) );
  XNOR2_X1 U8526 ( .A(n8641), .B(n6919), .ZN(n6906) );
  XNOR2_X1 U8527 ( .A(n6905), .B(n6906), .ZN(n8380) );
  NAND2_X1 U8528 ( .A1(n8380), .A2(n8622), .ZN(n6909) );
  INV_X1 U8529 ( .A(n6905), .ZN(n6907) );
  NAND2_X1 U8530 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8531 ( .A(n8749), .B(n6921), .ZN(n6911) );
  XNOR2_X1 U8532 ( .A(n8744), .B(n6919), .ZN(n6912) );
  NAND2_X1 U8533 ( .A1(n6912), .A2(n8621), .ZN(n6913) );
  NAND2_X1 U8534 ( .A1(n6914), .A2(n6913), .ZN(n8322) );
  XNOR2_X1 U8535 ( .A(n8603), .B(n6919), .ZN(n6915) );
  NAND2_X1 U8536 ( .A1(n8322), .A2(n8323), .ZN(n6918) );
  INV_X1 U8537 ( .A(n6915), .ZN(n6916) );
  NAND2_X1 U8538 ( .A1(n6916), .A2(n8611), .ZN(n6917) );
  XNOR2_X1 U8539 ( .A(n8803), .B(n6919), .ZN(n6920) );
  NAND2_X1 U8540 ( .A1(n6920), .A2(n8568), .ZN(n8259) );
  XNOR2_X1 U8541 ( .A(n8735), .B(n6921), .ZN(n6922) );
  NAND2_X1 U8542 ( .A1(n6922), .A2(n7493), .ZN(n8257) );
  OAI21_X1 U8543 ( .B1(n6922), .B2(n7493), .A(n8257), .ZN(n8258) );
  INV_X1 U8544 ( .A(n6923), .ZN(n6924) );
  NAND2_X1 U8545 ( .A1(n6931), .A2(n6924), .ZN(n6927) );
  INV_X1 U8546 ( .A(n6940), .ZN(n6925) );
  NAND2_X1 U8547 ( .A1(n6951), .A2(n6925), .ZN(n6926) );
  AOI21_X1 U8548 ( .B1(n6928), .B2(n8258), .A(n8403), .ZN(n6930) );
  NAND2_X1 U8549 ( .A1(n6930), .A2(n6929), .ZN(n6958) );
  NAND2_X1 U8550 ( .A1(n6931), .A2(n10308), .ZN(n6933) );
  NAND2_X1 U8551 ( .A1(n6933), .A2(n8712), .ZN(n8400) );
  INV_X1 U8552 ( .A(n8400), .ZN(n8419) );
  NOR2_X1 U8553 ( .A1(n4725), .A2(n8419), .ZN(n6956) );
  INV_X1 U8554 ( .A(n6934), .ZN(n6935) );
  AND3_X1 U8555 ( .A1(n6935), .A2(n7169), .A3(n6960), .ZN(n6939) );
  NAND2_X1 U8556 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  OAI211_X1 U8557 ( .C1(n6944), .C2(n6940), .A(n6939), .B(n6938), .ZN(n6941)
         );
  NAND2_X1 U8558 ( .A1(n6941), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6946) );
  INV_X1 U8559 ( .A(n6942), .ZN(n6943) );
  OR2_X1 U8560 ( .A1(n6944), .A2(n6943), .ZN(n6945) );
  NOR2_X1 U8561 ( .A1(n6949), .A2(n6948), .ZN(n6947) );
  NAND2_X1 U8562 ( .A1(n6951), .A2(n6947), .ZN(n8412) );
  INV_X1 U8563 ( .A(n6948), .ZN(n7297) );
  AND2_X1 U8564 ( .A1(n6949), .A2(n7297), .ZN(n6950) );
  AOI22_X1 U8565 ( .A1(n8410), .A2(n8422), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6952) );
  OAI21_X1 U8566 ( .B1(n8568), .B2(n8412), .A(n6952), .ZN(n6953) );
  AOI21_X1 U8567 ( .B1(n8580), .B2(n8415), .A(n6953), .ZN(n6954) );
  NAND2_X1 U8568 ( .A1(n6958), .A2(n6957), .ZN(P2_U3154) );
  NAND2_X1 U8569 ( .A1(n7169), .A2(n6959), .ZN(n6961) );
  NAND2_X1 U8570 ( .A1(n6961), .A2(n6960), .ZN(n7139) );
  NAND2_X1 U8571 ( .A1(n7139), .A2(n6962), .ZN(n6963) );
  NAND2_X1 U8572 ( .A1(n6963), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U8573 ( .A1(n6379), .A2(n8274), .ZN(n6964) );
  AND2_X2 U8574 ( .A1(n6964), .A2(n6982), .ZN(P1_U3973) );
  INV_X1 U8575 ( .A(n6965), .ZN(n6966) );
  INV_X2 U8576 ( .A(n8492), .ZN(P2_U3893) );
  XNOR2_X1 U8577 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8578 ( .A(n9013), .B(n6967), .S(P1_U3086), .Z(n6968) );
  INV_X1 U8579 ( .A(n6968), .ZN(P1_U3355) );
  NOR2_X1 U8580 ( .A1(n5065), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9697) );
  OAI222_X1 U8581 ( .A1(n8277), .A2(n6969), .B1(n8275), .B2(n6970), .C1(n8274), 
        .C2(n7096), .ZN(P1_U3353) );
  NOR2_X1 U8582 ( .A1(n5065), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8289) );
  INV_X2 U8583 ( .A(n8289), .ZN(n8848) );
  AND2_X1 U8584 ( .A1(n5065), .A2(P2_U3151), .ZN(n8288) );
  INV_X1 U8585 ( .A(n9038), .ZN(n7098) );
  OAI222_X1 U8586 ( .A1(n8277), .A2(n6972), .B1(n8275), .B2(n6973), .C1(n8274), 
        .C2(n7098), .ZN(P1_U3352) );
  OAI222_X1 U8587 ( .A1(n8848), .A2(n4559), .B1(n8851), .B2(n6973), .C1(n7158), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  OAI222_X1 U8588 ( .A1(n8275), .A2(n6978), .B1(n9807), .B2(P1_U3086), .C1(
        n5037), .C2(n8277), .ZN(P1_U3354) );
  INV_X1 U8589 ( .A(n7099), .ZN(n9820) );
  INV_X1 U8590 ( .A(n8277), .ZN(n7239) );
  AOI22_X1 U8591 ( .A1(n9835), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n7239), .ZN(n6977) );
  OAI21_X1 U8592 ( .B1(n6992), .B2(n8275), .A(n6977), .ZN(P1_U3350) );
  OAI222_X1 U8593 ( .A1(n8848), .A2(n6979), .B1(n8851), .B2(n6978), .C1(
        P2_U3151), .C2(n10118), .ZN(P2_U3294) );
  NAND2_X1 U8594 ( .A1(n8023), .A2(n6980), .ZN(n6989) );
  NAND2_X1 U8595 ( .A1(n6982), .A2(n6981), .ZN(n6984) );
  NAND2_X1 U8596 ( .A1(n6984), .A2(n6983), .ZN(n6988) );
  INV_X1 U8597 ( .A(n6988), .ZN(n6985) );
  NAND2_X1 U8598 ( .A1(n6989), .A2(n6985), .ZN(n7090) );
  OAI21_X1 U8599 ( .B1(n4451), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9009), .ZN(
        n9014) );
  AOI21_X1 U8600 ( .B1(n4451), .B2(n6986), .A(n9014), .ZN(n6987) );
  XNOR2_X1 U8601 ( .A(n6987), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6991) );
  AND2_X1 U8602 ( .A1(n6989), .A2(n6988), .ZN(n9811) );
  AOI22_X1 U8603 ( .A1(n9811), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6990) );
  OAI21_X1 U8604 ( .B1(n7090), .B2(n6991), .A(n6990), .ZN(P1_U3243) );
  OAI222_X1 U8605 ( .A1(n7389), .A2(P2_U3151), .B1(n8851), .B2(n6992), .C1(
        n9356), .C2(n8848), .ZN(P2_U3290) );
  NOR2_X1 U8606 ( .A1(n9811), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U8607 ( .A1(n6993), .A2(P1_U3973), .ZN(n6994) );
  OAI21_X1 U8608 ( .B1(P1_U3973), .B2(n5903), .A(n6994), .ZN(P1_U3585) );
  NAND2_X1 U8609 ( .A1(n7272), .A2(P1_U3973), .ZN(n6995) );
  OAI21_X1 U8610 ( .B1(P1_U3973), .B2(n5048), .A(n6995), .ZN(P1_U3554) );
  OAI222_X1 U8611 ( .A1(n7391), .A2(P2_U3151), .B1(n8851), .B2(n6996), .C1(
        n7000), .C2(n8848), .ZN(P2_U3289) );
  INV_X1 U8612 ( .A(n9845), .ZN(n7101) );
  OAI222_X1 U8613 ( .A1(n8277), .A2(n6997), .B1(n8275), .B2(n6996), .C1(n8274), 
        .C2(n7101), .ZN(P1_U3349) );
  AOI22_X1 U8614 ( .A1(n9716), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7239), .ZN(n6998) );
  OAI21_X1 U8615 ( .B1(n7006), .B2(n8275), .A(n6998), .ZN(P1_U3348) );
  MUX2_X1 U8616 ( .A(n7033), .B(n7544), .S(P1_U3973), .Z(n6999) );
  INV_X1 U8617 ( .A(n6999), .ZN(P1_U3563) );
  MUX2_X1 U8618 ( .A(n7000), .B(n7475), .S(P1_U3973), .Z(n7001) );
  INV_X1 U8619 ( .A(n7001), .ZN(P1_U3560) );
  MUX2_X1 U8620 ( .A(n7054), .B(n7709), .S(P1_U3973), .Z(n7002) );
  INV_X1 U8621 ( .A(n7002), .ZN(P1_U3565) );
  MUX2_X1 U8622 ( .A(n9356), .B(n7118), .S(P1_U3973), .Z(n7003) );
  INV_X1 U8623 ( .A(n7003), .ZN(P1_U3559) );
  MUX2_X1 U8624 ( .A(n7011), .B(n7476), .S(P1_U3973), .Z(n7004) );
  INV_X1 U8625 ( .A(n7004), .ZN(P1_U3562) );
  OAI222_X1 U8626 ( .A1(n7396), .A2(P2_U3151), .B1(n8851), .B2(n7006), .C1(
        n7005), .C2(n8848), .ZN(P2_U3288) );
  INV_X1 U8627 ( .A(n7007), .ZN(n7012) );
  AOI22_X1 U8628 ( .A1(n9731), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7239), .ZN(n7008) );
  OAI21_X1 U8629 ( .B1(n7012), .B2(n8275), .A(n7008), .ZN(P1_U3347) );
  AND2_X1 U8630 ( .A1(n7010), .A2(n7009), .ZN(n7038) );
  NOR2_X1 U8631 ( .A1(n7038), .A2(n9414), .ZN(P2_U3255) );
  NOR2_X1 U8632 ( .A1(n7038), .A2(n9327), .ZN(P2_U3257) );
  NOR2_X1 U8633 ( .A1(n7038), .A2(n9411), .ZN(P2_U3239) );
  INV_X1 U8634 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n9341) );
  NOR2_X1 U8635 ( .A1(n7038), .A2(n9341), .ZN(P2_U3248) );
  NOR2_X1 U8636 ( .A1(n7038), .A2(n9518), .ZN(P2_U3236) );
  INV_X1 U8637 ( .A(n8447), .ZN(n7638) );
  OAI222_X1 U8638 ( .A1(n7638), .A2(P2_U3151), .B1(n8851), .B2(n7012), .C1(
        n7011), .C2(n8848), .ZN(P2_U3287) );
  INV_X2 U8639 ( .A(n10109), .ZN(n10111) );
  INV_X1 U8640 ( .A(n7014), .ZN(n7016) );
  OR2_X1 U8641 ( .A1(n7937), .A2(n5880), .ZN(n7015) );
  NAND2_X1 U8642 ( .A1(n7016), .A2(n7015), .ZN(n9947) );
  NAND2_X1 U8643 ( .A1(n7018), .A2(n7017), .ZN(n7019) );
  NAND2_X1 U8644 ( .A1(n7313), .A2(n7019), .ZN(n7021) );
  OR2_X1 U8645 ( .A1(n7021), .A2(n7020), .ZN(n9960) );
  OR2_X1 U8646 ( .A1(n7023), .A2(n7022), .ZN(n10085) );
  NAND2_X1 U8647 ( .A1(n9960), .A2(n10085), .ZN(n10080) );
  OAI21_X1 U8648 ( .B1(n9947), .B2(n10080), .A(n7315), .ZN(n7024) );
  INV_X1 U8649 ( .A(n8972), .ZN(n8924) );
  NAND2_X1 U8650 ( .A1(n4440), .A2(n8924), .ZN(n7316) );
  OAI211_X1 U8651 ( .C1(n7313), .C2(n9976), .A(n7024), .B(n7316), .ZN(n7026)
         );
  NAND2_X1 U8652 ( .A1(n7026), .A2(n10111), .ZN(n7025) );
  OAI21_X1 U8653 ( .B1(n10111), .B2(n6986), .A(n7025), .ZN(P1_U3522) );
  INV_X1 U8654 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7028) );
  NAND2_X1 U8655 ( .A1(n7026), .A2(n10092), .ZN(n7027) );
  OAI21_X1 U8656 ( .B1(n10092), .B2(n7028), .A(n7027), .ZN(P1_U3453) );
  INV_X1 U8657 ( .A(n7029), .ZN(n7034) );
  AOI22_X1 U8658 ( .A1(n7434), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n7239), .ZN(n7030) );
  OAI21_X1 U8659 ( .B1(n7034), .B2(n8275), .A(n7030), .ZN(P1_U3346) );
  INV_X1 U8660 ( .A(n7031), .ZN(n7037) );
  AOI22_X1 U8661 ( .A1(n9712), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7239), .ZN(n7032) );
  OAI21_X1 U8662 ( .B1(n7037), .B2(n8275), .A(n7032), .ZN(P1_U3345) );
  INV_X1 U8663 ( .A(n7700), .ZN(n7659) );
  OAI222_X1 U8664 ( .A1(P2_U3151), .A2(n7659), .B1(n8851), .B2(n7034), .C1(
        n7033), .C2(n8848), .ZN(P2_U3286) );
  INV_X1 U8665 ( .A(n7038), .ZN(n7035) );
  AND2_X1 U8666 ( .A1(n7035), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8667 ( .A1(n7035), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8668 ( .A1(n7035), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8669 ( .A1(n7035), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8670 ( .A1(n7035), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8671 ( .A1(n7035), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8672 ( .A1(n7035), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8673 ( .A1(n7035), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8674 ( .A1(n7035), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  INV_X1 U8675 ( .A(n7728), .ZN(n7735) );
  OAI222_X1 U8676 ( .A1(P2_U3151), .A2(n7735), .B1(n8851), .B2(n7037), .C1(
        n7036), .C2(n8848), .ZN(P2_U3285) );
  INV_X1 U8677 ( .A(n8287), .ZN(n7039) );
  NOR4_X1 U8678 ( .A1(n7040), .A2(n7039), .A3(n7168), .A4(P2_U3151), .ZN(n7041) );
  AOI21_X1 U8679 ( .B1(n7035), .B2(n5600), .A(n7041), .ZN(P2_U3376) );
  NAND2_X1 U8680 ( .A1(n5625), .A2(P2_U3893), .ZN(n7042) );
  OAI21_X1 U8681 ( .B1(P2_U3893), .B2(n5034), .A(n7042), .ZN(P2_U3491) );
  AND2_X1 U8682 ( .A1(n7035), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8683 ( .A1(n7035), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8684 ( .A1(n7035), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8685 ( .A1(n7035), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8686 ( .A1(n7035), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8687 ( .A1(n7035), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8688 ( .A1(n7035), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8689 ( .A1(n7035), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8690 ( .A1(n7035), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8691 ( .A1(n7035), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8692 ( .A1(n7035), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8693 ( .A1(n7035), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8694 ( .A1(n7035), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8695 ( .A1(n7035), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8696 ( .A1(n7035), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8697 ( .A1(n7035), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  XOR2_X1 U8698 ( .A(n7043), .B(n7044), .Z(n7048) );
  NAND2_X1 U8699 ( .A1(n7045), .A2(n7268), .ZN(n7061) );
  INV_X1 U8700 ( .A(n8988), .ZN(n9786) );
  INV_X1 U8701 ( .A(n4438), .ZN(n8927) );
  INV_X1 U8702 ( .A(n9140), .ZN(n8948) );
  AOI22_X1 U8703 ( .A1(n8948), .A2(n4440), .B1(n9006), .B2(n8924), .ZN(n7277)
         );
  OAI22_X1 U8704 ( .A1(n7287), .A2(n9786), .B1(n8927), .B2(n7277), .ZN(n7046)
         );
  AOI21_X1 U8705 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7061), .A(n7046), .ZN(
        n7047) );
  OAI21_X1 U8706 ( .B1(n7048), .B2(n9791), .A(n7047), .ZN(P1_U3237) );
  XNOR2_X1 U8707 ( .A(n7050), .B(n7049), .ZN(n9010) );
  OAI22_X1 U8708 ( .A1(n9786), .A2(n9976), .B1(n8927), .B2(n7316), .ZN(n7051)
         );
  AOI21_X1 U8709 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7061), .A(n7051), .ZN(
        n7052) );
  OAI21_X1 U8710 ( .B1(n9791), .B2(n9010), .A(n7052), .ZN(P1_U3232) );
  INV_X1 U8711 ( .A(n7835), .ZN(n7840) );
  INV_X1 U8712 ( .A(n7053), .ZN(n7055) );
  OAI222_X1 U8713 ( .A1(n7840), .A2(P2_U3151), .B1(n8851), .B2(n7055), .C1(
        n7054), .C2(n8848), .ZN(P2_U3284) );
  INV_X1 U8714 ( .A(n9862), .ZN(n7432) );
  OAI222_X1 U8715 ( .A1(n8277), .A2(n9332), .B1(n8275), .B2(n7055), .C1(n8274), 
        .C2(n7432), .ZN(P1_U3344) );
  XOR2_X1 U8716 ( .A(n7057), .B(n7056), .Z(n7060) );
  INV_X1 U8717 ( .A(n9007), .ZN(n7067) );
  OAI22_X1 U8718 ( .A1(n7067), .A2(n9140), .B1(n7358), .B2(n8972), .ZN(n9946)
         );
  AOI22_X1 U8719 ( .A1(n9946), .A2(n4438), .B1(n8988), .B2(n6403), .ZN(n7059)
         );
  MUX2_X1 U8720 ( .A(n9796), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7058) );
  OAI211_X1 U8721 ( .C1(n7060), .C2(n9791), .A(n7059), .B(n7058), .ZN(P1_U3218) );
  INV_X1 U8722 ( .A(n7061), .ZN(n7071) );
  INV_X1 U8723 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7070) );
  OAI21_X1 U8724 ( .B1(n7062), .B2(n7064), .A(n7063), .ZN(n7065) );
  NAND2_X1 U8725 ( .A1(n7065), .A2(n8968), .ZN(n7069) );
  OAI22_X1 U8726 ( .A1(n7067), .A2(n8972), .B1(n7066), .B2(n9140), .ZN(n9966)
         );
  AOI22_X1 U8727 ( .A1(n9966), .A2(n4438), .B1(n8988), .B2(n7273), .ZN(n7068)
         );
  OAI211_X1 U8728 ( .C1(n7071), .C2(n7070), .A(n7069), .B(n7068), .ZN(P1_U3222) );
  INV_X1 U8729 ( .A(n7072), .ZN(n7113) );
  AOI22_X1 U8730 ( .A1(n9062), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7239), .ZN(n7073) );
  OAI21_X1 U8731 ( .B1(n7113), .B2(n8275), .A(n7073), .ZN(P1_U3343) );
  INV_X1 U8732 ( .A(n7434), .ZN(n7112) );
  OR2_X1 U8733 ( .A1(n7090), .A2(n9009), .ZN(n9821) );
  OR2_X1 U8734 ( .A1(n7090), .A2(n7074), .ZN(n9910) );
  INV_X1 U8735 ( .A(n9910), .ZN(n9861) );
  XNOR2_X1 U8736 ( .A(n7096), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U8737 ( .A1(n7092), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7077) );
  OR2_X1 U8738 ( .A1(n7092), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7075) );
  NAND2_X1 U8739 ( .A1(n7075), .A2(n7077), .ZN(n9799) );
  NOR3_X1 U8740 ( .A1(n9013), .A2(n6986), .A3(n9799), .ZN(n9797) );
  INV_X1 U8741 ( .A(n9797), .ZN(n7076) );
  NAND2_X1 U8742 ( .A1(n7077), .A2(n7076), .ZN(n9024) );
  NAND2_X1 U8743 ( .A1(n9023), .A2(n9024), .ZN(n9028) );
  INV_X1 U8744 ( .A(n7096), .ZN(n9031) );
  NAND2_X1 U8745 ( .A1(n9031), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7078) );
  NAND2_X1 U8746 ( .A1(n9028), .A2(n7078), .ZN(n9040) );
  XNOR2_X1 U8747 ( .A(n9038), .B(n10095), .ZN(n9041) );
  NAND2_X1 U8748 ( .A1(n9040), .A2(n9041), .ZN(n9039) );
  NAND2_X1 U8749 ( .A1(n9038), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U8750 ( .A1(n9039), .A2(n7079), .ZN(n9813) );
  INV_X1 U8751 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10097) );
  MUX2_X1 U8752 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10097), .S(n7099), .Z(n9814)
         );
  NAND2_X1 U8753 ( .A1(n9813), .A2(n9814), .ZN(n9812) );
  NAND2_X1 U8754 ( .A1(n7099), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U8755 ( .A1(n9812), .A2(n7080), .ZN(n9827) );
  MUX2_X1 U8756 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6121), .S(n9835), .Z(n9828)
         );
  NAND2_X1 U8757 ( .A1(n9827), .A2(n9828), .ZN(n9826) );
  NAND2_X1 U8758 ( .A1(n9835), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n7081) );
  AND2_X1 U8759 ( .A1(n9826), .A2(n7081), .ZN(n9842) );
  INV_X1 U8760 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7082) );
  MUX2_X1 U8761 ( .A(n7082), .B(P1_REG1_REG_6__SCAN_IN), .S(n9845), .Z(n9841)
         );
  NOR2_X1 U8762 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  AOI21_X1 U8763 ( .B1(n9845), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9840), .ZN(
        n9718) );
  OR2_X1 U8764 ( .A1(n9716), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7084) );
  NAND2_X1 U8765 ( .A1(n9716), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7083) );
  NAND2_X1 U8766 ( .A1(n7084), .A2(n7083), .ZN(n9719) );
  NOR2_X1 U8767 ( .A1(n9718), .A2(n9719), .ZN(n9717) );
  AOI21_X1 U8768 ( .B1(n9716), .B2(P1_REG1_REG_7__SCAN_IN), .A(n9717), .ZN(
        n9734) );
  OR2_X1 U8769 ( .A1(n9731), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7086) );
  NAND2_X1 U8770 ( .A1(n9731), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7085) );
  NAND2_X1 U8771 ( .A1(n7086), .A2(n7085), .ZN(n9733) );
  NOR2_X1 U8772 ( .A1(n9734), .A2(n9733), .ZN(n9732) );
  AOI21_X1 U8773 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9731), .A(n9732), .ZN(
        n7089) );
  MUX2_X1 U8774 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n7087), .S(n7434), .Z(n7088)
         );
  NAND2_X1 U8775 ( .A1(n7088), .A2(n7089), .ZN(n7436) );
  OAI21_X1 U8776 ( .B1(n7089), .B2(n7088), .A(n7436), .ZN(n7108) );
  INV_X1 U8777 ( .A(n7090), .ZN(n7091) );
  AND2_X1 U8778 ( .A1(n7091), .A2(n9012), .ZN(n9913) );
  XOR2_X1 U8779 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9038), .Z(n9044) );
  MUX2_X1 U8780 ( .A(n7095), .B(P1_REG2_REG_2__SCAN_IN), .S(n7096), .Z(n9017)
         );
  NAND2_X1 U8781 ( .A1(n7092), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U8782 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9802) );
  NOR2_X1 U8783 ( .A1(n9803), .A2(n9802), .ZN(n9801) );
  INV_X1 U8784 ( .A(n9801), .ZN(n7093) );
  NAND2_X1 U8785 ( .A1(n7094), .A2(n7093), .ZN(n9018) );
  NAND2_X1 U8786 ( .A1(n9017), .A2(n9018), .ZN(n9022) );
  OAI21_X1 U8787 ( .B1(n7096), .B2(n7095), .A(n9022), .ZN(n9043) );
  NAND2_X1 U8788 ( .A1(n9044), .A2(n9043), .ZN(n9042) );
  MUX2_X1 U8789 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n7333), .S(n7099), .Z(n9817)
         );
  NAND2_X1 U8790 ( .A1(n9835), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n7100) );
  OAI21_X1 U8791 ( .B1(n9835), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7100), .ZN(
        n9831) );
  NOR2_X1 U8792 ( .A1(n9832), .A2(n9831), .ZN(n9830) );
  AOI21_X1 U8793 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n9835), .A(n9830), .ZN(
        n9847) );
  AOI22_X1 U8794 ( .A1(n9845), .A2(n7350), .B1(P1_REG2_REG_6__SCAN_IN), .B2(
        n7101), .ZN(n9848) );
  NOR2_X1 U8795 ( .A1(n9847), .A2(n9848), .ZN(n9846) );
  AOI21_X1 U8796 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n9845), .A(n9846), .ZN(
        n9722) );
  NAND2_X1 U8797 ( .A1(n9716), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7102) );
  OAI21_X1 U8798 ( .B1(n9716), .B2(P1_REG2_REG_7__SCAN_IN), .A(n7102), .ZN(
        n9723) );
  NOR2_X1 U8799 ( .A1(n9722), .A2(n9723), .ZN(n9721) );
  NAND2_X1 U8800 ( .A1(n9731), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7103) );
  OAI21_X1 U8801 ( .B1(n9731), .B2(P1_REG2_REG_8__SCAN_IN), .A(n7103), .ZN(
        n9738) );
  MUX2_X1 U8802 ( .A(n7460), .B(P1_REG2_REG_9__SCAN_IN), .S(n7434), .Z(n7104)
         );
  INV_X1 U8803 ( .A(n7104), .ZN(n7105) );
  OAI21_X1 U8804 ( .B1(n7106), .B2(n7105), .A(n7431), .ZN(n7107) );
  AOI22_X1 U8805 ( .A1(n9861), .A2(n7108), .B1(n9913), .B2(n7107), .ZN(n7111)
         );
  NAND2_X1 U8806 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7781) );
  INV_X1 U8807 ( .A(n7781), .ZN(n7109) );
  AOI21_X1 U8808 ( .B1(n9811), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7109), .ZN(
        n7110) );
  OAI211_X1 U8809 ( .C1(n7112), .C2(n9821), .A(n7111), .B(n7110), .ZN(P1_U3252) );
  INV_X1 U8810 ( .A(n8504), .ZN(n7114) );
  OAI222_X1 U8811 ( .A1(P2_U3151), .A2(n7114), .B1(n8851), .B2(n7113), .C1(
        n9449), .C2(n8848), .ZN(P2_U3283) );
  AOI211_X1 U8812 ( .C1(n7117), .C2(n7115), .A(n9791), .B(n7116), .ZN(n7124)
         );
  OR2_X1 U8813 ( .A1(n7118), .A2(n8972), .ZN(n7120) );
  NAND2_X1 U8814 ( .A1(n9006), .A2(n8948), .ZN(n7119) );
  NAND2_X1 U8815 ( .A1(n7120), .A2(n7119), .ZN(n7331) );
  AOI22_X1 U8816 ( .A1(n4438), .A2(n7331), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3086), .ZN(n7122) );
  NAND2_X1 U8817 ( .A1(n8988), .A2(n10014), .ZN(n7121) );
  OAI211_X1 U8818 ( .C1(n9796), .C2(n7336), .A(n7122), .B(n7121), .ZN(n7123)
         );
  OR2_X1 U8819 ( .A1(n7124), .A2(n7123), .ZN(P1_U3230) );
  NAND2_X1 U8820 ( .A1(n8390), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7235) );
  NAND2_X1 U8821 ( .A1(n7235), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7127) );
  AOI22_X1 U8822 ( .A1(n7125), .A2(n8400), .B1(n8410), .B2(n6849), .ZN(n7126)
         );
  OAI211_X1 U8823 ( .C1(n8403), .C2(n8783), .A(n7127), .B(n7126), .ZN(P2_U3172) );
  NOR2_X1 U8824 ( .A1(n7642), .A2(P2_U3151), .ZN(n8232) );
  AND2_X1 U8825 ( .A1(n7139), .A2(n8232), .ZN(n7128) );
  MUX2_X1 U8826 ( .A(P2_U3893), .B(n7128), .S(n7138), .Z(n10232) );
  INV_X1 U8827 ( .A(n10232), .ZN(n7397) );
  MUX2_X1 U8828 ( .A(n7302), .B(n7129), .S(n7642), .Z(n7177) );
  NAND2_X1 U8829 ( .A1(n7177), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U8830 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7642), .Z(n7130) );
  INV_X1 U8831 ( .A(n7130), .ZN(n7131) );
  OAI22_X1 U8832 ( .A1(n7187), .A2(n7186), .B1(n7202), .B2(n7131), .ZN(n7206)
         );
  MUX2_X1 U8833 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n7642), .Z(n7132) );
  XNOR2_X1 U8834 ( .A(n7132), .B(n7158), .ZN(n7207) );
  NOR2_X1 U8835 ( .A1(n7132), .A2(n7158), .ZN(n7135) );
  MUX2_X1 U8836 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n7642), .Z(n7371) );
  XNOR2_X1 U8837 ( .A(n7371), .B(n7385), .ZN(n7134) );
  NOR3_X1 U8838 ( .A1(n7205), .A2(n7135), .A3(n7134), .ZN(n7370) );
  INV_X1 U8839 ( .A(n7370), .ZN(n7137) );
  OR2_X1 U8840 ( .A1(n8492), .A2(n7133), .ZN(n10159) );
  INV_X1 U8841 ( .A(n10159), .ZN(n10240) );
  OAI21_X1 U8842 ( .B1(n7205), .B2(n7135), .A(n7134), .ZN(n7136) );
  NAND3_X1 U8843 ( .A1(n7137), .A2(n10240), .A3(n7136), .ZN(n7176) );
  NOR2_X1 U8844 ( .A1(n7138), .A2(P2_U3151), .ZN(n8235) );
  AND2_X1 U8845 ( .A1(n7139), .A2(n8235), .ZN(n7154) );
  AND2_X1 U8846 ( .A1(n7154), .A2(n7642), .ZN(n10241) );
  MUX2_X1 U8847 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n7140), .S(n7385), .Z(n7153)
         );
  NAND2_X1 U8848 ( .A1(n7142), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U8849 ( .A1(n10118), .A2(n7146), .ZN(n7145) );
  NAND2_X1 U8850 ( .A1(n7178), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7143) );
  OR2_X1 U8851 ( .A1(n7143), .A2(n7142), .ZN(n7144) );
  NAND2_X1 U8852 ( .A1(n7145), .A2(n7144), .ZN(n10115) );
  NAND2_X1 U8853 ( .A1(n10115), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7147) );
  NAND2_X1 U8854 ( .A1(n7147), .A2(n7146), .ZN(n7194) );
  INV_X1 U8855 ( .A(n7158), .ZN(n7219) );
  XNOR2_X1 U8856 ( .A(n7149), .B(n7219), .ZN(n7208) );
  NAND2_X1 U8857 ( .A1(n7208), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7151) );
  NAND2_X1 U8858 ( .A1(n7149), .A2(n7158), .ZN(n7150) );
  NAND2_X1 U8859 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  NAND2_X1 U8860 ( .A1(n7152), .A2(n7153), .ZN(n7368) );
  OAI21_X1 U8861 ( .B1(n7153), .B2(n7152), .A(n7368), .ZN(n7174) );
  INV_X1 U8862 ( .A(n7154), .ZN(n7181) );
  OR2_X1 U8863 ( .A1(n7181), .A2(n7642), .ZN(n10246) );
  INV_X1 U8864 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7582) );
  AND2_X1 U8865 ( .A1(n7178), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8866 ( .A1(n7142), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7156) );
  OAI21_X1 U8867 ( .B1(n10118), .B2(n7155), .A(n7156), .ZN(n10112) );
  OR2_X1 U8868 ( .A1(n10112), .A2(n5017), .ZN(n10114) );
  NAND2_X1 U8869 ( .A1(n10114), .A2(n7156), .ZN(n7190) );
  NAND2_X1 U8870 ( .A1(n7191), .A2(n7190), .ZN(n7189) );
  NAND2_X1 U8871 ( .A1(n7189), .A2(n7157), .ZN(n7159) );
  NAND2_X1 U8872 ( .A1(n7159), .A2(n7158), .ZN(n7163) );
  OR2_X1 U8873 ( .A1(n7159), .A2(n7158), .ZN(n7160) );
  NAND2_X1 U8874 ( .A1(n7213), .A2(n7163), .ZN(n7161) );
  INV_X1 U8875 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7625) );
  XNOR2_X1 U8876 ( .A(n7385), .B(n7625), .ZN(n7162) );
  NAND2_X1 U8877 ( .A1(n7161), .A2(n7162), .ZN(n7387) );
  INV_X1 U8878 ( .A(n7162), .ZN(n7164) );
  NAND3_X1 U8879 ( .A1(n7213), .A2(n7164), .A3(n7163), .ZN(n7165) );
  AND2_X1 U8880 ( .A1(n7387), .A2(n7165), .ZN(n7167) );
  INV_X1 U8881 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9345) );
  NOR2_X1 U8882 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9345), .ZN(n7488) );
  INV_X1 U8883 ( .A(n7488), .ZN(n7166) );
  OAI21_X1 U8884 ( .B1(n10246), .B2(n7167), .A(n7166), .ZN(n7173) );
  NOR2_X1 U8885 ( .A1(n7169), .A2(n7168), .ZN(n7170) );
  OR2_X1 U8886 ( .A1(P2_U3150), .A2(n7170), .ZN(n10163) );
  INV_X1 U8887 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7171) );
  NOR2_X1 U8888 ( .A1(n10163), .A2(n7171), .ZN(n7172) );
  AOI211_X1 U8889 ( .C1(n10241), .C2(n7174), .A(n7173), .B(n7172), .ZN(n7175)
         );
  OAI211_X1 U8890 ( .C1(n7397), .C2(n7385), .A(n7176), .B(n7175), .ZN(P2_U3186) );
  INV_X1 U8891 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7185) );
  INV_X1 U8892 ( .A(n7177), .ZN(n7179) );
  NAND2_X1 U8893 ( .A1(n7179), .A2(n7178), .ZN(n7180) );
  AOI22_X1 U8894 ( .A1(n7181), .A2(n10159), .B1(n10123), .B2(n7180), .ZN(n7182) );
  AOI21_X1 U8895 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n7182), .ZN(
        n7184) );
  NAND2_X1 U8896 ( .A1(n10232), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7183) );
  OAI211_X1 U8897 ( .C1(n10163), .C2(n7185), .A(n7184), .B(n7183), .ZN(
        P2_U3182) );
  XNOR2_X1 U8898 ( .A(n7187), .B(n7186), .ZN(n7204) );
  INV_X1 U8899 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7188) );
  NOR2_X1 U8900 ( .A1(n10163), .A2(n7188), .ZN(n7201) );
  OAI21_X1 U8901 ( .B1(n7191), .B2(n7190), .A(n7189), .ZN(n7192) );
  INV_X1 U8902 ( .A(n7192), .ZN(n7199) );
  OAI21_X1 U8903 ( .B1(n7195), .B2(n7194), .A(n7193), .ZN(n7196) );
  NAND2_X1 U8904 ( .A1(n10241), .A2(n7196), .ZN(n7198) );
  NAND2_X1 U8905 ( .A1(P2_U3151), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7197) );
  OAI211_X1 U8906 ( .C1(n7199), .C2(n10246), .A(n7198), .B(n7197), .ZN(n7200)
         );
  AOI211_X1 U8907 ( .C1(n10232), .C2(n7202), .A(n7201), .B(n7200), .ZN(n7203)
         );
  OAI21_X1 U8908 ( .B1(n7204), .B2(n10159), .A(n7203), .ZN(P2_U3184) );
  AOI21_X1 U8909 ( .B1(n7207), .B2(n7206), .A(n7205), .ZN(n7221) );
  INV_X1 U8910 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7217) );
  XNOR2_X1 U8911 ( .A(n7208), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n7215) );
  INV_X1 U8912 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7209) );
  NOR2_X1 U8913 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7209), .ZN(n7261) );
  INV_X1 U8914 ( .A(n7210), .ZN(n7211) );
  NAND2_X1 U8915 ( .A1(n7211), .A2(n5074), .ZN(n7212) );
  AOI21_X1 U8916 ( .B1(n7213), .B2(n7212), .A(n10246), .ZN(n7214) );
  AOI211_X1 U8917 ( .C1(n10241), .C2(n7215), .A(n7261), .B(n7214), .ZN(n7216)
         );
  OAI21_X1 U8918 ( .B1(n7217), .B2(n10163), .A(n7216), .ZN(n7218) );
  AOI21_X1 U8919 ( .B1(n7219), .B2(n10232), .A(n7218), .ZN(n7220) );
  OAI21_X1 U8920 ( .B1(n7221), .B2(n10159), .A(n7220), .ZN(P2_U3185) );
  INV_X1 U8921 ( .A(n10165), .ZN(n8506) );
  INV_X1 U8922 ( .A(n7222), .ZN(n7223) );
  INV_X1 U8923 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9425) );
  OAI222_X1 U8924 ( .A1(n8506), .A2(P2_U3151), .B1(n8851), .B2(n7223), .C1(
        n9425), .C2(n8848), .ZN(P2_U3282) );
  INV_X1 U8925 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7224) );
  INV_X1 U8926 ( .A(n9881), .ZN(n9060) );
  OAI222_X1 U8927 ( .A1(n8277), .A2(n7224), .B1(n8275), .B2(n7223), .C1(n8274), 
        .C2(n9060), .ZN(P1_U3342) );
  XOR2_X1 U8928 ( .A(n7226), .B(n7225), .Z(n7230) );
  INV_X1 U8929 ( .A(n8412), .ZN(n8387) );
  AOI22_X1 U8930 ( .A1(n8387), .A2(n5625), .B1(n8410), .B2(n8438), .ZN(n7227)
         );
  OAI21_X1 U8931 ( .B1(n6848), .B2(n8419), .A(n7227), .ZN(n7228) );
  AOI21_X1 U8932 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7235), .A(n7228), .ZN(
        n7229) );
  OAI21_X1 U8933 ( .B1(n8403), .B2(n7230), .A(n7229), .ZN(P2_U3162) );
  XOR2_X1 U8934 ( .A(n7232), .B(n7231), .Z(n7237) );
  AOI22_X1 U8935 ( .A1(n8387), .A2(n6849), .B1(n8410), .B2(n4444), .ZN(n7233)
         );
  OAI21_X1 U8936 ( .B1(n10256), .B2(n8419), .A(n7233), .ZN(n7234) );
  AOI21_X1 U8937 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7235), .A(n7234), .ZN(
        n7236) );
  OAI21_X1 U8938 ( .B1(n7237), .B2(n8403), .A(n7236), .ZN(P2_U3177) );
  INV_X1 U8939 ( .A(n7238), .ZN(n7255) );
  AOI22_X1 U8940 ( .A1(n9893), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7239), .ZN(n7240) );
  OAI21_X1 U8941 ( .B1(n7255), .B2(n8275), .A(n7240), .ZN(P1_U3341) );
  INV_X1 U8942 ( .A(n7241), .ZN(n7243) );
  NAND2_X1 U8943 ( .A1(n7243), .A2(n7242), .ZN(n7245) );
  XNOR2_X1 U8944 ( .A(n7245), .B(n7244), .ZN(n7252) );
  OR2_X1 U8945 ( .A1(n7475), .A2(n8972), .ZN(n7247) );
  NAND2_X1 U8946 ( .A1(n9005), .A2(n8948), .ZN(n7246) );
  NAND2_X1 U8947 ( .A1(n7247), .A2(n7246), .ZN(n9931) );
  NOR2_X1 U8948 ( .A1(n7248), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9836) );
  AOI21_X1 U8949 ( .B1(n4438), .B2(n9931), .A(n9836), .ZN(n7250) );
  NAND2_X1 U8950 ( .A1(n8988), .A2(n7361), .ZN(n7249) );
  OAI211_X1 U8951 ( .C1(n9796), .C2(n9933), .A(n7250), .B(n7249), .ZN(n7251)
         );
  AOI21_X1 U8952 ( .B1(n7252), .B2(n8968), .A(n7251), .ZN(n7253) );
  INV_X1 U8953 ( .A(n7253), .ZN(P1_U3227) );
  INV_X1 U8954 ( .A(n10182), .ZN(n8499) );
  INV_X1 U8955 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7254) );
  OAI222_X1 U8956 ( .A1(n8499), .A2(P2_U3151), .B1(n8851), .B2(n7255), .C1(
        n7254), .C2(n8848), .ZN(P2_U3281) );
  INV_X1 U8957 ( .A(P1_U3973), .ZN(n9008) );
  NAND2_X1 U8958 ( .A1(n9008), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7256) );
  OAI21_X1 U8959 ( .B1(n7257), .B2(n9008), .A(n7256), .ZN(P1_U3583) );
  INV_X1 U8960 ( .A(n8403), .ZN(n8407) );
  OAI211_X1 U8961 ( .C1(n7260), .C2(n7259), .A(n7258), .B(n8407), .ZN(n7265)
         );
  INV_X1 U8962 ( .A(n8410), .ZN(n8397) );
  AOI21_X1 U8963 ( .B1(n8387), .B2(n8438), .A(n7261), .ZN(n7262) );
  OAI21_X1 U8964 ( .B1(n7608), .B2(n8397), .A(n7262), .ZN(n7263) );
  AOI21_X1 U8965 ( .B1(n10260), .B2(n8400), .A(n7263), .ZN(n7264) );
  OAI211_X1 U8966 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8390), .A(n7265), .B(
        n7264), .ZN(P2_U3158) );
  INV_X1 U8967 ( .A(n7266), .ZN(n7269) );
  NAND3_X1 U8968 ( .A1(n7269), .A2(n7268), .A3(n7267), .ZN(n7284) );
  AND2_X1 U8969 ( .A1(n9972), .A2(n9960), .ZN(n7270) );
  AND2_X1 U8970 ( .A1(n7272), .A2(n7271), .ZN(n9961) );
  XNOR2_X1 U8971 ( .A(n7325), .B(n7323), .ZN(n10002) );
  OAI21_X1 U8972 ( .B1(n7323), .B2(n7276), .A(n7275), .ZN(n7279) );
  INV_X1 U8973 ( .A(n7277), .ZN(n7278) );
  AOI21_X1 U8974 ( .B1(n7279), .B2(n9947), .A(n7278), .ZN(n10001) );
  INV_X1 U8975 ( .A(n10001), .ZN(n7289) );
  INV_X1 U8976 ( .A(n7280), .ZN(n7281) );
  NAND2_X1 U8977 ( .A1(n9974), .A2(n4447), .ZN(n7282) );
  NAND2_X1 U8978 ( .A1(n7282), .A2(n9975), .ZN(n7283) );
  NOR2_X1 U8979 ( .A1(n9955), .A2(n7283), .ZN(n9998) );
  OR2_X1 U8980 ( .A1(n7284), .A2(n6376), .ZN(n9585) );
  INV_X1 U8981 ( .A(n9585), .ZN(n9978) );
  INV_X1 U8982 ( .A(n9949), .ZN(n9967) );
  AOI22_X1 U8983 ( .A1(n9998), .A2(n9978), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9967), .ZN(n7286) );
  NAND2_X1 U8984 ( .A1(n9968), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7285) );
  OAI211_X1 U8985 ( .C1(n7287), .C2(n9970), .A(n7286), .B(n7285), .ZN(n7288)
         );
  AOI21_X1 U8986 ( .B1(n7289), .B2(n9588), .A(n7288), .ZN(n7290) );
  OAI21_X1 U8987 ( .B1(n9623), .B2(n10002), .A(n7290), .ZN(P1_U3291) );
  INV_X1 U8988 ( .A(n8846), .ZN(n7291) );
  NAND2_X1 U8989 ( .A1(n7292), .A2(n7291), .ZN(n7296) );
  NAND4_X1 U8990 ( .A1(n7296), .A2(n7295), .A3(n7294), .A4(n7293), .ZN(n7300)
         );
  OR2_X1 U8991 ( .A1(n7300), .A2(n8608), .ZN(n8714) );
  INV_X1 U8992 ( .A(n8712), .ZN(n8671) );
  NAND2_X1 U8993 ( .A1(n6849), .A2(n8694), .ZN(n8786) );
  INV_X1 U8994 ( .A(n8786), .ZN(n7299) );
  NOR3_X1 U8995 ( .A1(n8783), .A2(n10308), .A3(n7297), .ZN(n7298) );
  AOI211_X1 U8996 ( .C1(n8671), .C2(P2_REG3_REG_0__SCAN_IN), .A(n7299), .B(
        n7298), .ZN(n7301) );
  MUX2_X1 U8997 ( .A(n7302), .B(n7301), .S(n8700), .Z(n7303) );
  OAI21_X1 U8998 ( .B1(n8714), .B2(n8784), .A(n7303), .ZN(P2_U3233) );
  OAI21_X1 U8999 ( .B1(n7306), .B2(n7305), .A(n7304), .ZN(n7307) );
  NAND2_X1 U9000 ( .A1(n7307), .A2(n8968), .ZN(n7312) );
  INV_X1 U9001 ( .A(n7349), .ZN(n7310) );
  INV_X1 U9002 ( .A(n9796), .ZN(n8925) );
  AOI22_X1 U9003 ( .A1(n7362), .A2(n8948), .B1(n8924), .B2(n9004), .ZN(n7345)
         );
  INV_X1 U9004 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7308) );
  OAI22_X1 U9005 ( .A1(n7345), .A2(n8927), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7308), .ZN(n7309) );
  AOI21_X1 U9006 ( .B1(n7310), .B2(n8925), .A(n7309), .ZN(n7311) );
  OAI211_X1 U9007 ( .C1(n10028), .C2(n9786), .A(n7312), .B(n7311), .ZN(
        P1_U3239) );
  AOI21_X1 U9008 ( .B1(n9978), .B2(n9975), .A(n9599), .ZN(n7322) );
  INV_X1 U9009 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7318) );
  NAND3_X1 U9010 ( .A1(n7315), .A2(n7314), .A3(n7313), .ZN(n7317) );
  OAI211_X1 U9011 ( .C1(n9949), .C2(n7318), .A(n7317), .B(n7316), .ZN(n7320)
         );
  NOR2_X1 U9012 ( .A1(n9588), .A2(n6083), .ZN(n7319) );
  AOI21_X1 U9013 ( .B1(n9588), .B2(n7320), .A(n7319), .ZN(n7321) );
  OAI21_X1 U9014 ( .B1(n7322), .B2(n9976), .A(n7321), .ZN(P1_U3293) );
  INV_X1 U9015 ( .A(n7323), .ZN(n7324) );
  OR2_X1 U9016 ( .A1(n9007), .A2(n4447), .ZN(n7326) );
  NAND2_X1 U9017 ( .A1(n9953), .A2(n9954), .ZN(n7329) );
  NAND2_X1 U9018 ( .A1(n7327), .A2(n10007), .ZN(n7328) );
  NAND2_X1 U9019 ( .A1(n7329), .A2(n7328), .ZN(n7356) );
  XNOR2_X1 U9020 ( .A(n7356), .B(n7330), .ZN(n10017) );
  INV_X1 U9021 ( .A(n7330), .ZN(n7355) );
  XNOR2_X1 U9022 ( .A(n9928), .B(n7355), .ZN(n7332) );
  AOI21_X1 U9023 ( .B1(n7332), .B2(n9947), .A(n7331), .ZN(n10015) );
  MUX2_X1 U9024 ( .A(n10015), .B(n7333), .S(n9968), .Z(n7339) );
  INV_X1 U9025 ( .A(n7335), .ZN(n9940) );
  AOI211_X1 U9026 ( .C1(n10014), .C2(n7334), .A(n9612), .B(n9940), .ZN(n10013)
         );
  OAI22_X1 U9027 ( .A1(n9970), .A2(n7357), .B1(n9949), .B2(n7336), .ZN(n7337)
         );
  AOI21_X1 U9028 ( .B1(n10013), .B2(n9978), .A(n7337), .ZN(n7338) );
  OAI211_X1 U9029 ( .C1(n10017), .C2(n9623), .A(n7339), .B(n7338), .ZN(
        P1_U3289) );
  INV_X1 U9030 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7341) );
  INV_X1 U9031 ( .A(n7340), .ZN(n7343) );
  INV_X1 U9032 ( .A(n9905), .ZN(n9066) );
  OAI222_X1 U9033 ( .A1(n8277), .A2(n7341), .B1(n8275), .B2(n7343), .C1(n8274), 
        .C2(n9066), .ZN(P1_U3340) );
  INV_X1 U9034 ( .A(n10198), .ZN(n8510) );
  INV_X1 U9035 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7342) );
  OAI222_X1 U9036 ( .A1(n8510), .A2(P2_U3151), .B1(n8851), .B2(n7343), .C1(
        n7342), .C2(n8848), .ZN(P2_U3280) );
  INV_X1 U9037 ( .A(n9947), .ZN(n9963) );
  AOI21_X1 U9038 ( .B1(n7344), .B2(n7404), .A(n9963), .ZN(n7348) );
  INV_X1 U9039 ( .A(n7345), .ZN(n7346) );
  AOI21_X1 U9040 ( .B1(n7348), .B2(n7347), .A(n7346), .ZN(n10027) );
  INV_X1 U9041 ( .A(n9968), .ZN(n9588) );
  INV_X1 U9042 ( .A(n9588), .ZN(n9973) );
  OAI22_X1 U9043 ( .A1(n9588), .A2(n7350), .B1(n7349), .B2(n9949), .ZN(n7354)
         );
  NAND2_X1 U9044 ( .A1(n9939), .A2(n7407), .ZN(n7351) );
  NAND2_X1 U9045 ( .A1(n7351), .A2(n9975), .ZN(n7352) );
  OR2_X1 U9046 ( .A1(n7352), .A2(n7521), .ZN(n10026) );
  NOR2_X1 U9047 ( .A1(n10026), .A2(n9585), .ZN(n7353) );
  AOI211_X1 U9048 ( .C1(n9599), .C2(n7407), .A(n7354), .B(n7353), .ZN(n7366)
         );
  NAND2_X1 U9049 ( .A1(n7356), .A2(n7355), .ZN(n7360) );
  NAND2_X1 U9050 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  NAND2_X1 U9051 ( .A1(n7360), .A2(n7359), .ZN(n9937) );
  INV_X1 U9052 ( .A(n9929), .ZN(n9938) );
  NAND2_X1 U9053 ( .A1(n9937), .A2(n9938), .ZN(n7364) );
  OR2_X1 U9054 ( .A1(n7362), .A2(n7361), .ZN(n7363) );
  NAND2_X1 U9055 ( .A1(n7364), .A2(n7363), .ZN(n7405) );
  XNOR2_X1 U9056 ( .A(n7405), .B(n7404), .ZN(n10030) );
  NAND2_X1 U9057 ( .A1(n10030), .A2(n9957), .ZN(n7365) );
  OAI211_X1 U9058 ( .C1(n10027), .C2(n9973), .A(n7366), .B(n7365), .ZN(
        P1_U3287) );
  NAND2_X1 U9059 ( .A1(n7385), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7367) );
  NAND2_X1 U9060 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  MUX2_X1 U9061 ( .A(n7374), .B(P2_REG1_REG_6__SCAN_IN), .S(n7391), .Z(n10141)
         );
  INV_X1 U9062 ( .A(n7396), .ZN(n7655) );
  XNOR2_X1 U9063 ( .A(n7654), .B(n7655), .ZN(n7657) );
  XNOR2_X1 U9064 ( .A(n7657), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7402) );
  INV_X1 U9065 ( .A(n10241), .ZN(n10153) );
  AOI21_X1 U9066 ( .B1(n7371), .B2(n7385), .A(n7370), .ZN(n10135) );
  MUX2_X1 U9067 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n7642), .Z(n7372) );
  XNOR2_X1 U9068 ( .A(n7372), .B(n7389), .ZN(n10136) );
  INV_X1 U9069 ( .A(n7372), .ZN(n7373) );
  INV_X1 U9070 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7684) );
  MUX2_X1 U9071 ( .A(n7684), .B(n7374), .S(n7642), .Z(n7375) );
  INV_X1 U9072 ( .A(n7391), .ZN(n10151) );
  NAND2_X1 U9073 ( .A1(n7375), .A2(n10151), .ZN(n7376) );
  OAI21_X1 U9074 ( .B1(n7375), .B2(n10151), .A(n7376), .ZN(n10157) );
  INV_X1 U9075 ( .A(n7376), .ZN(n7382) );
  MUX2_X1 U9076 ( .A(n7377), .B(n7656), .S(n7642), .Z(n7378) );
  NAND2_X1 U9077 ( .A1(n7378), .A2(n7655), .ZN(n8440) );
  INV_X1 U9078 ( .A(n7378), .ZN(n7379) );
  NAND2_X1 U9079 ( .A1(n7379), .A2(n7396), .ZN(n7380) );
  AND2_X1 U9080 ( .A1(n8440), .A2(n7380), .ZN(n7381) );
  INV_X1 U9081 ( .A(n8441), .ZN(n7384) );
  NOR3_X1 U9082 ( .A1(n10156), .A2(n7382), .A3(n7381), .ZN(n7383) );
  OAI21_X1 U9083 ( .B1(n7384), .B2(n7383), .A(n10240), .ZN(n7401) );
  NAND2_X1 U9084 ( .A1(n7385), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7386) );
  NAND2_X1 U9085 ( .A1(n7387), .A2(n7386), .ZN(n7390) );
  INV_X1 U9086 ( .A(n7390), .ZN(n7388) );
  XNOR2_X1 U9087 ( .A(n7391), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n10145) );
  OAI21_X1 U9088 ( .B1(n7393), .B2(P2_REG2_REG_7__SCAN_IN), .A(n8453), .ZN(
        n7399) );
  INV_X1 U9089 ( .A(n10246), .ZN(n10175) );
  INV_X1 U9090 ( .A(n10163), .ZN(n10231) );
  INV_X1 U9091 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n7394) );
  NOR2_X1 U9092 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7394), .ZN(n7789) );
  AOI21_X1 U9093 ( .B1(n10231), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7789), .ZN(
        n7395) );
  OAI21_X1 U9094 ( .B1(n7397), .B2(n7396), .A(n7395), .ZN(n7398) );
  AOI21_X1 U9095 ( .B1(n7399), .B2(n10175), .A(n7398), .ZN(n7400) );
  OAI211_X1 U9096 ( .C1(n7402), .C2(n10153), .A(n7401), .B(n7400), .ZN(
        P2_U3189) );
  NAND2_X1 U9097 ( .A1(n9008), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7403) );
  OAI21_X1 U9098 ( .B1(n9167), .B2(n9008), .A(n7403), .ZN(P1_U3582) );
  NAND2_X1 U9099 ( .A1(n7405), .A2(n7404), .ZN(n7409) );
  INV_X1 U9100 ( .A(n7475), .ZN(n7406) );
  OR2_X1 U9101 ( .A1(n7407), .A2(n7406), .ZN(n7408) );
  NAND2_X1 U9102 ( .A1(n7409), .A2(n7408), .ZN(n7518) );
  INV_X1 U9103 ( .A(n7410), .ZN(n7519) );
  NAND2_X1 U9104 ( .A1(n7518), .A2(n7519), .ZN(n7413) );
  NAND2_X1 U9105 ( .A1(n10031), .A2(n7411), .ZN(n7412) );
  NAND2_X1 U9106 ( .A1(n7413), .A2(n7412), .ZN(n7464) );
  INV_X1 U9107 ( .A(n7449), .ZN(n7415) );
  OR2_X1 U9108 ( .A1(n7415), .A2(n7414), .ZN(n7463) );
  XNOR2_X1 U9109 ( .A(n7464), .B(n7463), .ZN(n10041) );
  INV_X1 U9110 ( .A(n10041), .ZN(n7429) );
  INV_X1 U9111 ( .A(n7463), .ZN(n7416) );
  XNOR2_X1 U9112 ( .A(n7417), .B(n7416), .ZN(n7418) );
  NAND2_X1 U9113 ( .A1(n7418), .A2(n9947), .ZN(n7422) );
  OR2_X1 U9114 ( .A1(n7544), .A2(n8972), .ZN(n7420) );
  NAND2_X1 U9115 ( .A1(n9004), .A2(n8948), .ZN(n7419) );
  NAND2_X1 U9116 ( .A1(n7420), .A2(n7419), .ZN(n9789) );
  INV_X1 U9117 ( .A(n9789), .ZN(n7421) );
  NAND2_X1 U9118 ( .A1(n7422), .A2(n7421), .ZN(n10046) );
  NAND2_X1 U9119 ( .A1(n10046), .A2(n9588), .ZN(n7428) );
  OAI22_X1 U9120 ( .A1(n9588), .A2(n7423), .B1(n9795), .B2(n9949), .ZN(n7426)
         );
  AOI21_X1 U9121 ( .B1(n7520), .B2(n7466), .A(n9612), .ZN(n7424) );
  NAND2_X1 U9122 ( .A1(n7424), .A2(n7454), .ZN(n10039) );
  NOR2_X1 U9123 ( .A1(n10039), .A2(n9585), .ZN(n7425) );
  AOI211_X1 U9124 ( .C1(n9599), .C2(n7466), .A(n7426), .B(n7425), .ZN(n7427)
         );
  OAI211_X1 U9125 ( .C1(n7429), .C2(n9623), .A(n7428), .B(n7427), .ZN(P1_U3285) );
  XNOR2_X1 U9126 ( .A(n9062), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U9127 ( .A1(n9712), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7430) );
  OAI21_X1 U9128 ( .B1(n9712), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7430), .ZN(
        n9709) );
  OAI21_X1 U9129 ( .B1(n7434), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7431), .ZN(
        n9708) );
  NOR2_X1 U9130 ( .A1(n9709), .A2(n9708), .ZN(n9707) );
  AOI22_X1 U9131 ( .A1(n9862), .A2(n6038), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n7432), .ZN(n9864) );
  XNOR2_X1 U9132 ( .A(n9064), .B(n9061), .ZN(n7448) );
  INV_X1 U9133 ( .A(n9913), .ZN(n9900) );
  OR2_X1 U9134 ( .A1(n9712), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7433) );
  NAND2_X1 U9135 ( .A1(n9712), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7437) );
  NAND2_X1 U9136 ( .A1(n7433), .A2(n7437), .ZN(n9705) );
  OR2_X1 U9137 ( .A1(n7434), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7435) );
  NAND2_X1 U9138 ( .A1(n7436), .A2(n7435), .ZN(n9706) );
  MUX2_X1 U9139 ( .A(n7438), .B(P1_REG1_REG_11__SCAN_IN), .S(n9862), .Z(n9856)
         );
  NOR2_X1 U9140 ( .A1(n9857), .A2(n9856), .ZN(n9858) );
  AOI21_X1 U9141 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9862), .A(n9858), .ZN(
        n7441) );
  MUX2_X1 U9142 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7439), .S(n9062), .Z(n7440)
         );
  NAND2_X1 U9143 ( .A1(n7440), .A2(n7441), .ZN(n9048) );
  OAI21_X1 U9144 ( .B1(n7441), .B2(n7440), .A(n9048), .ZN(n7446) );
  INV_X1 U9145 ( .A(n9062), .ZN(n7444) );
  NOR2_X1 U9146 ( .A1(n7442), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7985) );
  AOI21_X1 U9147 ( .B1(n9811), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7985), .ZN(
        n7443) );
  OAI21_X1 U9148 ( .B1(n7444), .B2(n9821), .A(n7443), .ZN(n7445) );
  AOI21_X1 U9149 ( .B1(n9861), .B2(n7446), .A(n7445), .ZN(n7447) );
  OAI21_X1 U9150 ( .B1(n7448), .B2(n9900), .A(n7447), .ZN(P1_U3255) );
  NAND2_X1 U9151 ( .A1(n4526), .A2(n7449), .ZN(n7452) );
  NAND2_X1 U9152 ( .A1(n7451), .A2(n7450), .ZN(n7542) );
  XNOR2_X1 U9153 ( .A(n7452), .B(n7542), .ZN(n7453) );
  NOR2_X1 U9154 ( .A1(n7476), .A2(n9140), .ZN(n7778) );
  AOI21_X1 U9155 ( .B1(n7453), .B2(n9947), .A(n7778), .ZN(n10054) );
  NAND2_X1 U9156 ( .A1(n7454), .A2(n10048), .ZN(n7455) );
  NAND2_X1 U9157 ( .A1(n7455), .A2(n9975), .ZN(n7456) );
  OR2_X1 U9158 ( .A1(n7456), .A2(n7539), .ZN(n7458) );
  NOR2_X1 U9159 ( .A1(n7565), .A2(n8972), .ZN(n7779) );
  INV_X1 U9160 ( .A(n7779), .ZN(n7457) );
  NAND2_X1 U9161 ( .A1(n7458), .A2(n7457), .ZN(n10050) );
  INV_X1 U9162 ( .A(n10048), .ZN(n7459) );
  NOR2_X1 U9163 ( .A1(n7459), .A2(n9970), .ZN(n7462) );
  OAI22_X1 U9164 ( .A1(n9588), .A2(n7460), .B1(n7782), .B2(n9949), .ZN(n7461)
         );
  AOI211_X1 U9165 ( .C1(n10050), .C2(n9978), .A(n7462), .B(n7461), .ZN(n7470)
         );
  NAND2_X1 U9166 ( .A1(n7464), .A2(n7463), .ZN(n7468) );
  INV_X1 U9167 ( .A(n7476), .ZN(n7465) );
  OR2_X1 U9168 ( .A1(n7466), .A2(n7465), .ZN(n7467) );
  NAND2_X1 U9169 ( .A1(n7468), .A2(n7467), .ZN(n7543) );
  XNOR2_X1 U9170 ( .A(n7543), .B(n7542), .ZN(n10051) );
  NAND2_X1 U9171 ( .A1(n10051), .A2(n9957), .ZN(n7469) );
  OAI211_X1 U9172 ( .C1(n10054), .C2(n9973), .A(n7470), .B(n7469), .ZN(
        P1_U3284) );
  XNOR2_X1 U9173 ( .A(n7473), .B(n7472), .ZN(n7474) );
  XNOR2_X1 U9174 ( .A(n7471), .B(n7474), .ZN(n7482) );
  NOR2_X1 U9175 ( .A1(n10031), .A2(n9786), .ZN(n7481) );
  OR2_X1 U9176 ( .A1(n7475), .A2(n9140), .ZN(n7478) );
  OR2_X1 U9177 ( .A1(n7476), .A2(n8972), .ZN(n7477) );
  NAND2_X1 U9178 ( .A1(n7478), .A2(n7477), .ZN(n7516) );
  AOI22_X1 U9179 ( .A1(n4438), .A2(n7516), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7479) );
  OAI21_X1 U9180 ( .B1(n9796), .B2(n7522), .A(n7479), .ZN(n7480) );
  AOI211_X1 U9181 ( .C1(n7482), .C2(n8968), .A(n7481), .B(n7480), .ZN(n7483)
         );
  INV_X1 U9182 ( .A(n7483), .ZN(P1_U3213) );
  AOI21_X1 U9183 ( .B1(n7485), .B2(n7484), .A(n4524), .ZN(n7492) );
  INV_X1 U9184 ( .A(n7486), .ZN(n7626) );
  NOR2_X1 U9185 ( .A1(n8412), .A2(n7622), .ZN(n7487) );
  AOI211_X1 U9186 ( .C1(n8410), .C2(n8436), .A(n7488), .B(n7487), .ZN(n7489)
         );
  OAI21_X1 U9187 ( .B1(n5632), .B2(n8419), .A(n7489), .ZN(n7490) );
  AOI21_X1 U9188 ( .B1(n7626), .B2(n8415), .A(n7490), .ZN(n7491) );
  OAI21_X1 U9189 ( .B1(n7492), .B2(n8403), .A(n7491), .ZN(P2_U3170) );
  NAND2_X1 U9190 ( .A1(n7493), .A2(P2_U3893), .ZN(n7494) );
  OAI21_X1 U9191 ( .B1(P2_U3893), .B2(n5827), .A(n7494), .ZN(P2_U3518) );
  INV_X1 U9192 ( .A(n10214), .ZN(n8498) );
  INV_X1 U9193 ( .A(n7495), .ZN(n7497) );
  INV_X1 U9194 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7496) );
  OAI222_X1 U9195 ( .A1(n8498), .A2(P2_U3151), .B1(n8851), .B2(n7497), .C1(
        n7496), .C2(n8848), .ZN(P2_U3279) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7498) );
  INV_X1 U9197 ( .A(n9084), .ZN(n9059) );
  OAI222_X1 U9198 ( .A1(n8277), .A2(n7498), .B1(n8275), .B2(n7497), .C1(n8274), 
        .C2(n9059), .ZN(P1_U3339) );
  AND2_X1 U9199 ( .A1(n7500), .A2(n7499), .ZN(n7574) );
  OR2_X1 U9200 ( .A1(n7944), .A2(n7574), .ZN(n7501) );
  NAND2_X1 U9201 ( .A1(n8700), .A2(n7501), .ZN(n8674) );
  INV_X1 U9202 ( .A(n8674), .ZN(n8727) );
  XNOR2_X1 U9203 ( .A(n7502), .B(n7505), .ZN(n10252) );
  OAI22_X1 U9204 ( .A1(n8714), .A2(n6848), .B1(n7503), .B2(n8712), .ZN(n7511)
         );
  OR2_X1 U9205 ( .A1(n8784), .A2(n8635), .ZN(n7504) );
  OAI21_X1 U9206 ( .B1(n7505), .B2(n7504), .A(n8718), .ZN(n7506) );
  NAND2_X1 U9207 ( .A1(n7506), .A2(n5625), .ZN(n7508) );
  NAND2_X1 U9208 ( .A1(n8438), .A2(n8694), .ZN(n7507) );
  OAI211_X1 U9209 ( .C1(n8635), .C2(n7509), .A(n7508), .B(n7507), .ZN(n10253)
         );
  MUX2_X1 U9210 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10253), .S(n8700), .Z(n7510)
         );
  AOI211_X1 U9211 ( .C1(n8727), .C2(n10252), .A(n7511), .B(n7510), .ZN(n7512)
         );
  INV_X1 U9212 ( .A(n7512), .ZN(P2_U3232) );
  NAND2_X1 U9213 ( .A1(n8492), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7513) );
  OAI21_X1 U9214 ( .B1(n7514), .B2(n8492), .A(n7513), .ZN(P2_U3521) );
  XNOR2_X1 U9215 ( .A(n7515), .B(n7519), .ZN(n7517) );
  AOI21_X1 U9216 ( .B1(n7517), .B2(n9947), .A(n7516), .ZN(n10037) );
  XNOR2_X1 U9217 ( .A(n7518), .B(n7519), .ZN(n10034) );
  OAI211_X1 U9218 ( .C1(n7521), .C2(n10031), .A(n9975), .B(n7520), .ZN(n10033)
         );
  OAI22_X1 U9219 ( .A1(n9588), .A2(n4661), .B1(n7522), .B2(n9949), .ZN(n7523)
         );
  AOI21_X1 U9220 ( .B1(n9599), .B2(n7524), .A(n7523), .ZN(n7525) );
  OAI21_X1 U9221 ( .B1(n10033), .B2(n9585), .A(n7525), .ZN(n7526) );
  AOI21_X1 U9222 ( .B1(n10034), .B2(n9957), .A(n7526), .ZN(n7527) );
  OAI21_X1 U9223 ( .B1(n10037), .B2(n9973), .A(n7527), .ZN(P1_U3286) );
  INV_X1 U9224 ( .A(n7528), .ZN(n7531) );
  INV_X1 U9225 ( .A(n9100), .ZN(n9089) );
  OAI222_X1 U9226 ( .A1(n8277), .A2(n7529), .B1(n8275), .B2(n7531), .C1(
        P1_U3086), .C2(n9089), .ZN(P1_U3338) );
  INV_X1 U9227 ( .A(n10233), .ZN(n8513) );
  OAI222_X1 U9228 ( .A1(n8513), .A2(P2_U3151), .B1(n8851), .B2(n7531), .C1(
        n7530), .C2(n8848), .ZN(P2_U3278) );
  OAI21_X1 U9229 ( .B1(n7547), .B2(n7533), .A(n7532), .ZN(n7536) );
  OR2_X1 U9230 ( .A1(n7544), .A2(n9140), .ZN(n7535) );
  OR2_X1 U9231 ( .A1(n7709), .A2(n8972), .ZN(n7534) );
  NAND2_X1 U9232 ( .A1(n7535), .A2(n7534), .ZN(n7957) );
  AOI21_X1 U9233 ( .B1(n7536), .B2(n9947), .A(n7957), .ZN(n10057) );
  OAI22_X1 U9234 ( .A1(n9588), .A2(n7537), .B1(n7959), .B2(n9949), .ZN(n7541)
         );
  INV_X1 U9235 ( .A(n7568), .ZN(n7538) );
  OAI211_X1 U9236 ( .C1(n10058), .C2(n7539), .A(n7538), .B(n9975), .ZN(n10056)
         );
  NOR2_X1 U9237 ( .A1(n10056), .A2(n9585), .ZN(n7540) );
  AOI211_X1 U9238 ( .C1(n9599), .C2(n7961), .A(n7541), .B(n7540), .ZN(n7549)
         );
  NAND2_X1 U9239 ( .A1(n7543), .A2(n7542), .ZN(n7546) );
  OR2_X1 U9240 ( .A1(n10048), .A2(n4828), .ZN(n7545) );
  NAND2_X1 U9241 ( .A1(n7546), .A2(n7545), .ZN(n7564) );
  INV_X1 U9242 ( .A(n7547), .ZN(n7563) );
  XNOR2_X1 U9243 ( .A(n7564), .B(n7563), .ZN(n10060) );
  NAND2_X1 U9244 ( .A1(n10060), .A2(n9957), .ZN(n7548) );
  OAI211_X1 U9245 ( .C1(n9968), .C2(n10057), .A(n7549), .B(n7548), .ZN(
        P1_U3283) );
  NAND2_X1 U9246 ( .A1(n7550), .A2(n7551), .ZN(n7552) );
  XOR2_X1 U9247 ( .A(n7554), .B(n7552), .Z(n7553) );
  AOI222_X1 U9248 ( .A1(n8781), .A2(n7553), .B1(n8437), .B2(n8694), .C1(n8438), 
        .C2(n8695), .ZN(n10263) );
  XNOR2_X1 U9249 ( .A(n7555), .B(n7554), .ZN(n10261) );
  NOR2_X1 U9250 ( .A1(n8700), .A2(n5074), .ZN(n7557) );
  OAI22_X1 U9251 ( .A1(n8714), .A2(n6846), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n8712), .ZN(n7556) );
  AOI211_X1 U9252 ( .C1(n10261), .C2(n8727), .A(n7557), .B(n7556), .ZN(n7558)
         );
  OAI21_X1 U9253 ( .B1(n10263), .B2(n8708), .A(n7558), .ZN(P2_U3230) );
  AOI21_X1 U9254 ( .B1(n7559), .B2(n7713), .A(n9963), .ZN(n7562) );
  OR2_X1 U9255 ( .A1(n7565), .A2(n9140), .ZN(n7560) );
  OAI21_X1 U9256 ( .B1(n7808), .B2(n8972), .A(n7560), .ZN(n8091) );
  AOI21_X1 U9257 ( .B1(n7562), .B2(n7561), .A(n8091), .ZN(n10063) );
  INV_X1 U9258 ( .A(n7565), .ZN(n9003) );
  OR2_X1 U9259 ( .A1(n7961), .A2(n9003), .ZN(n7566) );
  XNOR2_X1 U9260 ( .A(n7714), .B(n7713), .ZN(n10066) );
  NAND2_X1 U9261 ( .A1(n10066), .A2(n9957), .ZN(n7572) );
  OAI22_X1 U9262 ( .A1(n9588), .A2(n6038), .B1(n8093), .B2(n9949), .ZN(n7570)
         );
  OAI211_X1 U9263 ( .C1(n7568), .C2(n10064), .A(n9975), .B(n7567), .ZN(n10062)
         );
  NOR2_X1 U9264 ( .A1(n10062), .A2(n9585), .ZN(n7569) );
  AOI211_X1 U9265 ( .C1(n9599), .C2(n8095), .A(n7570), .B(n7569), .ZN(n7571)
         );
  OAI211_X1 U9266 ( .C1(n9968), .C2(n10063), .A(n7572), .B(n7571), .ZN(
        P1_U3282) );
  XNOR2_X1 U9267 ( .A(n7573), .B(n7576), .ZN(n10257) );
  NAND2_X1 U9268 ( .A1(n8700), .A2(n7574), .ZN(n8557) );
  INV_X1 U9269 ( .A(n7944), .ZN(n8251) );
  OAI21_X1 U9270 ( .B1(n7576), .B2(n7575), .A(n7550), .ZN(n7578) );
  OAI22_X1 U9271 ( .A1(n5051), .A2(n8718), .B1(n7622), .B2(n8720), .ZN(n7577)
         );
  AOI21_X1 U9272 ( .B1(n7578), .B2(n8781), .A(n7577), .ZN(n7579) );
  OAI21_X1 U9273 ( .B1(n10257), .B2(n8251), .A(n7579), .ZN(n10259) );
  OAI22_X1 U9274 ( .A1(n10256), .A2(n8608), .B1(n5054), .B2(n8712), .ZN(n7580)
         );
  NOR2_X1 U9275 ( .A1(n10259), .A2(n7580), .ZN(n7581) );
  MUX2_X1 U9276 ( .A(n7582), .B(n7581), .S(n8700), .Z(n7583) );
  OAI21_X1 U9277 ( .B1(n10257), .B2(n8557), .A(n7583), .ZN(P2_U3231) );
  INV_X1 U9278 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10335) );
  NOR2_X1 U9279 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(P2_ADDR_REG_17__SCAN_IN), 
        .ZN(n7584) );
  AOI21_X1 U9280 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n7584), .ZN(n10339) );
  NOR2_X1 U9281 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7585) );
  AOI21_X1 U9282 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7585), .ZN(n10342) );
  NOR2_X1 U9283 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7586) );
  AOI21_X1 U9284 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7586), .ZN(n10345) );
  NOR2_X1 U9285 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .ZN(n7587) );
  AOI21_X1 U9286 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n7587), .ZN(n10348) );
  NOR2_X1 U9287 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7588) );
  AOI21_X1 U9288 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n7588), .ZN(n10351) );
  NOR2_X1 U9289 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7589) );
  AOI21_X1 U9290 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7589), .ZN(n10354) );
  NOR2_X1 U9291 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7590) );
  AOI21_X1 U9292 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7590), .ZN(n10357) );
  NOR2_X1 U9293 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7591) );
  AOI21_X1 U9294 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7591), .ZN(n10360) );
  INV_X1 U9295 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7698) );
  INV_X1 U9296 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7592) );
  AOI22_X1 U9297 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P2_ADDR_REG_9__SCAN_IN), 
        .B1(n7698), .B2(n7592), .ZN(n10366) );
  NOR2_X1 U9298 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7593) );
  AOI21_X1 U9299 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7593), .ZN(n10375) );
  NOR2_X1 U9300 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7594) );
  AOI21_X1 U9301 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7594), .ZN(n10372) );
  NOR2_X1 U9302 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7595) );
  AOI21_X1 U9303 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7595), .ZN(n10369) );
  NOR2_X1 U9304 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7596) );
  AOI21_X1 U9305 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7596), .ZN(n10363) );
  INV_X1 U9306 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U9307 ( .A1(n10332), .A2(n7185), .ZN(n10331) );
  NOR2_X1 U9308 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10331), .ZN(n10327) );
  INV_X1 U9309 ( .A(n10327), .ZN(n10328) );
  INV_X1 U9310 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10330) );
  NAND3_X1 U9311 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U9312 ( .A1(n10330), .A2(n10329), .ZN(n10326) );
  NAND2_X1 U9313 ( .A1(n10328), .A2(n10326), .ZN(n10378) );
  NAND2_X1 U9314 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7597) );
  OAI21_X1 U9315 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7597), .ZN(n10377) );
  NOR2_X1 U9316 ( .A1(n10378), .A2(n10377), .ZN(n10376) );
  AOI21_X1 U9317 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10376), .ZN(n10381) );
  NAND2_X1 U9318 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7598) );
  OAI21_X1 U9319 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7598), .ZN(n10380) );
  NOR2_X1 U9320 ( .A1(n10381), .A2(n10380), .ZN(n10379) );
  AOI21_X1 U9321 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10379), .ZN(n10384) );
  NOR2_X1 U9322 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7599) );
  AOI21_X1 U9323 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7599), .ZN(n10383) );
  NAND2_X1 U9324 ( .A1(n10384), .A2(n10383), .ZN(n10382) );
  OAI21_X1 U9325 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10382), .ZN(n10362) );
  NAND2_X1 U9326 ( .A1(n10363), .A2(n10362), .ZN(n10361) );
  OAI21_X1 U9327 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10361), .ZN(n10368) );
  NAND2_X1 U9328 ( .A1(n10369), .A2(n10368), .ZN(n10367) );
  OAI21_X1 U9329 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10367), .ZN(n10371) );
  NAND2_X1 U9330 ( .A1(n10372), .A2(n10371), .ZN(n10370) );
  OAI21_X1 U9331 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10370), .ZN(n10374) );
  NAND2_X1 U9332 ( .A1(n10375), .A2(n10374), .ZN(n10373) );
  OAI21_X1 U9333 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10373), .ZN(n10365) );
  NAND2_X1 U9334 ( .A1(n10366), .A2(n10365), .ZN(n10364) );
  OAI21_X1 U9335 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n10364), .ZN(n10359) );
  NAND2_X1 U9336 ( .A1(n10360), .A2(n10359), .ZN(n10358) );
  OAI21_X1 U9337 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10358), .ZN(n10356) );
  NAND2_X1 U9338 ( .A1(n10357), .A2(n10356), .ZN(n10355) );
  OAI21_X1 U9339 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10355), .ZN(n10353) );
  NAND2_X1 U9340 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  OAI21_X1 U9341 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10352), .ZN(n10350) );
  NAND2_X1 U9342 ( .A1(n10351), .A2(n10350), .ZN(n10349) );
  OAI21_X1 U9343 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10349), .ZN(n10347) );
  NAND2_X1 U9344 ( .A1(n10348), .A2(n10347), .ZN(n10346) );
  OAI21_X1 U9345 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10346), .ZN(n10344) );
  NAND2_X1 U9346 ( .A1(n10345), .A2(n10344), .ZN(n10343) );
  OAI21_X1 U9347 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10343), .ZN(n10341) );
  NAND2_X1 U9348 ( .A1(n10342), .A2(n10341), .ZN(n10340) );
  OAI21_X1 U9349 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10340), .ZN(n10338) );
  NAND2_X1 U9350 ( .A1(n10339), .A2(n10338), .ZN(n10337) );
  OAI21_X1 U9351 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n10337), .ZN(n10334) );
  NAND2_X1 U9352 ( .A1(n10335), .A2(n10334), .ZN(n7600) );
  NOR2_X1 U9353 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  AOI21_X1 U9354 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7600), .A(n10333), .ZN(
        n7604) );
  NOR2_X1 U9355 ( .A1(n7602), .A2(n7601), .ZN(n7603) );
  XNOR2_X1 U9356 ( .A(n7604), .B(n7603), .ZN(ADD_1068_U4) );
  XOR2_X1 U9357 ( .A(n7606), .B(n7605), .Z(n7614) );
  INV_X1 U9358 ( .A(n7607), .ZN(n7757) );
  OAI22_X1 U9359 ( .A1(n8412), .A2(n7608), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10127), .ZN(n7609) );
  AOI21_X1 U9360 ( .B1(n8410), .B2(n8435), .A(n7609), .ZN(n7610) );
  OAI21_X1 U9361 ( .B1(n7611), .B2(n8419), .A(n7610), .ZN(n7612) );
  AOI21_X1 U9362 ( .B1(n7757), .B2(n8415), .A(n7612), .ZN(n7613) );
  OAI21_X1 U9363 ( .B1(n7614), .B2(n8403), .A(n7613), .ZN(P2_U3167) );
  NAND2_X1 U9364 ( .A1(n7616), .A2(n7615), .ZN(n7748) );
  INV_X1 U9365 ( .A(n7747), .ZN(n7619) );
  XNOR2_X1 U9366 ( .A(n7748), .B(n7619), .ZN(n10265) );
  AND2_X1 U9367 ( .A1(n7618), .A2(n7617), .ZN(n7620) );
  XNOR2_X1 U9368 ( .A(n7620), .B(n7619), .ZN(n7624) );
  NAND2_X1 U9369 ( .A1(n8436), .A2(n8694), .ZN(n7621) );
  OAI21_X1 U9370 ( .B1(n7622), .B2(n8718), .A(n7621), .ZN(n7623) );
  AOI21_X1 U9371 ( .B1(n7624), .B2(n8781), .A(n7623), .ZN(n10269) );
  MUX2_X1 U9372 ( .A(n7625), .B(n10269), .S(n8700), .Z(n7628) );
  AOI22_X1 U9373 ( .A1(n8702), .A2(n10266), .B1(n8671), .B2(n7626), .ZN(n7627)
         );
  OAI211_X1 U9374 ( .C1(n10265), .C2(n8674), .A(n7628), .B(n7627), .ZN(
        P2_U3229) );
  INV_X1 U9375 ( .A(n7629), .ZN(n7672) );
  INV_X1 U9376 ( .A(n8516), .ZN(n8523) );
  OAI222_X1 U9377 ( .A1(n8848), .A2(n7630), .B1(n8851), .B2(n7672), .C1(
        P2_U3151), .C2(n8523), .ZN(P2_U3277) );
  INV_X1 U9378 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7636) );
  MUX2_X1 U9379 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7636), .S(n8447), .Z(n8452)
         );
  AOI21_X1 U9380 ( .B1(n7631), .B2(n7700), .A(n7633), .ZN(n7632) );
  INV_X1 U9381 ( .A(n7632), .ZN(n7692) );
  AOI22_X1 U9382 ( .A1(P2_REG2_REG_10__SCAN_IN), .A2(n7728), .B1(n7735), .B2(
        n7949), .ZN(n7634) );
  AOI21_X1 U9383 ( .B1(n7635), .B2(n7634), .A(n7734), .ZN(n7671) );
  MUX2_X1 U9384 ( .A(n7636), .B(n7658), .S(n7642), .Z(n7637) );
  NAND2_X1 U9385 ( .A1(n7637), .A2(n8447), .ZN(n7641) );
  INV_X1 U9386 ( .A(n7637), .ZN(n7639) );
  NAND2_X1 U9387 ( .A1(n7639), .A2(n7638), .ZN(n7640) );
  NAND2_X1 U9388 ( .A1(n7641), .A2(n7640), .ZN(n8439) );
  INV_X1 U9389 ( .A(n7641), .ZN(n7695) );
  MUX2_X1 U9390 ( .A(n7872), .B(n7643), .S(n7642), .Z(n7644) );
  NAND2_X1 U9391 ( .A1(n7644), .A2(n7700), .ZN(n7652) );
  INV_X1 U9392 ( .A(n7644), .ZN(n7645) );
  NAND2_X1 U9393 ( .A1(n7645), .A2(n7659), .ZN(n7646) );
  AND2_X1 U9394 ( .A1(n7652), .A2(n7646), .ZN(n7694) );
  OAI21_X1 U9395 ( .B1(n8443), .B2(n7695), .A(n7694), .ZN(n7693) );
  MUX2_X1 U9396 ( .A(n7949), .B(n7647), .S(n7642), .Z(n7648) );
  NAND2_X1 U9397 ( .A1(n7648), .A2(n7728), .ZN(n7722) );
  INV_X1 U9398 ( .A(n7648), .ZN(n7649) );
  NAND2_X1 U9399 ( .A1(n7649), .A2(n7735), .ZN(n7650) );
  NAND2_X1 U9400 ( .A1(n7722), .A2(n7650), .ZN(n7651) );
  AND3_X1 U9401 ( .A1(n7693), .A2(n7652), .A3(n7651), .ZN(n7653) );
  OAI21_X1 U9402 ( .B1(n7724), .B2(n7653), .A(n10240), .ZN(n7670) );
  AOI22_X1 U9403 ( .A1(P2_REG1_REG_10__SCAN_IN), .A2(n7735), .B1(n7728), .B2(
        n7647), .ZN(n7663) );
  OAI22_X1 U9404 ( .A1(n7657), .A2(n7656), .B1(n7655), .B2(n7654), .ZN(n8449)
         );
  MUX2_X1 U9405 ( .A(n7658), .B(P2_REG1_REG_8__SCAN_IN), .S(n8447), .Z(n8450)
         );
  NAND2_X1 U9406 ( .A1(n8449), .A2(n8450), .ZN(n8448) );
  NAND2_X1 U9407 ( .A1(n7660), .A2(n7659), .ZN(n7661) );
  NAND2_X1 U9408 ( .A1(n7663), .A2(n7662), .ZN(n7727) );
  OAI21_X1 U9409 ( .B1(n7663), .B2(n7662), .A(n7727), .ZN(n7668) );
  INV_X1 U9410 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7666) );
  NAND2_X1 U9411 ( .A1(n10232), .A2(n7728), .ZN(n7665) );
  AND2_X1 U9412 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8120) );
  INV_X1 U9413 ( .A(n8120), .ZN(n7664) );
  OAI211_X1 U9414 ( .C1(n7666), .C2(n10163), .A(n7665), .B(n7664), .ZN(n7667)
         );
  AOI21_X1 U9415 ( .B1(n7668), .B2(n10241), .A(n7667), .ZN(n7669) );
  OAI211_X1 U9416 ( .C1(n7671), .C2(n10246), .A(n7670), .B(n7669), .ZN(
        P2_U3192) );
  INV_X1 U9417 ( .A(n9920), .ZN(n7673) );
  OAI222_X1 U9418 ( .A1(n8277), .A2(n9404), .B1(n7673), .B2(P1_U3086), .C1(
        n8275), .C2(n7672), .ZN(P1_U3337) );
  NAND2_X1 U9419 ( .A1(n7675), .A2(n7674), .ZN(n7677) );
  XNOR2_X1 U9420 ( .A(n7677), .B(n7676), .ZN(n10277) );
  XNOR2_X1 U9421 ( .A(n7679), .B(n7678), .ZN(n7683) );
  NAND2_X1 U9422 ( .A1(n8436), .A2(n8695), .ZN(n7680) );
  OAI21_X1 U9423 ( .B1(n7681), .B2(n8720), .A(n7680), .ZN(n7682) );
  AOI21_X1 U9424 ( .B1(n7683), .B2(n8781), .A(n7682), .ZN(n10279) );
  MUX2_X1 U9425 ( .A(n7684), .B(n10279), .S(n8700), .Z(n7688) );
  INV_X1 U9426 ( .A(n7685), .ZN(n7769) );
  AOI22_X1 U9427 ( .A1(n8702), .A2(n7686), .B1(n8671), .B2(n7769), .ZN(n7687)
         );
  OAI211_X1 U9428 ( .C1(n10277), .C2(n8674), .A(n7688), .B(n7687), .ZN(
        P2_U3227) );
  OAI21_X1 U9429 ( .B1(n7690), .B2(P2_REG1_REG_9__SCAN_IN), .A(n7689), .ZN(
        n7705) );
  AOI21_X1 U9430 ( .B1(n7692), .B2(n7872), .A(n7691), .ZN(n7703) );
  INV_X1 U9431 ( .A(n7693), .ZN(n7697) );
  NOR3_X1 U9432 ( .A1(n8443), .A2(n7695), .A3(n7694), .ZN(n7696) );
  OAI21_X1 U9433 ( .B1(n7697), .B2(n7696), .A(n10240), .ZN(n7702) );
  NOR2_X1 U9434 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9491), .ZN(n7879) );
  NOR2_X1 U9435 ( .A1(n10163), .A2(n7698), .ZN(n7699) );
  AOI211_X1 U9436 ( .C1(n10232), .C2(n7700), .A(n7879), .B(n7699), .ZN(n7701)
         );
  OAI211_X1 U9437 ( .C1(n7703), .C2(n10246), .A(n7702), .B(n7701), .ZN(n7704)
         );
  AOI21_X1 U9438 ( .B1(n10241), .B2(n7705), .A(n7704), .ZN(n7706) );
  INV_X1 U9439 ( .A(n7706), .ZN(P2_U3191) );
  XNOR2_X1 U9440 ( .A(n7708), .B(n7814), .ZN(n7712) );
  OR2_X1 U9441 ( .A1(n7709), .A2(n9140), .ZN(n7710) );
  OAI21_X1 U9442 ( .B1(n7711), .B2(n8972), .A(n7710), .ZN(n7986) );
  AOI21_X1 U9443 ( .B1(n7712), .B2(n9947), .A(n7986), .ZN(n10069) );
  XNOR2_X1 U9444 ( .A(n7815), .B(n7814), .ZN(n10072) );
  NAND2_X1 U9445 ( .A1(n10072), .A2(n9957), .ZN(n7721) );
  OAI22_X1 U9446 ( .A1(n9588), .A2(n7716), .B1(n7988), .B2(n9949), .ZN(n7719)
         );
  INV_X1 U9447 ( .A(n7567), .ZN(n7717) );
  OAI211_X1 U9448 ( .C1(n7717), .C2(n10070), .A(n9975), .B(n7810), .ZN(n10068)
         );
  NOR2_X1 U9449 ( .A1(n10068), .A2(n9585), .ZN(n7718) );
  AOI211_X1 U9450 ( .C1(n9599), .C2(n7990), .A(n7719), .B(n7718), .ZN(n7720)
         );
  OAI211_X1 U9451 ( .C1(n9968), .C2(n10069), .A(n7721), .B(n7720), .ZN(
        P1_U3281) );
  INV_X1 U9452 ( .A(n7722), .ZN(n7723) );
  NOR2_X1 U9453 ( .A1(n7724), .A2(n7723), .ZN(n7726) );
  MUX2_X1 U9454 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n7642), .Z(n7832) );
  XNOR2_X1 U9455 ( .A(n7832), .B(n7840), .ZN(n7725) );
  NOR2_X1 U9456 ( .A1(n7726), .A2(n7725), .ZN(n7833) );
  AOI21_X1 U9457 ( .B1(n7726), .B2(n7725), .A(n7833), .ZN(n7742) );
  OAI21_X1 U9458 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n7729), .A(n7841), .ZN(
        n7740) );
  INV_X1 U9459 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U9460 ( .A1(n10232), .A2(n7835), .ZN(n7732) );
  INV_X1 U9461 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7730) );
  NOR2_X1 U9462 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7730), .ZN(n8180) );
  INV_X1 U9463 ( .A(n8180), .ZN(n7731) );
  OAI211_X1 U9464 ( .C1(n7733), .C2(n10163), .A(n7732), .B(n7731), .ZN(n7739)
         );
  AOI21_X1 U9465 ( .B1(n5256), .B2(n7736), .A(n7827), .ZN(n7737) );
  NOR2_X1 U9466 ( .A1(n7737), .A2(n10246), .ZN(n7738) );
  AOI211_X1 U9467 ( .C1(n10241), .C2(n7740), .A(n7739), .B(n7738), .ZN(n7741)
         );
  OAI21_X1 U9468 ( .B1(n7742), .B2(n10159), .A(n7741), .ZN(P2_U3193) );
  INV_X1 U9469 ( .A(n7743), .ZN(n7746) );
  OAI222_X1 U9470 ( .A1(n8277), .A2(n7744), .B1(n8275), .B2(n7746), .C1(
        P1_U3086), .C2(n5880), .ZN(P1_U3336) );
  OAI222_X1 U9471 ( .A1(n8526), .A2(P2_U3151), .B1(n8851), .B2(n7746), .C1(
        n7745), .C2(n8848), .ZN(P2_U3276) );
  NAND2_X1 U9472 ( .A1(n7748), .A2(n7747), .ZN(n7750) );
  NAND2_X1 U9473 ( .A1(n7750), .A2(n7749), .ZN(n7751) );
  XNOR2_X1 U9474 ( .A(n7751), .B(n7753), .ZN(n10273) );
  INV_X1 U9475 ( .A(n10273), .ZN(n7760) );
  XNOR2_X1 U9476 ( .A(n7752), .B(n7753), .ZN(n7755) );
  AOI22_X1 U9477 ( .A1(n8437), .A2(n8695), .B1(n8694), .B2(n8435), .ZN(n7754)
         );
  OAI21_X1 U9478 ( .B1(n7755), .B2(n8635), .A(n7754), .ZN(n7756) );
  AOI21_X1 U9479 ( .B1(n7944), .B2(n10273), .A(n7756), .ZN(n10275) );
  MUX2_X1 U9480 ( .A(n4791), .B(n10275), .S(n8700), .Z(n7759) );
  AOI22_X1 U9481 ( .A1(n8702), .A2(n10271), .B1(n8671), .B2(n7757), .ZN(n7758)
         );
  OAI211_X1 U9482 ( .C1(n7760), .C2(n8557), .A(n7759), .B(n7758), .ZN(P2_U3228) );
  INV_X1 U9483 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9361) );
  NOR2_X1 U9484 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9361), .ZN(n10150) );
  NOR2_X1 U9485 ( .A1(n8412), .A2(n7761), .ZN(n7762) );
  AOI211_X1 U9486 ( .C1(n8410), .C2(n8434), .A(n10150), .B(n7762), .ZN(n7763)
         );
  OAI21_X1 U9487 ( .B1(n10276), .B2(n8419), .A(n7763), .ZN(n7768) );
  AOI211_X1 U9488 ( .C1(n7766), .C2(n7765), .A(n8403), .B(n7764), .ZN(n7767)
         );
  AOI211_X1 U9489 ( .C1(n7769), .C2(n8415), .A(n7768), .B(n7767), .ZN(n7770)
         );
  INV_X1 U9490 ( .A(n7770), .ZN(P2_U3179) );
  NAND2_X1 U9491 ( .A1(n7820), .A2(n9697), .ZN(n7772) );
  OAI211_X1 U9492 ( .C1(n7773), .C2(n8277), .A(n7772), .B(n7771), .ZN(P1_U3335) );
  NOR2_X1 U9493 ( .A1(n7776), .A2(n4877), .ZN(n7777) );
  XNOR2_X1 U9494 ( .A(n7774), .B(n7777), .ZN(n7785) );
  OAI21_X1 U9495 ( .B1(n7779), .B2(n7778), .A(n4438), .ZN(n7780) );
  OAI211_X1 U9496 ( .C1(n9796), .C2(n7782), .A(n7781), .B(n7780), .ZN(n7783)
         );
  AOI21_X1 U9497 ( .B1(n10048), .B2(n8988), .A(n7783), .ZN(n7784) );
  OAI21_X1 U9498 ( .B1(n7785), .B2(n9791), .A(n7784), .ZN(P1_U3231) );
  OAI21_X1 U9499 ( .B1(n7788), .B2(n7787), .A(n7786), .ZN(n7794) );
  NOR2_X1 U9500 ( .A1(n8419), .A2(n10281), .ZN(n7793) );
  AOI21_X1 U9501 ( .B1(n8387), .B2(n8435), .A(n7789), .ZN(n7791) );
  NAND2_X1 U9502 ( .A1(n8410), .A2(n8433), .ZN(n7790) );
  OAI211_X1 U9503 ( .C1(n8252), .C2(n8390), .A(n7791), .B(n7790), .ZN(n7792)
         );
  AOI211_X1 U9504 ( .C1(n7794), .C2(n8407), .A(n7793), .B(n7792), .ZN(n7795)
         );
  INV_X1 U9505 ( .A(n7795), .ZN(P2_U3153) );
  NAND2_X1 U9506 ( .A1(n8247), .A2(n7796), .ZN(n7798) );
  NAND2_X1 U9507 ( .A1(n7798), .A2(n7797), .ZN(n7864) );
  XNOR2_X1 U9508 ( .A(n6638), .B(n7864), .ZN(n7799) );
  AOI222_X1 U9509 ( .A1(n8781), .A2(n7799), .B1(n5211), .B2(n8694), .C1(n8434), 
        .C2(n8695), .ZN(n10290) );
  NAND2_X1 U9510 ( .A1(n8244), .A2(n7800), .ZN(n7801) );
  XNOR2_X1 U9511 ( .A(n7801), .B(n7863), .ZN(n10288) );
  NOR2_X1 U9512 ( .A1(n8714), .A2(n7802), .ZN(n7804) );
  OAI22_X1 U9513 ( .A1(n8700), .A2(n7636), .B1(n4464), .B2(n8712), .ZN(n7803)
         );
  AOI211_X1 U9514 ( .C1(n10288), .C2(n8727), .A(n7804), .B(n7803), .ZN(n7805)
         );
  OAI21_X1 U9515 ( .B1(n10290), .B2(n8708), .A(n7805), .ZN(P2_U3225) );
  XNOR2_X1 U9516 ( .A(n7806), .B(n7887), .ZN(n7809) );
  OR2_X1 U9517 ( .A1(n7908), .A2(n8972), .ZN(n7807) );
  OAI21_X1 U9518 ( .B1(n7808), .B2(n9140), .A(n7807), .ZN(n8063) );
  AOI21_X1 U9519 ( .B1(n7809), .B2(n9947), .A(n8063), .ZN(n10075) );
  OAI22_X1 U9520 ( .A1(n9588), .A2(n6025), .B1(n8065), .B2(n9949), .ZN(n7813)
         );
  INV_X1 U9521 ( .A(n7810), .ZN(n7811) );
  OAI211_X1 U9522 ( .C1(n10077), .C2(n7811), .A(n4521), .B(n9975), .ZN(n10074)
         );
  NOR2_X1 U9523 ( .A1(n10074), .A2(n9585), .ZN(n7812) );
  AOI211_X1 U9524 ( .C1(n9599), .C2(n8067), .A(n7813), .B(n7812), .ZN(n7819)
         );
  NAND2_X1 U9525 ( .A1(n7815), .A2(n7814), .ZN(n7817) );
  OR2_X1 U9526 ( .A1(n7990), .A2(n9002), .ZN(n7816) );
  NAND2_X1 U9527 ( .A1(n7817), .A2(n7816), .ZN(n7888) );
  XNOR2_X1 U9528 ( .A(n7888), .B(n7887), .ZN(n10079) );
  NAND2_X1 U9529 ( .A1(n10079), .A2(n9957), .ZN(n7818) );
  OAI211_X1 U9530 ( .C1(n9968), .C2(n10075), .A(n7819), .B(n7818), .ZN(
        P1_U3280) );
  INV_X1 U9531 ( .A(n7820), .ZN(n7822) );
  OAI222_X1 U9532 ( .A1(n7823), .A2(P2_U3151), .B1(n8851), .B2(n7822), .C1(
        n7821), .C2(n8848), .ZN(P2_U3275) );
  INV_X1 U9533 ( .A(n7824), .ZN(n7852) );
  OAI222_X1 U9534 ( .A1(n8275), .A2(n7852), .B1(n7826), .B2(P1_U3086), .C1(
        n7825), .C2(n8277), .ZN(P1_U3334) );
  NOR2_X1 U9535 ( .A1(n7835), .A2(n4469), .ZN(n7828) );
  NOR2_X1 U9536 ( .A1(n7828), .A2(n7827), .ZN(n7831) );
  INV_X1 U9537 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8462) );
  MUX2_X1 U9538 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n8462), .S(n8504), .Z(n7830)
         );
  INV_X1 U9539 ( .A(n8464), .ZN(n7829) );
  AOI21_X1 U9540 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n7850) );
  INV_X1 U9541 ( .A(n7832), .ZN(n7834) );
  MUX2_X1 U9542 ( .A(n8462), .B(n8503), .S(n7642), .Z(n7836) );
  NOR2_X1 U9543 ( .A1(n7836), .A2(n8504), .ZN(n8482) );
  NOR2_X1 U9544 ( .A1(n8482), .A2(n4528), .ZN(n7838) );
  NAND2_X1 U9545 ( .A1(n4522), .A2(n7838), .ZN(n7837) );
  OAI211_X1 U9546 ( .C1(n4522), .C2(n7838), .A(n10240), .B(n7837), .ZN(n7849)
         );
  NAND2_X1 U9547 ( .A1(n7840), .A2(n7839), .ZN(n7842) );
  XNOR2_X1 U9548 ( .A(n8504), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8500) );
  XNOR2_X1 U9549 ( .A(n8501), .B(n8500), .ZN(n7847) );
  INV_X1 U9550 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U9551 ( .A1(n10232), .A2(n8504), .ZN(n7844) );
  INV_X1 U9552 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9368) );
  NOR2_X1 U9553 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9368), .ZN(n8132) );
  INV_X1 U9554 ( .A(n8132), .ZN(n7843) );
  OAI211_X1 U9555 ( .C1(n7845), .C2(n10163), .A(n7844), .B(n7843), .ZN(n7846)
         );
  AOI21_X1 U9556 ( .B1(n7847), .B2(n10241), .A(n7846), .ZN(n7848) );
  OAI211_X1 U9557 ( .C1(n7850), .C2(n10246), .A(n7849), .B(n7848), .ZN(
        P2_U3194) );
  OAI222_X1 U9558 ( .A1(P2_U3151), .A2(n7853), .B1(n8851), .B2(n7852), .C1(
        n7851), .C2(n8848), .ZN(P2_U3274) );
  XOR2_X1 U9559 ( .A(n7855), .B(n7854), .Z(n7860) );
  AND2_X1 U9560 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8446) );
  AOI21_X1 U9561 ( .B1(n8387), .B2(n8434), .A(n8446), .ZN(n7857) );
  NAND2_X1 U9562 ( .A1(n8410), .A2(n5211), .ZN(n7856) );
  OAI211_X1 U9563 ( .C1(n4464), .C2(n8390), .A(n7857), .B(n7856), .ZN(n7858)
         );
  AOI21_X1 U9564 ( .B1(n10286), .B2(n8400), .A(n7858), .ZN(n7859) );
  OAI21_X1 U9565 ( .B1(n7860), .B2(n8403), .A(n7859), .ZN(P2_U3161) );
  OAI21_X1 U9566 ( .B1(n7862), .B2(n7867), .A(n7861), .ZN(n10293) );
  AOI22_X1 U9567 ( .A1(n8432), .A2(n8694), .B1(n8695), .B2(n8433), .ZN(n7871)
         );
  NAND2_X1 U9568 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  NAND2_X1 U9569 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  XNOR2_X1 U9570 ( .A(n7868), .B(n7867), .ZN(n7869) );
  NAND2_X1 U9571 ( .A1(n7869), .A2(n8781), .ZN(n7870) );
  OAI211_X1 U9572 ( .C1(n10293), .C2(n8251), .A(n7871), .B(n7870), .ZN(n10295)
         );
  NAND2_X1 U9574 ( .A1(n10295), .A2(n8700), .ZN(n7875) );
  OAI22_X1 U9575 ( .A1(n8700), .A2(n7872), .B1(n7882), .B2(n8712), .ZN(n7873)
         );
  AOI21_X1 U9576 ( .B1(n8702), .B2(n7884), .A(n7873), .ZN(n7874) );
  OAI211_X1 U9577 ( .C1(n10293), .C2(n8557), .A(n7875), .B(n7874), .ZN(
        P2_U3224) );
  OAI211_X1 U9578 ( .C1(n7878), .C2(n7877), .A(n7876), .B(n8407), .ZN(n7886)
         );
  AOI21_X1 U9579 ( .B1(n8387), .B2(n8433), .A(n7879), .ZN(n7881) );
  NAND2_X1 U9580 ( .A1(n8410), .A2(n8432), .ZN(n7880) );
  OAI211_X1 U9581 ( .C1(n7882), .C2(n8390), .A(n7881), .B(n7880), .ZN(n7883)
         );
  AOI21_X1 U9582 ( .B1(n7884), .B2(n8400), .A(n7883), .ZN(n7885) );
  NAND2_X1 U9583 ( .A1(n7886), .A2(n7885), .ZN(P2_U3171) );
  NAND2_X1 U9584 ( .A1(n7888), .A2(n7887), .ZN(n7890) );
  OR2_X1 U9585 ( .A1(n8067), .A2(n9001), .ZN(n7889) );
  NAND2_X1 U9586 ( .A1(n7890), .A2(n7889), .ZN(n7917) );
  XNOR2_X1 U9587 ( .A(n7917), .B(n7891), .ZN(n10086) );
  NAND2_X1 U9588 ( .A1(n7904), .A2(n9947), .ZN(n7897) );
  AOI21_X1 U9589 ( .B1(n7893), .B2(n7892), .A(n7891), .ZN(n7896) );
  OR2_X1 U9590 ( .A1(n7968), .A2(n8972), .ZN(n7895) );
  NAND2_X1 U9591 ( .A1(n9001), .A2(n8948), .ZN(n7894) );
  AND2_X1 U9592 ( .A1(n7895), .A2(n7894), .ZN(n8212) );
  OAI21_X1 U9593 ( .B1(n7897), .B2(n7896), .A(n8212), .ZN(n10081) );
  INV_X1 U9594 ( .A(n7898), .ZN(n7913) );
  AOI211_X1 U9595 ( .C1(n6021), .C2(n4521), .A(n9612), .B(n7913), .ZN(n10082)
         );
  NAND2_X1 U9596 ( .A1(n10082), .A2(n9978), .ZN(n7901) );
  INV_X1 U9597 ( .A(n7899), .ZN(n8214) );
  AOI22_X1 U9598 ( .A1(n9968), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8214), .B2(
        n9967), .ZN(n7900) );
  OAI211_X1 U9599 ( .C1(n8217), .C2(n9970), .A(n7901), .B(n7900), .ZN(n7902)
         );
  AOI21_X1 U9600 ( .B1(n9588), .B2(n10081), .A(n7902), .ZN(n7903) );
  OAI21_X1 U9601 ( .B1(n10086), .B2(n9623), .A(n7903), .ZN(P1_U3279) );
  INV_X1 U9602 ( .A(n7904), .ZN(n7906) );
  OAI21_X1 U9603 ( .B1(n7906), .B2(n7905), .A(n7972), .ZN(n7907) );
  AOI21_X1 U9604 ( .B1(n7907), .B2(n7965), .A(n9963), .ZN(n7911) );
  OR2_X1 U9605 ( .A1(n8071), .A2(n8972), .ZN(n7910) );
  OR2_X1 U9606 ( .A1(n7908), .A2(n9140), .ZN(n7909) );
  NAND2_X1 U9607 ( .A1(n7910), .A2(n7909), .ZN(n8984) );
  NOR2_X1 U9608 ( .A1(n7911), .A2(n8984), .ZN(n9768) );
  OAI22_X1 U9609 ( .A1(n9588), .A2(n7912), .B1(n8986), .B2(n9949), .ZN(n7915)
         );
  OAI211_X1 U9610 ( .C1(n7913), .C2(n9769), .A(n9975), .B(n4993), .ZN(n9767)
         );
  NOR2_X1 U9611 ( .A1(n9767), .A2(n9585), .ZN(n7914) );
  AOI211_X1 U9612 ( .C1(n9599), .C2(n8989), .A(n7915), .B(n7914), .ZN(n7921)
         );
  NAND2_X1 U9613 ( .A1(n7917), .A2(n7916), .ZN(n7919) );
  OR2_X1 U9614 ( .A1(n6021), .A2(n9000), .ZN(n7918) );
  NAND2_X1 U9615 ( .A1(n7919), .A2(n7918), .ZN(n7973) );
  XNOR2_X1 U9616 ( .A(n7973), .B(n7972), .ZN(n9771) );
  NAND2_X1 U9617 ( .A1(n9771), .A2(n9957), .ZN(n7920) );
  OAI211_X1 U9618 ( .C1(n9768), .C2(n9973), .A(n7921), .B(n7920), .ZN(P1_U3278) );
  OR2_X1 U9619 ( .A1(n7922), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U9620 ( .A1(n7925), .A2(n7924), .ZN(n7927) );
  XNOR2_X1 U9621 ( .A(n7927), .B(n7926), .ZN(n10304) );
  XNOR2_X1 U9622 ( .A(n7928), .B(n7929), .ZN(n7930) );
  OAI222_X1 U9623 ( .A1(n8720), .A2(n7932), .B1(n8718), .B2(n7931), .C1(n8635), 
        .C2(n7930), .ZN(n10305) );
  NOR2_X1 U9624 ( .A1(n8712), .A2(n8183), .ZN(n7933) );
  OAI21_X1 U9625 ( .B1(n10305), .B2(n7933), .A(n8700), .ZN(n7935) );
  AOI22_X1 U9626 ( .A1(n10307), .A2(n8702), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n8708), .ZN(n7934) );
  OAI211_X1 U9627 ( .C1(n8674), .C2(n10304), .A(n7935), .B(n7934), .ZN(
        P2_U3222) );
  INV_X1 U9628 ( .A(n7936), .ZN(n7940) );
  OAI222_X1 U9629 ( .A1(n8277), .A2(n7938), .B1(n8275), .B2(n7940), .C1(n8274), 
        .C2(n7937), .ZN(P1_U3333) );
  OAI222_X1 U9630 ( .A1(n7941), .A2(P2_U3151), .B1(n8851), .B2(n7940), .C1(
        n7939), .C2(n8848), .ZN(P2_U3273) );
  XOR2_X1 U9631 ( .A(n7922), .B(n7943), .Z(n10298) );
  XNOR2_X1 U9632 ( .A(n7942), .B(n7943), .ZN(n7948) );
  INV_X1 U9633 ( .A(n10298), .ZN(n7945) );
  NAND2_X1 U9634 ( .A1(n7945), .A2(n7944), .ZN(n7947) );
  AOI22_X1 U9635 ( .A1(n8695), .A2(n5211), .B1(n8431), .B2(n8694), .ZN(n7946)
         );
  OAI211_X1 U9636 ( .C1(n8635), .C2(n7948), .A(n7947), .B(n7946), .ZN(n10300)
         );
  NAND2_X1 U9637 ( .A1(n10300), .A2(n8700), .ZN(n7952) );
  OAI22_X1 U9638 ( .A1(n8700), .A2(n7949), .B1(n8123), .B2(n8712), .ZN(n7950)
         );
  AOI21_X1 U9639 ( .B1(n8702), .B2(n10301), .A(n7950), .ZN(n7951) );
  OAI211_X1 U9640 ( .C1(n10298), .C2(n8557), .A(n7952), .B(n7951), .ZN(
        P2_U3223) );
  XNOR2_X1 U9641 ( .A(n7953), .B(n8086), .ZN(n7956) );
  INV_X1 U9642 ( .A(n7954), .ZN(n7955) );
  NOR2_X1 U9643 ( .A1(n7956), .A2(n7955), .ZN(n8085) );
  AOI21_X1 U9644 ( .B1(n7956), .B2(n7955), .A(n8085), .ZN(n7963) );
  AOI22_X1 U9645 ( .A1(n4438), .A2(n7957), .B1(P1_REG3_REG_10__SCAN_IN), .B2(
        P1_U3086), .ZN(n7958) );
  OAI21_X1 U9646 ( .B1(n9796), .B2(n7959), .A(n7958), .ZN(n7960) );
  AOI21_X1 U9647 ( .B1(n7961), .B2(n8988), .A(n7960), .ZN(n7962) );
  OAI21_X1 U9648 ( .B1(n7963), .B2(n9791), .A(n7962), .ZN(P1_U3217) );
  AND2_X1 U9649 ( .A1(n7965), .A2(n7964), .ZN(n7967) );
  OAI211_X1 U9650 ( .C1(n7967), .C2(n4996), .A(n9947), .B(n7966), .ZN(n7971)
         );
  OR2_X1 U9651 ( .A1(n8143), .A2(n8972), .ZN(n7970) );
  OR2_X1 U9652 ( .A1(n7968), .A2(n9140), .ZN(n7969) );
  AND2_X1 U9653 ( .A1(n7970), .A2(n7969), .ZN(n8911) );
  NAND2_X1 U9654 ( .A1(n7971), .A2(n8911), .ZN(n9762) );
  INV_X1 U9655 ( .A(n9762), .ZN(n7982) );
  OR2_X1 U9656 ( .A1(n8989), .A2(n8999), .ZN(n7974) );
  NAND2_X1 U9657 ( .A1(n7976), .A2(n4996), .ZN(n9764) );
  NAND3_X1 U9658 ( .A1(n8074), .A2(n9764), .A3(n9957), .ZN(n7981) );
  AOI211_X1 U9659 ( .C1(n9763), .C2(n4993), .A(n9612), .B(n8079), .ZN(n9761)
         );
  AOI22_X1 U9660 ( .A1(n9968), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8909), .B2(
        n9967), .ZN(n7977) );
  OAI21_X1 U9661 ( .B1(n7978), .B2(n9970), .A(n7977), .ZN(n7979) );
  AOI21_X1 U9662 ( .B1(n9761), .B2(n9978), .A(n7979), .ZN(n7980) );
  OAI211_X1 U9663 ( .C1(n9968), .C2(n7982), .A(n7981), .B(n7980), .ZN(P1_U3277) );
  XOR2_X1 U9664 ( .A(n7983), .B(n7984), .Z(n7992) );
  AOI21_X1 U9665 ( .B1(n7986), .B2(n4438), .A(n7985), .ZN(n7987) );
  OAI21_X1 U9666 ( .B1(n9796), .B2(n7988), .A(n7987), .ZN(n7989) );
  AOI21_X1 U9667 ( .B1(n7990), .B2(n8988), .A(n7989), .ZN(n7991) );
  OAI21_X1 U9668 ( .B1(n7992), .B2(n9791), .A(n7991), .ZN(P1_U3224) );
  OR2_X1 U9669 ( .A1(n7922), .A2(n7993), .ZN(n7995) );
  AND2_X1 U9670 ( .A1(n7995), .A2(n7994), .ZN(n7996) );
  XNOR2_X1 U9671 ( .A(n7996), .B(n8000), .ZN(n8018) );
  INV_X1 U9672 ( .A(n8377), .ZN(n8006) );
  NOR2_X1 U9673 ( .A1(n7928), .A2(n7997), .ZN(n7999) );
  NOR2_X1 U9674 ( .A1(n7999), .A2(n7998), .ZN(n8002) );
  INV_X1 U9675 ( .A(n8000), .ZN(n8001) );
  XNOR2_X1 U9676 ( .A(n8002), .B(n8001), .ZN(n8005) );
  NAND2_X1 U9677 ( .A1(n8430), .A2(n8695), .ZN(n8003) );
  OAI21_X1 U9678 ( .B1(n8413), .B2(n8720), .A(n8003), .ZN(n8004) );
  AOI21_X1 U9679 ( .B1(n8005), .B2(n8781), .A(n8004), .ZN(n8014) );
  OAI21_X1 U9680 ( .B1(n8006), .B2(n8608), .A(n8014), .ZN(n8007) );
  NAND2_X1 U9681 ( .A1(n8007), .A2(n8700), .ZN(n8010) );
  INV_X1 U9682 ( .A(n8375), .ZN(n8008) );
  AOI22_X1 U9683 ( .A1(n8708), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n8671), .B2(
        n8008), .ZN(n8009) );
  OAI211_X1 U9684 ( .C1(n8018), .C2(n8674), .A(n8010), .B(n8009), .ZN(P2_U3220) );
  MUX2_X1 U9685 ( .A(n8011), .B(n8014), .S(n10325), .Z(n8013) );
  NAND2_X1 U9686 ( .A1(n8377), .A2(n8762), .ZN(n8012) );
  OAI211_X1 U9687 ( .C1(n8018), .C2(n8778), .A(n8013), .B(n8012), .ZN(P2_U3472) );
  INV_X1 U9688 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8015) );
  MUX2_X1 U9689 ( .A(n8015), .B(n8014), .S(n10309), .Z(n8017) );
  NAND2_X1 U9690 ( .A1(n8377), .A2(n6371), .ZN(n8016) );
  OAI211_X1 U9691 ( .C1(n8018), .C2(n8841), .A(n8017), .B(n8016), .ZN(P2_U3429) );
  NAND2_X1 U9692 ( .A1(n8022), .A2(n8288), .ZN(n8020) );
  OAI211_X1 U9693 ( .C1(n8021), .C2(n8848), .A(n8020), .B(n8019), .ZN(P2_U3272) );
  NAND2_X1 U9694 ( .A1(n8022), .A2(n9697), .ZN(n8024) );
  OAI211_X1 U9695 ( .C1(n9354), .C2(n8277), .A(n8024), .B(n8023), .ZN(P1_U3332) );
  OR2_X1 U9696 ( .A1(n7922), .A2(n8025), .ZN(n8028) );
  AND2_X1 U9697 ( .A1(n8028), .A2(n8026), .ZN(n8030) );
  NAND2_X1 U9698 ( .A1(n8028), .A2(n8027), .ZN(n8029) );
  OAI21_X1 U9699 ( .B1(n8030), .B2(n8035), .A(n8029), .ZN(n8103) );
  OR2_X1 U9700 ( .A1(n7928), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U9701 ( .A1(n8033), .A2(n8032), .ZN(n8034) );
  XOR2_X1 U9702 ( .A(n8035), .B(n8034), .Z(n8036) );
  OAI222_X1 U9703 ( .A1(n8720), .A2(n8037), .B1(n8718), .B2(n8134), .C1(n8635), 
        .C2(n8036), .ZN(n8098) );
  NOR2_X1 U9704 ( .A1(n8712), .A2(n8131), .ZN(n8038) );
  OAI21_X1 U9705 ( .B1(n8098), .B2(n8038), .A(n8700), .ZN(n8040) );
  AOI22_X1 U9706 ( .A1(n8127), .A2(n8702), .B1(P2_REG2_REG_12__SCAN_IN), .B2(
        n8708), .ZN(n8039) );
  OAI211_X1 U9707 ( .C1(n8103), .C2(n8674), .A(n8040), .B(n8039), .ZN(P2_U3221) );
  OR2_X1 U9708 ( .A1(n7922), .A2(n8041), .ZN(n8043) );
  AND2_X1 U9709 ( .A1(n8043), .A2(n8042), .ZN(n8045) );
  XNOR2_X1 U9710 ( .A(n8045), .B(n8044), .ZN(n8060) );
  XNOR2_X1 U9711 ( .A(n8047), .B(n8046), .ZN(n8048) );
  AOI222_X1 U9712 ( .A1(n8781), .A2(n8048), .B1(n8427), .B2(n8694), .C1(n8429), 
        .C2(n8695), .ZN(n8054) );
  MUX2_X1 U9713 ( .A(n8508), .B(n8054), .S(n10325), .Z(n8050) );
  NAND2_X1 U9714 ( .A1(n8300), .A2(n8762), .ZN(n8049) );
  OAI211_X1 U9715 ( .C1(n8060), .C2(n8778), .A(n8050), .B(n8049), .ZN(P2_U3473) );
  INV_X1 U9716 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8051) );
  MUX2_X1 U9717 ( .A(n8051), .B(n8054), .S(n10309), .Z(n8053) );
  NAND2_X1 U9718 ( .A1(n8300), .A2(n6371), .ZN(n8052) );
  OAI211_X1 U9719 ( .C1(n8060), .C2(n8841), .A(n8053), .B(n8052), .ZN(P2_U3432) );
  INV_X1 U9720 ( .A(n8054), .ZN(n8057) );
  INV_X1 U9721 ( .A(n8300), .ZN(n8055) );
  OAI22_X1 U9722 ( .A1(n8055), .A2(n8608), .B1(n8298), .B2(n8712), .ZN(n8056)
         );
  OAI21_X1 U9723 ( .B1(n8057), .B2(n8056), .A(n8700), .ZN(n8059) );
  NAND2_X1 U9724 ( .A1(n8708), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8058) );
  OAI211_X1 U9725 ( .C1(n8060), .C2(n8674), .A(n8059), .B(n8058), .ZN(P2_U3219) );
  XOR2_X1 U9726 ( .A(n8061), .B(n8062), .Z(n8069) );
  AOI22_X1 U9727 ( .A1(n4438), .A2(n8063), .B1(P1_REG3_REG_13__SCAN_IN), .B2(
        P1_U3086), .ZN(n8064) );
  OAI21_X1 U9728 ( .B1(n9796), .B2(n8065), .A(n8064), .ZN(n8066) );
  AOI21_X1 U9729 ( .B1(n8067), .B2(n8988), .A(n8066), .ZN(n8068) );
  OAI21_X1 U9730 ( .B1(n8069), .B2(n9791), .A(n8068), .ZN(P1_U3234) );
  XNOR2_X1 U9731 ( .A(n8070), .B(n8075), .ZN(n8072) );
  INV_X1 U9732 ( .A(n8071), .ZN(n8998) );
  AOI22_X1 U9733 ( .A1(n8996), .A2(n8924), .B1(n8948), .B2(n8998), .ZN(n8919)
         );
  OAI21_X1 U9734 ( .B1(n8072), .B2(n9963), .A(n8919), .ZN(n9759) );
  INV_X1 U9735 ( .A(n9759), .ZN(n8084) );
  NAND2_X1 U9736 ( .A1(n9763), .A2(n8998), .ZN(n8073) );
  NAND2_X1 U9737 ( .A1(n8074), .A2(n8073), .ZN(n8076) );
  INV_X1 U9738 ( .A(n8076), .ZN(n8078) );
  INV_X1 U9739 ( .A(n8075), .ZN(n8077) );
  OAI21_X1 U9740 ( .B1(n8078), .B2(n8077), .A(n4462), .ZN(n9760) );
  OAI211_X1 U9741 ( .C1(n9757), .C2(n8079), .A(n9975), .B(n8146), .ZN(n9756)
         );
  AOI22_X1 U9742 ( .A1(n9973), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n8917), .B2(
        n9967), .ZN(n8081) );
  NAND2_X1 U9743 ( .A1(n8921), .A2(n9599), .ZN(n8080) );
  OAI211_X1 U9744 ( .C1(n9756), .C2(n9585), .A(n8081), .B(n8080), .ZN(n8082)
         );
  AOI21_X1 U9745 ( .B1(n9760), .B2(n9957), .A(n8082), .ZN(n8083) );
  OAI21_X1 U9746 ( .B1(n9973), .B2(n8084), .A(n8083), .ZN(P1_U3276) );
  AOI21_X1 U9747 ( .B1(n8086), .B2(n7953), .A(n8085), .ZN(n8090) );
  XNOR2_X1 U9748 ( .A(n8088), .B(n8087), .ZN(n8089) );
  XNOR2_X1 U9749 ( .A(n8090), .B(n8089), .ZN(n8097) );
  AOI22_X1 U9750 ( .A1(n8091), .A2(n4438), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n8092) );
  OAI21_X1 U9751 ( .B1(n9796), .B2(n8093), .A(n8092), .ZN(n8094) );
  AOI21_X1 U9752 ( .B1(n8095), .B2(n8988), .A(n8094), .ZN(n8096) );
  OAI21_X1 U9753 ( .B1(n8097), .B2(n9791), .A(n8096), .ZN(P1_U3236) );
  AOI21_X1 U9754 ( .B1(n10308), .B2(n8127), .A(n8098), .ZN(n8100) );
  MUX2_X1 U9755 ( .A(n8503), .B(n8100), .S(n10325), .Z(n8099) );
  OAI21_X1 U9756 ( .B1(n8778), .B2(n8103), .A(n8099), .ZN(P2_U3471) );
  MUX2_X1 U9757 ( .A(n8101), .B(n8100), .S(n10309), .Z(n8102) );
  OAI21_X1 U9758 ( .B1(n8103), .B2(n8841), .A(n8102), .ZN(P2_U3426) );
  XNOR2_X1 U9759 ( .A(n8105), .B(n8104), .ZN(n8119) );
  XNOR2_X1 U9760 ( .A(n8107), .B(n8106), .ZN(n8108) );
  AOI222_X1 U9761 ( .A1(n8781), .A2(n8108), .B1(n8426), .B2(n8694), .C1(n8428), 
        .C2(n8695), .ZN(n8115) );
  MUX2_X1 U9762 ( .A(n10207), .B(n8115), .S(n8700), .Z(n8111) );
  INV_X1 U9763 ( .A(n8109), .ZN(n8416) );
  AOI22_X1 U9764 ( .A1(n8405), .A2(n8702), .B1(n8671), .B2(n8416), .ZN(n8110)
         );
  OAI211_X1 U9765 ( .C1(n8119), .C2(n8674), .A(n8111), .B(n8110), .ZN(P2_U3218) );
  MUX2_X1 U9766 ( .A(n8112), .B(n8115), .S(n10325), .Z(n8114) );
  NAND2_X1 U9767 ( .A1(n8405), .A2(n8762), .ZN(n8113) );
  OAI211_X1 U9768 ( .C1(n8778), .C2(n8119), .A(n8114), .B(n8113), .ZN(P2_U3474) );
  INV_X1 U9769 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8116) );
  MUX2_X1 U9770 ( .A(n8116), .B(n8115), .S(n10309), .Z(n8118) );
  NAND2_X1 U9771 ( .A1(n8405), .A2(n6371), .ZN(n8117) );
  OAI211_X1 U9772 ( .C1(n8119), .C2(n8841), .A(n8118), .B(n8117), .ZN(P2_U3435) );
  XNOR2_X1 U9773 ( .A(n8175), .B(n8432), .ZN(n8177) );
  XOR2_X1 U9774 ( .A(n8176), .B(n8177), .Z(n8126) );
  AOI21_X1 U9775 ( .B1(n8387), .B2(n5211), .A(n8120), .ZN(n8122) );
  NAND2_X1 U9776 ( .A1(n8410), .A2(n8431), .ZN(n8121) );
  OAI211_X1 U9777 ( .C1(n8123), .C2(n8390), .A(n8122), .B(n8121), .ZN(n8124)
         );
  AOI21_X1 U9778 ( .B1(n10301), .B2(n8400), .A(n8124), .ZN(n8125) );
  OAI21_X1 U9779 ( .B1(n8126), .B2(n8403), .A(n8125), .ZN(P2_U3157) );
  INV_X1 U9780 ( .A(n8127), .ZN(n8139) );
  OAI211_X1 U9781 ( .C1(n8130), .C2(n8129), .A(n8128), .B(n8407), .ZN(n8138)
         );
  INV_X1 U9782 ( .A(n8131), .ZN(n8136) );
  AOI21_X1 U9783 ( .B1(n8410), .B2(n8429), .A(n8132), .ZN(n8133) );
  OAI21_X1 U9784 ( .B1(n8134), .B2(n8412), .A(n8133), .ZN(n8135) );
  AOI21_X1 U9785 ( .B1(n8136), .B2(n8415), .A(n8135), .ZN(n8137) );
  OAI211_X1 U9786 ( .C1(n8139), .C2(n8419), .A(n8138), .B(n8137), .ZN(P2_U3164) );
  NAND2_X1 U9787 ( .A1(n8195), .A2(n8140), .ZN(n8141) );
  NAND2_X1 U9788 ( .A1(n8188), .A2(n8141), .ZN(n8142) );
  OAI22_X1 U9789 ( .A1(n8937), .A2(n8972), .B1(n8143), .B2(n9140), .ZN(n8964)
         );
  AOI21_X1 U9790 ( .B1(n8142), .B2(n9947), .A(n8964), .ZN(n9752) );
  INV_X1 U9791 ( .A(n8143), .ZN(n8997) );
  OR2_X1 U9792 ( .A1(n8921), .A2(n8997), .ZN(n8144) );
  XNOR2_X1 U9793 ( .A(n8196), .B(n8195), .ZN(n9755) );
  NAND2_X1 U9794 ( .A1(n9755), .A2(n9957), .ZN(n8151) );
  INV_X1 U9795 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8145) );
  OAI22_X1 U9796 ( .A1(n9588), .A2(n8145), .B1(n8961), .B2(n9949), .ZN(n8149)
         );
  INV_X1 U9797 ( .A(n8146), .ZN(n8147) );
  OAI211_X1 U9798 ( .C1(n8147), .C2(n9753), .A(n9975), .B(n8200), .ZN(n9751)
         );
  NOR2_X1 U9799 ( .A1(n9751), .A2(n9585), .ZN(n8148) );
  AOI211_X1 U9800 ( .C1(n9599), .C2(n8197), .A(n8149), .B(n8148), .ZN(n8150)
         );
  OAI211_X1 U9801 ( .C1(n9968), .C2(n9752), .A(n8151), .B(n8150), .ZN(P1_U3275) );
  INV_X1 U9802 ( .A(n8152), .ZN(n8286) );
  OAI222_X1 U9803 ( .A1(n8277), .A2(n8153), .B1(n5876), .B2(P1_U3086), .C1(
        n8275), .C2(n8286), .ZN(P1_U3331) );
  NAND2_X1 U9804 ( .A1(n8155), .A2(n8154), .ZN(n8156) );
  XNOR2_X1 U9805 ( .A(n8156), .B(n8157), .ZN(n8174) );
  NAND2_X1 U9806 ( .A1(n8158), .A2(n8157), .ZN(n8159) );
  NAND3_X1 U9807 ( .A1(n8160), .A2(n8781), .A3(n8159), .ZN(n8164) );
  OAI22_X1 U9808 ( .A1(n8161), .A2(n8718), .B1(n8334), .B2(n8720), .ZN(n8162)
         );
  INV_X1 U9809 ( .A(n8162), .ZN(n8163) );
  AND2_X1 U9810 ( .A1(n8164), .A2(n8163), .ZN(n8170) );
  MUX2_X1 U9811 ( .A(n8512), .B(n8170), .S(n10325), .Z(n8166) );
  NAND2_X1 U9812 ( .A1(n8339), .A2(n8762), .ZN(n8165) );
  OAI211_X1 U9813 ( .C1(n8174), .C2(n8778), .A(n8166), .B(n8165), .ZN(P2_U3475) );
  INV_X1 U9814 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8167) );
  MUX2_X1 U9815 ( .A(n8170), .B(n8167), .S(n10311), .Z(n8169) );
  NAND2_X1 U9816 ( .A1(n8339), .A2(n6371), .ZN(n8168) );
  OAI211_X1 U9817 ( .C1(n8174), .C2(n8841), .A(n8169), .B(n8168), .ZN(P2_U3438) );
  MUX2_X1 U9818 ( .A(n8170), .B(n8472), .S(n8708), .Z(n8173) );
  AOI22_X1 U9819 ( .A1(n8339), .A2(n8702), .B1(n8671), .B2(n8171), .ZN(n8172)
         );
  OAI211_X1 U9820 ( .C1(n8174), .C2(n8674), .A(n8173), .B(n8172), .ZN(P2_U3217) );
  OAI22_X1 U9821 ( .A1(n8177), .A2(n8176), .B1(n8432), .B2(n8175), .ZN(n8178)
         );
  XOR2_X1 U9822 ( .A(n8179), .B(n8178), .Z(n8186) );
  AOI21_X1 U9823 ( .B1(n8387), .B2(n8432), .A(n8180), .ZN(n8182) );
  NAND2_X1 U9824 ( .A1(n8410), .A2(n8430), .ZN(n8181) );
  OAI211_X1 U9825 ( .C1(n8183), .C2(n8390), .A(n8182), .B(n8181), .ZN(n8184)
         );
  AOI21_X1 U9826 ( .B1(n10307), .B2(n8400), .A(n8184), .ZN(n8185) );
  OAI21_X1 U9827 ( .B1(n8186), .B2(n8403), .A(n8185), .ZN(P2_U3176) );
  NAND3_X1 U9828 ( .A1(n8188), .A2(n8187), .A3(n8199), .ZN(n8189) );
  NAND2_X1 U9829 ( .A1(n8190), .A2(n8189), .ZN(n8194) );
  OR2_X1 U9830 ( .A1(n8889), .A2(n8972), .ZN(n8192) );
  NAND2_X1 U9831 ( .A1(n8996), .A2(n8948), .ZN(n8191) );
  AND2_X1 U9832 ( .A1(n8192), .A2(n8191), .ZN(n8881) );
  INV_X1 U9833 ( .A(n8881), .ZN(n8193) );
  AOI21_X1 U9834 ( .B1(n8194), .B2(n9947), .A(n8193), .ZN(n9747) );
  OR2_X1 U9835 ( .A1(n8197), .A2(n8996), .ZN(n8198) );
  XNOR2_X1 U9836 ( .A(n9144), .B(n8199), .ZN(n9750) );
  NAND2_X1 U9837 ( .A1(n9750), .A2(n9957), .ZN(n8206) );
  INV_X1 U9838 ( .A(n9146), .ZN(n9748) );
  INV_X1 U9839 ( .A(n8200), .ZN(n8201) );
  OAI211_X1 U9840 ( .C1(n9748), .C2(n8201), .A(n4460), .B(n9975), .ZN(n9746)
         );
  INV_X1 U9841 ( .A(n9746), .ZN(n8204) );
  AOI22_X1 U9842 ( .A1(n8879), .A2(n9967), .B1(n9968), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n8202) );
  OAI21_X1 U9843 ( .B1(n9748), .B2(n9970), .A(n8202), .ZN(n8203) );
  AOI21_X1 U9844 ( .B1(n8204), .B2(n9978), .A(n8203), .ZN(n8205) );
  OAI211_X1 U9845 ( .C1(n9968), .C2(n9747), .A(n8206), .B(n8205), .ZN(P1_U3274) );
  OAI21_X1 U9846 ( .B1(n8209), .B2(n8208), .A(n8207), .ZN(n8210) );
  NAND2_X1 U9847 ( .A1(n8210), .A2(n8968), .ZN(n8216) );
  INV_X1 U9848 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8211) );
  AOI21_X1 U9849 ( .B1(n8214), .B2(n8925), .A(n8213), .ZN(n8215) );
  OAI211_X1 U9850 ( .C1(n8217), .C2(n9786), .A(n8216), .B(n8215), .ZN(P1_U3215) );
  INV_X1 U9851 ( .A(n8218), .ZN(n8221) );
  INV_X1 U9852 ( .A(n8219), .ZN(n8222) );
  OAI222_X1 U9853 ( .A1(n8221), .A2(P2_U3151), .B1(n8851), .B2(n8222), .C1(
        n8220), .C2(n8848), .ZN(P2_U3270) );
  OAI222_X1 U9854 ( .A1(n8277), .A2(n8224), .B1(n8223), .B2(P1_U3086), .C1(
        n8275), .C2(n8222), .ZN(P1_U3330) );
  INV_X1 U9855 ( .A(n8225), .ZN(n8228) );
  OAI222_X1 U9856 ( .A1(n8227), .A2(P2_U3151), .B1(n8851), .B2(n8228), .C1(
        n8226), .C2(n8848), .ZN(P2_U3269) );
  OAI222_X1 U9857 ( .A1(n8277), .A2(n8230), .B1(n8229), .B2(P1_U3086), .C1(
        n8275), .C2(n8228), .ZN(P1_U3329) );
  INV_X1 U9858 ( .A(n8231), .ZN(n8240) );
  AOI21_X1 U9859 ( .B1(n8289), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8232), .ZN(
        n8233) );
  OAI21_X1 U9860 ( .B1(n8240), .B2(n8851), .A(n8233), .ZN(P2_U3268) );
  INV_X1 U9861 ( .A(n8234), .ZN(n8239) );
  AOI21_X1 U9862 ( .B1(n8289), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8235), .ZN(
        n8236) );
  OAI21_X1 U9863 ( .B1(n8239), .B2(n8851), .A(n8236), .ZN(P2_U3267) );
  OAI222_X1 U9864 ( .A1(n8275), .A2(n8239), .B1(n8238), .B2(P1_U3086), .C1(
        n8237), .C2(n8277), .ZN(P1_U3327) );
  OAI222_X1 U9865 ( .A1(n4451), .A2(P1_U3086), .B1(n8275), .B2(n8240), .C1(
        n8277), .C2(n5827), .ZN(P1_U3328) );
  INV_X1 U9866 ( .A(n6351), .ZN(n9702) );
  OAI222_X1 U9867 ( .A1(P2_U3151), .A2(n8242), .B1(n8851), .B2(n9702), .C1(
        n8241), .C2(n8848), .ZN(P2_U3266) );
  OAI21_X1 U9868 ( .B1(n8245), .B2(n8246), .A(n8244), .ZN(n10282) );
  AOI22_X1 U9869 ( .A1(n8694), .A2(n8433), .B1(n8435), .B2(n8695), .ZN(n8250)
         );
  XNOR2_X1 U9870 ( .A(n8247), .B(n8246), .ZN(n8248) );
  NAND2_X1 U9871 ( .A1(n8248), .A2(n8781), .ZN(n8249) );
  OAI211_X1 U9872 ( .C1(n10282), .C2(n8251), .A(n8250), .B(n8249), .ZN(n10284)
         );
  NAND2_X1 U9873 ( .A1(n10284), .A2(n8700), .ZN(n8256) );
  OAI22_X1 U9874 ( .A1(n8700), .A2(n7377), .B1(n8252), .B2(n8712), .ZN(n8253)
         );
  AOI21_X1 U9875 ( .B1(n8702), .B2(n8254), .A(n8253), .ZN(n8255) );
  OAI211_X1 U9876 ( .C1(n10282), .C2(n8557), .A(n8256), .B(n8255), .ZN(
        P2_U3226) );
  AND2_X1 U9877 ( .A1(n8395), .A2(n8257), .ZN(n8263) );
  INV_X1 U9878 ( .A(n8257), .ZN(n8262) );
  INV_X1 U9879 ( .A(n8258), .ZN(n8260) );
  AND2_X1 U9880 ( .A1(n8260), .A2(n8259), .ZN(n8261) );
  XNOR2_X1 U9881 ( .A(n8264), .B(n6851), .ZN(n8265) );
  XNOR2_X1 U9882 ( .A(n8266), .B(n8265), .ZN(n8271) );
  NOR2_X1 U9883 ( .A1(n8390), .A2(n8560), .ZN(n8269) );
  AOI22_X1 U9884 ( .A1(n8410), .A2(n8421), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8267) );
  OAI21_X1 U9885 ( .B1(n8589), .B2(n8412), .A(n8267), .ZN(n8268) );
  AOI211_X1 U9886 ( .C1(n8563), .C2(n8400), .A(n8269), .B(n8268), .ZN(n8270)
         );
  OAI21_X1 U9887 ( .B1(n8271), .B2(n8403), .A(n8270), .ZN(P2_U3160) );
  INV_X1 U9888 ( .A(n8272), .ZN(n8850) );
  OAI222_X1 U9889 ( .A1(n8277), .A2(n8276), .B1(n8275), .B2(n8850), .C1(n8274), 
        .C2(n8273), .ZN(P1_U3325) );
  XOR2_X1 U9890 ( .A(n8279), .B(n8278), .Z(n8284) );
  NAND2_X1 U9891 ( .A1(n8415), .A2(n8661), .ZN(n8281) );
  AOI22_X1 U9892 ( .A1(n8387), .A2(n8657), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8280) );
  OAI211_X1 U9893 ( .C1(n8622), .C2(n8397), .A(n8281), .B(n8280), .ZN(n8282)
         );
  AOI21_X1 U9894 ( .B1(n5444), .B2(n8400), .A(n8282), .ZN(n8283) );
  OAI21_X1 U9895 ( .B1(n8284), .B2(n8403), .A(n8283), .ZN(P2_U3163) );
  OAI222_X1 U9896 ( .A1(n8287), .A2(P2_U3151), .B1(n8851), .B2(n8286), .C1(
        n8285), .C2(n8848), .ZN(P2_U3271) );
  NAND3_X1 U9897 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_STATE_REG_SCAN_IN), .A3(
        n5011), .ZN(n8292) );
  NAND2_X1 U9898 ( .A1(n9698), .A2(n8288), .ZN(n8291) );
  NAND2_X1 U9899 ( .A1(n8289), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8290) );
  OAI211_X1 U9900 ( .C1(n8293), .C2(n8292), .A(n8291), .B(n8290), .ZN(P2_U3264) );
  XOR2_X1 U9901 ( .A(n8295), .B(n8294), .Z(n8302) );
  AOI22_X1 U9902 ( .A1(n8410), .A2(n8427), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8297) );
  NAND2_X1 U9903 ( .A1(n8387), .A2(n8429), .ZN(n8296) );
  OAI211_X1 U9904 ( .C1(n8390), .C2(n8298), .A(n8297), .B(n8296), .ZN(n8299)
         );
  AOI21_X1 U9905 ( .B1(n8300), .B2(n8400), .A(n8299), .ZN(n8301) );
  OAI21_X1 U9906 ( .B1(n8302), .B2(n8403), .A(n8301), .ZN(P2_U3155) );
  XNOR2_X1 U9907 ( .A(n8303), .B(n8424), .ZN(n8309) );
  INV_X1 U9908 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8304) );
  OAI22_X1 U9909 ( .A1(n8622), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8304), .ZN(n8306) );
  NOR2_X1 U9910 ( .A1(n8621), .A2(n8397), .ZN(n8305) );
  AOI211_X1 U9911 ( .C1(n8625), .C2(n8415), .A(n8306), .B(n8305), .ZN(n8308)
         );
  NAND2_X1 U9912 ( .A1(n8749), .A2(n8400), .ZN(n8307) );
  OAI211_X1 U9913 ( .C1(n8309), .C2(n8403), .A(n8308), .B(n8307), .ZN(P2_U3156) );
  NAND2_X1 U9914 ( .A1(n8310), .A2(n8386), .ZN(n8315) );
  NAND2_X1 U9915 ( .A1(n8315), .A2(n8311), .ZN(n8313) );
  AOI21_X1 U9916 ( .B1(n8313), .B2(n8312), .A(n8403), .ZN(n8317) );
  NAND2_X1 U9917 ( .A1(n8315), .A2(n8314), .ZN(n8316) );
  NAND2_X1 U9918 ( .A1(n8317), .A2(n8316), .ZN(n8321) );
  NAND2_X1 U9919 ( .A1(n8410), .A2(n8657), .ZN(n8318) );
  NAND2_X1 U9920 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8532) );
  OAI211_X1 U9921 ( .C1(n8721), .C2(n8412), .A(n8318), .B(n8532), .ZN(n8319)
         );
  AOI21_X1 U9922 ( .B1(n8682), .B2(n8415), .A(n8319), .ZN(n8320) );
  OAI211_X1 U9923 ( .C1(n8768), .C2(n8419), .A(n8321), .B(n8320), .ZN(P2_U3159) );
  XOR2_X1 U9924 ( .A(n8323), .B(n8322), .Z(n8329) );
  OAI22_X1 U9925 ( .A1(n8621), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8324), .ZN(n8326) );
  NOR2_X1 U9926 ( .A1(n8568), .A2(n8397), .ZN(n8325) );
  AOI211_X1 U9927 ( .C1(n8601), .C2(n8415), .A(n8326), .B(n8325), .ZN(n8328)
         );
  NAND2_X1 U9928 ( .A1(n8809), .A2(n8400), .ZN(n8327) );
  OAI211_X1 U9929 ( .C1(n8329), .C2(n8403), .A(n8328), .B(n8327), .ZN(P2_U3165) );
  NAND2_X1 U9930 ( .A1(n8331), .A2(n8330), .ZN(n8333) );
  XOR2_X1 U9931 ( .A(n8333), .B(n8332), .Z(n8341) );
  NAND2_X1 U9932 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n10228) );
  OAI21_X1 U9933 ( .B1(n8397), .B2(n8334), .A(n10228), .ZN(n8335) );
  AOI21_X1 U9934 ( .B1(n8387), .B2(n8427), .A(n8335), .ZN(n8336) );
  OAI21_X1 U9935 ( .B1(n8337), .B2(n8390), .A(n8336), .ZN(n8338) );
  AOI21_X1 U9936 ( .B1(n8339), .B2(n8400), .A(n8338), .ZN(n8340) );
  OAI21_X1 U9937 ( .B1(n8341), .B2(n8403), .A(n8340), .ZN(P2_U3166) );
  XOR2_X1 U9938 ( .A(n8343), .B(n8342), .Z(n8349) );
  OAI22_X1 U9939 ( .A1(n8397), .A2(n8721), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8344), .ZN(n8345) );
  AOI21_X1 U9940 ( .B1(n8387), .B2(n8426), .A(n8345), .ZN(n8346) );
  OAI21_X1 U9941 ( .B1(n8713), .B2(n8390), .A(n8346), .ZN(n8347) );
  AOI21_X1 U9942 ( .B1(n8711), .B2(n8400), .A(n8347), .ZN(n8348) );
  OAI21_X1 U9943 ( .B1(n8349), .B2(n8403), .A(n8348), .ZN(P2_U3168) );
  XOR2_X1 U9944 ( .A(n8351), .B(n8350), .Z(n8356) );
  AOI22_X1 U9945 ( .A1(n8424), .A2(n8387), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8353) );
  NAND2_X1 U9946 ( .A1(n8415), .A2(n8613), .ZN(n8352) );
  OAI211_X1 U9947 ( .C1(n8611), .C2(n8397), .A(n8353), .B(n8352), .ZN(n8354)
         );
  AOI21_X1 U9948 ( .B1(n8744), .B2(n8400), .A(n8354), .ZN(n8355) );
  OAI21_X1 U9949 ( .B1(n8356), .B2(n8403), .A(n8355), .ZN(P2_U3169) );
  NAND2_X1 U9950 ( .A1(n8310), .A2(n8357), .ZN(n8359) );
  AND2_X1 U9951 ( .A1(n8359), .A2(n8358), .ZN(n8360) );
  AOI21_X1 U9952 ( .B1(n8361), .B2(n8360), .A(n4994), .ZN(n8367) );
  NAND2_X1 U9953 ( .A1(n8415), .A2(n8670), .ZN(n8363) );
  AOI22_X1 U9954 ( .A1(n8667), .A2(n8410), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8362) );
  OAI211_X1 U9955 ( .C1(n8364), .C2(n8412), .A(n8363), .B(n8362), .ZN(n8365)
         );
  AOI21_X1 U9956 ( .B1(n8832), .B2(n8400), .A(n8365), .ZN(n8366) );
  OAI21_X1 U9957 ( .B1(n8367), .B2(n8403), .A(n8366), .ZN(P2_U3173) );
  INV_X1 U9958 ( .A(n8368), .ZN(n8369) );
  AOI21_X1 U9959 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8379) );
  OAI22_X1 U9960 ( .A1(n8397), .A2(n8413), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8372), .ZN(n8373) );
  AOI21_X1 U9961 ( .B1(n8387), .B2(n8430), .A(n8373), .ZN(n8374) );
  OAI21_X1 U9962 ( .B1(n8375), .B2(n8390), .A(n8374), .ZN(n8376) );
  AOI21_X1 U9963 ( .B1(n8377), .B2(n8400), .A(n8376), .ZN(n8378) );
  OAI21_X1 U9964 ( .B1(n8379), .B2(n8403), .A(n8378), .ZN(P2_U3174) );
  XNOR2_X1 U9965 ( .A(n8380), .B(n8658), .ZN(n8385) );
  NAND2_X1 U9966 ( .A1(n8415), .A2(n8642), .ZN(n8382) );
  AOI22_X1 U9967 ( .A1(n8387), .A2(n8667), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8381) );
  OAI211_X1 U9968 ( .C1(n8637), .C2(n8397), .A(n8382), .B(n8381), .ZN(n8383)
         );
  AOI21_X1 U9969 ( .B1(n8641), .B2(n8400), .A(n8383), .ZN(n8384) );
  OAI21_X1 U9970 ( .B1(n8385), .B2(n8403), .A(n8384), .ZN(P2_U3175) );
  XOR2_X1 U9971 ( .A(n8310), .B(n8386), .Z(n8393) );
  AOI22_X1 U9972 ( .A1(n8410), .A2(n8693), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8389) );
  NAND2_X1 U9973 ( .A1(n8387), .A2(n8696), .ZN(n8388) );
  OAI211_X1 U9974 ( .C1(n8390), .C2(n8699), .A(n8389), .B(n8388), .ZN(n8391)
         );
  AOI21_X1 U9975 ( .B1(n8703), .B2(n8400), .A(n8391), .ZN(n8392) );
  OAI21_X1 U9976 ( .B1(n8393), .B2(n8403), .A(n8392), .ZN(P2_U3178) );
  XNOR2_X1 U9977 ( .A(n8394), .B(n4925), .ZN(n8404) );
  OAI22_X1 U9978 ( .A1(n8611), .A2(n8412), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8396), .ZN(n8399) );
  NOR2_X1 U9979 ( .A1(n8589), .A2(n8397), .ZN(n8398) );
  AOI211_X1 U9980 ( .C1(n8592), .C2(n8415), .A(n8399), .B(n8398), .ZN(n8402)
         );
  NAND2_X1 U9981 ( .A1(n8803), .A2(n8400), .ZN(n8401) );
  OAI211_X1 U9982 ( .C1(n8404), .C2(n8403), .A(n8402), .B(n8401), .ZN(P2_U3180) );
  INV_X1 U9983 ( .A(n8405), .ZN(n8420) );
  OAI211_X1 U9984 ( .C1(n8406), .C2(n8409), .A(n8408), .B(n8407), .ZN(n8418)
         );
  AND2_X1 U9985 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10206) );
  AOI21_X1 U9986 ( .B1(n8410), .B2(n8426), .A(n10206), .ZN(n8411) );
  OAI21_X1 U9987 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  AOI21_X1 U9988 ( .B1(n8416), .B2(n8415), .A(n8414), .ZN(n8417) );
  OAI211_X1 U9989 ( .C1(n8420), .C2(n8419), .A(n8418), .B(n8417), .ZN(P2_U3181) );
  MUX2_X1 U9990 ( .A(n8544), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8492), .Z(
        P2_U3522) );
  MUX2_X1 U9991 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8421), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U9992 ( .A(n8422), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8492), .Z(
        P2_U3519) );
  MUX2_X1 U9993 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8598), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9994 ( .A(n8423), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8492), .Z(
        P2_U3516) );
  MUX2_X1 U9995 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8599), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9996 ( .A(n8424), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8492), .Z(
        P2_U3514) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8658), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9998 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8667), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9999 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8657), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10000 ( .A(n8693), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8492), .Z(
        P2_U3510) );
  MUX2_X1 U10001 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8425), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10002 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8696), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10003 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8426), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10004 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8427), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10005 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8428), .S(P2_U3893), .Z(
        P2_U3505) );
  MUX2_X1 U10006 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8429), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10007 ( .A(n8430), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8492), .Z(
        P2_U3503) );
  MUX2_X1 U10008 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8431), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10009 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8432), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10010 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n5211), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10011 ( .A(n8433), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8492), .Z(
        P2_U3499) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8434), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10013 ( .A(n8435), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8492), .Z(
        P2_U3497) );
  MUX2_X1 U10014 ( .A(n8436), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8492), .Z(
        P2_U3496) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8437), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n4444), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10017 ( .A(n8438), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8492), .Z(
        P2_U3493) );
  MUX2_X1 U10018 ( .A(n6849), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8492), .Z(
        P2_U3492) );
  AND3_X1 U10019 ( .A1(n8441), .A2(n8440), .A3(n8439), .ZN(n8442) );
  OAI21_X1 U10020 ( .B1(n8443), .B2(n8442), .A(n10240), .ZN(n8459) );
  INV_X1 U10021 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8444) );
  NOR2_X1 U10022 ( .A1(n10163), .A2(n8444), .ZN(n8445) );
  AOI211_X1 U10023 ( .C1(n10232), .C2(n8447), .A(n8446), .B(n8445), .ZN(n8458)
         );
  OAI21_X1 U10024 ( .B1(n8450), .B2(n8449), .A(n8448), .ZN(n8451) );
  NAND2_X1 U10025 ( .A1(n8451), .A2(n10241), .ZN(n8457) );
  AND3_X1 U10026 ( .A1(n8453), .A2(n8452), .A3(n4465), .ZN(n8454) );
  OAI21_X1 U10027 ( .B1(n8455), .B2(n8454), .A(n10175), .ZN(n8456) );
  NAND4_X1 U10028 ( .A1(n8459), .A2(n8458), .A3(n8457), .A4(n8456), .ZN(
        P2_U3190) );
  INV_X1 U10029 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8461) );
  NOR2_X1 U10030 ( .A1(n8523), .A2(n8461), .ZN(n8460) );
  AOI21_X1 U10031 ( .B1(n8461), .B2(n8523), .A(n8460), .ZN(n8477) );
  OR2_X1 U10032 ( .A1(n8504), .A2(n8462), .ZN(n8463) );
  INV_X1 U10033 ( .A(n8466), .ZN(n8465) );
  NOR2_X1 U10034 ( .A1(n10165), .A2(n8465), .ZN(n8468) );
  XNOR2_X1 U10035 ( .A(n10182), .B(n8469), .ZN(n10192) );
  XNOR2_X1 U10036 ( .A(n10198), .B(n8471), .ZN(n10208) );
  NOR2_X1 U10037 ( .A1(n8498), .A2(n8472), .ZN(n8473) );
  AOI21_X1 U10038 ( .B1(n8472), .B2(n8498), .A(n8473), .ZN(n10224) );
  NOR2_X1 U10039 ( .A1(n10233), .A2(n8475), .ZN(n8476) );
  AOI21_X1 U10040 ( .B1(n8477), .B2(n4476), .A(n8521), .ZN(n8520) );
  INV_X1 U10041 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8497) );
  MUX2_X1 U10042 ( .A(n8478), .B(n9447), .S(n7642), .Z(n8487) );
  XNOR2_X1 U10043 ( .A(n8487), .B(n8513), .ZN(n10238) );
  MUX2_X1 U10044 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n7642), .Z(n8479) );
  OR2_X1 U10045 ( .A1(n8479), .A2(n8498), .ZN(n8486) );
  XNOR2_X1 U10046 ( .A(n8479), .B(n10214), .ZN(n10220) );
  MUX2_X1 U10047 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n7642), .Z(n8480) );
  OR2_X1 U10048 ( .A1(n8480), .A2(n8510), .ZN(n8485) );
  XNOR2_X1 U10049 ( .A(n8480), .B(n10198), .ZN(n10203) );
  MUX2_X1 U10050 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n7642), .Z(n8481) );
  OR2_X1 U10051 ( .A1(n8481), .A2(n8499), .ZN(n8484) );
  XNOR2_X1 U10052 ( .A(n8481), .B(n10182), .ZN(n10188) );
  MUX2_X1 U10053 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n7642), .Z(n8483) );
  XNOR2_X1 U10054 ( .A(n8483), .B(n10165), .ZN(n10170) );
  NAND2_X1 U10055 ( .A1(n10188), .A2(n10187), .ZN(n10186) );
  NAND2_X1 U10056 ( .A1(n8486), .A2(n10218), .ZN(n10237) );
  MUX2_X1 U10057 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n7642), .Z(n8490) );
  INV_X1 U10058 ( .A(n8490), .ZN(n8488) );
  NAND2_X1 U10059 ( .A1(n8489), .A2(n8488), .ZN(n8528) );
  INV_X1 U10060 ( .A(n8528), .ZN(n8495) );
  NAND2_X1 U10061 ( .A1(n8491), .A2(n8490), .ZN(n8493) );
  NAND2_X1 U10062 ( .A1(n8493), .A2(n8516), .ZN(n8529) );
  INV_X1 U10063 ( .A(n8493), .ZN(n8494) );
  OAI211_X1 U10064 ( .C1(n8495), .C2(n8494), .A(n10240), .B(n8523), .ZN(n8496)
         );
  AOI22_X1 U10065 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8498), .B1(n10214), 
        .B2(n8512), .ZN(n10217) );
  AOI22_X1 U10066 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8499), .B1(n10182), 
        .B2(n8508), .ZN(n10185) );
  NAND2_X1 U10067 ( .A1(n8501), .A2(n8500), .ZN(n8502) );
  OAI21_X1 U10068 ( .B1(n8504), .B2(n8503), .A(n8502), .ZN(n8505) );
  NAND2_X1 U10069 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  XOR2_X1 U10070 ( .A(n8506), .B(n8505), .Z(n10167) );
  NAND2_X1 U10071 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10167), .ZN(n10166) );
  NAND2_X1 U10072 ( .A1(n8510), .A2(n8509), .ZN(n8511) );
  NAND2_X1 U10073 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10200), .ZN(n10199) );
  NAND2_X1 U10074 ( .A1(n8511), .A2(n10199), .ZN(n10216) );
  NAND2_X1 U10075 ( .A1(n10217), .A2(n10216), .ZN(n10215) );
  OAI21_X1 U10076 ( .B1(n10214), .B2(n8512), .A(n10215), .ZN(n8514) );
  NAND2_X1 U10077 ( .A1(n8513), .A2(n8514), .ZN(n8515) );
  XNOR2_X1 U10078 ( .A(n10233), .B(n8514), .ZN(n10235) );
  XNOR2_X1 U10079 ( .A(n8516), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8524) );
  XNOR2_X1 U10080 ( .A(n8525), .B(n8524), .ZN(n8517) );
  NAND2_X1 U10081 ( .A1(n8517), .A2(n10241), .ZN(n8518) );
  OAI211_X1 U10082 ( .C1(n8520), .C2(n10246), .A(n8519), .B(n8518), .ZN(
        P2_U3200) );
  MUX2_X1 U10083 ( .A(n8684), .B(P2_REG2_REG_19__SCAN_IN), .S(n8535), .Z(n8527) );
  XNOR2_X1 U10084 ( .A(n8522), .B(n8527), .ZN(n8541) );
  MUX2_X1 U10085 ( .A(n8527), .B(n4529), .S(n7642), .Z(n8531) );
  NAND2_X1 U10086 ( .A1(n8529), .A2(n8528), .ZN(n8530) );
  XOR2_X1 U10087 ( .A(n8531), .B(n8530), .Z(n8537) );
  INV_X1 U10088 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8533) );
  OAI21_X1 U10089 ( .B1(n10163), .B2(n8533), .A(n8532), .ZN(n8534) );
  AOI21_X1 U10090 ( .B1(n8535), .B2(n10232), .A(n8534), .ZN(n8536) );
  OAI21_X1 U10091 ( .B1(n8537), .B2(n10159), .A(n8536), .ZN(n8538) );
  AOI21_X1 U10092 ( .B1(n8539), .B2(n10241), .A(n8538), .ZN(n8540) );
  OAI21_X1 U10093 ( .B1(n8541), .B2(n10246), .A(n8540), .ZN(P2_U3201) );
  INV_X1 U10094 ( .A(n8542), .ZN(n8543) );
  AND2_X1 U10095 ( .A1(n8544), .A2(n8543), .ZN(n8790) );
  NOR2_X1 U10096 ( .A1(n8712), .A2(n8545), .ZN(n8554) );
  AOI21_X1 U10097 ( .B1(n8700), .B2(n8790), .A(n8554), .ZN(n8547) );
  NAND2_X1 U10098 ( .A1(n8708), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8546) );
  OAI211_X1 U10099 ( .C1(n8793), .C2(n8714), .A(n8547), .B(n8546), .ZN(
        P2_U3202) );
  NAND2_X1 U10100 ( .A1(n6657), .A2(n8702), .ZN(n8548) );
  OAI211_X1 U10101 ( .C1(n8700), .C2(n8549), .A(n8548), .B(n8547), .ZN(
        P2_U3203) );
  INV_X1 U10102 ( .A(n8550), .ZN(n8558) );
  NAND2_X1 U10103 ( .A1(n8551), .A2(n8700), .ZN(n8556) );
  NOR2_X1 U10104 ( .A1(n8552), .A2(n8714), .ZN(n8553) );
  AOI211_X1 U10105 ( .C1(n8708), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8554), .B(
        n8553), .ZN(n8555) );
  OAI211_X1 U10106 ( .C1(n8558), .C2(n8557), .A(n8556), .B(n8555), .ZN(
        P2_U3204) );
  NAND2_X1 U10107 ( .A1(n8559), .A2(n8700), .ZN(n8565) );
  OAI22_X1 U10108 ( .A1(n8700), .A2(n8561), .B1(n8560), .B2(n8712), .ZN(n8562)
         );
  AOI21_X1 U10109 ( .B1(n8563), .B2(n8702), .A(n8562), .ZN(n8564) );
  OAI211_X1 U10110 ( .C1(n8566), .C2(n8674), .A(n8565), .B(n8564), .ZN(
        P2_U3205) );
  XNOR2_X1 U10111 ( .A(n8567), .B(n8576), .ZN(n8573) );
  OAI22_X1 U10112 ( .A1(n8570), .A2(n8569), .B1(n8718), .B2(n8568), .ZN(n8571)
         );
  NAND2_X1 U10113 ( .A1(n8575), .A2(n8574), .ZN(n8577) );
  NAND2_X1 U10114 ( .A1(n8577), .A2(n8576), .ZN(n8578) );
  NAND2_X1 U10115 ( .A1(n8579), .A2(n8578), .ZN(n8800) );
  AOI22_X1 U10116 ( .A1(n8580), .A2(n8671), .B1(n8708), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8582) );
  NAND2_X1 U10117 ( .A1(n8735), .A2(n8702), .ZN(n8581) );
  OAI211_X1 U10118 ( .C1(n8800), .C2(n8674), .A(n8582), .B(n8581), .ZN(n8583)
         );
  AOI21_X1 U10119 ( .B1(n8734), .B2(n8700), .A(n8583), .ZN(n8584) );
  INV_X1 U10120 ( .A(n8584), .ZN(P2_U3206) );
  XNOR2_X1 U10121 ( .A(n8585), .B(n8586), .ZN(n8806) );
  XNOR2_X1 U10122 ( .A(n8588), .B(n8587), .ZN(n8591) );
  OAI22_X1 U10123 ( .A1(n8589), .A2(n8720), .B1(n8611), .B2(n8718), .ZN(n8590)
         );
  AOI21_X1 U10124 ( .B1(n8591), .B2(n8781), .A(n8590), .ZN(n8801) );
  MUX2_X1 U10125 ( .A(n9306), .B(n8801), .S(n8700), .Z(n8594) );
  AOI22_X1 U10126 ( .A1(n8803), .A2(n8702), .B1(n8671), .B2(n8592), .ZN(n8593)
         );
  OAI211_X1 U10127 ( .C1(n8806), .C2(n8674), .A(n8594), .B(n8593), .ZN(
        P2_U3207) );
  XNOR2_X1 U10128 ( .A(n8595), .B(n8596), .ZN(n8812) );
  XNOR2_X1 U10129 ( .A(n8597), .B(n8596), .ZN(n8600) );
  AOI222_X1 U10130 ( .A1(n8781), .A2(n8600), .B1(n8599), .B2(n8695), .C1(n8598), .C2(n8694), .ZN(n8807) );
  INV_X1 U10131 ( .A(n8807), .ZN(n8605) );
  INV_X1 U10132 ( .A(n8601), .ZN(n8602) );
  OAI22_X1 U10133 ( .A1(n8603), .A2(n8608), .B1(n8602), .B2(n8712), .ZN(n8604)
         );
  OAI21_X1 U10134 ( .B1(n8605), .B2(n8604), .A(n8700), .ZN(n8607) );
  NAND2_X1 U10135 ( .A1(n8708), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8606) );
  OAI211_X1 U10136 ( .C1(n8812), .C2(n8674), .A(n8607), .B(n8606), .ZN(
        P2_U3208) );
  INV_X1 U10137 ( .A(n8608), .ZN(n8612) );
  XOR2_X1 U10138 ( .A(n8615), .B(n8609), .Z(n8610) );
  OAI222_X1 U10139 ( .A1(n8718), .A2(n8637), .B1(n8720), .B2(n8611), .C1(n8635), .C2(n8610), .ZN(n8745) );
  AOI21_X1 U10140 ( .B1(n8612), .B2(n8744), .A(n8745), .ZN(n8618) );
  AOI22_X1 U10141 ( .A1(n8613), .A2(n8671), .B1(n8708), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8617) );
  XOR2_X1 U10142 ( .A(n8614), .B(n8615), .Z(n8746) );
  NAND2_X1 U10143 ( .A1(n8746), .A2(n8727), .ZN(n8616) );
  OAI211_X1 U10144 ( .C1(n8618), .C2(n8708), .A(n8617), .B(n8616), .ZN(
        P2_U3209) );
  XNOR2_X1 U10145 ( .A(n8619), .B(n8623), .ZN(n8620) );
  OAI222_X1 U10146 ( .A1(n8718), .A2(n8622), .B1(n8720), .B2(n8621), .C1(n8635), .C2(n8620), .ZN(n8748) );
  XNOR2_X1 U10147 ( .A(n8624), .B(n8623), .ZN(n8820) );
  AOI22_X1 U10148 ( .A1(n8708), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8625), .B2(
        n8671), .ZN(n8627) );
  NAND2_X1 U10149 ( .A1(n8749), .A2(n8702), .ZN(n8626) );
  OAI211_X1 U10150 ( .C1(n8820), .C2(n8674), .A(n8627), .B(n8626), .ZN(n8628)
         );
  AOI21_X1 U10151 ( .B1(n8748), .B2(n8700), .A(n8628), .ZN(n8629) );
  INV_X1 U10152 ( .A(n8629), .ZN(P2_U3210) );
  NAND3_X1 U10153 ( .A1(n8630), .A2(n8638), .A3(n8631), .ZN(n8632) );
  AND2_X1 U10154 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  OAI222_X1 U10155 ( .A1(n8720), .A2(n8637), .B1(n8718), .B2(n8636), .C1(n8635), .C2(n8634), .ZN(n8753) );
  NOR2_X1 U10156 ( .A1(n8639), .A2(n8638), .ZN(n8752) );
  INV_X1 U10157 ( .A(n8754), .ZN(n8640) );
  NOR3_X1 U10158 ( .A1(n8752), .A2(n8640), .A3(n8674), .ZN(n8645) );
  INV_X1 U10159 ( .A(n8641), .ZN(n8824) );
  AOI22_X1 U10160 ( .A1(n8708), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8671), .B2(
        n8642), .ZN(n8643) );
  OAI21_X1 U10161 ( .B1(n8824), .B2(n8714), .A(n8643), .ZN(n8644) );
  AOI211_X1 U10162 ( .C1(n8753), .C2(n8700), .A(n8645), .B(n8644), .ZN(n8647)
         );
  INV_X1 U10163 ( .A(n8647), .ZN(P2_U3211) );
  NAND2_X1 U10164 ( .A1(n8648), .A2(n8649), .ZN(n8651) );
  NAND2_X1 U10165 ( .A1(n8651), .A2(n8650), .ZN(n8653) );
  XNOR2_X1 U10166 ( .A(n8653), .B(n8652), .ZN(n8829) );
  INV_X1 U10167 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8660) );
  NAND3_X1 U10168 ( .A1(n8664), .A2(n8655), .A3(n8654), .ZN(n8656) );
  NAND2_X1 U10169 ( .A1(n8630), .A2(n8656), .ZN(n8659) );
  AOI222_X1 U10170 ( .A1(n8781), .A2(n8659), .B1(n8658), .B2(n8694), .C1(n8657), .C2(n8695), .ZN(n8825) );
  MUX2_X1 U10171 ( .A(n8660), .B(n8825), .S(n8700), .Z(n8663) );
  AOI22_X1 U10172 ( .A1(n5444), .A2(n8702), .B1(n8671), .B2(n8661), .ZN(n8662)
         );
  OAI211_X1 U10173 ( .C1(n8829), .C2(n8674), .A(n8663), .B(n8662), .ZN(
        P2_U3212) );
  XNOR2_X1 U10174 ( .A(n8648), .B(n8665), .ZN(n8835) );
  INV_X1 U10175 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8669) );
  OAI21_X1 U10176 ( .B1(n8666), .B2(n8665), .A(n8664), .ZN(n8668) );
  AOI222_X1 U10177 ( .A1(n8781), .A2(n8668), .B1(n8693), .B2(n8695), .C1(n8667), .C2(n8694), .ZN(n8830) );
  MUX2_X1 U10178 ( .A(n8669), .B(n8830), .S(n8700), .Z(n8673) );
  AOI22_X1 U10179 ( .A1(n8832), .A2(n8702), .B1(n8671), .B2(n8670), .ZN(n8672)
         );
  OAI211_X1 U10180 ( .C1(n8835), .C2(n8674), .A(n8673), .B(n8672), .ZN(
        P2_U3213) );
  XNOR2_X1 U10181 ( .A(n8676), .B(n8675), .ZN(n8677) );
  NAND2_X1 U10182 ( .A1(n8677), .A2(n8781), .ZN(n8681) );
  OAI22_X1 U10183 ( .A1(n8678), .A2(n8720), .B1(n8721), .B2(n8718), .ZN(n8679)
         );
  INV_X1 U10184 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U10185 ( .A1(n8681), .A2(n8680), .ZN(n8770) );
  INV_X1 U10186 ( .A(n8770), .ZN(n8690) );
  INV_X1 U10187 ( .A(n8682), .ZN(n8683) );
  OAI22_X1 U10188 ( .A1(n8700), .A2(n8684), .B1(n8683), .B2(n8712), .ZN(n8685)
         );
  AOI21_X1 U10189 ( .B1(n8686), .B2(n8702), .A(n8685), .ZN(n8689) );
  NAND2_X1 U10190 ( .A1(n4516), .A2(n8687), .ZN(n8766) );
  NAND3_X1 U10191 ( .A1(n8766), .A2(n8727), .A3(n8765), .ZN(n8688) );
  OAI211_X1 U10192 ( .C1(n8690), .C2(n8708), .A(n8689), .B(n8688), .ZN(
        P2_U3214) );
  XNOR2_X1 U10193 ( .A(n8691), .B(n5648), .ZN(n8692) );
  NAND2_X1 U10194 ( .A1(n8692), .A2(n8781), .ZN(n8698) );
  AOI22_X1 U10195 ( .A1(n8696), .A2(n8695), .B1(n8694), .B2(n8693), .ZN(n8697)
         );
  NAND2_X1 U10196 ( .A1(n8698), .A2(n8697), .ZN(n8776) );
  INV_X1 U10197 ( .A(n8776), .ZN(n8709) );
  OAI22_X1 U10198 ( .A1(n8700), .A2(n8461), .B1(n8699), .B2(n8712), .ZN(n8701)
         );
  AOI21_X1 U10199 ( .B1(n8703), .B2(n8702), .A(n8701), .ZN(n8707) );
  NAND2_X1 U10200 ( .A1(n8705), .A2(n8704), .ZN(n8771) );
  NAND3_X1 U10201 ( .A1(n8772), .A2(n8771), .A3(n8727), .ZN(n8706) );
  OAI211_X1 U10202 ( .C1(n8709), .C2(n8708), .A(n8707), .B(n8706), .ZN(
        P2_U3215) );
  XNOR2_X1 U10203 ( .A(n8710), .B(n8717), .ZN(n8842) );
  INV_X1 U10204 ( .A(n8842), .ZN(n8728) );
  INV_X1 U10205 ( .A(n8711), .ZN(n8840) );
  OAI22_X1 U10206 ( .A1(n8840), .A2(n8714), .B1(n8713), .B2(n8712), .ZN(n8726)
         );
  OAI211_X1 U10207 ( .C1(n8717), .C2(n8716), .A(n8715), .B(n8781), .ZN(n8724)
         );
  OAI22_X1 U10208 ( .A1(n8721), .A2(n8720), .B1(n8719), .B2(n8718), .ZN(n8722)
         );
  INV_X1 U10209 ( .A(n8722), .ZN(n8723) );
  NAND2_X1 U10210 ( .A1(n8724), .A2(n8723), .ZN(n8838) );
  MUX2_X1 U10211 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8838), .S(n8700), .Z(n8725) );
  AOI211_X1 U10212 ( .C1(n8728), .C2(n8727), .A(n8726), .B(n8725), .ZN(n8729)
         );
  INV_X1 U10213 ( .A(n8729), .ZN(P2_U3216) );
  NAND2_X1 U10214 ( .A1(n8730), .A2(n8762), .ZN(n8731) );
  NAND2_X1 U10215 ( .A1(n10325), .A2(n8790), .ZN(n8732) );
  OAI211_X1 U10216 ( .C1(n10325), .C2(n6619), .A(n8731), .B(n8732), .ZN(
        P2_U3490) );
  NAND2_X1 U10217 ( .A1(n6657), .A2(n8762), .ZN(n8733) );
  OAI211_X1 U10218 ( .C1(n10325), .C2(n9335), .A(n8733), .B(n8732), .ZN(
        P2_U3489) );
  AOI21_X1 U10219 ( .B1(n10308), .B2(n8735), .A(n8734), .ZN(n8797) );
  MUX2_X1 U10220 ( .A(n8736), .B(n8797), .S(n10325), .Z(n8737) );
  OAI21_X1 U10221 ( .B1(n8778), .B2(n8800), .A(n8737), .ZN(P2_U3486) );
  INV_X1 U10222 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8738) );
  MUX2_X1 U10223 ( .A(n8738), .B(n8801), .S(n10325), .Z(n8740) );
  NAND2_X1 U10224 ( .A1(n8803), .A2(n8762), .ZN(n8739) );
  OAI211_X1 U10225 ( .C1(n8806), .C2(n8778), .A(n8740), .B(n8739), .ZN(
        P2_U3485) );
  MUX2_X1 U10226 ( .A(n8741), .B(n8807), .S(n10325), .Z(n8743) );
  NAND2_X1 U10227 ( .A1(n8809), .A2(n8762), .ZN(n8742) );
  OAI211_X1 U10228 ( .C1(n8812), .C2(n8778), .A(n8743), .B(n8742), .ZN(
        P2_U3484) );
  INV_X1 U10229 ( .A(n8744), .ZN(n8816) );
  AOI21_X1 U10230 ( .B1(n8746), .B2(n10287), .A(n8745), .ZN(n8813) );
  MUX2_X1 U10231 ( .A(n9427), .B(n8813), .S(n10325), .Z(n8747) );
  OAI21_X1 U10232 ( .B1(n8816), .B2(n8777), .A(n8747), .ZN(P2_U3483) );
  AOI21_X1 U10233 ( .B1(n10308), .B2(n8749), .A(n8748), .ZN(n8817) );
  MUX2_X1 U10234 ( .A(n8750), .B(n8817), .S(n10325), .Z(n8751) );
  OAI21_X1 U10235 ( .B1(n8820), .B2(n8778), .A(n8751), .ZN(P2_U3482) );
  INV_X1 U10236 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8756) );
  NOR2_X1 U10237 ( .A1(n8752), .A2(n10303), .ZN(n8755) );
  AOI21_X1 U10238 ( .B1(n8755), .B2(n8754), .A(n8753), .ZN(n8821) );
  MUX2_X1 U10239 ( .A(n8756), .B(n8821), .S(n10325), .Z(n8757) );
  OAI21_X1 U10240 ( .B1(n8824), .B2(n8777), .A(n8757), .ZN(P2_U3481) );
  INV_X1 U10241 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8758) );
  MUX2_X1 U10242 ( .A(n8758), .B(n8825), .S(n10325), .Z(n8760) );
  NAND2_X1 U10243 ( .A1(n5444), .A2(n8762), .ZN(n8759) );
  OAI211_X1 U10244 ( .C1(n8778), .C2(n8829), .A(n8760), .B(n8759), .ZN(
        P2_U3480) );
  INV_X1 U10245 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U10246 ( .A(n8761), .B(n8830), .S(n10325), .Z(n8764) );
  NAND2_X1 U10247 ( .A1(n8832), .A2(n8762), .ZN(n8763) );
  OAI211_X1 U10248 ( .C1(n8835), .C2(n8778), .A(n8764), .B(n8763), .ZN(
        P2_U3479) );
  NAND3_X1 U10249 ( .A1(n8766), .A2(n8765), .A3(n10287), .ZN(n8767) );
  OAI21_X1 U10250 ( .B1(n8768), .B2(n10291), .A(n8767), .ZN(n8769) );
  MUX2_X1 U10251 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8836), .S(n10325), .Z(
        P2_U3478) );
  NAND3_X1 U10252 ( .A1(n8772), .A2(n10287), .A3(n8771), .ZN(n8773) );
  OAI21_X1 U10253 ( .B1(n8774), .B2(n10291), .A(n8773), .ZN(n8775) );
  MUX2_X1 U10254 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8837), .S(n10325), .Z(
        P2_U3477) );
  MUX2_X1 U10255 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8838), .S(n10325), .Z(
        n8780) );
  OAI22_X1 U10256 ( .A1(n8842), .A2(n8778), .B1(n8840), .B2(n8777), .ZN(n8779)
         );
  OR2_X1 U10257 ( .A1(n8780), .A2(n8779), .ZN(P2_U3476) );
  NOR2_X1 U10258 ( .A1(n10287), .A2(n8781), .ZN(n8782) );
  OR2_X1 U10259 ( .A1(n8783), .A2(n8782), .ZN(n8788) );
  OR2_X1 U10260 ( .A1(n8784), .A2(n10291), .ZN(n8785) );
  AND2_X1 U10261 ( .A1(n8786), .A2(n8785), .ZN(n8787) );
  AND2_X1 U10262 ( .A1(n8788), .A2(n8787), .ZN(n10251) );
  INV_X1 U10263 ( .A(n10251), .ZN(n8789) );
  MUX2_X1 U10264 ( .A(n8789), .B(P2_REG1_REG_0__SCAN_IN), .S(n10323), .Z(
        P2_U3459) );
  INV_X1 U10265 ( .A(n8790), .ZN(n8791) );
  NOR2_X1 U10266 ( .A1(n10311), .A2(n8791), .ZN(n8794) );
  AOI21_X1 U10267 ( .B1(n10311), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8794), .ZN(
        n8792) );
  OAI21_X1 U10268 ( .B1(n8793), .B2(n8839), .A(n8792), .ZN(P2_U3458) );
  NAND2_X1 U10269 ( .A1(n6657), .A2(n6371), .ZN(n8796) );
  INV_X1 U10270 ( .A(n8794), .ZN(n8795) );
  OAI211_X1 U10271 ( .C1(n6357), .C2(n10309), .A(n8796), .B(n8795), .ZN(
        P2_U3457) );
  INV_X1 U10272 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8798) );
  MUX2_X1 U10273 ( .A(n8798), .B(n8797), .S(n10309), .Z(n8799) );
  OAI21_X1 U10274 ( .B1(n8800), .B2(n8841), .A(n8799), .ZN(P2_U3454) );
  INV_X1 U10275 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10276 ( .A(n8802), .B(n8801), .S(n10309), .Z(n8805) );
  NAND2_X1 U10277 ( .A1(n8803), .A2(n6371), .ZN(n8804) );
  OAI211_X1 U10278 ( .C1(n8806), .C2(n8841), .A(n8805), .B(n8804), .ZN(
        P2_U3453) );
  INV_X1 U10279 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8808) );
  MUX2_X1 U10280 ( .A(n8808), .B(n8807), .S(n10309), .Z(n8811) );
  NAND2_X1 U10281 ( .A1(n8809), .A2(n6371), .ZN(n8810) );
  OAI211_X1 U10282 ( .C1(n8812), .C2(n8841), .A(n8811), .B(n8810), .ZN(
        P2_U3452) );
  INV_X1 U10283 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8814) );
  MUX2_X1 U10284 ( .A(n8814), .B(n8813), .S(n10309), .Z(n8815) );
  OAI21_X1 U10285 ( .B1(n8816), .B2(n8839), .A(n8815), .ZN(P2_U3451) );
  INV_X1 U10286 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8818) );
  MUX2_X1 U10287 ( .A(n8818), .B(n8817), .S(n10309), .Z(n8819) );
  OAI21_X1 U10288 ( .B1(n8820), .B2(n8841), .A(n8819), .ZN(P2_U3450) );
  INV_X1 U10289 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8822) );
  MUX2_X1 U10290 ( .A(n8822), .B(n8821), .S(n10309), .Z(n8823) );
  OAI21_X1 U10291 ( .B1(n8824), .B2(n8839), .A(n8823), .ZN(P2_U3449) );
  INV_X1 U10292 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8826) );
  MUX2_X1 U10293 ( .A(n8826), .B(n8825), .S(n10309), .Z(n8828) );
  NAND2_X1 U10294 ( .A1(n5444), .A2(n6371), .ZN(n8827) );
  OAI211_X1 U10295 ( .C1(n8829), .C2(n8841), .A(n8828), .B(n8827), .ZN(
        P2_U3448) );
  INV_X1 U10296 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8831) );
  MUX2_X1 U10297 ( .A(n8831), .B(n8830), .S(n10309), .Z(n8834) );
  NAND2_X1 U10298 ( .A1(n8832), .A2(n6371), .ZN(n8833) );
  OAI211_X1 U10299 ( .C1(n8835), .C2(n8841), .A(n8834), .B(n8833), .ZN(
        P2_U3447) );
  MUX2_X1 U10300 ( .A(n8836), .B(P2_REG0_REG_19__SCAN_IN), .S(n10311), .Z(
        P2_U3446) );
  MUX2_X1 U10301 ( .A(n8837), .B(P2_REG0_REG_18__SCAN_IN), .S(n10311), .Z(
        P2_U3444) );
  MUX2_X1 U10302 ( .A(n8838), .B(P2_REG0_REG_17__SCAN_IN), .S(n10311), .Z(
        n8844) );
  OAI22_X1 U10303 ( .A1(n8842), .A2(n8841), .B1(n8840), .B2(n8839), .ZN(n8843)
         );
  OR2_X1 U10304 ( .A1(n8844), .A2(n8843), .ZN(P2_U3441) );
  MUX2_X1 U10305 ( .A(n8846), .B(P2_D_REG_1__SCAN_IN), .S(n8845), .Z(P2_U3377)
         );
  OAI222_X1 U10306 ( .A1(n8847), .A2(P2_U3151), .B1(n8851), .B2(n8850), .C1(
        n8849), .C2(n8848), .ZN(P2_U3265) );
  INV_X1 U10307 ( .A(n8852), .ZN(n8853) );
  MUX2_X1 U10308 ( .A(n8853), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U10309 ( .B1(n8967), .B2(n8855), .A(n8854), .ZN(n8856) );
  OAI21_X1 U10310 ( .B1(n8857), .B2(n8856), .A(n8968), .ZN(n8863) );
  OR2_X1 U10311 ( .A1(n9167), .A2(n8972), .ZN(n8859) );
  OR2_X1 U10312 ( .A1(n8994), .A2(n9140), .ZN(n8858) );
  NAND2_X1 U10313 ( .A1(n8859), .A2(n8858), .ZN(n9199) );
  AOI22_X1 U10314 ( .A1(n4438), .A2(n9199), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n8860) );
  OAI21_X1 U10315 ( .B1(n9796), .B2(n9204), .A(n8860), .ZN(n8861) );
  AOI21_X1 U10316 ( .B1(n9640), .B2(n8988), .A(n8861), .ZN(n8862) );
  NAND2_X1 U10317 ( .A1(n8863), .A2(n8862), .ZN(P1_U3214) );
  INV_X1 U10318 ( .A(n8864), .ZN(n8866) );
  NOR3_X1 U10319 ( .A1(n4454), .A2(n8866), .A3(n8865), .ZN(n8869) );
  INV_X1 U10320 ( .A(n8867), .ZN(n8868) );
  OAI21_X1 U10321 ( .B1(n8869), .B2(n8868), .A(n8968), .ZN(n8874) );
  OAI22_X1 U10322 ( .A1(n8899), .A2(n8972), .B1(n8995), .B2(n9140), .ZN(n9569)
         );
  INV_X1 U10323 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8870) );
  OAI22_X1 U10324 ( .A1(n8871), .A2(n9796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8870), .ZN(n8872) );
  AOI21_X1 U10325 ( .B1(n9569), .B2(n4438), .A(n8872), .ZN(n8873) );
  OAI211_X1 U10326 ( .C1(n9564), .C2(n9786), .A(n8874), .B(n8873), .ZN(
        P1_U3216) );
  XNOR2_X1 U10327 ( .A(n8876), .B(n8875), .ZN(n8877) );
  XNOR2_X1 U10328 ( .A(n8878), .B(n8877), .ZN(n8884) );
  NAND2_X1 U10329 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U10330 ( .A1(n8925), .A2(n8879), .ZN(n8880) );
  OAI211_X1 U10331 ( .C1(n8881), .C2(n8927), .A(n9110), .B(n8880), .ZN(n8882)
         );
  AOI21_X1 U10332 ( .B1(n9146), .B2(n8988), .A(n8882), .ZN(n8883) );
  OAI21_X1 U10333 ( .B1(n8884), .B2(n9791), .A(n8883), .ZN(P1_U3219) );
  OAI21_X1 U10334 ( .B1(n8887), .B2(n8886), .A(n8885), .ZN(n8888) );
  NAND2_X1 U10335 ( .A1(n8888), .A2(n8968), .ZN(n8893) );
  OAI22_X1 U10336 ( .A1(n8995), .A2(n8972), .B1(n8889), .B2(n9140), .ZN(n9596)
         );
  OAI22_X1 U10337 ( .A1(n9602), .A2(n9796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8890), .ZN(n8891) );
  AOI21_X1 U10338 ( .B1(n9596), .B2(n4438), .A(n8891), .ZN(n8892) );
  OAI211_X1 U10339 ( .C1(n8894), .C2(n9786), .A(n8893), .B(n8892), .ZN(
        P1_U3223) );
  OAI21_X1 U10340 ( .B1(n8897), .B2(n8895), .A(n8896), .ZN(n8898) );
  NAND2_X1 U10341 ( .A1(n8898), .A2(n8968), .ZN(n8902) );
  OAI22_X1 U10342 ( .A1(n8899), .A2(n9140), .B1(n8994), .B2(n8972), .ZN(n9234)
         );
  INV_X1 U10343 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9436) );
  OAI22_X1 U10344 ( .A1(n9796), .A2(n9227), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9436), .ZN(n8900) );
  AOI21_X1 U10345 ( .B1(n9234), .B2(n4438), .A(n8900), .ZN(n8901) );
  OAI211_X1 U10346 ( .C1(n9230), .C2(n9786), .A(n8902), .B(n8901), .ZN(
        P1_U3225) );
  XNOR2_X1 U10347 ( .A(n8903), .B(n8904), .ZN(n8982) );
  NOR2_X1 U10348 ( .A1(n8982), .A2(n8981), .ZN(n8980) );
  AOI21_X1 U10349 ( .B1(n8904), .B2(n8903), .A(n8980), .ZN(n8908) );
  XNOR2_X1 U10350 ( .A(n8906), .B(n8905), .ZN(n8907) );
  XNOR2_X1 U10351 ( .A(n8908), .B(n8907), .ZN(n8914) );
  NAND2_X1 U10352 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9058) );
  NAND2_X1 U10353 ( .A1(n8925), .A2(n8909), .ZN(n8910) );
  OAI211_X1 U10354 ( .C1(n8911), .C2(n8927), .A(n9058), .B(n8910), .ZN(n8912)
         );
  AOI21_X1 U10355 ( .B1(n9763), .B2(n8988), .A(n8912), .ZN(n8913) );
  OAI21_X1 U10356 ( .B1(n8914), .B2(n9791), .A(n8913), .ZN(P1_U3226) );
  XOR2_X1 U10357 ( .A(n8915), .B(n8916), .Z(n8923) );
  NAND2_X1 U10358 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9088) );
  NAND2_X1 U10359 ( .A1(n8925), .A2(n8917), .ZN(n8918) );
  OAI211_X1 U10360 ( .C1(n8919), .C2(n8927), .A(n9088), .B(n8918), .ZN(n8920)
         );
  AOI21_X1 U10361 ( .B1(n8921), .B2(n8988), .A(n8920), .ZN(n8922) );
  OAI21_X1 U10362 ( .B1(n8923), .B2(n9791), .A(n8922), .ZN(P1_U3228) );
  INV_X1 U10363 ( .A(n8947), .ZN(n9155) );
  INV_X1 U10364 ( .A(n8971), .ZN(n9159) );
  AOI22_X1 U10365 ( .A1(n9155), .A2(n8948), .B1(n8924), .B2(n9159), .ZN(n9542)
         );
  AOI22_X1 U10366 ( .A1(n9547), .A2(n8925), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8926) );
  OAI21_X1 U10367 ( .B1(n9542), .B2(n8927), .A(n8926), .ZN(n8933) );
  NAND3_X1 U10368 ( .A1(n8867), .A2(n8930), .A3(n4893), .ZN(n8931) );
  AOI21_X1 U10369 ( .B1(n8928), .B2(n8931), .A(n9791), .ZN(n8932) );
  AOI211_X1 U10370 ( .C1(n9655), .C2(n8988), .A(n8933), .B(n8932), .ZN(n8934)
         );
  INV_X1 U10371 ( .A(n8934), .ZN(P1_U3229) );
  AOI21_X1 U10372 ( .B1(n8935), .B2(n8936), .A(n4487), .ZN(n8944) );
  OAI22_X1 U10373 ( .A1(n8938), .A2(n8972), .B1(n8937), .B2(n9140), .ZN(n9618)
         );
  INV_X1 U10374 ( .A(n9613), .ZN(n8940) );
  OAI22_X1 U10375 ( .A1(n8940), .A2(n9796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8939), .ZN(n8942) );
  NOR2_X1 U10376 ( .A1(n9615), .A2(n9786), .ZN(n8941) );
  AOI211_X1 U10377 ( .C1(n4438), .C2(n9618), .A(n8942), .B(n8941), .ZN(n8943)
         );
  OAI21_X1 U10378 ( .B1(n8944), .B2(n9791), .A(n8943), .ZN(P1_U3233) );
  AOI21_X1 U10379 ( .B1(n8946), .B2(n8945), .A(n4454), .ZN(n8955) );
  OR2_X1 U10380 ( .A1(n8947), .A2(n8972), .ZN(n8950) );
  NAND2_X1 U10381 ( .A1(n9151), .A2(n8948), .ZN(n8949) );
  NAND2_X1 U10382 ( .A1(n8950), .A2(n8949), .ZN(n9580) );
  INV_X1 U10383 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9410) );
  OAI22_X1 U10384 ( .A1(n9582), .A2(n9796), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9410), .ZN(n8953) );
  NOR2_X1 U10385 ( .A1(n8951), .A2(n9786), .ZN(n8952) );
  AOI211_X1 U10386 ( .C1(n4438), .C2(n9580), .A(n8953), .B(n8952), .ZN(n8954)
         );
  OAI21_X1 U10387 ( .B1(n8955), .B2(n9791), .A(n8954), .ZN(P1_U3235) );
  XNOR2_X1 U10388 ( .A(n8958), .B(n8957), .ZN(n8959) );
  XNOR2_X1 U10389 ( .A(n8956), .B(n8959), .ZN(n8966) );
  OAI22_X1 U10390 ( .A1(n9796), .A2(n8961), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8960), .ZN(n8963) );
  NOR2_X1 U10391 ( .A1(n9753), .A2(n9786), .ZN(n8962) );
  AOI211_X1 U10392 ( .C1(n4438), .C2(n8964), .A(n8963), .B(n8962), .ZN(n8965)
         );
  OAI21_X1 U10393 ( .B1(n8966), .B2(n9791), .A(n8965), .ZN(P1_U3238) );
  NAND2_X1 U10394 ( .A1(n8967), .A2(n8968), .ZN(n8979) );
  AOI21_X1 U10395 ( .B1(n8896), .B2(n8970), .A(n8969), .ZN(n8978) );
  OR2_X1 U10396 ( .A1(n8971), .A2(n9140), .ZN(n8974) );
  OR2_X1 U10397 ( .A1(n8993), .A2(n8972), .ZN(n8973) );
  NAND2_X1 U10398 ( .A1(n8974), .A2(n8973), .ZN(n9211) );
  AOI22_X1 U10399 ( .A1(n4438), .A2(n9211), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8975) );
  OAI21_X1 U10400 ( .B1(n9796), .B2(n9219), .A(n8975), .ZN(n8976) );
  AOI21_X1 U10401 ( .B1(n9643), .B2(n8988), .A(n8976), .ZN(n8977) );
  OAI21_X1 U10402 ( .B1(n8979), .B2(n8978), .A(n8977), .ZN(P1_U3240) );
  AOI21_X1 U10403 ( .B1(n8982), .B2(n8981), .A(n8980), .ZN(n8991) );
  AOI22_X1 U10404 ( .A1(n8984), .A2(n4438), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n8985) );
  OAI21_X1 U10405 ( .B1(n8986), .B2(n9796), .A(n8985), .ZN(n8987) );
  AOI21_X1 U10406 ( .B1(n8989), .B2(n8988), .A(n8987), .ZN(n8990) );
  OAI21_X1 U10407 ( .B1(n8991), .B2(n9791), .A(n8990), .ZN(P1_U3241) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8992), .S(P1_U3973), .Z(
        P1_U3584) );
  INV_X1 U10409 ( .A(n8993), .ZN(n9165) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9165), .S(P1_U3973), .Z(
        P1_U3581) );
  INV_X1 U10411 ( .A(n8994), .ZN(n9163) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9163), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9159), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9156), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9155), .S(P1_U3973), .Z(
        P1_U3577) );
  INV_X1 U10416 ( .A(n8995), .ZN(n9153) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9153), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9151), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9149), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9145), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n8996), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n8997), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n8998), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8999), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9000), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9001), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9002), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9003), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10429 ( .A(n9004), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9008), .Z(
        P1_U3561) );
  MUX2_X1 U10430 ( .A(n9005), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9008), .Z(
        P1_U3558) );
  MUX2_X1 U10431 ( .A(n9006), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9008), .Z(
        P1_U3557) );
  MUX2_X1 U10432 ( .A(n9007), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9008), .Z(
        P1_U3556) );
  MUX2_X1 U10433 ( .A(n4440), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9008), .Z(
        P1_U3555) );
  NAND3_X1 U10434 ( .A1(n9010), .A2(n9009), .A3(n4451), .ZN(n9016) );
  INV_X1 U10435 ( .A(n9802), .ZN(n9011) );
  AOI22_X1 U10436 ( .A1(n9014), .A2(n9013), .B1(n9012), .B2(n9011), .ZN(n9015)
         );
  NAND3_X1 U10437 ( .A1(n9016), .A2(P1_U3973), .A3(n9015), .ZN(n9823) );
  AOI22_X1 U10438 ( .A1(n9811), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n9034) );
  INV_X1 U10439 ( .A(n9017), .ZN(n9020) );
  INV_X1 U10440 ( .A(n9018), .ZN(n9019) );
  NAND2_X1 U10441 ( .A1(n9020), .A2(n9019), .ZN(n9021) );
  NAND3_X1 U10442 ( .A1(n9913), .A2(n9022), .A3(n9021), .ZN(n9030) );
  INV_X1 U10443 ( .A(n9023), .ZN(n9026) );
  INV_X1 U10444 ( .A(n9024), .ZN(n9025) );
  NAND2_X1 U10445 ( .A1(n9026), .A2(n9025), .ZN(n9027) );
  NAND3_X1 U10446 ( .A1(n9861), .A2(n9028), .A3(n9027), .ZN(n9029) );
  AND2_X1 U10447 ( .A1(n9030), .A2(n9029), .ZN(n9033) );
  INV_X1 U10448 ( .A(n9821), .ZN(n9921) );
  NAND2_X1 U10449 ( .A1(n9921), .A2(n9031), .ZN(n9032) );
  NAND4_X1 U10450 ( .A1(n9823), .A2(n9034), .A3(n9033), .A4(n9032), .ZN(
        P1_U3245) );
  INV_X1 U10451 ( .A(n9811), .ZN(n9924) );
  INV_X1 U10452 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9036) );
  NAND2_X1 U10453 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9035) );
  OAI21_X1 U10454 ( .B1(n9924), .B2(n9036), .A(n9035), .ZN(n9037) );
  AOI21_X1 U10455 ( .B1(n9038), .B2(n9921), .A(n9037), .ZN(n9047) );
  OAI211_X1 U10456 ( .C1(n9041), .C2(n9040), .A(n9861), .B(n9039), .ZN(n9046)
         );
  OAI211_X1 U10457 ( .C1(n9044), .C2(n9043), .A(n9913), .B(n9042), .ZN(n9045)
         );
  NAND3_X1 U10458 ( .A1(n9047), .A2(n9046), .A3(n9045), .ZN(P1_U3246) );
  OAI21_X1 U10459 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n9062), .A(n9048), .ZN(
        n9877) );
  INV_X1 U10460 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9049) );
  MUX2_X1 U10461 ( .A(n9049), .B(P1_REG1_REG_13__SCAN_IN), .S(n9881), .Z(n9878) );
  NOR2_X1 U10462 ( .A1(n9877), .A2(n9878), .ZN(n9876) );
  AOI21_X1 U10463 ( .B1(n9881), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9876), .ZN(
        n9890) );
  MUX2_X1 U10464 ( .A(n9050), .B(P1_REG1_REG_14__SCAN_IN), .S(n9893), .Z(n9889) );
  NOR2_X1 U10465 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  AOI21_X1 U10466 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n9893), .A(n9888), .ZN(
        n9051) );
  NOR2_X1 U10467 ( .A1(n9051), .A2(n9066), .ZN(n9052) );
  INV_X1 U10468 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9898) );
  XNOR2_X1 U10469 ( .A(n9066), .B(n9051), .ZN(n9899) );
  NOR2_X1 U10470 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  NOR2_X1 U10471 ( .A1(n9052), .A2(n9897), .ZN(n9056) );
  NOR2_X1 U10472 ( .A1(n9059), .A2(n9053), .ZN(n9054) );
  AOI21_X1 U10473 ( .B1(n9053), .B2(n9059), .A(n9054), .ZN(n9055) );
  NAND2_X1 U10474 ( .A1(n9056), .A2(n9055), .ZN(n9083) );
  OAI21_X1 U10475 ( .B1(n9056), .B2(n9055), .A(n9083), .ZN(n9074) );
  NAND2_X1 U10476 ( .A1(n9811), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n9057) );
  OAI211_X1 U10477 ( .C1(n9821), .C2(n9059), .A(n9058), .B(n9057), .ZN(n9073)
         );
  AOI22_X1 U10478 ( .A1(n9881), .A2(n6025), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n9060), .ZN(n9875) );
  OAI22_X1 U10479 ( .A1(n9064), .A2(n9063), .B1(P1_REG2_REG_12__SCAN_IN), .B2(
        n9062), .ZN(n9874) );
  NOR2_X1 U10480 ( .A1(n9875), .A2(n9874), .ZN(n9873) );
  NAND2_X1 U10481 ( .A1(n9893), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9065) );
  OAI21_X1 U10482 ( .B1(n9893), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9065), .ZN(
        n9886) );
  NOR2_X1 U10483 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  NOR2_X1 U10484 ( .A1(n7912), .A2(n9902), .ZN(n9901) );
  NOR2_X1 U10485 ( .A1(n9068), .A2(n9901), .ZN(n9071) );
  XNOR2_X1 U10486 ( .A(n9084), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9070) );
  INV_X1 U10487 ( .A(n9078), .ZN(n9069) );
  AOI211_X1 U10488 ( .C1(n9071), .C2(n9070), .A(n9900), .B(n9069), .ZN(n9072)
         );
  AOI211_X1 U10489 ( .C1(n9861), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9075)
         );
  INV_X1 U10490 ( .A(n9075), .ZN(P1_U3259) );
  OR2_X1 U10491 ( .A1(n9100), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U10492 ( .A1(n9100), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9076) );
  AND2_X1 U10493 ( .A1(n9094), .A2(n9076), .ZN(n9079) );
  NAND2_X1 U10494 ( .A1(n9084), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9077) );
  OAI21_X1 U10495 ( .B1(n9079), .B2(n4520), .A(n9095), .ZN(n9080) );
  NAND2_X1 U10496 ( .A1(n9080), .A2(n9913), .ZN(n9093) );
  NOR2_X1 U10497 ( .A1(n9089), .A2(n9081), .ZN(n9082) );
  AOI21_X1 U10498 ( .B1(n9081), .B2(n9089), .A(n9082), .ZN(n9086) );
  OAI21_X1 U10499 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(n9084), .A(n9083), .ZN(
        n9085) );
  NAND2_X1 U10500 ( .A1(n9085), .A2(n9086), .ZN(n9099) );
  OAI21_X1 U10501 ( .B1(n9086), .B2(n9085), .A(n9099), .ZN(n9091) );
  NAND2_X1 U10502 ( .A1(n9811), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9087) );
  OAI211_X1 U10503 ( .C1(n9821), .C2(n9089), .A(n9088), .B(n9087), .ZN(n9090)
         );
  AOI21_X1 U10504 ( .B1(n9091), .B2(n9861), .A(n9090), .ZN(n9092) );
  NAND2_X1 U10505 ( .A1(n9093), .A2(n9092), .ZN(P1_U3260) );
  INV_X1 U10506 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U10507 ( .A1(n9920), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9097) );
  OR2_X1 U10508 ( .A1(n9920), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9096) );
  AND2_X1 U10509 ( .A1(n9097), .A2(n9096), .ZN(n9915) );
  NAND2_X1 U10510 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  NAND2_X1 U10511 ( .A1(n9914), .A2(n9097), .ZN(n9098) );
  XNOR2_X1 U10512 ( .A(n9098), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9107) );
  INV_X1 U10513 ( .A(n9107), .ZN(n9104) );
  OAI21_X1 U10514 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9100), .A(n9099), .ZN(
        n9911) );
  NOR2_X1 U10515 ( .A1(n9920), .A2(n9101), .ZN(n9102) );
  AOI21_X1 U10516 ( .B1(n9920), .B2(n9101), .A(n9102), .ZN(n9912) );
  NOR2_X1 U10517 ( .A1(n9911), .A2(n9912), .ZN(n9909) );
  AOI21_X1 U10518 ( .B1(n9920), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9909), .ZN(
        n9103) );
  XNOR2_X1 U10519 ( .A(n9103), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9105) );
  AOI22_X1 U10520 ( .A1(n9104), .A2(n9913), .B1(n9861), .B2(n9105), .ZN(n9109)
         );
  OAI21_X1 U10521 ( .B1(n9105), .B2(n9910), .A(n9821), .ZN(n9106) );
  AOI21_X1 U10522 ( .B1(n9107), .B2(n9913), .A(n9106), .ZN(n9108) );
  MUX2_X1 U10523 ( .A(n9109), .B(n9108), .S(n6376), .Z(n9111) );
  OAI211_X1 U10524 ( .C1(n9112), .C2(n9924), .A(n9111), .B(n9110), .ZN(
        P1_U3262) );
  XNOR2_X1 U10525 ( .A(n9113), .B(n6138), .ZN(n9114) );
  NAND2_X1 U10526 ( .A1(n9114), .A2(n9975), .ZN(n9625) );
  NOR2_X1 U10527 ( .A1(n9588), .A2(n9115), .ZN(n9116) );
  NOR2_X1 U10528 ( .A1(n9973), .A2(n9624), .ZN(n9119) );
  AOI211_X1 U10529 ( .C1(n6138), .C2(n9599), .A(n9116), .B(n9119), .ZN(n9117)
         );
  OAI21_X1 U10530 ( .B1(n9625), .B2(n9585), .A(n9117), .ZN(P1_U3263) );
  NOR2_X1 U10531 ( .A1(n4636), .A2(n9970), .ZN(n9118) );
  AOI211_X1 U10532 ( .C1(n9968), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9119), .B(
        n9118), .ZN(n9120) );
  OAI21_X1 U10533 ( .B1(n9585), .B2(n9121), .A(n9120), .ZN(P1_U3264) );
  NAND2_X1 U10534 ( .A1(n9567), .A2(n9565), .ZN(n9126) );
  OAI21_X1 U10535 ( .B1(n9577), .B2(n9126), .A(n9125), .ZN(n9539) );
  NOR2_X1 U10536 ( .A1(n9539), .A2(n4622), .ZN(n9543) );
  INV_X1 U10537 ( .A(n9127), .ZN(n9128) );
  NOR2_X1 U10538 ( .A1(n9543), .A2(n9128), .ZN(n9233) );
  INV_X1 U10539 ( .A(n9130), .ZN(n9131) );
  INV_X1 U10540 ( .A(n9132), .ZN(n9133) );
  OAI21_X1 U10541 ( .B1(n9180), .B2(n9188), .A(n9136), .ZN(n9137) );
  XNOR2_X1 U10542 ( .A(n9137), .B(n4638), .ZN(n9142) );
  OAI22_X1 U10543 ( .A1(n9167), .A2(n9140), .B1(n9139), .B2(n9138), .ZN(n9141)
         );
  NOR2_X1 U10544 ( .A1(n9146), .A2(n9145), .ZN(n9143) );
  NAND2_X1 U10545 ( .A1(n9146), .A2(n9145), .ZN(n9147) );
  OR2_X1 U10546 ( .A1(n9674), .A2(n9149), .ZN(n9150) );
  INV_X1 U10547 ( .A(n9594), .ZN(n9604) );
  NAND2_X1 U10548 ( .A1(n9605), .A2(n9604), .ZN(n9603) );
  OR2_X1 U10549 ( .A1(n9669), .A2(n9151), .ZN(n9152) );
  NAND2_X1 U10550 ( .A1(n9603), .A2(n9152), .ZN(n9575) );
  OR2_X1 U10551 ( .A1(n9664), .A2(n9153), .ZN(n9154) );
  INV_X1 U10552 ( .A(n9567), .ZN(n9556) );
  NOR2_X1 U10553 ( .A1(n9655), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U10554 ( .A1(n9655), .A2(n9156), .ZN(n9157) );
  OR2_X1 U10555 ( .A1(n9649), .A2(n9159), .ZN(n9160) );
  NAND2_X1 U10556 ( .A1(n9643), .A2(n9163), .ZN(n9164) );
  OR2_X1 U10557 ( .A1(n9640), .A2(n9165), .ZN(n9166) );
  NAND2_X1 U10558 ( .A1(n9968), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9170) );
  OAI21_X1 U10559 ( .B1(n9949), .B2(n9171), .A(n9170), .ZN(n9172) );
  AOI21_X1 U10560 ( .B1(n5918), .B2(n9599), .A(n9172), .ZN(n9177) );
  AOI21_X1 U10561 ( .B1(n5918), .B2(n9183), .A(n9612), .ZN(n9175) );
  NAND2_X1 U10562 ( .A1(n9628), .A2(n9978), .ZN(n9176) );
  OAI211_X1 U10563 ( .C1(n9631), .C2(n9623), .A(n9177), .B(n9176), .ZN(n9178)
         );
  INV_X1 U10564 ( .A(n9178), .ZN(n9179) );
  OAI21_X1 U10565 ( .B1(n9630), .B2(n9973), .A(n9179), .ZN(P1_U3356) );
  XNOR2_X1 U10566 ( .A(n9180), .B(n9188), .ZN(n9182) );
  AOI21_X1 U10567 ( .B1(n9182), .B2(n9947), .A(n9181), .ZN(n9637) );
  AOI211_X1 U10568 ( .C1(n9633), .C2(n9202), .A(n9612), .B(n9173), .ZN(n9632)
         );
  NOR2_X1 U10569 ( .A1(n4674), .A2(n9970), .ZN(n9187) );
  OAI22_X1 U10570 ( .A1(n9588), .A2(n9185), .B1(n9184), .B2(n9949), .ZN(n9186)
         );
  AOI211_X1 U10571 ( .C1(n9632), .C2(n9978), .A(n9187), .B(n9186), .ZN(n9192)
         );
  NAND3_X1 U10572 ( .A1(n9634), .A2(n9957), .A3(n9190), .ZN(n9191) );
  OAI211_X1 U10573 ( .C1(n9637), .C2(n9973), .A(n9192), .B(n9191), .ZN(
        P1_U3265) );
  OAI21_X1 U10574 ( .B1(n9194), .B2(n9197), .A(n9193), .ZN(n9195) );
  INV_X1 U10575 ( .A(n9195), .ZN(n9641) );
  AOI21_X1 U10576 ( .B1(n9198), .B2(n9197), .A(n9196), .ZN(n9201) );
  INV_X1 U10577 ( .A(n9199), .ZN(n9200) );
  NAND2_X1 U10578 ( .A1(n9638), .A2(n9588), .ZN(n9209) );
  AOI211_X1 U10579 ( .C1(n9640), .C2(n9213), .A(n9612), .B(n4676), .ZN(n9639)
         );
  INV_X1 U10580 ( .A(n9640), .ZN(n9203) );
  NOR2_X1 U10581 ( .A1(n9203), .A2(n9970), .ZN(n9207) );
  OAI22_X1 U10582 ( .A1(n9588), .A2(n9205), .B1(n9204), .B2(n9949), .ZN(n9206)
         );
  AOI211_X1 U10583 ( .C1(n9639), .C2(n9978), .A(n9207), .B(n9206), .ZN(n9208)
         );
  OAI211_X1 U10584 ( .C1(n9641), .C2(n9623), .A(n9209), .B(n9208), .ZN(
        P1_U3266) );
  XNOR2_X1 U10585 ( .A(n9210), .B(n9216), .ZN(n9212) );
  AOI21_X1 U10586 ( .B1(n9212), .B2(n9947), .A(n9211), .ZN(n9647) );
  OAI211_X1 U10587 ( .C1(n9214), .C2(n9226), .A(n9975), .B(n9213), .ZN(n9645)
         );
  NAND2_X1 U10588 ( .A1(n9217), .A2(n9216), .ZN(n9642) );
  NAND3_X1 U10589 ( .A1(n9215), .A2(n9642), .A3(n9957), .ZN(n9222) );
  NAND2_X1 U10590 ( .A1(n9968), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9218) );
  OAI21_X1 U10591 ( .B1(n9949), .B2(n9219), .A(n9218), .ZN(n9220) );
  AOI21_X1 U10592 ( .B1(n9643), .B2(n9599), .A(n9220), .ZN(n9221) );
  OAI211_X1 U10593 ( .C1(n9645), .C2(n9585), .A(n9222), .B(n9221), .ZN(n9223)
         );
  INV_X1 U10594 ( .A(n9223), .ZN(n9224) );
  OAI21_X1 U10595 ( .B1(n9647), .B2(n9973), .A(n9224), .ZN(P1_U3267) );
  XNOR2_X1 U10596 ( .A(n9225), .B(n9232), .ZN(n9652) );
  AOI211_X1 U10597 ( .C1(n9649), .C2(n9545), .A(n9612), .B(n9226), .ZN(n9648)
         );
  INV_X1 U10598 ( .A(n9227), .ZN(n9228) );
  AOI22_X1 U10599 ( .A1(n9968), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9228), .B2(
        n9967), .ZN(n9229) );
  OAI21_X1 U10600 ( .B1(n9230), .B2(n9970), .A(n9229), .ZN(n9237) );
  AOI211_X1 U10601 ( .C1(n9233), .C2(n9232), .A(n9963), .B(n9231), .ZN(n9235)
         );
  NOR2_X1 U10602 ( .A1(n9235), .A2(n9234), .ZN(n9651) );
  NOR2_X1 U10603 ( .A1(n9651), .A2(n9973), .ZN(n9236) );
  AOI211_X1 U10604 ( .C1(n9648), .C2(n9978), .A(n9237), .B(n9236), .ZN(n9238)
         );
  OAI21_X1 U10605 ( .B1(n9623), .B2(n9652), .A(n9238), .ZN(P1_U3268) );
  NAND2_X1 U10606 ( .A1(keyinput121), .A2(keyinput14), .ZN(n9239) );
  NOR3_X1 U10607 ( .A1(keyinput9), .A2(keyinput50), .A3(n9239), .ZN(n9240) );
  NAND3_X1 U10608 ( .A1(keyinput34), .A2(keyinput72), .A3(n9240), .ZN(n9252)
         );
  NOR2_X1 U10609 ( .A1(keyinput53), .A2(keyinput104), .ZN(n9241) );
  NAND3_X1 U10610 ( .A1(keyinput101), .A2(keyinput85), .A3(n9241), .ZN(n9242)
         );
  NOR3_X1 U10611 ( .A1(keyinput39), .A2(keyinput118), .A3(n9242), .ZN(n9250)
         );
  NOR3_X1 U10612 ( .A1(keyinput35), .A2(keyinput81), .A3(keyinput80), .ZN(
        n9243) );
  NAND2_X1 U10613 ( .A1(keyinput51), .A2(n9243), .ZN(n9248) );
  NAND4_X1 U10614 ( .A1(keyinput1), .A2(keyinput89), .A3(keyinput12), .A4(
        keyinput106), .ZN(n9247) );
  OR4_X1 U10615 ( .A1(keyinput26), .A2(keyinput111), .A3(keyinput94), .A4(
        keyinput19), .ZN(n9246) );
  INV_X1 U10616 ( .A(keyinput82), .ZN(n9244) );
  NAND4_X1 U10617 ( .A1(keyinput87), .A2(keyinput44), .A3(keyinput97), .A4(
        n9244), .ZN(n9245) );
  NOR4_X1 U10618 ( .A1(n9248), .A2(n9247), .A3(n9246), .A4(n9245), .ZN(n9249)
         );
  NAND4_X1 U10619 ( .A1(keyinput24), .A2(keyinput33), .A3(n9250), .A4(n9249), 
        .ZN(n9251) );
  NOR4_X1 U10620 ( .A1(keyinput47), .A2(keyinput32), .A3(n9252), .A4(n9251), 
        .ZN(n9282) );
  INV_X1 U10621 ( .A(keyinput117), .ZN(n9253) );
  NAND4_X1 U10622 ( .A1(keyinput115), .A2(keyinput45), .A3(keyinput49), .A4(
        n9253), .ZN(n9262) );
  NOR2_X1 U10623 ( .A1(keyinput98), .A2(keyinput55), .ZN(n9254) );
  NAND3_X1 U10624 ( .A1(keyinput5), .A2(keyinput13), .A3(n9254), .ZN(n9261) );
  NOR4_X1 U10625 ( .A1(keyinput6), .A2(keyinput57), .A3(keyinput52), .A4(
        keyinput70), .ZN(n9259) );
  INV_X1 U10626 ( .A(keyinput23), .ZN(n9255) );
  NOR4_X1 U10627 ( .A1(keyinput86), .A2(keyinput21), .A3(keyinput41), .A4(
        n9255), .ZN(n9258) );
  NOR4_X1 U10628 ( .A1(keyinput103), .A2(keyinput25), .A3(keyinput99), .A4(
        keyinput58), .ZN(n9257) );
  NOR4_X1 U10629 ( .A1(keyinput18), .A2(keyinput120), .A3(keyinput127), .A4(
        keyinput76), .ZN(n9256) );
  NAND4_X1 U10630 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n9260)
         );
  NOR3_X1 U10631 ( .A1(n9262), .A2(n9261), .A3(n9260), .ZN(n9281) );
  NAND4_X1 U10632 ( .A1(keyinput74), .A2(keyinput10), .A3(keyinput67), .A4(
        keyinput122), .ZN(n9263) );
  NOR3_X1 U10633 ( .A1(keyinput114), .A2(keyinput2), .A3(n9263), .ZN(n9271) );
  INV_X1 U10634 ( .A(keyinput59), .ZN(n9520) );
  NAND4_X1 U10635 ( .A1(keyinput123), .A2(keyinput126), .A3(keyinput65), .A4(
        n9520), .ZN(n9269) );
  NAND4_X1 U10636 ( .A1(keyinput100), .A2(keyinput28), .A3(keyinput43), .A4(
        keyinput27), .ZN(n9268) );
  NOR2_X1 U10637 ( .A1(keyinput38), .A2(keyinput61), .ZN(n9264) );
  NAND3_X1 U10638 ( .A1(keyinput3), .A2(keyinput78), .A3(n9264), .ZN(n9267) );
  INV_X1 U10639 ( .A(keyinput102), .ZN(n9265) );
  NAND4_X1 U10640 ( .A1(keyinput75), .A2(keyinput22), .A3(keyinput77), .A4(
        n9265), .ZN(n9266) );
  NOR4_X1 U10641 ( .A1(n9269), .A2(n9268), .A3(n9267), .A4(n9266), .ZN(n9270)
         );
  AND4_X1 U10642 ( .A1(keyinput31), .A2(keyinput7), .A3(n9271), .A4(n9270), 
        .ZN(n9280) );
  INV_X1 U10643 ( .A(keyinput16), .ZN(n9272) );
  NOR4_X1 U10644 ( .A1(keyinput88), .A2(keyinput37), .A3(keyinput29), .A4(
        n9272), .ZN(n9278) );
  NAND2_X1 U10645 ( .A1(keyinput90), .A2(keyinput8), .ZN(n9273) );
  NOR3_X1 U10646 ( .A1(keyinput11), .A2(keyinput109), .A3(n9273), .ZN(n9277)
         );
  NOR4_X1 U10647 ( .A1(keyinput68), .A2(keyinput107), .A3(keyinput4), .A4(
        keyinput91), .ZN(n9276) );
  NAND2_X1 U10648 ( .A1(keyinput64), .A2(keyinput83), .ZN(n9274) );
  NOR3_X1 U10649 ( .A1(keyinput60), .A2(keyinput54), .A3(n9274), .ZN(n9275) );
  AND4_X1 U10650 ( .A1(n9278), .A2(n9277), .A3(n9276), .A4(n9275), .ZN(n9279)
         );
  AND4_X1 U10651 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(n9537)
         );
  NOR4_X1 U10652 ( .A1(keyinput42), .A2(keyinput0), .A3(keyinput46), .A4(
        keyinput95), .ZN(n9283) );
  NAND3_X1 U10653 ( .A1(keyinput84), .A2(keyinput62), .A3(n9283), .ZN(n9296)
         );
  NOR2_X1 U10654 ( .A1(keyinput48), .A2(keyinput112), .ZN(n9284) );
  NAND3_X1 U10655 ( .A1(keyinput105), .A2(keyinput30), .A3(n9284), .ZN(n9285)
         );
  NOR3_X1 U10656 ( .A1(keyinput119), .A2(keyinput116), .A3(n9285), .ZN(n9294)
         );
  NOR2_X1 U10657 ( .A1(keyinput73), .A2(keyinput20), .ZN(n9286) );
  NAND3_X1 U10658 ( .A1(keyinput124), .A2(keyinput71), .A3(n9286), .ZN(n9292)
         );
  INV_X1 U10659 ( .A(keyinput66), .ZN(n9287) );
  NAND4_X1 U10660 ( .A1(keyinput69), .A2(keyinput56), .A3(keyinput108), .A4(
        n9287), .ZN(n9291) );
  OR4_X1 U10661 ( .A1(keyinput92), .A2(keyinput17), .A3(keyinput15), .A4(
        keyinput79), .ZN(n9290) );
  INV_X1 U10662 ( .A(keyinput36), .ZN(n9288) );
  NAND4_X1 U10663 ( .A1(keyinput93), .A2(keyinput113), .A3(keyinput63), .A4(
        n9288), .ZN(n9289) );
  NOR4_X1 U10664 ( .A1(n9292), .A2(n9291), .A3(n9290), .A4(n9289), .ZN(n9293)
         );
  NAND4_X1 U10665 ( .A1(keyinput40), .A2(keyinput125), .A3(n9294), .A4(n9293), 
        .ZN(n9295) );
  NOR4_X1 U10666 ( .A1(keyinput110), .A2(keyinput96), .A3(n9296), .A4(n9295), 
        .ZN(n9536) );
  INV_X1 U10667 ( .A(SI_18_), .ZN(n9299) );
  AOI22_X1 U10668 ( .A1(n9299), .A2(keyinput82), .B1(keyinput87), .B2(n9298), 
        .ZN(n9297) );
  OAI221_X1 U10669 ( .B1(n9299), .B2(keyinput82), .C1(n9298), .C2(keyinput87), 
        .A(n9297), .ZN(n9311) );
  AOI22_X1 U10670 ( .A1(n9301), .A2(keyinput26), .B1(keyinput111), .B2(n5256), 
        .ZN(n9300) );
  OAI221_X1 U10671 ( .B1(n9301), .B2(keyinput26), .C1(n5256), .C2(keyinput111), 
        .A(n9300), .ZN(n9310) );
  INV_X1 U10672 ( .A(keyinput44), .ZN(n9304) );
  INV_X1 U10673 ( .A(keyinput97), .ZN(n9303) );
  AOI22_X1 U10674 ( .A1(n9304), .A2(P1_ADDR_REG_9__SCAN_IN), .B1(
        P1_ADDR_REG_13__SCAN_IN), .B2(n9303), .ZN(n9302) );
  OAI221_X1 U10675 ( .B1(n9304), .B2(P1_ADDR_REG_9__SCAN_IN), .C1(n9303), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n9302), .ZN(n9309) );
  INV_X1 U10676 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9306) );
  AOI22_X1 U10677 ( .A1(n9307), .A2(keyinput94), .B1(keyinput19), .B2(n9306), 
        .ZN(n9305) );
  OAI221_X1 U10678 ( .B1(n9307), .B2(keyinput94), .C1(n9306), .C2(keyinput19), 
        .A(n9305), .ZN(n9308) );
  NOR4_X1 U10679 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), .ZN(n9325)
         );
  INV_X1 U10680 ( .A(SI_7_), .ZN(n9313) );
  INV_X1 U10681 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U10682 ( .A1(n9313), .A2(keyinput18), .B1(n9987), .B2(keyinput120), 
        .ZN(n9312) );
  OAI221_X1 U10683 ( .B1(n9313), .B2(keyinput18), .C1(n9987), .C2(keyinput120), 
        .A(n9312), .ZN(n9323) );
  INV_X1 U10684 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9316) );
  INV_X1 U10685 ( .A(keyinput76), .ZN(n9315) );
  AOI22_X1 U10686 ( .A1(n9316), .A2(keyinput127), .B1(P1_ADDR_REG_17__SCAN_IN), 
        .B2(n9315), .ZN(n9314) );
  OAI221_X1 U10687 ( .B1(n9316), .B2(keyinput127), .C1(n9315), .C2(
        P1_ADDR_REG_17__SCAN_IN), .A(n9314), .ZN(n9322) );
  AOI22_X1 U10688 ( .A1(n9318), .A2(keyinput103), .B1(keyinput25), .B2(n4685), 
        .ZN(n9317) );
  OAI221_X1 U10689 ( .B1(n9318), .B2(keyinput103), .C1(n4685), .C2(keyinput25), 
        .A(n9317), .ZN(n9321) );
  INV_X1 U10690 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10061) );
  INV_X1 U10691 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n9989) );
  AOI22_X1 U10692 ( .A1(n10061), .A2(keyinput99), .B1(n9989), .B2(keyinput58), 
        .ZN(n9319) );
  OAI221_X1 U10693 ( .B1(n10061), .B2(keyinput99), .C1(n9989), .C2(keyinput58), 
        .A(n9319), .ZN(n9320) );
  NOR4_X1 U10694 ( .A1(n9323), .A2(n9322), .A3(n9321), .A4(n9320), .ZN(n9324)
         );
  NAND2_X1 U10695 ( .A1(n9325), .A2(n9324), .ZN(n9535) );
  INV_X1 U10696 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U10697 ( .A1(n9327), .A2(keyinput16), .B1(n9776), .B2(keyinput29), 
        .ZN(n9326) );
  OAI221_X1 U10698 ( .B1(n9327), .B2(keyinput16), .C1(n9776), .C2(keyinput29), 
        .A(n9326), .ZN(n9339) );
  AOI22_X1 U10699 ( .A1(n9329), .A2(keyinput88), .B1(n5559), .B2(keyinput37), 
        .ZN(n9328) );
  OAI221_X1 U10700 ( .B1(n9329), .B2(keyinput88), .C1(n5559), .C2(keyinput37), 
        .A(n9328), .ZN(n9338) );
  AOI22_X1 U10701 ( .A1(n9332), .A2(keyinput11), .B1(keyinput90), .B2(n9331), 
        .ZN(n9330) );
  OAI221_X1 U10702 ( .B1(n9332), .B2(keyinput11), .C1(n9331), .C2(keyinput90), 
        .A(n9330), .ZN(n9337) );
  INV_X1 U10703 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9334) );
  AOI22_X1 U10704 ( .A1(n9335), .A2(keyinput8), .B1(n9334), .B2(keyinput109), 
        .ZN(n9333) );
  OAI221_X1 U10705 ( .B1(n9335), .B2(keyinput8), .C1(n9334), .C2(keyinput109), 
        .A(n9333), .ZN(n9336) );
  NOR4_X1 U10706 ( .A1(n9339), .A2(n9338), .A3(n9337), .A4(n9336), .ZN(n9351)
         );
  AOI22_X1 U10707 ( .A1(n9341), .A2(keyinput39), .B1(n5858), .B2(keyinput118), 
        .ZN(n9340) );
  OAI221_X1 U10708 ( .B1(n9341), .B2(keyinput39), .C1(n5858), .C2(keyinput118), 
        .A(n9340), .ZN(n9349) );
  AOI22_X1 U10709 ( .A1(n5054), .A2(keyinput101), .B1(n6121), .B2(keyinput53), 
        .ZN(n9342) );
  OAI221_X1 U10710 ( .B1(n5054), .B2(keyinput101), .C1(n6121), .C2(keyinput53), 
        .A(n9342), .ZN(n9348) );
  AOI22_X1 U10711 ( .A1(n5011), .A2(keyinput24), .B1(keyinput33), .B2(n5018), 
        .ZN(n9343) );
  OAI221_X1 U10712 ( .B1(n5011), .B2(keyinput24), .C1(n5018), .C2(keyinput33), 
        .A(n9343), .ZN(n9347) );
  AOI22_X1 U10713 ( .A1(n4683), .A2(keyinput85), .B1(keyinput104), .B2(n9345), 
        .ZN(n9344) );
  OAI221_X1 U10714 ( .B1(n4683), .B2(keyinput85), .C1(n9345), .C2(keyinput104), 
        .A(n9344), .ZN(n9346) );
  NOR4_X1 U10715 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n9350)
         );
  AND2_X1 U10716 ( .A1(n9351), .A2(n9350), .ZN(n9533) );
  INV_X1 U10717 ( .A(keyinput77), .ZN(n9353) );
  AOI22_X1 U10718 ( .A1(n9354), .A2(keyinput102), .B1(P1_ADDR_REG_4__SCAN_IN), 
        .B2(n9353), .ZN(n9352) );
  OAI221_X1 U10719 ( .B1(n9354), .B2(keyinput102), .C1(n9353), .C2(
        P1_ADDR_REG_4__SCAN_IN), .A(n9352), .ZN(n9365) );
  INV_X1 U10720 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U10721 ( .A1(n9986), .A2(keyinput22), .B1(keyinput75), .B2(n9356), 
        .ZN(n9355) );
  OAI221_X1 U10722 ( .B1(n9986), .B2(keyinput22), .C1(n9356), .C2(keyinput75), 
        .A(n9355), .ZN(n9364) );
  INV_X1 U10723 ( .A(keyinput38), .ZN(n9358) );
  AOI22_X1 U10724 ( .A1(n5838), .A2(keyinput78), .B1(P2_ADDR_REG_13__SCAN_IN), 
        .B2(n9358), .ZN(n9357) );
  OAI221_X1 U10725 ( .B1(n5838), .B2(keyinput78), .C1(n9358), .C2(
        P2_ADDR_REG_13__SCAN_IN), .A(n9357), .ZN(n9363) );
  AOI22_X1 U10726 ( .A1(n9361), .A2(keyinput3), .B1(n9360), .B2(keyinput61), 
        .ZN(n9359) );
  OAI221_X1 U10727 ( .B1(n9361), .B2(keyinput3), .C1(n9360), .C2(keyinput61), 
        .A(n9359), .ZN(n9362) );
  NOR4_X1 U10728 ( .A1(n9365), .A2(n9364), .A3(n9363), .A4(n9362), .ZN(n9532)
         );
  INV_X1 U10729 ( .A(keyinput125), .ZN(n9367) );
  AOI22_X1 U10730 ( .A1(n9368), .A2(keyinput40), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9367), .ZN(n9366) );
  OAI221_X1 U10731 ( .B1(n9368), .B2(keyinput40), .C1(n9367), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9366), .ZN(n9373) );
  INV_X1 U10732 ( .A(keyinput105), .ZN(n9370) );
  AOI22_X1 U10733 ( .A1(n9371), .A2(keyinput48), .B1(P2_ADDR_REG_0__SCAN_IN), 
        .B2(n9370), .ZN(n9369) );
  OAI221_X1 U10734 ( .B1(n9371), .B2(keyinput48), .C1(n9370), .C2(
        P2_ADDR_REG_0__SCAN_IN), .A(n9369), .ZN(n9372) );
  NOR2_X1 U10735 ( .A1(n9373), .A2(n9372), .ZN(n9397) );
  INV_X1 U10736 ( .A(keyinput28), .ZN(n9375) );
  AOI22_X1 U10737 ( .A1(n9376), .A2(keyinput100), .B1(P2_ADDR_REG_10__SCAN_IN), 
        .B2(n9375), .ZN(n9374) );
  OAI221_X1 U10738 ( .B1(n9376), .B2(keyinput100), .C1(n9375), .C2(
        P2_ADDR_REG_10__SCAN_IN), .A(n9374), .ZN(n9381) );
  INV_X1 U10739 ( .A(keyinput50), .ZN(n9378) );
  NOR2_X1 U10740 ( .A1(n9381), .A2(n9380), .ZN(n9396) );
  INV_X1 U10741 ( .A(keyinput81), .ZN(n9383) );
  AOI22_X1 U10742 ( .A1(n7350), .A2(keyinput35), .B1(P1_ADDR_REG_0__SCAN_IN), 
        .B2(n9383), .ZN(n9382) );
  OAI221_X1 U10743 ( .B1(n7350), .B2(keyinput35), .C1(n9383), .C2(
        P1_ADDR_REG_0__SCAN_IN), .A(n9382), .ZN(n9388) );
  INV_X1 U10744 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9386) );
  INV_X1 U10745 ( .A(keyinput13), .ZN(n9385) );
  AOI22_X1 U10746 ( .A1(n9386), .A2(keyinput55), .B1(P1_ADDR_REG_2__SCAN_IN), 
        .B2(n9385), .ZN(n9384) );
  OAI221_X1 U10747 ( .B1(n9386), .B2(keyinput55), .C1(n9385), .C2(
        P1_ADDR_REG_2__SCAN_IN), .A(n9384), .ZN(n9387) );
  NOR2_X1 U10748 ( .A1(n9388), .A2(n9387), .ZN(n9395) );
  INV_X1 U10749 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n9982) );
  AOI22_X1 U10750 ( .A1(n9390), .A2(keyinput6), .B1(n9982), .B2(keyinput57), 
        .ZN(n9389) );
  OAI221_X1 U10751 ( .B1(n9390), .B2(keyinput6), .C1(n9982), .C2(keyinput57), 
        .A(n9389), .ZN(n9393) );
  INV_X1 U10752 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9778) );
  INV_X1 U10753 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9983) );
  AOI22_X1 U10754 ( .A1(n9778), .A2(keyinput23), .B1(n9983), .B2(keyinput21), 
        .ZN(n9391) );
  OAI221_X1 U10755 ( .B1(n9778), .B2(keyinput23), .C1(n9983), .C2(keyinput21), 
        .A(n9391), .ZN(n9392) );
  NOR2_X1 U10756 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND4_X1 U10757 ( .A1(n9397), .A2(n9396), .A3(n9395), .A4(n9394), .ZN(n9423)
         );
  INV_X1 U10758 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9399) );
  INV_X1 U10759 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9985) );
  AOI22_X1 U10760 ( .A1(n9399), .A2(keyinput20), .B1(n9985), .B2(keyinput71), 
        .ZN(n9398) );
  OAI221_X1 U10761 ( .B1(n9399), .B2(keyinput20), .C1(n9985), .C2(keyinput71), 
        .A(n9398), .ZN(n9402) );
  INV_X1 U10762 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U10763 ( .A1(n7636), .A2(keyinput45), .B1(n10073), .B2(keyinput49), 
        .ZN(n9400) );
  OAI221_X1 U10764 ( .B1(n7636), .B2(keyinput45), .C1(n10073), .C2(keyinput49), 
        .A(n9400), .ZN(n9401) );
  NOR2_X1 U10765 ( .A1(n9402), .A2(n9401), .ZN(n9421) );
  AOI22_X1 U10766 ( .A1(n7082), .A2(keyinput15), .B1(n9404), .B2(keyinput79), 
        .ZN(n9403) );
  OAI221_X1 U10767 ( .B1(n7082), .B2(keyinput15), .C1(n9404), .C2(keyinput79), 
        .A(n9403), .ZN(n9408) );
  AOI22_X1 U10768 ( .A1(n7439), .A2(keyinput112), .B1(keyinput30), .B2(n9406), 
        .ZN(n9405) );
  OAI221_X1 U10769 ( .B1(n7439), .B2(keyinput112), .C1(n9406), .C2(keyinput30), 
        .A(n9405), .ZN(n9407) );
  NOR2_X1 U10770 ( .A1(n9408), .A2(n9407), .ZN(n9420) );
  AOI22_X1 U10771 ( .A1(n9411), .A2(keyinput36), .B1(n9410), .B2(keyinput63), 
        .ZN(n9409) );
  OAI221_X1 U10772 ( .B1(n9411), .B2(keyinput36), .C1(n9410), .C2(keyinput63), 
        .A(n9409), .ZN(n9416) );
  AOI22_X1 U10773 ( .A1(n9414), .A2(keyinput46), .B1(keyinput95), .B2(n9413), 
        .ZN(n9412) );
  OAI221_X1 U10774 ( .B1(n9414), .B2(keyinput46), .C1(n9413), .C2(keyinput95), 
        .A(n9412), .ZN(n9415) );
  NOR2_X1 U10775 ( .A1(n9416), .A2(n9415), .ZN(n9419) );
  INV_X1 U10776 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9984) );
  INV_X1 U10777 ( .A(keyinput41), .ZN(n9417) );
  XNOR2_X1 U10778 ( .A(n9984), .B(n9417), .ZN(n9418) );
  NAND4_X1 U10779 ( .A1(n9421), .A2(n9420), .A3(n9419), .A4(n9418), .ZN(n9422)
         );
  NOR2_X1 U10780 ( .A1(n9423), .A2(n9422), .ZN(n9531) );
  AOI22_X1 U10781 ( .A1(n9425), .A2(keyinput108), .B1(keyinput66), .B2(n7949), 
        .ZN(n9424) );
  OAI221_X1 U10782 ( .B1(n9425), .B2(keyinput108), .C1(n7949), .C2(keyinput66), 
        .A(n9424), .ZN(n9434) );
  AOI22_X1 U10783 ( .A1(n9428), .A2(keyinput114), .B1(keyinput2), .B2(n9427), 
        .ZN(n9426) );
  OAI221_X1 U10784 ( .B1(n9428), .B2(keyinput114), .C1(n9427), .C2(keyinput2), 
        .A(n9426), .ZN(n9433) );
  AOI22_X1 U10785 ( .A1(n9431), .A2(keyinput60), .B1(keyinput83), .B2(n9430), 
        .ZN(n9429) );
  OAI221_X1 U10786 ( .B1(n9431), .B2(keyinput60), .C1(n9430), .C2(keyinput83), 
        .A(n9429), .ZN(n9432) );
  NOR3_X1 U10787 ( .A1(n9434), .A2(n9433), .A3(n9432), .ZN(n9486) );
  AOI22_X1 U10788 ( .A1(n9436), .A2(keyinput92), .B1(keyinput17), .B2(n6025), 
        .ZN(n9435) );
  OAI221_X1 U10789 ( .B1(n9436), .B2(keyinput92), .C1(n6025), .C2(keyinput17), 
        .A(n9435), .ZN(n9445) );
  INV_X1 U10790 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9439) );
  AOI22_X1 U10791 ( .A1(n9439), .A2(keyinput126), .B1(keyinput65), .B2(n9438), 
        .ZN(n9437) );
  OAI221_X1 U10792 ( .B1(n9439), .B2(keyinput126), .C1(n9438), .C2(keyinput65), 
        .A(n9437), .ZN(n9444) );
  AOI22_X1 U10793 ( .A1(n9442), .A2(keyinput56), .B1(keyinput69), .B2(n9441), 
        .ZN(n9440) );
  OAI221_X1 U10794 ( .B1(n9442), .B2(keyinput56), .C1(n9441), .C2(keyinput69), 
        .A(n9440), .ZN(n9443) );
  NOR3_X1 U10795 ( .A1(n9445), .A2(n9444), .A3(n9443), .ZN(n9485) );
  INV_X1 U10796 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U10797 ( .A1(n10296), .A2(keyinput31), .B1(n9447), .B2(keyinput7), 
        .ZN(n9446) );
  OAI221_X1 U10798 ( .B1(n10296), .B2(keyinput31), .C1(n9447), .C2(keyinput7), 
        .A(n9446), .ZN(n9460) );
  AOI22_X1 U10799 ( .A1(n5758), .A2(keyinput47), .B1(keyinput32), .B2(n9449), 
        .ZN(n9448) );
  OAI221_X1 U10800 ( .B1(n5758), .B2(keyinput47), .C1(n9449), .C2(keyinput32), 
        .A(n9448), .ZN(n9459) );
  XNOR2_X1 U10801 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput106), .ZN(n9453) );
  XNOR2_X1 U10802 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput14), .ZN(n9452) );
  XNOR2_X1 U10803 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput119), .ZN(n9451) );
  XNOR2_X1 U10804 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput73), .ZN(n9450) );
  AND4_X1 U10805 ( .A1(n9453), .A2(n9452), .A3(n9451), .A4(n9450), .ZN(n9457)
         );
  XNOR2_X1 U10806 ( .A(keyinput43), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9456) );
  XNOR2_X1 U10807 ( .A(SI_9_), .B(keyinput93), .ZN(n9455) );
  XNOR2_X1 U10808 ( .A(SI_3_), .B(keyinput113), .ZN(n9454) );
  NAND4_X1 U10809 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .ZN(n9458)
         );
  NOR3_X1 U10810 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(n9484) );
  XNOR2_X1 U10811 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput124), .ZN(n9464) );
  XNOR2_X1 U10812 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput10), .ZN(n9463) );
  XNOR2_X1 U10813 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput86), .ZN(n9462) );
  XNOR2_X1 U10814 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput68), .ZN(n9461) );
  NAND4_X1 U10815 ( .A1(n9464), .A2(n9463), .A3(n9462), .A4(n9461), .ZN(n9470)
         );
  XNOR2_X1 U10816 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(keyinput74), .ZN(n9468)
         );
  XNOR2_X1 U10817 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput80), .ZN(n9467) );
  XNOR2_X1 U10818 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput0), .ZN(n9466) );
  XNOR2_X1 U10819 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput9), .ZN(n9465) );
  NAND4_X1 U10820 ( .A1(n9468), .A2(n9467), .A3(n9466), .A4(n9465), .ZN(n9469)
         );
  NOR2_X1 U10821 ( .A1(n9470), .A2(n9469), .ZN(n9482) );
  XNOR2_X1 U10822 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput12), .ZN(n9474) );
  XNOR2_X1 U10823 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput27), .ZN(n9473) );
  XNOR2_X1 U10824 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput115), .ZN(n9472) );
  XNOR2_X1 U10825 ( .A(P2_REG2_REG_1__SCAN_IN), .B(keyinput4), .ZN(n9471) );
  NAND4_X1 U10826 ( .A1(n9474), .A2(n9473), .A3(n9472), .A4(n9471), .ZN(n9480)
         );
  XNOR2_X1 U10827 ( .A(keyinput117), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n9478)
         );
  XNOR2_X1 U10828 ( .A(keyinput107), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9477) );
  XNOR2_X1 U10829 ( .A(keyinput116), .B(P1_REG2_REG_20__SCAN_IN), .ZN(n9476)
         );
  XNOR2_X1 U10830 ( .A(keyinput51), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n9475) );
  NAND4_X1 U10831 ( .A1(n9478), .A2(n9477), .A3(n9476), .A4(n9475), .ZN(n9479)
         );
  NOR2_X1 U10832 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  AND2_X1 U10833 ( .A1(n9482), .A2(n9481), .ZN(n9483) );
  NAND4_X1 U10834 ( .A1(n9486), .A2(n9485), .A3(n9484), .A4(n9483), .ZN(n9529)
         );
  INV_X1 U10835 ( .A(SI_5_), .ZN(n9488) );
  AOI22_X1 U10836 ( .A1(n9488), .A2(keyinput52), .B1(keyinput70), .B2(n5034), 
        .ZN(n9487) );
  OAI221_X1 U10837 ( .B1(n9488), .B2(keyinput52), .C1(n5034), .C2(keyinput70), 
        .A(n9487), .ZN(n9497) );
  AOI22_X1 U10838 ( .A1(n9491), .A2(keyinput67), .B1(keyinput122), .B2(n9490), 
        .ZN(n9489) );
  OAI221_X1 U10839 ( .B1(n9491), .B2(keyinput67), .C1(n9490), .C2(keyinput122), 
        .A(n9489), .ZN(n9496) );
  AOI22_X1 U10840 ( .A1(n9494), .A2(keyinput34), .B1(n9493), .B2(keyinput72), 
        .ZN(n9492) );
  OAI221_X1 U10841 ( .B1(n9494), .B2(keyinput34), .C1(n9493), .C2(keyinput72), 
        .A(n9492), .ZN(n9495) );
  NOR3_X1 U10842 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(n9527) );
  INV_X1 U10843 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9499) );
  AOI22_X1 U10844 ( .A1(n9500), .A2(keyinput98), .B1(keyinput5), .B2(n9499), 
        .ZN(n9498) );
  OAI221_X1 U10845 ( .B1(n9500), .B2(keyinput98), .C1(n9499), .C2(keyinput5), 
        .A(n9498), .ZN(n9505) );
  INV_X1 U10846 ( .A(keyinput64), .ZN(n9502) );
  AOI22_X1 U10847 ( .A1(n9503), .A2(keyinput54), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n9502), .ZN(n9501) );
  OAI221_X1 U10848 ( .B1(n9503), .B2(keyinput54), .C1(n9502), .C2(
        P2_ADDR_REG_15__SCAN_IN), .A(n9501), .ZN(n9504) );
  NOR2_X1 U10849 ( .A1(n9505), .A2(n9504), .ZN(n9526) );
  AOI22_X1 U10850 ( .A1(n9508), .A2(keyinput110), .B1(n9507), .B2(keyinput96), 
        .ZN(n9506) );
  OAI221_X1 U10851 ( .B1(n9508), .B2(keyinput110), .C1(n9507), .C2(keyinput96), 
        .A(n9506), .ZN(n9509) );
  INV_X1 U10852 ( .A(n9509), .ZN(n9513) );
  XNOR2_X1 U10853 ( .A(keyinput91), .B(n8561), .ZN(n9511) );
  XNOR2_X1 U10854 ( .A(keyinput42), .B(n5580), .ZN(n9510) );
  NOR2_X1 U10855 ( .A1(n9511), .A2(n9510), .ZN(n9512) );
  NAND2_X1 U10856 ( .A1(n9513), .A2(n9512), .ZN(n9516) );
  NOR2_X1 U10857 ( .A1(n9516), .A2(n9515), .ZN(n9525) );
  INV_X1 U10858 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U10859 ( .A1(n9518), .A2(keyinput84), .B1(keyinput62), .B2(n10310), 
        .ZN(n9517) );
  OAI221_X1 U10860 ( .B1(n9518), .B2(keyinput84), .C1(n10310), .C2(keyinput62), 
        .A(n9517), .ZN(n9523) );
  INV_X1 U10861 ( .A(SI_16_), .ZN(n9521) );
  AOI22_X1 U10862 ( .A1(n9521), .A2(keyinput123), .B1(P2_ADDR_REG_16__SCAN_IN), 
        .B2(n9520), .ZN(n9519) );
  OAI221_X1 U10863 ( .B1(n9521), .B2(keyinput123), .C1(n9520), .C2(
        P2_ADDR_REG_16__SCAN_IN), .A(n9519), .ZN(n9522) );
  NOR2_X1 U10864 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  NAND4_X1 U10865 ( .A1(n9527), .A2(n9526), .A3(n9525), .A4(n9524), .ZN(n9528)
         );
  NOR2_X1 U10866 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NAND4_X1 U10867 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n9534)
         );
  AOI211_X1 U10868 ( .C1(n9537), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9554)
         );
  XNOR2_X1 U10869 ( .A(n9538), .B(n9540), .ZN(n9657) );
  INV_X1 U10870 ( .A(n9539), .ZN(n9541) );
  OAI21_X1 U10871 ( .B1(n9541), .B2(n9540), .A(n9947), .ZN(n9544) );
  OAI21_X1 U10872 ( .B1(n9544), .B2(n9543), .A(n9542), .ZN(n9653) );
  INV_X1 U10873 ( .A(n9655), .ZN(n9550) );
  INV_X1 U10874 ( .A(n9545), .ZN(n9546) );
  AOI211_X1 U10875 ( .C1(n9655), .C2(n9559), .A(n9612), .B(n9546), .ZN(n9654)
         );
  NAND2_X1 U10876 ( .A1(n9654), .A2(n9978), .ZN(n9549) );
  AOI22_X1 U10877 ( .A1(n9547), .A2(n9967), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9973), .ZN(n9548) );
  OAI211_X1 U10878 ( .C1(n9550), .C2(n9970), .A(n9549), .B(n9548), .ZN(n9551)
         );
  AOI21_X1 U10879 ( .B1(n9588), .B2(n9653), .A(n9551), .ZN(n9552) );
  OAI21_X1 U10880 ( .B1(n9657), .B2(n9623), .A(n9552), .ZN(n9553) );
  XOR2_X1 U10881 ( .A(n9554), .B(n9553), .Z(P1_U3269) );
  OAI21_X1 U10882 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9558) );
  INV_X1 U10883 ( .A(n9558), .ZN(n9662) );
  INV_X1 U10884 ( .A(n9583), .ZN(n9561) );
  INV_X1 U10885 ( .A(n9559), .ZN(n9560) );
  AOI211_X1 U10886 ( .C1(n9659), .C2(n9561), .A(n9612), .B(n9560), .ZN(n9658)
         );
  AOI22_X1 U10887 ( .A1(n9562), .A2(n9967), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9973), .ZN(n9563) );
  OAI21_X1 U10888 ( .B1(n9564), .B2(n9970), .A(n9563), .ZN(n9572) );
  INV_X1 U10889 ( .A(n9565), .ZN(n9566) );
  NOR2_X1 U10890 ( .A1(n9577), .A2(n9566), .ZN(n9568) );
  XNOR2_X1 U10891 ( .A(n9568), .B(n9567), .ZN(n9570) );
  AOI21_X1 U10892 ( .B1(n9570), .B2(n9947), .A(n9569), .ZN(n9661) );
  NOR2_X1 U10893 ( .A1(n9661), .A2(n9973), .ZN(n9571) );
  AOI211_X1 U10894 ( .C1(n9658), .C2(n9978), .A(n9572), .B(n9571), .ZN(n9573)
         );
  OAI21_X1 U10895 ( .B1(n9662), .B2(n9623), .A(n9573), .ZN(P1_U3270) );
  OAI21_X1 U10896 ( .B1(n9575), .B2(n9579), .A(n9574), .ZN(n9576) );
  INV_X1 U10897 ( .A(n9576), .ZN(n9667) );
  AOI211_X1 U10898 ( .C1(n9579), .C2(n9578), .A(n9963), .B(n9577), .ZN(n9581)
         );
  NOR2_X1 U10899 ( .A1(n9581), .A2(n9580), .ZN(n9666) );
  OAI21_X1 U10900 ( .B1(n9582), .B2(n9949), .A(n9666), .ZN(n9589) );
  AOI211_X1 U10901 ( .C1(n9664), .C2(n4518), .A(n9612), .B(n9583), .ZN(n9663)
         );
  INV_X1 U10902 ( .A(n9663), .ZN(n9586) );
  AOI22_X1 U10903 ( .A1(n9664), .A2(n9599), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9973), .ZN(n9584) );
  OAI21_X1 U10904 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9587) );
  AOI21_X1 U10905 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(n9590) );
  OAI21_X1 U10906 ( .B1(n9667), .B2(n9623), .A(n9590), .ZN(P1_U3271) );
  INV_X1 U10907 ( .A(n9591), .ZN(n9592) );
  AOI21_X1 U10908 ( .B1(n9617), .B2(n9593), .A(n9592), .ZN(n9595) );
  XNOR2_X1 U10909 ( .A(n9595), .B(n9594), .ZN(n9597) );
  AOI21_X1 U10910 ( .B1(n9597), .B2(n9947), .A(n9596), .ZN(n9671) );
  AOI21_X1 U10911 ( .B1(n9669), .B2(n9611), .A(n9612), .ZN(n9598) );
  AND2_X1 U10912 ( .A1(n9598), .A2(n4518), .ZN(n9668) );
  NAND2_X1 U10913 ( .A1(n9669), .A2(n9599), .ZN(n9601) );
  NAND2_X1 U10914 ( .A1(n9968), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9600) );
  OAI211_X1 U10915 ( .C1(n9949), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9608)
         );
  OAI21_X1 U10916 ( .B1(n9605), .B2(n9604), .A(n9603), .ZN(n9606) );
  INV_X1 U10917 ( .A(n9606), .ZN(n9672) );
  NOR2_X1 U10918 ( .A1(n9672), .A2(n9623), .ZN(n9607) );
  AOI211_X1 U10919 ( .C1(n9668), .C2(n9978), .A(n9608), .B(n9607), .ZN(n9609)
         );
  OAI21_X1 U10920 ( .B1(n9968), .B2(n9671), .A(n9609), .ZN(P1_U3272) );
  XNOR2_X1 U10921 ( .A(n9610), .B(n9616), .ZN(n9677) );
  AOI211_X1 U10922 ( .C1(n9674), .C2(n4460), .A(n9612), .B(n4680), .ZN(n9673)
         );
  AOI22_X1 U10923 ( .A1(n9613), .A2(n9967), .B1(n9968), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9614) );
  OAI21_X1 U10924 ( .B1(n9615), .B2(n9970), .A(n9614), .ZN(n9621) );
  XNOR2_X1 U10925 ( .A(n9617), .B(n9616), .ZN(n9619) );
  AOI21_X1 U10926 ( .B1(n9619), .B2(n9947), .A(n9618), .ZN(n9676) );
  NOR2_X1 U10927 ( .A1(n9676), .A2(n9973), .ZN(n9620) );
  AOI211_X1 U10928 ( .C1(n9673), .C2(n9978), .A(n9621), .B(n9620), .ZN(n9622)
         );
  OAI21_X1 U10929 ( .B1(n9623), .B2(n9677), .A(n9622), .ZN(P1_U3273) );
  INV_X1 U10930 ( .A(n6138), .ZN(n9626) );
  OAI211_X1 U10931 ( .C1(n9626), .C2(n10076), .A(n9625), .B(n9624), .ZN(n9678)
         );
  MUX2_X1 U10932 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9678), .S(n10111), .Z(
        P1_U3553) );
  MUX2_X1 U10933 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9627), .S(n10111), .Z(
        P1_U3552) );
  INV_X1 U10934 ( .A(n10080), .ZN(n10018) );
  INV_X1 U10935 ( .A(n10076), .ZN(n10083) );
  AOI21_X1 U10936 ( .B1(n10083), .B2(n5918), .A(n9628), .ZN(n9629) );
  OAI211_X1 U10937 ( .C1(n9631), .C2(n10018), .A(n9630), .B(n9629), .ZN(n9679)
         );
  MUX2_X1 U10938 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9679), .S(n10111), .Z(
        P1_U3551) );
  AOI21_X1 U10939 ( .B1(n10083), .B2(n9633), .A(n9632), .ZN(n9636) );
  NAND3_X1 U10940 ( .A1(n9634), .A2(n9190), .A3(n10080), .ZN(n9635) );
  NAND3_X1 U10941 ( .A1(n9637), .A2(n9636), .A3(n9635), .ZN(n9680) );
  MUX2_X1 U10942 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9680), .S(n10111), .Z(
        P1_U3550) );
  MUX2_X1 U10943 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9681), .S(n10111), .Z(
        P1_U3549) );
  NAND3_X1 U10944 ( .A1(n9215), .A2(n10080), .A3(n9642), .ZN(n9646) );
  NAND2_X1 U10945 ( .A1(n9643), .A2(n10083), .ZN(n9644) );
  NAND4_X1 U10946 ( .A1(n9647), .A2(n9646), .A3(n9645), .A4(n9644), .ZN(n9682)
         );
  MUX2_X1 U10947 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9682), .S(n10111), .Z(
        P1_U3548) );
  AOI21_X1 U10948 ( .B1(n10083), .B2(n9649), .A(n9648), .ZN(n9650) );
  OAI211_X1 U10949 ( .C1(n10018), .C2(n9652), .A(n9651), .B(n9650), .ZN(n9683)
         );
  MUX2_X1 U10950 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9683), .S(n10111), .Z(
        P1_U3547) );
  AOI211_X1 U10951 ( .C1(n10083), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9656)
         );
  OAI21_X1 U10952 ( .B1(n10018), .B2(n9657), .A(n9656), .ZN(n9684) );
  MUX2_X1 U10953 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9684), .S(n10111), .Z(
        P1_U3546) );
  AOI21_X1 U10954 ( .B1(n10083), .B2(n9659), .A(n9658), .ZN(n9660) );
  OAI211_X1 U10955 ( .C1(n9662), .C2(n10018), .A(n9661), .B(n9660), .ZN(n9685)
         );
  MUX2_X1 U10956 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9685), .S(n10111), .Z(
        P1_U3545) );
  AOI21_X1 U10957 ( .B1(n10083), .B2(n9664), .A(n9663), .ZN(n9665) );
  OAI211_X1 U10958 ( .C1(n10018), .C2(n9667), .A(n9666), .B(n9665), .ZN(n9686)
         );
  MUX2_X1 U10959 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9686), .S(n10111), .Z(
        P1_U3544) );
  AOI21_X1 U10960 ( .B1(n10083), .B2(n9669), .A(n9668), .ZN(n9670) );
  OAI211_X1 U10961 ( .C1(n9672), .C2(n10018), .A(n9671), .B(n9670), .ZN(n9687)
         );
  MUX2_X1 U10962 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9687), .S(n10111), .Z(
        P1_U3543) );
  AOI21_X1 U10963 ( .B1(n10083), .B2(n9674), .A(n9673), .ZN(n9675) );
  OAI211_X1 U10964 ( .C1(n9677), .C2(n10018), .A(n9676), .B(n9675), .ZN(n9688)
         );
  MUX2_X1 U10965 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9688), .S(n10111), .Z(
        P1_U3542) );
  MUX2_X1 U10966 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9678), .S(n10092), .Z(
        P1_U3521) );
  MUX2_X1 U10967 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9679), .S(n10092), .Z(
        P1_U3519) );
  MUX2_X1 U10968 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9680), .S(n10092), .Z(
        P1_U3518) );
  MUX2_X1 U10969 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9682), .S(n10092), .Z(
        P1_U3516) );
  MUX2_X1 U10970 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9683), .S(n10092), .Z(
        P1_U3515) );
  MUX2_X1 U10971 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9684), .S(n10092), .Z(
        P1_U3514) );
  MUX2_X1 U10972 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9685), .S(n10092), .Z(
        P1_U3513) );
  MUX2_X1 U10973 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9686), .S(n10092), .Z(
        P1_U3512) );
  MUX2_X1 U10974 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9687), .S(n10092), .Z(
        P1_U3511) );
  MUX2_X1 U10975 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9688), .S(n10092), .Z(
        P1_U3510) );
  AND2_X1 U10976 ( .A1(n9690), .A2(n9689), .ZN(n9990) );
  MUX2_X1 U10977 ( .A(P1_D_REG_1__SCAN_IN), .B(n9691), .S(n9990), .Z(P1_U3440)
         );
  MUX2_X1 U10978 ( .A(P1_D_REG_0__SCAN_IN), .B(n9692), .S(n9990), .Z(P1_U3439)
         );
  NAND3_X1 U10979 ( .A1(n9386), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9695) );
  OAI22_X1 U10980 ( .A1(n9693), .A2(n9695), .B1(n9694), .B2(n8277), .ZN(n9696)
         );
  AOI21_X1 U10981 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9699) );
  INV_X1 U10982 ( .A(n9699), .ZN(P1_U3324) );
  OAI222_X1 U10983 ( .A1(n8275), .A2(n9702), .B1(n9701), .B2(P1_U3086), .C1(
        n9700), .C2(n8277), .ZN(P1_U3326) );
  INV_X1 U10984 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9715) );
  INV_X1 U10985 ( .A(n9703), .ZN(n9704) );
  AOI211_X1 U10986 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n9910), .ZN(n9711)
         );
  AOI211_X1 U10987 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n9900), .ZN(n9710)
         );
  AOI211_X1 U10988 ( .C1(n9921), .C2(n9712), .A(n9711), .B(n9710), .ZN(n9714)
         );
  NAND2_X1 U10989 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9713) );
  OAI211_X1 U10990 ( .C1(n9924), .C2(n9715), .A(n9714), .B(n9713), .ZN(
        P1_U3253) );
  INV_X1 U10991 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9730) );
  AOI21_X1 U10992 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9720) );
  NAND2_X1 U10993 ( .A1(n9861), .A2(n9720), .ZN(n9726) );
  AOI21_X1 U10994 ( .B1(n9723), .B2(n9722), .A(n9721), .ZN(n9724) );
  NAND2_X1 U10995 ( .A1(n9913), .A2(n9724), .ZN(n9725) );
  OAI211_X1 U10996 ( .C1(n9821), .C2(n4662), .A(n9726), .B(n9725), .ZN(n9727)
         );
  INV_X1 U10997 ( .A(n9727), .ZN(n9729) );
  NAND2_X1 U10998 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9728) );
  OAI211_X1 U10999 ( .C1(n9924), .C2(n9730), .A(n9729), .B(n9728), .ZN(
        P1_U3250) );
  INV_X1 U11000 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9745) );
  INV_X1 U11001 ( .A(n9731), .ZN(n9742) );
  AOI21_X1 U11002 ( .B1(n9734), .B2(n9733), .A(n9732), .ZN(n9735) );
  NAND2_X1 U11003 ( .A1(n9861), .A2(n9735), .ZN(n9741) );
  AOI21_X1 U11004 ( .B1(n9738), .B2(n9737), .A(n9736), .ZN(n9739) );
  NAND2_X1 U11005 ( .A1(n9913), .A2(n9739), .ZN(n9740) );
  OAI211_X1 U11006 ( .C1(n9821), .C2(n9742), .A(n9741), .B(n9740), .ZN(n9743)
         );
  INV_X1 U11007 ( .A(n9743), .ZN(n9744) );
  NAND2_X1 U11008 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9785) );
  OAI211_X1 U11009 ( .C1(n9924), .C2(n9745), .A(n9744), .B(n9785), .ZN(
        P1_U3251) );
  OAI211_X1 U11010 ( .C1(n9748), .C2(n10076), .A(n9747), .B(n9746), .ZN(n9749)
         );
  AOI21_X1 U11011 ( .B1(n9750), .B2(n10080), .A(n9749), .ZN(n9773) );
  AOI22_X1 U11012 ( .A1(n10111), .A2(n9773), .B1(n5987), .B2(n10109), .ZN(
        P1_U3541) );
  OAI211_X1 U11013 ( .C1(n9753), .C2(n10076), .A(n9752), .B(n9751), .ZN(n9754)
         );
  AOI21_X1 U11014 ( .B1(n9755), .B2(n10080), .A(n9754), .ZN(n9775) );
  AOI22_X1 U11015 ( .A1(n10111), .A2(n9775), .B1(n9101), .B2(n10109), .ZN(
        P1_U3540) );
  OAI21_X1 U11016 ( .B1(n9757), .B2(n10076), .A(n9756), .ZN(n9758) );
  AOI211_X1 U11017 ( .C1(n9760), .C2(n10080), .A(n9759), .B(n9758), .ZN(n9777)
         );
  AOI22_X1 U11018 ( .A1(n10111), .A2(n9777), .B1(n9081), .B2(n10109), .ZN(
        P1_U3539) );
  AOI211_X1 U11019 ( .C1(n10083), .C2(n9763), .A(n9762), .B(n9761), .ZN(n9766)
         );
  NAND3_X1 U11020 ( .A1(n8074), .A2(n9764), .A3(n10080), .ZN(n9765) );
  AND2_X1 U11021 ( .A1(n9766), .A2(n9765), .ZN(n9779) );
  AOI22_X1 U11022 ( .A1(n10111), .A2(n9779), .B1(n9053), .B2(n10109), .ZN(
        P1_U3538) );
  OAI211_X1 U11023 ( .C1(n9769), .C2(n10076), .A(n9768), .B(n9767), .ZN(n9770)
         );
  AOI21_X1 U11024 ( .B1(n10080), .B2(n9771), .A(n9770), .ZN(n9781) );
  AOI22_X1 U11025 ( .A1(n10111), .A2(n9781), .B1(n9898), .B2(n10109), .ZN(
        P1_U3537) );
  INV_X1 U11026 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U11027 ( .A1(n10092), .A2(n9773), .B1(n9772), .B2(n10090), .ZN(
        P1_U3509) );
  INV_X1 U11028 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U11029 ( .A1(n10092), .A2(n9775), .B1(n9774), .B2(n10090), .ZN(
        P1_U3507) );
  AOI22_X1 U11030 ( .A1(n10092), .A2(n9777), .B1(n9776), .B2(n10090), .ZN(
        P1_U3504) );
  AOI22_X1 U11031 ( .A1(n10092), .A2(n9779), .B1(n9778), .B2(n10090), .ZN(
        P1_U3501) );
  INV_X1 U11032 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U11033 ( .A1(n10092), .A2(n9781), .B1(n9780), .B2(n10090), .ZN(
        P1_U3498) );
  XNOR2_X1 U11034 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI21_X1 U11035 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9792) );
  INV_X1 U11036 ( .A(n9785), .ZN(n9788) );
  NOR2_X1 U11037 ( .A1(n10040), .A2(n9786), .ZN(n9787) );
  AOI211_X1 U11038 ( .C1(n4438), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9790)
         );
  OAI21_X1 U11039 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9793) );
  INV_X1 U11040 ( .A(n9793), .ZN(n9794) );
  OAI21_X1 U11041 ( .B1(n9796), .B2(n9795), .A(n9794), .ZN(P1_U3221) );
  AOI22_X1 U11042 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9811), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9810) );
  NAND2_X1 U11043 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9798) );
  AOI21_X1 U11044 ( .B1(n9799), .B2(n9798), .A(n9797), .ZN(n9800) );
  NAND2_X1 U11045 ( .A1(n9861), .A2(n9800), .ZN(n9806) );
  AOI21_X1 U11046 ( .B1(n9803), .B2(n9802), .A(n9801), .ZN(n9804) );
  NAND2_X1 U11047 ( .A1(n9913), .A2(n9804), .ZN(n9805) );
  OAI211_X1 U11048 ( .C1(n9821), .C2(n9807), .A(n9806), .B(n9805), .ZN(n9808)
         );
  INV_X1 U11049 ( .A(n9808), .ZN(n9809) );
  NAND2_X1 U11050 ( .A1(n9810), .A2(n9809), .ZN(P1_U3244) );
  AOI22_X1 U11051 ( .A1(n9811), .A2(P1_ADDR_REG_4__SCAN_IN), .B1(
        P1_REG3_REG_4__SCAN_IN), .B2(P1_U3086), .ZN(n9825) );
  OAI211_X1 U11052 ( .C1(n9814), .C2(n9813), .A(n9861), .B(n9812), .ZN(n9819)
         );
  OAI211_X1 U11053 ( .C1(n9817), .C2(n9816), .A(n9913), .B(n9815), .ZN(n9818)
         );
  OAI211_X1 U11054 ( .C1(n9821), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9822)
         );
  INV_X1 U11055 ( .A(n9822), .ZN(n9824) );
  NAND3_X1 U11056 ( .A1(n9825), .A2(n9824), .A3(n9823), .ZN(P1_U3247) );
  INV_X1 U11057 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9839) );
  OAI211_X1 U11058 ( .C1(n9828), .C2(n9827), .A(n9861), .B(n9826), .ZN(n9829)
         );
  INV_X1 U11059 ( .A(n9829), .ZN(n9834) );
  AOI211_X1 U11060 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9900), .ZN(n9833)
         );
  AOI211_X1 U11061 ( .C1(n9921), .C2(n9835), .A(n9834), .B(n9833), .ZN(n9838)
         );
  INV_X1 U11062 ( .A(n9836), .ZN(n9837) );
  OAI211_X1 U11063 ( .C1(n9924), .C2(n9839), .A(n9838), .B(n9837), .ZN(
        P1_U3248) );
  INV_X1 U11064 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9855) );
  INV_X1 U11065 ( .A(n9840), .ZN(n9844) );
  NAND2_X1 U11066 ( .A1(n9842), .A2(n9841), .ZN(n9843) );
  NAND3_X1 U11067 ( .A1(n9861), .A2(n9844), .A3(n9843), .ZN(n9852) );
  NAND2_X1 U11068 ( .A1(n9921), .A2(n9845), .ZN(n9851) );
  AOI21_X1 U11069 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9849) );
  NAND2_X1 U11070 ( .A1(n9913), .A2(n9849), .ZN(n9850) );
  AND3_X1 U11071 ( .A1(n9852), .A2(n9851), .A3(n9850), .ZN(n9854) );
  NAND2_X1 U11072 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9853) );
  OAI211_X1 U11073 ( .C1(n9924), .C2(n9855), .A(n9854), .B(n9853), .ZN(
        P1_U3249) );
  INV_X1 U11074 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U11075 ( .A1(n9857), .A2(n9856), .ZN(n9860) );
  INV_X1 U11076 ( .A(n9858), .ZN(n9859) );
  NAND3_X1 U11077 ( .A1(n9861), .A2(n9860), .A3(n9859), .ZN(n9869) );
  NAND2_X1 U11078 ( .A1(n9921), .A2(n9862), .ZN(n9868) );
  AOI21_X1 U11079 ( .B1(n9865), .B2(n9864), .A(n9863), .ZN(n9866) );
  NAND2_X1 U11080 ( .A1(n9913), .A2(n9866), .ZN(n9867) );
  AND3_X1 U11081 ( .A1(n9869), .A2(n9868), .A3(n9867), .ZN(n9871) );
  NAND2_X1 U11082 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9870) );
  OAI211_X1 U11083 ( .C1(n9924), .C2(n9872), .A(n9871), .B(n9870), .ZN(
        P1_U3254) );
  INV_X1 U11084 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9884) );
  AOI211_X1 U11085 ( .C1(n9875), .C2(n9874), .A(n9873), .B(n9900), .ZN(n9880)
         );
  AOI211_X1 U11086 ( .C1(n9878), .C2(n9877), .A(n9910), .B(n9876), .ZN(n9879)
         );
  AOI211_X1 U11087 ( .C1(n9921), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9883)
         );
  NAND2_X1 U11088 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9882) );
  OAI211_X1 U11089 ( .C1(n9884), .C2(n9924), .A(n9883), .B(n9882), .ZN(
        P1_U3256) );
  INV_X1 U11090 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9896) );
  AOI211_X1 U11091 ( .C1(n9887), .C2(n9886), .A(n9885), .B(n9900), .ZN(n9892)
         );
  AOI211_X1 U11092 ( .C1(n9890), .C2(n9889), .A(n9888), .B(n9910), .ZN(n9891)
         );
  AOI211_X1 U11093 ( .C1(n9921), .C2(n9893), .A(n9892), .B(n9891), .ZN(n9895)
         );
  NAND2_X1 U11094 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9894) );
  OAI211_X1 U11095 ( .C1(n9896), .C2(n9924), .A(n9895), .B(n9894), .ZN(
        P1_U3257) );
  INV_X1 U11096 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9908) );
  AOI211_X1 U11097 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9910), .ZN(n9904)
         );
  AOI211_X1 U11098 ( .C1(n9902), .C2(n7912), .A(n9901), .B(n9900), .ZN(n9903)
         );
  AOI211_X1 U11099 ( .C1(n9921), .C2(n9905), .A(n9904), .B(n9903), .ZN(n9907)
         );
  NAND2_X1 U11100 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n9906) );
  OAI211_X1 U11101 ( .C1(n9924), .C2(n9908), .A(n9907), .B(n9906), .ZN(
        P1_U3258) );
  AOI211_X1 U11102 ( .C1(n9912), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9919)
         );
  OAI211_X1 U11103 ( .C1(n9916), .C2(n9915), .A(n9914), .B(n9913), .ZN(n9917)
         );
  INV_X1 U11104 ( .A(n9917), .ZN(n9918) );
  AOI211_X1 U11105 ( .C1(n9921), .C2(n9920), .A(n9919), .B(n9918), .ZN(n9923)
         );
  NAND2_X1 U11106 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n9922) );
  OAI211_X1 U11107 ( .C1(n9924), .C2(n10335), .A(n9923), .B(n9922), .ZN(
        P1_U3261) );
  INV_X1 U11108 ( .A(n9925), .ZN(n9927) );
  OAI21_X1 U11109 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9930) );
  XNOR2_X1 U11110 ( .A(n9930), .B(n9929), .ZN(n9932) );
  AOI21_X1 U11111 ( .B1(n9932), .B2(n9947), .A(n9931), .ZN(n10021) );
  NOR2_X1 U11112 ( .A1(n9949), .A2(n9933), .ZN(n9934) );
  AOI21_X1 U11113 ( .B1(n9968), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9934), .ZN(
        n9935) );
  OAI21_X1 U11114 ( .B1(n9970), .B2(n4557), .A(n9935), .ZN(n9936) );
  INV_X1 U11115 ( .A(n9936), .ZN(n9943) );
  XNOR2_X1 U11116 ( .A(n9938), .B(n9937), .ZN(n10024) );
  OAI211_X1 U11117 ( .C1(n9940), .C2(n4557), .A(n9975), .B(n9939), .ZN(n10020)
         );
  INV_X1 U11118 ( .A(n10020), .ZN(n9941) );
  AOI22_X1 U11119 ( .A1(n10024), .A2(n9957), .B1(n9978), .B2(n9941), .ZN(n9942) );
  OAI211_X1 U11120 ( .C1(n9973), .C2(n10021), .A(n9943), .B(n9942), .ZN(
        P1_U3288) );
  XNOR2_X1 U11121 ( .A(n9945), .B(n9944), .ZN(n9948) );
  AOI21_X1 U11122 ( .B1(n9948), .B2(n9947), .A(n9946), .ZN(n10008) );
  NOR2_X1 U11123 ( .A1(n9949), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9950) );
  AOI21_X1 U11124 ( .B1(n9968), .B2(P1_REG2_REG_3__SCAN_IN), .A(n9950), .ZN(
        n9951) );
  OAI21_X1 U11125 ( .B1(n9970), .B2(n10007), .A(n9951), .ZN(n9952) );
  INV_X1 U11126 ( .A(n9952), .ZN(n9959) );
  XNOR2_X1 U11127 ( .A(n9954), .B(n9953), .ZN(n10011) );
  OAI211_X1 U11128 ( .C1(n9955), .C2(n10007), .A(n7334), .B(n9975), .ZN(n10006) );
  INV_X1 U11129 ( .A(n10006), .ZN(n9956) );
  AOI22_X1 U11130 ( .A1(n10011), .A2(n9957), .B1(n9978), .B2(n9956), .ZN(n9958) );
  OAI211_X1 U11131 ( .C1(n9973), .C2(n10008), .A(n9959), .B(n9958), .ZN(
        P1_U3290) );
  INV_X1 U11132 ( .A(n9960), .ZN(n10089) );
  XNOR2_X1 U11133 ( .A(n7274), .B(n9961), .ZN(n9996) );
  XNOR2_X1 U11134 ( .A(n9962), .B(n7274), .ZN(n9964) );
  NOR2_X1 U11135 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  AOI211_X1 U11136 ( .C1(n10089), .C2(n9996), .A(n9966), .B(n9965), .ZN(n9993)
         );
  AOI22_X1 U11137 ( .A1(n9968), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9967), .ZN(n9969) );
  OAI21_X1 U11138 ( .B1(n9970), .B2(n9992), .A(n9969), .ZN(n9971) );
  INV_X1 U11139 ( .A(n9971), .ZN(n9981) );
  NOR2_X1 U11140 ( .A1(n9973), .A2(n9972), .ZN(n9979) );
  OAI211_X1 U11141 ( .C1(n9992), .C2(n9976), .A(n9975), .B(n9974), .ZN(n9991)
         );
  INV_X1 U11142 ( .A(n9991), .ZN(n9977) );
  AOI22_X1 U11143 ( .A1(n9996), .A2(n9979), .B1(n9978), .B2(n9977), .ZN(n9980)
         );
  OAI211_X1 U11144 ( .C1(n9973), .C2(n9993), .A(n9981), .B(n9980), .ZN(
        P1_U3292) );
  NOR2_X1 U11145 ( .A1(n9990), .A2(n9982), .ZN(P1_U3294) );
  INV_X1 U11146 ( .A(n9990), .ZN(n9988) );
  AND2_X1 U11147 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9988), .ZN(P1_U3295) );
  AND2_X1 U11148 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9988), .ZN(P1_U3296) );
  AND2_X1 U11149 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9988), .ZN(P1_U3297) );
  AND2_X1 U11150 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9988), .ZN(P1_U3298) );
  AND2_X1 U11151 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9988), .ZN(P1_U3299) );
  AND2_X1 U11152 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9988), .ZN(P1_U3300) );
  NOR2_X1 U11153 ( .A1(n9990), .A2(n9983), .ZN(P1_U3301) );
  AND2_X1 U11154 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9988), .ZN(P1_U3302) );
  AND2_X1 U11155 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9988), .ZN(P1_U3303) );
  AND2_X1 U11156 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9988), .ZN(P1_U3304) );
  NOR2_X1 U11157 ( .A1(n9990), .A2(n9984), .ZN(P1_U3305) );
  AND2_X1 U11158 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9988), .ZN(P1_U3306) );
  AND2_X1 U11159 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9988), .ZN(P1_U3307) );
  NOR2_X1 U11160 ( .A1(n9990), .A2(n9985), .ZN(P1_U3308) );
  AND2_X1 U11161 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9988), .ZN(P1_U3309) );
  NOR2_X1 U11162 ( .A1(n9990), .A2(n9986), .ZN(P1_U3310) );
  AND2_X1 U11163 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9988), .ZN(P1_U3311) );
  AND2_X1 U11164 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9988), .ZN(P1_U3312) );
  AND2_X1 U11165 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9988), .ZN(P1_U3313) );
  AND2_X1 U11166 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9988), .ZN(P1_U3314) );
  AND2_X1 U11167 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9988), .ZN(P1_U3315) );
  AND2_X1 U11168 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9988), .ZN(P1_U3316) );
  AND2_X1 U11169 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9988), .ZN(P1_U3317) );
  AND2_X1 U11170 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9988), .ZN(P1_U3318) );
  AND2_X1 U11171 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9988), .ZN(P1_U3319) );
  AND2_X1 U11172 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9988), .ZN(P1_U3320) );
  NOR2_X1 U11173 ( .A1(n9990), .A2(n9987), .ZN(P1_U3321) );
  AND2_X1 U11174 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9988), .ZN(P1_U3322) );
  NOR2_X1 U11175 ( .A1(n9990), .A2(n9989), .ZN(P1_U3323) );
  INV_X1 U11176 ( .A(n10085), .ZN(n10042) );
  OAI21_X1 U11177 ( .B1(n9992), .B2(n10076), .A(n9991), .ZN(n9995) );
  INV_X1 U11178 ( .A(n9993), .ZN(n9994) );
  AOI211_X1 U11179 ( .C1(n10042), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10093) );
  INV_X1 U11180 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9997) );
  AOI22_X1 U11181 ( .A1(n10092), .A2(n10093), .B1(n9997), .B2(n10090), .ZN(
        P1_U3456) );
  INV_X1 U11182 ( .A(n10002), .ZN(n10004) );
  AOI21_X1 U11183 ( .B1(n10083), .B2(n4447), .A(n9998), .ZN(n10000) );
  OAI211_X1 U11184 ( .C1(n10085), .C2(n10002), .A(n10001), .B(n10000), .ZN(
        n10003) );
  AOI21_X1 U11185 ( .B1(n10089), .B2(n10004), .A(n10003), .ZN(n10094) );
  INV_X1 U11186 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U11187 ( .A1(n10092), .A2(n10094), .B1(n10005), .B2(n10090), .ZN(
        P1_U3459) );
  OAI21_X1 U11188 ( .B1(n10007), .B2(n10076), .A(n10006), .ZN(n10010) );
  INV_X1 U11189 ( .A(n10008), .ZN(n10009) );
  AOI211_X1 U11190 ( .C1(n10080), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10096) );
  INV_X1 U11191 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10012) );
  AOI22_X1 U11192 ( .A1(n10092), .A2(n10096), .B1(n10012), .B2(n10090), .ZN(
        P1_U3462) );
  AOI21_X1 U11193 ( .B1(n10083), .B2(n10014), .A(n10013), .ZN(n10016) );
  OAI211_X1 U11194 ( .C1(n10018), .C2(n10017), .A(n10016), .B(n10015), .ZN(
        n10019) );
  INV_X1 U11195 ( .A(n10019), .ZN(n10098) );
  AOI22_X1 U11196 ( .A1(n10092), .A2(n10098), .B1(n6109), .B2(n10090), .ZN(
        P1_U3465) );
  OAI21_X1 U11197 ( .B1(n4557), .B2(n10076), .A(n10020), .ZN(n10023) );
  INV_X1 U11198 ( .A(n10021), .ZN(n10022) );
  AOI211_X1 U11199 ( .C1(n10024), .C2(n10080), .A(n10023), .B(n10022), .ZN(
        n10099) );
  INV_X1 U11200 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10025) );
  AOI22_X1 U11201 ( .A1(n10092), .A2(n10099), .B1(n10025), .B2(n10090), .ZN(
        P1_U3468) );
  OAI211_X1 U11202 ( .C1(n10028), .C2(n10076), .A(n10027), .B(n10026), .ZN(
        n10029) );
  AOI21_X1 U11203 ( .B1(n10080), .B2(n10030), .A(n10029), .ZN(n10100) );
  AOI22_X1 U11204 ( .A1(n10092), .A2(n10100), .B1(n6074), .B2(n10090), .ZN(
        P1_U3471) );
  OR2_X1 U11205 ( .A1(n10031), .A2(n10076), .ZN(n10032) );
  AND2_X1 U11206 ( .A1(n10033), .A2(n10032), .ZN(n10036) );
  NAND2_X1 U11207 ( .A1(n10034), .A2(n10080), .ZN(n10035) );
  AND3_X1 U11208 ( .A1(n10037), .A2(n10036), .A3(n10035), .ZN(n10102) );
  INV_X1 U11209 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U11210 ( .A1(n10092), .A2(n10102), .B1(n10038), .B2(n10090), .ZN(
        P1_U3474) );
  OAI21_X1 U11211 ( .B1(n10040), .B2(n10076), .A(n10039), .ZN(n10045) );
  OAI21_X1 U11212 ( .B1(n10089), .B2(n10042), .A(n10041), .ZN(n10043) );
  INV_X1 U11213 ( .A(n10043), .ZN(n10044) );
  NOR3_X1 U11214 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10103) );
  INV_X1 U11215 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10047) );
  AOI22_X1 U11216 ( .A1(n10092), .A2(n10103), .B1(n10047), .B2(n10090), .ZN(
        P1_U3477) );
  AND2_X1 U11217 ( .A1(n10048), .A2(n10083), .ZN(n10049) );
  NOR2_X1 U11218 ( .A1(n10050), .A2(n10049), .ZN(n10053) );
  NAND2_X1 U11219 ( .A1(n10051), .A2(n10080), .ZN(n10052) );
  AND3_X1 U11220 ( .A1(n10054), .A2(n10053), .A3(n10052), .ZN(n10104) );
  INV_X1 U11221 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11222 ( .A1(n10092), .A2(n10104), .B1(n10055), .B2(n10090), .ZN(
        P1_U3480) );
  OAI211_X1 U11223 ( .C1(n10058), .C2(n10076), .A(n10057), .B(n10056), .ZN(
        n10059) );
  AOI21_X1 U11224 ( .B1(n10060), .B2(n10080), .A(n10059), .ZN(n10105) );
  AOI22_X1 U11225 ( .A1(n10092), .A2(n10105), .B1(n10061), .B2(n10090), .ZN(
        P1_U3483) );
  OAI211_X1 U11226 ( .C1(n10064), .C2(n10076), .A(n10063), .B(n10062), .ZN(
        n10065) );
  AOI21_X1 U11227 ( .B1(n10080), .B2(n10066), .A(n10065), .ZN(n10106) );
  INV_X1 U11228 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10067) );
  AOI22_X1 U11229 ( .A1(n10092), .A2(n10106), .B1(n10067), .B2(n10090), .ZN(
        P1_U3486) );
  OAI211_X1 U11230 ( .C1(n10070), .C2(n10076), .A(n10069), .B(n10068), .ZN(
        n10071) );
  AOI21_X1 U11231 ( .B1(n10080), .B2(n10072), .A(n10071), .ZN(n10107) );
  AOI22_X1 U11232 ( .A1(n10092), .A2(n10107), .B1(n10073), .B2(n10090), .ZN(
        P1_U3489) );
  OAI211_X1 U11233 ( .C1(n10077), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10078) );
  AOI21_X1 U11234 ( .B1(n10080), .B2(n10079), .A(n10078), .ZN(n10108) );
  AOI22_X1 U11235 ( .A1(n10092), .A2(n10108), .B1(n6022), .B2(n10090), .ZN(
        P1_U3492) );
  INV_X1 U11236 ( .A(n10086), .ZN(n10088) );
  AOI211_X1 U11237 ( .C1(n10083), .C2(n6021), .A(n10082), .B(n10081), .ZN(
        n10084) );
  OAI21_X1 U11238 ( .B1(n10086), .B2(n10085), .A(n10084), .ZN(n10087) );
  AOI21_X1 U11239 ( .B1(n10089), .B2(n10088), .A(n10087), .ZN(n10110) );
  INV_X1 U11240 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U11241 ( .A1(n10092), .A2(n10110), .B1(n10091), .B2(n10090), .ZN(
        P1_U3495) );
  AOI22_X1 U11242 ( .A1(n10111), .A2(n10093), .B1(n6094), .B2(n10109), .ZN(
        P1_U3523) );
  AOI22_X1 U11243 ( .A1(n10111), .A2(n10094), .B1(n6100), .B2(n10109), .ZN(
        P1_U3524) );
  INV_X1 U11244 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U11245 ( .A1(n10111), .A2(n10096), .B1(n10095), .B2(n10109), .ZN(
        P1_U3525) );
  AOI22_X1 U11246 ( .A1(n10111), .A2(n10098), .B1(n10097), .B2(n10109), .ZN(
        P1_U3526) );
  AOI22_X1 U11247 ( .A1(n10111), .A2(n10099), .B1(n6121), .B2(n10109), .ZN(
        P1_U3527) );
  AOI22_X1 U11248 ( .A1(n10111), .A2(n10100), .B1(n7082), .B2(n10109), .ZN(
        P1_U3528) );
  INV_X1 U11249 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11250 ( .A1(n10111), .A2(n10102), .B1(n10101), .B2(n10109), .ZN(
        P1_U3529) );
  AOI22_X1 U11251 ( .A1(n10111), .A2(n10103), .B1(n6050), .B2(n10109), .ZN(
        P1_U3530) );
  AOI22_X1 U11252 ( .A1(n10111), .A2(n10104), .B1(n7087), .B2(n10109), .ZN(
        P1_U3531) );
  AOI22_X1 U11253 ( .A1(n10111), .A2(n10105), .B1(n6066), .B2(n10109), .ZN(
        P1_U3532) );
  AOI22_X1 U11254 ( .A1(n10111), .A2(n10106), .B1(n7438), .B2(n10109), .ZN(
        P1_U3533) );
  AOI22_X1 U11255 ( .A1(n10111), .A2(n10107), .B1(n7439), .B2(n10109), .ZN(
        P1_U3534) );
  AOI22_X1 U11256 ( .A1(n10111), .A2(n10108), .B1(n9049), .B2(n10109), .ZN(
        P1_U3535) );
  AOI22_X1 U11257 ( .A1(n10111), .A2(n10110), .B1(n9050), .B2(n10109), .ZN(
        P1_U3536) );
  NAND2_X1 U11258 ( .A1(n10112), .A2(n5017), .ZN(n10113) );
  NAND2_X1 U11259 ( .A1(n10114), .A2(n10113), .ZN(n10117) );
  XNOR2_X1 U11260 ( .A(n10115), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U11261 ( .A1(n10175), .A2(n10117), .B1(n10241), .B2(n10116), .ZN(
        n10120) );
  NAND2_X1 U11262 ( .A1(n10232), .A2(n4584), .ZN(n10119) );
  OAI211_X1 U11263 ( .C1(n10330), .C2(n10163), .A(n10120), .B(n10119), .ZN(
        n10121) );
  INV_X1 U11264 ( .A(n10121), .ZN(n10126) );
  XOR2_X1 U11265 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND2_X1 U11266 ( .A1(n10124), .A2(n10240), .ZN(n10125) );
  OAI211_X1 U11267 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7503), .A(n10126), .B(
        n10125), .ZN(P2_U3183) );
  INV_X1 U11268 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10140) );
  OAI21_X1 U11269 ( .B1(n4531), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10146), .ZN(
        n10129) );
  NOR2_X1 U11270 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10127), .ZN(n10128) );
  AOI21_X1 U11271 ( .B1(n10175), .B2(n10129), .A(n10128), .ZN(n10134) );
  NAND2_X1 U11272 ( .A1(n10232), .A2(n4789), .ZN(n10133) );
  XNOR2_X1 U11273 ( .A(n10130), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n10131) );
  NAND2_X1 U11274 ( .A1(n10241), .A2(n10131), .ZN(n10132) );
  AND3_X1 U11275 ( .A1(n10134), .A2(n10133), .A3(n10132), .ZN(n10139) );
  XOR2_X1 U11276 ( .A(n10136), .B(n10135), .Z(n10137) );
  NAND2_X1 U11277 ( .A1(n10137), .A2(n10240), .ZN(n10138) );
  OAI211_X1 U11278 ( .C1(n10140), .C2(n10163), .A(n10139), .B(n10138), .ZN(
        P2_U3187) );
  INV_X1 U11279 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10164) );
  AOI21_X1 U11280 ( .B1(n10142), .B2(n10141), .A(n4532), .ZN(n10154) );
  INV_X1 U11281 ( .A(n10143), .ZN(n10148) );
  NAND3_X1 U11282 ( .A1(n10146), .A2(n10145), .A3(n10144), .ZN(n10147) );
  AOI21_X1 U11283 ( .B1(n10148), .B2(n10147), .A(n10246), .ZN(n10149) );
  AOI211_X1 U11284 ( .C1(n10232), .C2(n10151), .A(n10150), .B(n10149), .ZN(
        n10152) );
  OAI21_X1 U11285 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10155) );
  INV_X1 U11286 ( .A(n10155), .ZN(n10162) );
  AOI21_X1 U11287 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10160) );
  OR2_X1 U11288 ( .A1(n10160), .A2(n10159), .ZN(n10161) );
  OAI211_X1 U11289 ( .C1(n10164), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        P2_U3188) );
  AOI22_X1 U11290 ( .A1(n10165), .A2(n10232), .B1(P2_ADDR_REG_13__SCAN_IN), 
        .B2(n10231), .ZN(n10181) );
  OAI21_X1 U11291 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10167), .A(n10166), 
        .ZN(n10172) );
  OAI21_X1 U11292 ( .B1(n10170), .B2(n10169), .A(n10168), .ZN(n10171) );
  AOI22_X1 U11293 ( .A1(n10172), .A2(n10241), .B1(n10240), .B2(n10171), .ZN(
        n10180) );
  NAND2_X1 U11294 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n10179)
         );
  INV_X1 U11295 ( .A(n10173), .ZN(n10174) );
  NOR2_X1 U11296 ( .A1(n10174), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10177) );
  OAI21_X1 U11297 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(n10178) );
  NAND4_X1 U11298 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        P2_U3195) );
  AOI22_X1 U11299 ( .A1(n10182), .A2(n10232), .B1(n10231), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n10197) );
  OAI21_X1 U11300 ( .B1(n10185), .B2(n10184), .A(n10183), .ZN(n10190) );
  OAI21_X1 U11301 ( .B1(n10188), .B2(n10187), .A(n10186), .ZN(n10189) );
  AOI22_X1 U11302 ( .A1(n10190), .A2(n10241), .B1(n10240), .B2(n10189), .ZN(
        n10196) );
  NAND2_X1 U11303 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n10195)
         );
  AOI21_X1 U11304 ( .B1(n4512), .B2(n10192), .A(n10191), .ZN(n10193) );
  OR2_X1 U11305 ( .A1(n10193), .A2(n10246), .ZN(n10194) );
  NAND4_X1 U11306 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        P2_U3196) );
  AOI22_X1 U11307 ( .A1(n10198), .A2(n10232), .B1(P2_ADDR_REG_15__SCAN_IN), 
        .B2(n10231), .ZN(n10213) );
  OAI21_X1 U11308 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10200), .A(n10199), 
        .ZN(n10205) );
  OAI21_X1 U11309 ( .B1(n10203), .B2(n10202), .A(n10201), .ZN(n10204) );
  AOI22_X1 U11310 ( .A1(n10205), .A2(n10241), .B1(n10240), .B2(n10204), .ZN(
        n10212) );
  INV_X1 U11311 ( .A(n10206), .ZN(n10211) );
  OR2_X1 U11312 ( .A1(n10209), .A2(n10246), .ZN(n10210) );
  NAND4_X1 U11313 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        P2_U3197) );
  AOI22_X1 U11314 ( .A1(n10214), .A2(n10232), .B1(P2_ADDR_REG_16__SCAN_IN), 
        .B2(n10231), .ZN(n10230) );
  OAI21_X1 U11315 ( .B1(n10217), .B2(n10216), .A(n10215), .ZN(n10222) );
  OAI21_X1 U11316 ( .B1(n10220), .B2(n10219), .A(n10218), .ZN(n10221) );
  AOI22_X1 U11317 ( .A1(n10222), .A2(n10241), .B1(n10240), .B2(n10221), .ZN(
        n10229) );
  AOI21_X1 U11318 ( .B1(n10225), .B2(n10224), .A(n10223), .ZN(n10226) );
  OR2_X1 U11319 ( .A1(n10226), .A2(n10246), .ZN(n10227) );
  NAND4_X1 U11320 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        P2_U3198) );
  AOI22_X1 U11321 ( .A1(n10233), .A2(n10232), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n10231), .ZN(n10250) );
  OAI21_X1 U11322 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10235), .A(n10234), 
        .ZN(n10242) );
  OAI21_X1 U11323 ( .B1(n10238), .B2(n10237), .A(n10236), .ZN(n10239) );
  AOI22_X1 U11324 ( .A1(n10242), .A2(n10241), .B1(n10240), .B2(n10239), .ZN(
        n10249) );
  NAND2_X1 U11325 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10248)
         );
  AOI21_X1 U11326 ( .B1(n10244), .B2(n8478), .A(n10243), .ZN(n10245) );
  OR2_X1 U11327 ( .A1(n10246), .A2(n10245), .ZN(n10247) );
  NAND4_X1 U11328 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        P2_U3199) );
  AOI22_X1 U11329 ( .A1(n10311), .A2(n5042), .B1(n10251), .B2(n10309), .ZN(
        P2_U3390) );
  AND2_X1 U11330 ( .A1(n10252), .A2(n10287), .ZN(n10255) );
  NOR2_X1 U11331 ( .A1(n6848), .A2(n10291), .ZN(n10254) );
  NOR3_X1 U11332 ( .A1(n10255), .A2(n10254), .A3(n10253), .ZN(n10312) );
  AOI22_X1 U11333 ( .A1(n10311), .A2(n5018), .B1(n10312), .B2(n10309), .ZN(
        P2_U3393) );
  OAI22_X1 U11334 ( .A1(n10257), .A2(n10297), .B1(n10256), .B2(n10291), .ZN(
        n10258) );
  NOR2_X1 U11335 ( .A1(n10259), .A2(n10258), .ZN(n10313) );
  AOI22_X1 U11336 ( .A1(n10311), .A2(n5053), .B1(n10313), .B2(n10309), .ZN(
        P2_U3396) );
  INV_X1 U11337 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U11338 ( .A1(n10261), .A2(n10287), .B1(n10308), .B2(n10260), .ZN(
        n10262) );
  AND2_X1 U11339 ( .A1(n10263), .A2(n10262), .ZN(n10314) );
  AOI22_X1 U11340 ( .A1(n10311), .A2(n10264), .B1(n10314), .B2(n10309), .ZN(
        P2_U3399) );
  OR2_X1 U11341 ( .A1(n10265), .A2(n10303), .ZN(n10268) );
  NAND2_X1 U11342 ( .A1(n10266), .A2(n10308), .ZN(n10267) );
  AND2_X1 U11343 ( .A1(n10268), .A2(n10267), .ZN(n10270) );
  AND2_X1 U11344 ( .A1(n10270), .A2(n10269), .ZN(n10315) );
  AOI22_X1 U11345 ( .A1(n10311), .A2(n5092), .B1(n10315), .B2(n10309), .ZN(
        P2_U3402) );
  AOI22_X1 U11346 ( .A1(n10273), .A2(n10272), .B1(n10308), .B2(n10271), .ZN(
        n10274) );
  AND2_X1 U11347 ( .A1(n10275), .A2(n10274), .ZN(n10317) );
  AOI22_X1 U11348 ( .A1(n10311), .A2(n5114), .B1(n10317), .B2(n10309), .ZN(
        P2_U3405) );
  OAI22_X1 U11349 ( .A1(n10277), .A2(n10303), .B1(n10276), .B2(n10291), .ZN(
        n10278) );
  INV_X1 U11350 ( .A(n10278), .ZN(n10280) );
  AND2_X1 U11351 ( .A1(n10280), .A2(n10279), .ZN(n10318) );
  AOI22_X1 U11352 ( .A1(n10311), .A2(n5140), .B1(n10318), .B2(n10309), .ZN(
        P2_U3408) );
  INV_X1 U11353 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10285) );
  OAI22_X1 U11354 ( .A1(n10282), .A2(n10297), .B1(n10281), .B2(n10291), .ZN(
        n10283) );
  NOR2_X1 U11355 ( .A1(n10284), .A2(n10283), .ZN(n10319) );
  AOI22_X1 U11356 ( .A1(n10311), .A2(n10285), .B1(n10319), .B2(n10309), .ZN(
        P2_U3411) );
  AOI22_X1 U11357 ( .A1(n10288), .A2(n10287), .B1(n10308), .B2(n10286), .ZN(
        n10289) );
  AND2_X1 U11358 ( .A1(n10290), .A2(n10289), .ZN(n10320) );
  AOI22_X1 U11359 ( .A1(n10311), .A2(n5200), .B1(n10320), .B2(n10309), .ZN(
        P2_U3414) );
  OAI22_X1 U11360 ( .A1(n10293), .A2(n10297), .B1(n10292), .B2(n10291), .ZN(
        n10294) );
  NOR2_X1 U11361 ( .A1(n10295), .A2(n10294), .ZN(n10321) );
  AOI22_X1 U11362 ( .A1(n10311), .A2(n10296), .B1(n10321), .B2(n10309), .ZN(
        P2_U3417) );
  INV_X1 U11363 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10302) );
  NOR2_X1 U11364 ( .A1(n10298), .A2(n10297), .ZN(n10299) );
  AOI211_X1 U11365 ( .C1(n10308), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10322) );
  AOI22_X1 U11366 ( .A1(n10311), .A2(n10302), .B1(n10322), .B2(n10309), .ZN(
        P2_U3420) );
  NOR2_X1 U11367 ( .A1(n10304), .A2(n10303), .ZN(n10306) );
  AOI211_X1 U11368 ( .C1(n10308), .C2(n10307), .A(n10306), .B(n10305), .ZN(
        n10324) );
  AOI22_X1 U11369 ( .A1(n10311), .A2(n10310), .B1(n10324), .B2(n10309), .ZN(
        P2_U3423) );
  AOI22_X1 U11370 ( .A1(n10325), .A2(n10312), .B1(n5021), .B2(n10323), .ZN(
        P2_U3460) );
  AOI22_X1 U11371 ( .A1(n10325), .A2(n10313), .B1(n7141), .B2(n10323), .ZN(
        P2_U3461) );
  AOI22_X1 U11372 ( .A1(n10325), .A2(n10314), .B1(n5075), .B2(n10323), .ZN(
        P2_U3462) );
  AOI22_X1 U11373 ( .A1(n10325), .A2(n10315), .B1(n7140), .B2(n10323), .ZN(
        P2_U3463) );
  INV_X1 U11374 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U11375 ( .A1(n10325), .A2(n10317), .B1(n10316), .B2(n10323), .ZN(
        P2_U3464) );
  AOI22_X1 U11376 ( .A1(n10325), .A2(n10318), .B1(n7374), .B2(n10323), .ZN(
        P2_U3465) );
  AOI22_X1 U11377 ( .A1(n10325), .A2(n10319), .B1(n7656), .B2(n10323), .ZN(
        P2_U3466) );
  AOI22_X1 U11378 ( .A1(n10325), .A2(n10320), .B1(n7658), .B2(n10323), .ZN(
        P2_U3467) );
  AOI22_X1 U11379 ( .A1(n10325), .A2(n10321), .B1(n7643), .B2(n10323), .ZN(
        P2_U3468) );
  AOI22_X1 U11380 ( .A1(n10325), .A2(n10322), .B1(n7647), .B2(n10323), .ZN(
        P2_U3469) );
  AOI22_X1 U11381 ( .A1(n10325), .A2(n10324), .B1(n5255), .B2(n10323), .ZN(
        P2_U3470) );
  OAI222_X1 U11382 ( .A1(n10330), .A2(n10329), .B1(n10330), .B2(n10328), .C1(
        n10327), .C2(n10326), .ZN(ADD_1068_U5) );
  AOI21_X1 U11383 ( .B1(n10332), .B2(n7185), .A(n10331), .ZN(ADD_1068_U46) );
  AOI21_X1 U11384 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(n10336) );
  XOR2_X1 U11385 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10336), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11386 ( .B1(n10339), .B2(n10338), .A(n10337), .ZN(ADD_1068_U56) );
  OAI21_X1 U11387 ( .B1(n10342), .B2(n10341), .A(n10340), .ZN(ADD_1068_U57) );
  OAI21_X1 U11388 ( .B1(n10345), .B2(n10344), .A(n10343), .ZN(ADD_1068_U58) );
  OAI21_X1 U11389 ( .B1(n10348), .B2(n10347), .A(n10346), .ZN(ADD_1068_U59) );
  OAI21_X1 U11390 ( .B1(n10351), .B2(n10350), .A(n10349), .ZN(ADD_1068_U60) );
  OAI21_X1 U11391 ( .B1(n10354), .B2(n10353), .A(n10352), .ZN(ADD_1068_U61) );
  OAI21_X1 U11392 ( .B1(n10357), .B2(n10356), .A(n10355), .ZN(ADD_1068_U62) );
  OAI21_X1 U11393 ( .B1(n10360), .B2(n10359), .A(n10358), .ZN(ADD_1068_U63) );
  OAI21_X1 U11394 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(ADD_1068_U51) );
  OAI21_X1 U11395 ( .B1(n10366), .B2(n10365), .A(n10364), .ZN(ADD_1068_U47) );
  OAI21_X1 U11396 ( .B1(n10369), .B2(n10368), .A(n10367), .ZN(ADD_1068_U50) );
  OAI21_X1 U11397 ( .B1(n10372), .B2(n10371), .A(n10370), .ZN(ADD_1068_U49) );
  OAI21_X1 U11398 ( .B1(n10375), .B2(n10374), .A(n10373), .ZN(ADD_1068_U48) );
  AOI21_X1 U11399 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(ADD_1068_U54) );
  AOI21_X1 U11400 ( .B1(n10381), .B2(n10380), .A(n10379), .ZN(ADD_1068_U53) );
  OAI21_X1 U11401 ( .B1(n10384), .B2(n10383), .A(n10382), .ZN(ADD_1068_U52) );
  NOR2_X1 U7318 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5699) );
  OAI22_X1 U4945 ( .A1(n8212), .A2(n8927), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8211), .ZN(n8213) );
  CLKBUF_X1 U4951 ( .A(n4904), .Z(n4903) );
  NOR2_X1 U4959 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5705) );
  CLKBUF_X2 U4989 ( .A(n5819), .Z(n4443) );
  NAND2_X1 U6108 ( .A1(n8293), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5012) );
  INV_X2 U7324 ( .A(n8708), .ZN(n8700) );
endmodule

