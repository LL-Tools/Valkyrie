

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4420, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616;

  NAND2_X1 U4926 ( .A1(n9655), .A2(n9653), .ZN(n9689) );
  INV_X1 U4927 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10311) );
  AND2_X1 U4928 ( .A1(n5903), .A2(n5902), .ZN(n9431) );
  AND2_X1 U4929 ( .A1(n10339), .A2(n10347), .ZN(n5186) );
  INV_X1 U4930 ( .A(n8066), .ZN(n10230) );
  INV_X1 U4931 ( .A(n9791), .ZN(n9792) );
  NAND2_X2 U4932 ( .A1(n5624), .A2(n5623), .ZN(n8026) );
  INV_X1 U4933 ( .A(n9370), .ZN(n10245) );
  CLKBUF_X1 U4934 ( .A(n6287), .Z(n6545) );
  INV_X1 U4935 ( .A(n5582), .ZN(n6919) );
  INV_X1 U4936 ( .A(n7876), .ZN(n5815) );
  CLKBUF_X1 U4937 ( .A(n5509), .Z(n4439) );
  AND3_X1 U4938 ( .A1(n6249), .A2(n4468), .A3(n6250), .ZN(n7958) );
  XNOR2_X1 U4939 ( .A(n5501), .B(n5500), .ZN(n7106) );
  AND2_X1 U4940 ( .A1(n5434), .A2(n10322), .ZN(n5509) );
  CLKBUF_X2 U4941 ( .A(n6286), .Z(n4430) );
  AND2_X1 U4942 ( .A1(n6164), .A2(n6165), .ZN(n6287) );
  AND2_X1 U4943 ( .A1(n6244), .A2(n4431), .ZN(n6553) );
  NAND2_X1 U4944 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5554) );
  AND2_X1 U4945 ( .A1(n6022), .A2(n4540), .ZN(n10310) );
  INV_X2 U4946 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10312) );
  CLKBUF_X1 U4948 ( .A(n9805), .Z(n4420) );
  NOR2_X1 U4949 ( .A1(n6085), .A2(n8005), .ZN(n9805) );
  AND2_X1 U4950 ( .A1(n5201), .A2(n9705), .ZN(n7917) );
  OAI21_X1 U4951 ( .B1(n5331), .B2(n6073), .A(n5012), .ZN(n5201) );
  INV_X1 U4954 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4955 ( .A(n7888), .ZN(n9660) );
  NOR2_X1 U4956 ( .A1(n7524), .A2(n5336), .ZN(n5335) );
  INV_X1 U4957 ( .A(n9345), .ZN(n8141) );
  OR2_X1 U4958 ( .A1(n5965), .A2(n9539), .ZN(n5986) );
  INV_X1 U4959 ( .A(n6453), .ZN(n6557) );
  NAND2_X1 U4960 ( .A1(n7597), .A2(n6612), .ZN(n7659) );
  INV_X1 U4961 ( .A(n7963), .ZN(n6803) );
  INV_X2 U4962 ( .A(n5508), .ZN(n6081) );
  INV_X1 U4963 ( .A(n9406), .ZN(n7920) );
  OR2_X1 U4964 ( .A1(n10036), .A2(n5905), .ZN(n4955) );
  INV_X1 U4965 ( .A(n7808), .ZN(n10439) );
  CLKBUF_X3 U4966 ( .A(n6428), .Z(n6453) );
  NAND2_X1 U4968 ( .A1(n5589), .A2(n5588), .ZN(n7528) );
  NAND2_X1 U4969 ( .A1(n4611), .A2(n5408), .ZN(n9477) );
  INV_X1 U4970 ( .A(n4438), .ZN(n5625) );
  AND2_X1 U4971 ( .A1(n6001), .A2(n5987), .ZN(n10002) );
  INV_X1 U4972 ( .A(n7375), .ZN(n6694) );
  AOI21_X2 U4973 ( .B1(n10002), .B2(n6083), .A(n5991), .ZN(n9538) );
  NAND4_X2 U4974 ( .A1(n5487), .A2(n4472), .A3(n5486), .A4(n5403), .ZN(n9838)
         );
  BUF_X1 U4975 ( .A(n6286), .Z(n4429) );
  AND3_X1 U4976 ( .A1(n4642), .A2(n4641), .A3(n9608), .ZN(n4424) );
  OAI21_X2 U4977 ( .B1(n9477), .B2(n5054), .A(n5052), .ZN(n4610) );
  NOR2_X2 U4978 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n6102) );
  XNOR2_X2 U4979 ( .A(n6141), .B(n6158), .ZN(n6676) );
  XNOR2_X2 U4980 ( .A(n5542), .B(SI_4_), .ZN(n5540) );
  OAI211_X1 U4981 ( .C1(n4731), .C2(n4730), .A(n4728), .B(n4726), .ZN(n6859)
         );
  NAND2_X1 U4982 ( .A1(n8814), .A2(n8815), .ZN(n4731) );
  OR2_X2 U4983 ( .A1(n5576), .A2(n5485), .ZN(n5403) );
  NAND2_X2 U4984 ( .A1(n5323), .A2(n5321), .ZN(n7480) );
  NAND2_X2 U4985 ( .A1(n8165), .A2(n9345), .ZN(n7198) );
  BUF_X8 U4986 ( .A(n6889), .Z(n6142) );
  BUF_X8 U4987 ( .A(n6142), .Z(n4956) );
  BUF_X1 U4988 ( .A(n9196), .Z(n4425) );
  OAI21_X2 U4989 ( .B1(n5020), .B2(n5021), .A(n6391), .ZN(n6418) );
  AOI22_X2 U4990 ( .A1(n8421), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n8420), .B2(
        n8419), .ZN(n8441) );
  OAI211_X2 U4991 ( .C1(n9656), .C2(n9716), .A(n9707), .B(n9791), .ZN(n9657)
         );
  OR2_X2 U4992 ( .A1(n5786), .A2(n4973), .ZN(n4967) );
  OAI222_X1 U4994 ( .A1(P1_U3086), .A2(n7106), .B1(n10335), .B2(n6899), .C1(
        n6896), .C2(n10332), .ZN(P1_U3353) );
  NAND2_X4 U4995 ( .A1(n4658), .A2(n5816), .ZN(n10206) );
  OR2_X2 U4996 ( .A1(n10027), .A2(n10026), .ZN(n10182) );
  NAND2_X1 U4997 ( .A1(n4433), .A2(n4431), .ZN(n4426) );
  NAND2_X2 U4998 ( .A1(n4433), .A2(n4431), .ZN(n7876) );
  AND2_X2 U4999 ( .A1(n4943), .A2(n4942), .ZN(n7849) );
  OAI21_X2 U5000 ( .B1(n6731), .B2(n8335), .A(n8245), .ZN(n8299) );
  AOI21_X2 U5001 ( .B1(n5636), .B2(n4441), .A(n5023), .ZN(n5022) );
  XNOR2_X2 U5002 ( .A(n5455), .B(n5454), .ZN(n6972) );
  NOR2_X2 U5003 ( .A1(n7917), .A2(n9689), .ZN(n7916) );
  NAND2_X2 U5004 ( .A1(n9296), .A2(n6164), .ZN(n6428) );
  OAI211_X2 U5005 ( .C1(n5498), .C2(n5497), .A(n5496), .B(n5495), .ZN(n5520)
         );
  BUF_X4 U5006 ( .A(n5552), .Z(n4436) );
  OAI21_X2 U5007 ( .B1(n7916), .B2(n5375), .A(n5378), .ZN(n7891) );
  AOI22_X2 U5008 ( .A1(n8465), .A2(n8464), .B1(n8463), .B2(n8462), .ZN(n8490)
         );
  AND3_X1 U5009 ( .A1(n6857), .A2(n6860), .A3(n10548), .ZN(n4769) );
  AND3_X1 U5010 ( .A1(n6857), .A2(n6860), .A3(n10557), .ZN(n4890) );
  OAI21_X1 U5011 ( .B1(n6859), .B2(n9069), .A(n6855), .ZN(n6856) );
  AND2_X1 U5012 ( .A1(n7536), .A2(n7535), .ZN(n9364) );
  NOR2_X2 U5013 ( .A1(n9005), .A2(n9022), .ZN(n6592) );
  NAND2_X1 U5014 ( .A1(n7799), .A2(n9571), .ZN(n7645) );
  NAND2_X1 U5015 ( .A1(n6621), .A2(n6370), .ZN(n9005) );
  NAND2_X1 U5016 ( .A1(n7704), .A2(n7703), .ZN(n7702) );
  NAND2_X1 U5017 ( .A1(n9571), .A2(n9746), .ZN(n7798) );
  CLKBUF_X2 U5018 ( .A(n4599), .Z(n4428) );
  INV_X1 U5019 ( .A(n6886), .ZN(n4599) );
  NAND2_X1 U5020 ( .A1(n6694), .A2(n10533), .ZN(n6581) );
  CLKBUF_X2 U5021 ( .A(n6684), .Z(n4435) );
  INV_X2 U5022 ( .A(n7958), .ZN(n8339) );
  INV_X1 U5023 ( .A(n9063), .ZN(n7595) );
  INV_X2 U5024 ( .A(n9838), .ZN(n7201) );
  INV_X2 U5025 ( .A(n5421), .ZN(n8108) );
  CLKBUF_X2 U5026 ( .A(n5509), .Z(n4438) );
  INV_X1 U5027 ( .A(n9784), .ZN(n4613) );
  NAND2_X2 U5028 ( .A1(n5582), .A2(n4956), .ZN(n5587) );
  INV_X2 U5029 ( .A(n9991), .ZN(n9800) );
  NOR2_X1 U5030 ( .A1(n6671), .A2(n6670), .ZN(n7869) );
  AND2_X1 U5031 ( .A1(n4859), .A2(n4834), .ZN(n4524) );
  OR2_X1 U5032 ( .A1(n5068), .A2(n6656), .ZN(n4835) );
  AOI211_X1 U5033 ( .C1(n6090), .C2(n7920), .A(n7929), .B(n7930), .ZN(n7923)
         );
  AND2_X1 U5034 ( .A1(n7884), .A2(n6011), .ZN(n7992) );
  NAND2_X1 U5035 ( .A1(n4731), .A2(n4727), .ZN(n4726) );
  NAND2_X1 U5036 ( .A1(n9397), .A2(n9398), .ZN(n9531) );
  OR2_X1 U5037 ( .A1(n10177), .A2(n10164), .ZN(n4941) );
  XNOR2_X1 U5038 ( .A(n10006), .B(n10005), .ZN(n10177) );
  NAND2_X1 U5039 ( .A1(n5244), .A2(n6009), .ZN(n7884) );
  OAI21_X1 U5040 ( .B1(n8186), .B2(n8188), .A(n8253), .ZN(n8189) );
  NAND2_X1 U5041 ( .A1(n9428), .A2(n8149), .ZN(n9397) );
  INV_X1 U5042 ( .A(n5414), .ZN(n4730) );
  AOI21_X1 U5043 ( .B1(n8859), .B2(n9061), .A(n4881), .ZN(n9208) );
  OR2_X1 U5044 ( .A1(n10044), .A2(n6073), .ZN(n5016) );
  NOR2_X1 U5045 ( .A1(n5009), .A2(n4512), .ZN(n5008) );
  AND2_X1 U5046 ( .A1(n7878), .A2(n7877), .ZN(n10166) );
  NAND2_X1 U5047 ( .A1(n6144), .A2(n6143), .ZN(n9177) );
  OR2_X1 U5048 ( .A1(n7886), .A2(n7885), .ZN(n9698) );
  NAND2_X1 U5049 ( .A1(n6741), .A2(n6740), .ZN(n8275) );
  NAND2_X1 U5050 ( .A1(n7874), .A2(n7873), .ZN(n9730) );
  AND2_X1 U5051 ( .A1(n4717), .A2(n5144), .ZN(n8833) );
  NAND2_X1 U5052 ( .A1(n9379), .A2(n4612), .ZN(n4611) );
  OR2_X1 U5053 ( .A1(n6834), .A2(n4550), .ZN(n4717) );
  XNOR2_X1 U5054 ( .A(n6132), .B(n6131), .ZN(n9291) );
  OAI21_X1 U5055 ( .B1(n6552), .B2(n6551), .A(n6129), .ZN(n6132) );
  AND2_X1 U5056 ( .A1(n10014), .A2(n5397), .ZN(n7899) );
  AOI21_X1 U5057 ( .B1(n5314), .B2(n5317), .A(n5312), .ZN(n5311) );
  AND2_X1 U5058 ( .A1(n5279), .A2(n6644), .ZN(n5278) );
  NOR2_X1 U5059 ( .A1(n9941), .A2(n4567), .ZN(n9956) );
  NAND2_X1 U5060 ( .A1(n4700), .A2(n4492), .ZN(n8917) );
  NAND2_X1 U5061 ( .A1(n10133), .A2(n6064), .ZN(n10122) );
  XNOR2_X1 U5062 ( .A(n6115), .B(n6114), .ZN(n8004) );
  NOR2_X1 U5063 ( .A1(n8452), .A2(n8453), .ZN(n8472) );
  NAND2_X1 U5064 ( .A1(n5160), .A2(n5162), .ZN(n8924) );
  AND2_X1 U5065 ( .A1(n4981), .A2(n4571), .ZN(n8772) );
  NAND2_X1 U5066 ( .A1(n9463), .A2(n5344), .ZN(n5343) );
  INV_X1 U5067 ( .A(n5342), .ZN(n5341) );
  OR2_X1 U5068 ( .A1(n8116), .A2(n9376), .ZN(n5408) );
  NAND2_X1 U5069 ( .A1(n5996), .A2(n5995), .ZN(n6115) );
  NAND2_X1 U5070 ( .A1(n5913), .A2(n5912), .ZN(n6074) );
  NAND2_X1 U5071 ( .A1(n5978), .A2(n5977), .ZN(n5994) );
  NAND2_X1 U5072 ( .A1(n5906), .A2(n5892), .ZN(n7865) );
  NAND2_X1 U5073 ( .A1(n5957), .A2(n5956), .ZN(n5976) );
  AND2_X1 U5074 ( .A1(n4946), .A2(n4945), .ZN(n7817) );
  NAND2_X1 U5075 ( .A1(n4854), .A2(n4853), .ZN(n7819) );
  NAND2_X1 U5076 ( .A1(n7684), .A2(n7683), .ZN(n7682) );
  NAND2_X1 U5077 ( .A1(n4443), .A2(n5046), .ZN(n5044) );
  NAND2_X1 U5078 ( .A1(n5846), .A2(n5845), .ZN(n10194) );
  AND2_X1 U5079 ( .A1(n9769), .A2(n9771), .ZN(n10093) );
  NAND2_X1 U5080 ( .A1(n5870), .A2(n5869), .ZN(n9562) );
  NAND2_X1 U5081 ( .A1(n9768), .A2(n9625), .ZN(n10101) );
  AOI21_X1 U5082 ( .B1(n4916), .B2(n4919), .A(n4914), .ZN(n4913) );
  NAND2_X1 U5083 ( .A1(n6456), .A2(n6455), .ZN(n9238) );
  NAND2_X1 U5084 ( .A1(n5790), .A2(n5789), .ZN(n6067) );
  NOR2_X1 U5085 ( .A1(n6376), .A2(n4428), .ZN(n4808) );
  NAND2_X1 U5086 ( .A1(n5733), .A2(n5732), .ZN(n10225) );
  AND2_X1 U5087 ( .A1(n5035), .A2(n4533), .ZN(n7293) );
  OR2_X1 U5088 ( .A1(n10230), .A2(n5389), .ZN(n5388) );
  NAND2_X1 U5089 ( .A1(n10349), .A2(n10474), .ZN(n7822) );
  XNOR2_X1 U5090 ( .A(n9276), .B(n9046), .ZN(n9020) );
  OR2_X1 U5091 ( .A1(n10235), .A2(n8062), .ZN(n9758) );
  NAND2_X1 U5092 ( .A1(n8039), .A2(n8037), .ZN(n9594) );
  AND2_X1 U5093 ( .A1(n5004), .A2(n5003), .ZN(n7624) );
  OR2_X2 U5094 ( .A1(n10240), .A2(n9605), .ZN(n9590) );
  AND3_X1 U5095 ( .A1(n5109), .A2(n9575), .A3(n4536), .ZN(n4895) );
  NAND2_X1 U5096 ( .A1(n4934), .A2(n5642), .ZN(n8039) );
  NAND2_X1 U5097 ( .A1(n5663), .A2(n5662), .ZN(n9603) );
  AND2_X1 U5098 ( .A1(n9581), .A2(n9591), .ZN(n9678) );
  AND2_X2 U5099 ( .A1(n7341), .A2(n9087), .ZN(n8981) );
  NAND2_X1 U5100 ( .A1(n6210), .A2(n6209), .ZN(n9155) );
  NAND2_X1 U5101 ( .A1(n5698), .A2(n5697), .ZN(n10235) );
  NAND2_X2 U5102 ( .A1(n5680), .A2(n5679), .ZN(n10240) );
  NAND2_X1 U5103 ( .A1(n4629), .A2(n4627), .ZN(n5786) );
  OR2_X1 U5104 ( .A1(n7681), .A2(n7655), .ZN(n9034) );
  XNOR2_X1 U5105 ( .A(n5726), .B(n5724), .ZN(n7132) );
  AND2_X1 U5106 ( .A1(n9583), .A2(n9584), .ZN(n7782) );
  AND2_X1 U5107 ( .A1(n4809), .A2(n4600), .ZN(n6270) );
  NAND2_X1 U5108 ( .A1(n5896), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5914) );
  OAI211_X1 U5109 ( .C1(n5636), .C2(n4657), .A(n4656), .B(n4654), .ZN(n6934)
         );
  NOR2_X2 U5110 ( .A1(n10367), .A2(n9527), .ZN(n10368) );
  NAND2_X1 U5111 ( .A1(n7702), .A2(n5197), .ZN(n9570) );
  OR2_X1 U5112 ( .A1(n9076), .A2(n7595), .ZN(n9032) );
  XNOR2_X1 U5113 ( .A(n5022), .B(n4517), .ZN(n6947) );
  BUF_X4 U5114 ( .A(n6693), .Z(n7967) );
  NAND2_X1 U5115 ( .A1(n6324), .A2(n6323), .ZN(n9076) );
  NAND2_X1 U5116 ( .A1(n4796), .A2(n10439), .ZN(n10367) );
  NAND2_X1 U5117 ( .A1(n5634), .A2(n5633), .ZN(n5636) );
  INV_X1 U5118 ( .A(n7528), .ZN(n10455) );
  NOR2_X1 U5119 ( .A1(n7559), .A2(n7560), .ZN(n7621) );
  NAND2_X1 U5120 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  INV_X1 U5121 ( .A(n8137), .ZN(n8163) );
  AND2_X1 U5122 ( .A1(n5141), .A2(n7364), .ZN(n6804) );
  AND2_X1 U5123 ( .A1(n6052), .A2(n6053), .ZN(n5197) );
  NAND2_X1 U5124 ( .A1(n6803), .A2(n8340), .ZN(n6260) );
  INV_X2 U5125 ( .A(n8165), .ZN(n9342) );
  BUF_X1 U5126 ( .A(n6684), .Z(n4434) );
  CLKBUF_X1 U5127 ( .A(n9551), .Z(n9522) );
  INV_X1 U5128 ( .A(n7596), .ZN(n8337) );
  AND2_X1 U5129 ( .A1(n4686), .A2(n4685), .ZN(n7553) );
  NAND2_X1 U5130 ( .A1(n4529), .A2(n4449), .ZN(n9837) );
  AND4_X2 U5131 ( .A1(n6265), .A2(n6263), .A3(n6264), .A4(n6262), .ZN(n7375)
         );
  INV_X1 U5132 ( .A(n7203), .ZN(n10426) );
  INV_X1 U5133 ( .A(n6257), .ZN(n7352) );
  XNOR2_X1 U5134 ( .A(n6181), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6684) );
  CLKBUF_X1 U5135 ( .A(n6257), .Z(n8340) );
  NAND2_X1 U5136 ( .A1(n4471), .A2(n5561), .ZN(n9836) );
  NAND4_X1 U5137 ( .A1(n6331), .A2(n6330), .A3(n6329), .A4(n6328), .ZN(n9063)
         );
  NAND2_X1 U5138 ( .A1(n5507), .A2(n5506), .ZN(n7203) );
  AND4_X1 U5139 ( .A1(n5632), .A2(n5631), .A3(n5630), .A4(n5629), .ZN(n7668)
         );
  AND4_X1 U5140 ( .A1(n5581), .A2(n5580), .A3(n5579), .A4(n5578), .ZN(n7526)
         );
  NAND2_X1 U5141 ( .A1(n6180), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U5142 ( .A1(n5545), .A2(n5544), .ZN(n4625) );
  AND4_X1 U5143 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n7538)
         );
  AND3_X1 U5144 ( .A1(n6256), .A2(n6255), .A3(n6254), .ZN(n7357) );
  NAND4_X1 U5145 ( .A1(n6229), .A2(n6228), .A3(n6230), .A4(n6227), .ZN(n6257)
         );
  NAND2_X1 U5146 ( .A1(n7829), .A2(n8794), .ZN(n6685) );
  NAND2_X1 U5147 ( .A1(n6666), .A2(n6672), .ZN(n6682) );
  OAI211_X1 U5148 ( .C1(n6895), .C2(n4426), .A(n5456), .B(n5457), .ZN(n4772)
         );
  XNOR2_X1 U5149 ( .A(n6179), .B(n6178), .ZN(n7829) );
  AOI21_X2 U5150 ( .B1(n7066), .B2(n9806), .A(n7072), .ZN(n7067) );
  CLKBUF_X1 U5151 ( .A(n6275), .Z(n4768) );
  OR2_X1 U5152 ( .A1(n6275), .A2(n7312), .ZN(n6227) );
  CLKBUF_X1 U5153 ( .A(n5572), .Z(n6083) );
  NAND2_X1 U5154 ( .A1(n6111), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6179) );
  INV_X2 U5155 ( .A(n6306), .ZN(n6472) );
  INV_X1 U5156 ( .A(n4437), .ZN(n5576) );
  INV_X1 U5157 ( .A(n9787), .ZN(n9806) );
  NAND2_X1 U5158 ( .A1(n4897), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n6666) );
  OR2_X1 U5159 ( .A1(n5587), .A2(n6899), .ZN(n5479) );
  NAND2_X1 U5160 ( .A1(n6165), .A2(n9299), .ZN(n6286) );
  NAND2_X1 U5161 ( .A1(n6043), .A2(n6013), .ZN(n7066) );
  AOI21_X1 U5162 ( .B1(n5300), .B2(n4760), .A(n7186), .ZN(n7232) );
  NAND2_X1 U5163 ( .A1(n9784), .A2(n9800), .ZN(n9787) );
  XNOR2_X1 U5164 ( .A(n6112), .B(n6113), .ZN(n8794) );
  AND2_X1 U5165 ( .A1(n5434), .A2(n5433), .ZN(n5572) );
  OR3_X2 U5166 ( .A1(n10328), .A2(n10336), .A3(n10331), .ZN(n7205) );
  INV_X1 U5167 ( .A(n6244), .ZN(n6454) );
  CLKBUF_X1 U5168 ( .A(n6084), .Z(n8005) );
  XNOR2_X1 U5169 ( .A(n6029), .B(n6028), .ZN(n10328) );
  INV_X1 U5170 ( .A(n5654), .ZN(n5023) );
  OAI21_X1 U5171 ( .B1(n5432), .B2(P1_IR_REG_29__SCAN_IN), .A(n4694), .ZN(
        n10322) );
  NAND2_X1 U5172 ( .A1(n9292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5159) );
  INV_X1 U5173 ( .A(n5434), .ZN(n10318) );
  NAND2_X1 U5174 ( .A1(n6027), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6029) );
  NAND2_X1 U5175 ( .A1(n6027), .A2(n6021), .ZN(n10331) );
  NAND2_X1 U5176 ( .A1(n4713), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U5177 ( .A1(n5813), .A2(n5812), .ZN(n6016) );
  XNOR2_X1 U5178 ( .A(n5593), .B(SI_7_), .ZN(n5590) );
  NAND2_X1 U5179 ( .A1(n5449), .A2(n5448), .ZN(n6242) );
  OR2_X1 U5180 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U5181 ( .A1(n6020), .A2(n6019), .ZN(n6027) );
  NAND2_X2 U5182 ( .A1(n4431), .A2(P2_U3151), .ZN(n9307) );
  AND2_X1 U5183 ( .A1(n6022), .A2(n5128), .ZN(n5439) );
  NAND2_X1 U5184 ( .A1(n6140), .A2(n4745), .ZN(n4746) );
  AND2_X1 U5185 ( .A1(n6140), .A2(n6158), .ZN(n4712) );
  AND2_X1 U5186 ( .A1(n4513), .A2(n4699), .ZN(n6022) );
  NAND2_X1 U5187 ( .A1(n6253), .A2(n6252), .ZN(n7183) );
  NOR2_X1 U5188 ( .A1(n6105), .A2(n6106), .ZN(n6137) );
  AND4_X1 U5189 ( .A1(n6135), .A2(n6134), .A3(n6107), .A4(n6133), .ZN(n6136)
         );
  AND4_X1 U5190 ( .A1(n4604), .A2(n4603), .A3(n4602), .A4(n4601), .ZN(n5423)
         );
  NOR2_X1 U5191 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(n4469), .ZN(n5400) );
  AND2_X1 U5192 ( .A1(n5430), .A2(n5444), .ZN(n5130) );
  AND3_X1 U5193 ( .A1(n4751), .A2(n4978), .A3(n4931), .ZN(n4724) );
  NAND2_X1 U5194 ( .A1(n7743), .A2(n5328), .ZN(n5327) );
  NAND4_X1 U5195 ( .A1(n6379), .A2(n6102), .A3(n6101), .A4(n6216), .ZN(n6106)
         );
  AND2_X1 U5196 ( .A1(n8579), .A2(n6100), .ZN(n5277) );
  AND3_X2 U5197 ( .A1(n5601), .A2(n5330), .A3(n5513), .ZN(n5517) );
  INV_X1 U5198 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8579) );
  INV_X1 U5199 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5749) );
  INV_X4 U5200 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5201 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6404) );
  INV_X1 U5202 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8661) );
  INV_X1 U5203 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8578) );
  INV_X1 U5204 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6138) );
  INV_X1 U5205 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8573) );
  NOR2_X1 U5206 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5770) );
  NOR2_X1 U5207 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4604) );
  NOR2_X1 U5208 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4603) );
  NOR2_X1 U5209 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4602) );
  NOR2_X1 U5210 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4601) );
  INV_X1 U5211 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8556) );
  NOR2_X2 U5212 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5601) );
  AND2_X1 U5213 ( .A1(n5331), .A2(n4521), .ZN(n10044) );
  OR2_X2 U5214 ( .A1(n6444), .A2(n6443), .ZN(n5034) );
  INV_X1 U5215 ( .A(n10374), .ZN(n4846) );
  NOR2_X1 U5216 ( .A1(n6997), .A2(n6996), .ZN(n7028) );
  NAND2_X2 U5217 ( .A1(n5262), .A2(n5263), .ZN(n8914) );
  OR2_X1 U5218 ( .A1(n5601), .A2(n10312), .ZN(n5501) );
  OR2_X2 U5219 ( .A1(n9347), .A2(n7892), .ZN(n7888) );
  BUF_X4 U5220 ( .A(n8138), .Z(n4427) );
  INV_X1 U5221 ( .A(n5421), .ZN(n8138) );
  AND2_X1 U5222 ( .A1(n6248), .A2(n4844), .ZN(n4468) );
  AOI21_X2 U5223 ( .B1(n4846), .B2(n6054), .A(n4845), .ZN(n7799) );
  AOI21_X2 U5224 ( .B1(n8299), .B2(n4903), .A(n4900), .ZN(n4899) );
  NAND2_X2 U5225 ( .A1(n10355), .A2(n6056), .ZN(n9743) );
  NAND2_X2 U5226 ( .A1(n7645), .A2(n9746), .ZN(n10355) );
  NAND2_X2 U5227 ( .A1(n9296), .A2(n9299), .ZN(n6275) );
  INV_X1 U5228 ( .A(n6889), .ZN(n5449) );
  OAI222_X1 U5229 ( .A1(P2_U3151), .A2(n7317), .B1(n9307), .B2(n6911), .C1(
        n6910), .C2(n8134), .ZN(P2_U3294) );
  OAI222_X1 U5230 ( .A1(n10311), .A2(n6972), .B1(n10335), .B2(n6911), .C1(
        n6895), .C2(n10332), .ZN(P1_U3354) );
  XNOR2_X1 U5231 ( .A(n5451), .B(n5452), .ZN(n6911) );
  NAND2_X1 U5232 ( .A1(n6084), .A2(n6924), .ZN(n4432) );
  NAND2_X1 U5233 ( .A1(n6084), .A2(n6924), .ZN(n4433) );
  NAND2_X2 U5234 ( .A1(n6084), .A2(n6924), .ZN(n5582) );
  NAND2_X2 U5235 ( .A1(n10122), .A2(n6065), .ZN(n10125) );
  NAND2_X2 U5236 ( .A1(n4787), .A2(n7816), .ZN(n7818) );
  OAI222_X1 U5237 ( .A1(n10332), .A2(n10325), .B1(P1_U3086), .B2(n6924), .C1(
        n10335), .C2(n10324), .ZN(P1_U3328) );
  INV_X2 U5238 ( .A(n10414), .ZN(n5458) );
  XNOR2_X2 U5239 ( .A(n5617), .B(n5616), .ZN(n6912) );
  OR2_X1 U5240 ( .A1(n6428), .A2(n10496), .ZN(n6263) );
  BUF_X4 U5241 ( .A(n5552), .Z(n4437) );
  AND2_X2 U5242 ( .A1(n10322), .A2(n10318), .ZN(n5552) );
  INV_X1 U5243 ( .A(n5603), .ZN(n5605) );
  OR2_X1 U5244 ( .A1(n8287), .A2(n9066), .ZN(n6711) );
  OR2_X1 U5245 ( .A1(n6879), .A2(n6770), .ZN(n6789) );
  NOR2_X1 U5246 ( .A1(n9720), .A2(n6075), .ZN(n9996) );
  AND2_X1 U5247 ( .A1(n5013), .A2(n5014), .ZN(n5012) );
  NOR2_X1 U5248 ( .A1(n10025), .A2(n5015), .ZN(n5014) );
  NOR2_X1 U5249 ( .A1(n6774), .A2(n6758), .ZN(n6793) );
  INV_X1 U5250 ( .A(n6566), .ZN(n4579) );
  NAND2_X1 U5251 ( .A1(n6569), .A2(n7968), .ZN(n4578) );
  AND2_X1 U5252 ( .A1(n6177), .A2(n6176), .ZN(n6838) );
  INV_X1 U5253 ( .A(n4768), .ZN(n6534) );
  NAND2_X1 U5254 ( .A1(n5006), .A2(n5005), .ZN(n5004) );
  NAND2_X1 U5255 ( .A1(n7569), .A2(n7570), .ZN(n5005) );
  OAI22_X1 U5256 ( .A1(n8445), .A2(n8444), .B1(n8443), .B2(n8442), .ZN(n8465)
         );
  OAI21_X1 U5257 ( .B1(n8441), .B2(n5089), .A(n4564), .ZN(n5085) );
  NAND2_X1 U5258 ( .A1(n5090), .A2(n4563), .ZN(n5089) );
  NAND2_X1 U5259 ( .A1(n8127), .A2(n6533), .ZN(n8819) );
  XNOR2_X1 U5260 ( .A(n9192), .B(n8834), .ZN(n8823) );
  AND2_X1 U5261 ( .A1(n4428), .A2(n6853), .ZN(n9064) );
  INV_X1 U5262 ( .A(n9008), .ZN(n9065) );
  NAND2_X1 U5263 ( .A1(n4635), .A2(n4633), .ZN(n4632) );
  INV_X1 U5264 ( .A(n9730), .ZN(n10168) );
  NOR2_X1 U5265 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5812) );
  NOR2_X1 U5266 ( .A1(n9598), .A2(n5106), .ZN(n5105) );
  INV_X1 U5267 ( .A(n9596), .ZN(n5106) );
  AOI21_X1 U5268 ( .B1(n5179), .B2(n5177), .A(n6886), .ZN(n5021) );
  NAND2_X1 U5269 ( .A1(n6639), .A2(n6638), .ZN(n5033) );
  NAND2_X1 U5270 ( .A1(n6636), .A2(n6638), .ZN(n4581) );
  AOI21_X1 U5271 ( .B1(n6482), .B2(n4584), .A(n4583), .ZN(n4582) );
  NOR2_X1 U5272 ( .A1(n5761), .A2(n5373), .ZN(n5372) );
  NOR2_X1 U5273 ( .A1(n5760), .A2(SI_16_), .ZN(n5761) );
  INV_X1 U5274 ( .A(n5743), .ZN(n5373) );
  AOI211_X1 U5275 ( .C1(n8854), .C2(n6579), .A(n6508), .B(n6507), .ZN(n6509)
         );
  NAND2_X1 U5276 ( .A1(n8450), .A2(n8449), .ZN(n8451) );
  NOR2_X1 U5277 ( .A1(n5252), .A2(n5945), .ZN(n5251) );
  INV_X1 U5278 ( .A(n5921), .ZN(n5252) );
  NOR2_X1 U5279 ( .A1(n5368), .A2(n5724), .ZN(n5366) );
  INV_X1 U5280 ( .A(n5372), .ZN(n5368) );
  AND2_X1 U5281 ( .A1(n4977), .A2(n5707), .ZN(n4861) );
  INV_X1 U5282 ( .A(n7448), .ZN(n5324) );
  NAND2_X1 U5283 ( .A1(n7234), .A2(n4483), .ZN(n4756) );
  NAND2_X1 U5284 ( .A1(n7272), .A2(n4755), .ZN(n4754) );
  INV_X1 U5285 ( .A(n7274), .ZN(n4755) );
  NAND2_X1 U5286 ( .A1(n7621), .A2(n4494), .ZN(n4764) );
  NAND2_X1 U5287 ( .A1(n7560), .A2(n4767), .ZN(n4765) );
  AND2_X1 U5288 ( .A1(n5303), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5302) );
  NAND2_X1 U5289 ( .A1(n8389), .A2(n8390), .ZN(n4763) );
  INV_X1 U5290 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5291 ( .B1(n6822), .B2(n4723), .A(n6824), .ZN(n4722) );
  OR2_X1 U5292 ( .A1(n9204), .A2(n8314), .ZN(n6648) );
  AOI21_X1 U5293 ( .B1(n4735), .B2(n4738), .A(n4734), .ZN(n4733) );
  NAND2_X1 U5294 ( .A1(n6627), .A2(n4735), .ZN(n4732) );
  INV_X1 U5295 ( .A(n6630), .ZN(n4734) );
  OAI21_X1 U5296 ( .B1(n6620), .B2(n6226), .A(n6622), .ZN(n5275) );
  INV_X1 U5297 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4931) );
  NAND2_X1 U5298 ( .A1(n5974), .A2(n5973), .ZN(n5255) );
  OR2_X1 U5299 ( .A1(n10197), .A2(n6071), .ZN(n9699) );
  OR2_X1 U5300 ( .A1(n10206), .A2(n6070), .ZN(n9769) );
  NAND2_X1 U5301 ( .A1(n10160), .A2(n6061), .ZN(n5221) );
  AND2_X1 U5302 ( .A1(n7066), .A2(n7063), .ZN(n7059) );
  INV_X1 U5303 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U5304 ( .A1(n5948), .A2(n5946), .ZN(n5924) );
  NAND2_X1 U5305 ( .A1(n4967), .A2(n4966), .ZN(n5864) );
  NAND2_X1 U5306 ( .A1(n5826), .A2(n5807), .ZN(n5827) );
  OAI21_X1 U5307 ( .B1(n5786), .B2(n5785), .A(n5784), .ZN(n5804) );
  NAND2_X1 U5308 ( .A1(n5711), .A2(n5710), .ZN(n5726) );
  NAND2_X1 U5310 ( .A1(n4896), .A2(n8277), .ZN(n8186) );
  AND2_X1 U5311 ( .A1(n6717), .A2(n4917), .ZN(n4916) );
  OR2_X1 U5312 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  NAND2_X1 U5313 ( .A1(n6712), .A2(n4918), .ZN(n4917) );
  AND2_X1 U5314 ( .A1(n4856), .A2(n6654), .ZN(n5068) );
  NOR2_X1 U5315 ( .A1(n6655), .A2(n4858), .ZN(n4857) );
  NAND2_X1 U5316 ( .A1(n5297), .A2(n5298), .ZN(n5300) );
  AOI21_X1 U5317 ( .B1(n7268), .B2(n4684), .A(n4683), .ZN(n7552) );
  AND2_X1 U5318 ( .A1(n7269), .A2(n7270), .ZN(n4683) );
  OR2_X1 U5319 ( .A1(n7269), .A2(n7270), .ZN(n4684) );
  INV_X1 U5320 ( .A(n7625), .ZN(n5003) );
  OR2_X1 U5321 ( .A1(n8448), .A2(n9148), .ZN(n5103) );
  NAND2_X1 U5322 ( .A1(n4985), .A2(n4983), .ZN(n8773) );
  AND2_X1 U5323 ( .A1(n4987), .A2(n4984), .ZN(n4983) );
  NAND2_X1 U5324 ( .A1(n4580), .A2(n6155), .ZN(n6197) );
  INV_X1 U5325 ( .A(n5163), .ZN(n5162) );
  OAI21_X1 U5326 ( .B1(n6829), .B2(n5164), .A(n6828), .ZN(n5163) );
  OR2_X1 U5327 ( .A1(n8948), .A2(n8954), .ZN(n8927) );
  OAI211_X1 U5328 ( .C1(n6819), .C2(n4544), .A(n4706), .B(n6820), .ZN(n9004)
         );
  INV_X1 U5329 ( .A(n4544), .ZN(n4707) );
  NAND2_X1 U5330 ( .A1(n6606), .A2(n6605), .ZN(n7429) );
  NAND2_X1 U5331 ( .A1(n4921), .A2(n6944), .ZN(n4920) );
  NAND2_X1 U5332 ( .A1(n7869), .A2(n4922), .ZN(n4921) );
  NAND2_X1 U5333 ( .A1(n4715), .A2(n4714), .ZN(n8825) );
  AOI21_X1 U5334 ( .B1(n4716), .B2(n4550), .A(n4451), .ZN(n4714) );
  NAND2_X1 U5335 ( .A1(n6834), .A2(n4716), .ZN(n4715) );
  XNOR2_X1 U5336 ( .A(n6838), .B(n9198), .ZN(n6507) );
  NAND2_X1 U5337 ( .A1(n4532), .A2(n5149), .ZN(n5146) );
  AND2_X1 U5338 ( .A1(n6645), .A2(n6579), .ZN(n8856) );
  AOI21_X1 U5339 ( .B1(n4743), .B2(n6481), .A(n4741), .ZN(n4740) );
  NAND2_X1 U5340 ( .A1(n8914), .A2(n4743), .ZN(n4739) );
  INV_X1 U5341 ( .A(n6638), .ZN(n4741) );
  NAND2_X1 U5342 ( .A1(n7429), .A2(n6607), .ZN(n5285) );
  AND2_X1 U5343 ( .A1(n6674), .A2(n6885), .ZN(n6787) );
  OR2_X1 U5344 ( .A1(n6887), .A2(n6680), .ZN(n6674) );
  NAND2_X1 U5345 ( .A1(n4746), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6141) );
  NOR2_X1 U5346 ( .A1(n4464), .A2(n5409), .ZN(n5041) );
  INV_X1 U5347 ( .A(n7064), .ZN(n4614) );
  AND2_X1 U5348 ( .A1(n9796), .A2(n6076), .ZN(n9735) );
  AND4_X1 U5349 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n8062)
         );
  NOR2_X1 U5350 ( .A1(n9347), .A2(n5398), .ZN(n5397) );
  INV_X1 U5351 ( .A(n5399), .ZN(n5398) );
  AND2_X1 U5352 ( .A1(n10001), .A2(n10000), .ZN(n10173) );
  NOR2_X1 U5353 ( .A1(n5203), .A2(n9645), .ZN(n5202) );
  NOR2_X1 U5354 ( .A1(n9689), .A2(n9705), .ZN(n5203) );
  NOR2_X1 U5355 ( .A1(n4485), .A2(n5242), .ZN(n5241) );
  INV_X1 U5356 ( .A(n5797), .ZN(n5242) );
  NAND2_X1 U5357 ( .A1(n5212), .A2(n5211), .ZN(n10115) );
  AOI21_X1 U5358 ( .B1(n5214), .B2(n5216), .A(n4506), .ZN(n5211) );
  NAND2_X1 U5359 ( .A1(n7849), .A2(n5214), .ZN(n5212) );
  INV_X1 U5360 ( .A(n5217), .ZN(n5216) );
  OR2_X1 U5361 ( .A1(n10240), .A2(n9829), .ZN(n4944) );
  INV_X1 U5362 ( .A(n7059), .ZN(n10254) );
  AND2_X1 U5363 ( .A1(n6031), .A2(n6030), .ZN(n7056) );
  NAND2_X1 U5364 ( .A1(n5924), .A2(n4551), .ZN(n5906) );
  XNOR2_X1 U5365 ( .A(n6045), .B(n6044), .ZN(n7866) );
  NAND2_X1 U5366 ( .A1(n6014), .A2(n5365), .ZN(n5364) );
  NAND2_X1 U5367 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .ZN(n5365) );
  INV_X1 U5368 ( .A(n5363), .ZN(n5362) );
  OAI21_X1 U5369 ( .B1(n5364), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5363) );
  AOI21_X1 U5370 ( .B1(n5811), .B2(n5810), .A(n5809), .ZN(n5814) );
  NAND2_X1 U5371 ( .A1(n6782), .A2(n9087), .ZN(n8316) );
  NAND2_X1 U5372 ( .A1(n5061), .A2(n6539), .ZN(n8826) );
  NAND2_X1 U5373 ( .A1(n8819), .A2(n6534), .ZN(n5061) );
  INV_X1 U5374 ( .A(n6838), .ZN(n8841) );
  INV_X1 U5375 ( .A(n8314), .ZN(n8858) );
  NAND2_X1 U5376 ( .A1(n6252), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4680) );
  OR2_X1 U5377 ( .A1(P2_U3150), .A2(n4589), .ZN(n8778) );
  INV_X1 U5378 ( .A(n9087), .ZN(n10518) );
  INV_X1 U5379 ( .A(n5175), .ZN(n5172) );
  AOI21_X1 U5380 ( .B1(n8817), .B2(n9065), .A(n5176), .ZN(n5175) );
  NAND2_X1 U5381 ( .A1(n6521), .A2(n6520), .ZN(n9192) );
  OR2_X1 U5382 ( .A1(n4432), .A2(n6972), .ZN(n5456) );
  NAND2_X1 U5383 ( .A1(n5972), .A2(n5971), .ZN(n9816) );
  INV_X1 U5384 ( .A(n10164), .ZN(n10393) );
  INV_X1 U5385 ( .A(n9579), .ZN(n5110) );
  NAND2_X1 U5386 ( .A1(n9582), .A2(n9791), .ZN(n4814) );
  NAND2_X1 U5387 ( .A1(n4816), .A2(n9792), .ZN(n4815) );
  INV_X1 U5388 ( .A(n9581), .ZN(n4816) );
  AOI211_X1 U5389 ( .C1(n10374), .C2(n9568), .A(n9574), .B(n9566), .ZN(n9580)
         );
  AND2_X1 U5390 ( .A1(n6582), .A2(n4599), .ZN(n4701) );
  NAND2_X1 U5391 ( .A1(n4644), .A2(n4424), .ZN(n9615) );
  NOR2_X1 U5392 ( .A1(n4646), .A2(n9792), .ZN(n4645) );
  OAI21_X1 U5393 ( .B1(n6269), .B2(n6268), .A(n4500), .ZN(n6273) );
  AOI21_X1 U5394 ( .B1(n9620), .B2(n5112), .A(n10123), .ZN(n4660) );
  AOI21_X1 U5395 ( .B1(n9617), .B2(n5114), .A(n5113), .ZN(n5112) );
  AND2_X1 U5396 ( .A1(n9768), .A2(n10099), .ZN(n5111) );
  NOR2_X1 U5397 ( .A1(n5033), .A2(n4523), .ZN(n5030) );
  OAI21_X1 U5398 ( .B1(n5033), .B2(n4520), .A(n8850), .ZN(n5028) );
  NAND2_X1 U5399 ( .A1(n4446), .A2(n5032), .ZN(n5031) );
  NAND2_X1 U5400 ( .A1(n9590), .A2(n9589), .ZN(n9599) );
  AOI21_X1 U5401 ( .B1(n5155), .B2(n5153), .A(n6496), .ZN(n6511) );
  NOR2_X1 U5402 ( .A1(n5157), .A2(n5156), .ZN(n5155) );
  NAND2_X1 U5403 ( .A1(n4826), .A2(n4823), .ZN(n4822) );
  INV_X1 U5404 ( .A(n8892), .ZN(n4826) );
  NOR2_X1 U5405 ( .A1(n8915), .A2(n4824), .ZN(n4823) );
  AND2_X1 U5406 ( .A1(n6591), .A2(n4818), .ZN(n6594) );
  AND2_X1 U5407 ( .A1(n6592), .A2(n4819), .ZN(n4818) );
  NAND2_X1 U5408 ( .A1(n9702), .A2(n9563), .ZN(n5121) );
  NOR2_X1 U5409 ( .A1(n5827), .A2(n5358), .ZN(n5357) );
  INV_X1 U5410 ( .A(n5802), .ZN(n5358) );
  NOR2_X1 U5411 ( .A1(n6747), .A2(n5319), .ZN(n5318) );
  INV_X1 U5412 ( .A(n8277), .ZN(n5319) );
  AND2_X1 U5413 ( .A1(n8469), .A2(n4456), .ZN(n4752) );
  INV_X1 U5414 ( .A(n9625), .ZN(n5192) );
  NAND2_X1 U5415 ( .A1(n9746), .A2(n7643), .ZN(n9574) );
  NAND2_X1 U5416 ( .A1(n7077), .A2(n10414), .ZN(n9745) );
  NAND2_X1 U5417 ( .A1(n5805), .A2(n8513), .ZN(n5826) );
  INV_X1 U5418 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5655) );
  INV_X1 U5419 ( .A(n5549), .ZN(n5350) );
  AND2_X1 U5420 ( .A1(n9177), .A2(n8808), .ZN(n6575) );
  NAND2_X1 U5421 ( .A1(n4828), .A2(n4827), .ZN(n6657) );
  AND2_X1 U5422 ( .A1(n6598), .A2(n4829), .ZN(n4828) );
  INV_X1 U5423 ( .A(n6655), .ZN(n4827) );
  OR2_X1 U5424 ( .A1(n8451), .A2(n5101), .ZN(n4863) );
  NOR2_X1 U5425 ( .A1(n5087), .A2(n8480), .ZN(n5086) );
  INV_X1 U5426 ( .A(n5091), .ZN(n5087) );
  NOR2_X1 U5427 ( .A1(n8479), .A2(n9141), .ZN(n5093) );
  NAND2_X1 U5428 ( .A1(n8483), .A2(n8767), .ZN(n8485) );
  INV_X1 U5429 ( .A(n8826), .ZN(n7968) );
  NOR2_X1 U5430 ( .A1(n6465), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6464) );
  AND2_X1 U5431 ( .A1(n6153), .A2(n5071), .ZN(n5070) );
  INV_X1 U5432 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5071) );
  AND2_X1 U5433 ( .A1(n6152), .A2(n8738), .ZN(n6425) );
  AND2_X1 U5434 ( .A1(n6150), .A2(n5074), .ZN(n5073) );
  INV_X1 U5435 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5074) );
  INV_X1 U5436 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6150) );
  INV_X1 U5437 ( .A(n6385), .ZN(n6151) );
  NAND2_X1 U5438 ( .A1(n6287), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n4844) );
  OAI21_X1 U5439 ( .B1(n4597), .B2(n4515), .A(n4746), .ZN(n6677) );
  AOI21_X1 U5440 ( .B1(n5287), .B2(P2_IR_REG_31__SCAN_IN), .A(n4598), .ZN(
        n4597) );
  AND2_X1 U5441 ( .A1(n5144), .A2(n4541), .ZN(n4716) );
  NAND2_X1 U5442 ( .A1(n9210), .A2(n8871), .ZN(n5149) );
  OR2_X1 U5443 ( .A1(n8282), .A2(n8213), .ZN(n8852) );
  OR2_X1 U5444 ( .A1(n9226), .A2(n8882), .ZN(n8850) );
  OR2_X1 U5445 ( .A1(n9232), .A2(n8204), .ZN(n6637) );
  OR2_X1 U5446 ( .A1(n9253), .A2(n8327), .ZN(n6631) );
  NAND2_X1 U5447 ( .A1(n5404), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U5448 ( .A1(n6665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4898) );
  INV_X1 U5449 ( .A(n7292), .ZN(n5333) );
  AND2_X1 U5450 ( .A1(n8120), .A2(n5057), .ZN(n5056) );
  NAND2_X1 U5451 ( .A1(n5058), .A2(n4458), .ZN(n5057) );
  INV_X1 U5452 ( .A(n4458), .ZN(n5053) );
  INV_X1 U5453 ( .A(n9836), .ZN(n7463) );
  NOR2_X1 U5454 ( .A1(n9562), .A2(n5392), .ZN(n5391) );
  NAND2_X1 U5455 ( .A1(n10059), .A2(n5393), .ZN(n5392) );
  INV_X1 U5456 ( .A(n4876), .ZN(n5777) );
  INV_X1 U5457 ( .A(n5019), .ZN(n5195) );
  NAND2_X1 U5458 ( .A1(n6934), .A2(n5637), .ZN(n4934) );
  NAND2_X1 U5459 ( .A1(n4934), .A2(n4932), .ZN(n9597) );
  NOR2_X1 U5460 ( .A1(n8037), .A2(n4933), .ZN(n4932) );
  INV_X1 U5461 ( .A(n5642), .ZN(n4933) );
  NOR2_X1 U5462 ( .A1(n10245), .A2(n7528), .ZN(n5396) );
  NAND2_X1 U5463 ( .A1(n9835), .A2(n10445), .ZN(n7643) );
  NAND2_X1 U5464 ( .A1(n7201), .A2(n7203), .ZN(n6053) );
  NAND2_X1 U5465 ( .A1(n10426), .A2(n9838), .ZN(n9567) );
  INV_X1 U5466 ( .A(n5251), .ZN(n5248) );
  NOR2_X1 U5467 ( .A1(n5249), .A2(n5922), .ZN(n5246) );
  NOR2_X1 U5468 ( .A1(n9996), .A2(n5257), .ZN(n5256) );
  INV_X1 U5469 ( .A(n5973), .ZN(n5257) );
  INV_X1 U5470 ( .A(n4951), .ZN(n4950) );
  AND2_X1 U5471 ( .A1(n5251), .A2(n4952), .ZN(n4951) );
  NAND2_X1 U5472 ( .A1(n4953), .A2(n5905), .ZN(n4952) );
  INV_X1 U5473 ( .A(n9825), .ZN(n8083) );
  OAI21_X1 U5474 ( .B1(n6542), .B2(n8701), .A(n6123), .ZN(n6552) );
  XNOR2_X1 U5475 ( .A(n6122), .B(n6121), .ZN(n6542) );
  AND2_X1 U5476 ( .A1(n5400), .A2(n5444), .ZN(n5128) );
  AND2_X1 U5477 ( .A1(n5977), .A2(n5962), .ZN(n5975) );
  AND2_X1 U5478 ( .A1(n5956), .A2(n5934), .ZN(n5950) );
  INV_X1 U5479 ( .A(n5829), .ZN(n5353) );
  INV_X1 U5480 ( .A(n5799), .ZN(n5803) );
  XNOR2_X1 U5481 ( .A(n5800), .B(SI_18_), .ZN(n5799) );
  NOR2_X1 U5482 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5769) );
  NOR2_X1 U5483 ( .A1(n4491), .A2(n4628), .ZN(n4627) );
  INV_X1 U5484 ( .A(n5367), .ZN(n4628) );
  NAND2_X1 U5485 ( .A1(n5784), .A2(n5766), .ZN(n5785) );
  XNOR2_X1 U5486 ( .A(n5709), .B(SI_13_), .ZN(n5706) );
  INV_X1 U5487 ( .A(n4965), .ZN(n5338) );
  OAI21_X1 U5488 ( .B1(n5339), .B2(n4441), .A(n5673), .ZN(n4965) );
  NAND2_X1 U5489 ( .A1(n4517), .A2(n5654), .ZN(n5339) );
  NOR2_X1 U5490 ( .A1(n5651), .A2(n5340), .ZN(n4655) );
  XNOR2_X1 U5491 ( .A(n5652), .B(SI_10_), .ZN(n5651) );
  INV_X1 U5492 ( .A(n5590), .ZN(n5591) );
  NAND2_X1 U5493 ( .A1(n5615), .A2(n5599), .ZN(n5616) );
  INV_X1 U5494 ( .A(SI_6_), .ZN(n8588) );
  OAI21_X1 U5495 ( .B1(n6142), .B2(n4783), .A(n4782), .ZN(n5586) );
  NAND2_X1 U5496 ( .A1(n6142), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4782) );
  INV_X1 U5497 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5446) );
  AND2_X1 U5498 ( .A1(n5306), .A2(n4904), .ZN(n4903) );
  OR2_X1 U5499 ( .A1(n8298), .A2(n4461), .ZN(n4904) );
  AND2_X1 U5500 ( .A1(n8259), .A2(n5307), .ZN(n5306) );
  OR2_X1 U5501 ( .A1(n8202), .A2(n5308), .ZN(n5307) );
  INV_X1 U5502 ( .A(n6735), .ZN(n5308) );
  INV_X1 U5503 ( .A(n6712), .ZN(n4919) );
  AOI21_X1 U5504 ( .B1(n4927), .B2(n4929), .A(n4925), .ZN(n4924) );
  INV_X1 U5505 ( .A(n8244), .ZN(n4925) );
  INV_X1 U5506 ( .A(n5323), .ZN(n7446) );
  OR2_X1 U5507 ( .A1(n9177), .A2(n8808), .ZN(n6578) );
  AND2_X1 U5508 ( .A1(n5065), .A2(n5066), .ZN(n4859) );
  NOR2_X1 U5509 ( .A1(n4478), .A2(n5067), .ZN(n5066) );
  AND2_X1 U5510 ( .A1(n6562), .A2(n6549), .ZN(n7976) );
  INV_X1 U5511 ( .A(n6287), .ZN(n6489) );
  OAI21_X1 U5512 ( .B1(n7317), .B2(n7180), .A(n7181), .ZN(n7310) );
  NOR2_X1 U5513 ( .A1(n7310), .A2(n7962), .ZN(n7309) );
  XNOR2_X1 U5514 ( .A(n7158), .B(n4679), .ZN(n7306) );
  OAI21_X1 U5515 ( .B1(n8770), .B2(n7962), .A(n4999), .ZN(n7158) );
  NAND2_X1 U5516 ( .A1(n8770), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4999) );
  INV_X1 U5517 ( .A(n7183), .ZN(n7175) );
  XNOR2_X1 U5518 ( .A(n7183), .B(n4682), .ZN(n7215) );
  XNOR2_X1 U5519 ( .A(n7183), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7218) );
  INV_X1 U5520 ( .A(n4760), .ZN(n4759) );
  NAND3_X1 U5521 ( .A1(n4756), .A2(n4754), .A3(n4504), .ZN(n4758) );
  NOR2_X1 U5522 ( .A1(n7624), .A2(n5002), .ZN(n7751) );
  AND2_X1 U5523 ( .A1(n7572), .A2(n7573), .ZN(n5002) );
  NAND2_X1 U5524 ( .A1(n7557), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4685) );
  INV_X1 U5525 ( .A(n4884), .ZN(n4766) );
  NOR2_X1 U5526 ( .A1(n7754), .A2(n4884), .ZN(n7756) );
  AND2_X1 U5527 ( .A1(n5301), .A2(n5302), .ZN(n8350) );
  OR2_X1 U5528 ( .A1(n8371), .A2(n8370), .ZN(n4779) );
  AOI21_X1 U5529 ( .B1(n8359), .B2(n8358), .A(n4691), .ZN(n8379) );
  NOR2_X1 U5530 ( .A1(n8367), .A2(n9165), .ZN(n4691) );
  AOI22_X1 U5531 ( .A1(n8385), .A2(n8384), .B1(n8382), .B2(n8383), .ZN(n8403)
         );
  NAND2_X1 U5532 ( .A1(n4763), .A2(n4499), .ZN(n5291) );
  AND2_X1 U5533 ( .A1(n8424), .A2(n4885), .ZN(n4761) );
  OAI22_X1 U5534 ( .A1(n8403), .A2(n8402), .B1(n8401), .B2(n8400), .ZN(n8426)
         );
  NAND2_X1 U5535 ( .A1(n8409), .A2(n8420), .ZN(n8431) );
  NAND2_X1 U5536 ( .A1(n5289), .A2(n8431), .ZN(n8433) );
  INV_X1 U5537 ( .A(n5290), .ZN(n5289) );
  NAND2_X1 U5538 ( .A1(n5292), .A2(n5296), .ZN(n5293) );
  INV_X1 U5539 ( .A(n8761), .ZN(n5292) );
  NAND2_X1 U5540 ( .A1(n8485), .A2(n5295), .ZN(n5294) );
  AND2_X1 U5541 ( .A1(n5296), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5295) );
  OAI21_X1 U5542 ( .B1(n8755), .B2(n4665), .A(n4674), .ZN(n4669) );
  NAND2_X1 U5543 ( .A1(n8799), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5544 ( .A1(n8800), .A2(n4879), .ZN(n4665) );
  NAND2_X1 U5545 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  AND2_X1 U5546 ( .A1(n8800), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4671) );
  INV_X1 U5547 ( .A(n8757), .ZN(n4672) );
  INV_X1 U5548 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5075) );
  OR2_X1 U5549 ( .A1(n6487), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6499) );
  AND2_X1 U5550 ( .A1(n6580), .A2(n6635), .ZN(n8930) );
  AOI21_X1 U5551 ( .B1(n4721), .B2(n4723), .A(n4489), .ZN(n4718) );
  NAND2_X1 U5552 ( .A1(n8989), .A2(n4721), .ZN(n4719) );
  NAND2_X1 U5553 ( .A1(n4576), .A2(n6149), .ZN(n6354) );
  INV_X1 U5554 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6149) );
  INV_X1 U5555 ( .A(n6327), .ZN(n4576) );
  NAND2_X1 U5556 ( .A1(n6148), .A2(n6147), .ZN(n6337) );
  INV_X1 U5557 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6147) );
  INV_X1 U5558 ( .A(n6335), .ZN(n6148) );
  OR2_X1 U5559 ( .A1(n6298), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U5560 ( .A1(n7958), .A2(n7357), .ZN(n7364) );
  AND2_X1 U5561 ( .A1(n6541), .A2(n6540), .ZN(n7970) );
  INV_X1 U5562 ( .A(n6553), .ZN(n6306) );
  AOI21_X1 U5563 ( .B1(n5271), .B2(n5273), .A(n5268), .ZN(n5267) );
  INV_X1 U5564 ( .A(n6651), .ZN(n5268) );
  XNOR2_X1 U5565 ( .A(n9186), .B(n8826), .ZN(n8815) );
  INV_X1 U5566 ( .A(n8794), .ZN(n6772) );
  NAND2_X1 U5567 ( .A1(n8924), .A2(n5417), .ZN(n4700) );
  AOI21_X1 U5568 ( .B1(n4474), .B2(n5266), .A(n6480), .ZN(n5263) );
  AND3_X1 U5569 ( .A1(n6441), .A2(n6440), .A3(n6439), .ZN(n8954) );
  OR2_X1 U5570 ( .A1(n6886), .A2(n6853), .ZN(n9008) );
  NAND2_X1 U5571 ( .A1(n6621), .A2(n4750), .ZN(n4748) );
  INV_X1 U5572 ( .A(n5275), .ZN(n5274) );
  NAND2_X1 U5573 ( .A1(n5276), .A2(n6620), .ZN(n9003) );
  INV_X1 U5574 ( .A(n9001), .ZN(n5276) );
  INV_X1 U5575 ( .A(n9020), .ZN(n9022) );
  AND2_X1 U5576 ( .A1(n9039), .A2(n4538), .ZN(n4708) );
  NOR2_X1 U5577 ( .A1(n5284), .A2(n5286), .ZN(n5283) );
  INV_X1 U5578 ( .A(n6611), .ZN(n5284) );
  INV_X1 U5579 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6158) );
  XNOR2_X1 U5580 ( .A(n6208), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U5581 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4692) );
  NAND2_X1 U5582 ( .A1(n4470), .A2(n8579), .ZN(n6252) );
  NAND2_X1 U5583 ( .A1(n5529), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5574) );
  NOR2_X1 U5584 ( .A1(n5060), .A2(n5059), .ZN(n5058) );
  INV_X1 U5585 ( .A(n9475), .ZN(n5059) );
  INV_X1 U5586 ( .A(n9474), .ZN(n5060) );
  INV_X1 U5587 ( .A(n9837), .ZN(n7291) );
  NAND2_X1 U5588 ( .A1(n5043), .A2(n4498), .ZN(n5042) );
  INV_X1 U5589 ( .A(n8102), .ZN(n5043) );
  INV_X1 U5590 ( .A(n9357), .ZN(n5049) );
  AND2_X1 U5591 ( .A1(n8149), .A2(n8148), .ZN(n9425) );
  NAND2_X1 U5592 ( .A1(n5051), .A2(n5056), .ZN(n8136) );
  NAND2_X1 U5593 ( .A1(n9477), .A2(n4458), .ZN(n5051) );
  INV_X1 U5594 ( .A(n9336), .ZN(n5039) );
  INV_X1 U5595 ( .A(n5042), .ZN(n4617) );
  OAI21_X1 U5596 ( .B1(n8028), .B2(n5047), .A(n4514), .ZN(n5046) );
  NAND2_X1 U5597 ( .A1(n4443), .A2(n8033), .ZN(n5045) );
  INV_X1 U5598 ( .A(n7125), .ZN(n4605) );
  AND2_X1 U5599 ( .A1(n10409), .A2(n7204), .ZN(n7608) );
  NOR2_X1 U5600 ( .A1(n6085), .A2(n7112), .ZN(n9551) );
  AND4_X1 U5601 ( .A1(n5722), .A2(n5721), .A3(n5720), .A4(n5719), .ZN(n8064)
         );
  AND4_X1 U5602 ( .A1(n5672), .A2(n5671), .A3(n5670), .A4(n5669), .ZN(n9601)
         );
  INV_X1 U5603 ( .A(n10166), .ZN(n9666) );
  NAND2_X1 U5604 ( .A1(n6078), .A2(n6002), .ZN(n9352) );
  NAND2_X1 U5605 ( .A1(n5985), .A2(n5984), .ZN(n10174) );
  INV_X1 U5606 ( .A(n4891), .ZN(n5938) );
  NAND2_X1 U5607 ( .A1(n10188), .A2(n9431), .ZN(n9702) );
  INV_X1 U5608 ( .A(n10058), .ZN(n5199) );
  NOR2_X1 U5609 ( .A1(n10086), .A2(n10197), .ZN(n10075) );
  NOR2_X1 U5610 ( .A1(n10101), .A2(n6068), .ZN(n6069) );
  OR2_X1 U5611 ( .A1(n10215), .A2(n9506), .ZN(n10099) );
  OR2_X1 U5612 ( .A1(n10230), .A2(n8064), .ZN(n10148) );
  NAND2_X1 U5613 ( .A1(n6060), .A2(n7818), .ZN(n5196) );
  AND2_X1 U5614 ( .A1(n10148), .A2(n9613), .ZN(n9685) );
  NAND2_X1 U5615 ( .A1(n10462), .A2(n7668), .ZN(n5237) );
  NAND2_X1 U5616 ( .A1(n5223), .A2(n5237), .ZN(n5230) );
  INV_X1 U5617 ( .A(n7787), .ZN(n5223) );
  NOR2_X1 U5618 ( .A1(n7782), .A2(n5109), .ZN(n5234) );
  OAI21_X1 U5619 ( .B1(n7782), .B2(n5239), .A(n5238), .ZN(n5233) );
  OR2_X1 U5620 ( .A1(n5587), .A2(n6893), .ZN(n5566) );
  NAND2_X1 U5621 ( .A1(n9998), .A2(n10377), .ZN(n5007) );
  AND2_X1 U5622 ( .A1(n9641), .A2(n9702), .ZN(n10047) );
  INV_X1 U5623 ( .A(n4939), .ZN(n4938) );
  OAI21_X1 U5624 ( .B1(n5241), .B2(n4440), .A(n5839), .ZN(n4939) );
  NAND2_X1 U5625 ( .A1(n10098), .A2(n5796), .ZN(n5798) );
  INV_X1 U5626 ( .A(n5215), .ZN(n5214) );
  OAI21_X1 U5627 ( .B1(n5218), .B2(n5216), .A(n10135), .ZN(n5215) );
  AND2_X1 U5628 ( .A1(n5221), .A2(n5723), .ZN(n5218) );
  NAND2_X1 U5629 ( .A1(n4531), .A2(n5221), .ZN(n5217) );
  NAND2_X1 U5630 ( .A1(n9473), .A2(n8062), .ZN(n4942) );
  NAND2_X1 U5631 ( .A1(n7093), .A2(n5637), .ZN(n5680) );
  INV_X1 U5632 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5431) );
  XNOR2_X1 U5633 ( .A(n6552), .B(n6551), .ZN(n9295) );
  INV_X1 U5634 ( .A(n5443), .ZN(n5129) );
  XNOR2_X1 U5635 ( .A(n5976), .B(n5975), .ZN(n7868) );
  NAND2_X1 U5636 ( .A1(n5038), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6020) );
  NOR2_X1 U5637 ( .A1(n5428), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5037) );
  XNOR2_X1 U5638 ( .A(n5935), .B(n5950), .ZN(n8133) );
  NAND2_X1 U5639 ( .A1(n5930), .A2(n5953), .ZN(n5935) );
  NAND2_X1 U5640 ( .A1(n5924), .A2(n5949), .ZN(n5930) );
  XNOR2_X1 U5641 ( .A(n5911), .B(n5910), .ZN(n9308) );
  NAND2_X1 U5642 ( .A1(n5906), .A2(n5925), .ZN(n5911) );
  NAND2_X1 U5643 ( .A1(n5887), .A2(n5886), .ZN(n5948) );
  INV_X1 U5644 ( .A(n5885), .ZN(n5886) );
  AOI21_X1 U5645 ( .B1(n6016), .B2(n5362), .A(n5360), .ZN(n5359) );
  NAND2_X1 U5646 ( .A1(n5361), .A2(n6012), .ZN(n5360) );
  NAND2_X1 U5647 ( .A1(n5362), .A2(n5364), .ZN(n5361) );
  INV_X1 U5648 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6014) );
  XNOR2_X1 U5649 ( .A(n5844), .B(n5843), .ZN(n7832) );
  OAI211_X1 U5650 ( .C1(n5354), .C2(n5353), .A(n5352), .B(n5351), .ZN(n7813)
         );
  NAND2_X1 U5651 ( .A1(n4970), .A2(n5829), .ZN(n5351) );
  NAND2_X1 U5652 ( .A1(n5354), .A2(n4480), .ZN(n5352) );
  NAND2_X1 U5653 ( .A1(n4968), .A2(n4972), .ZN(n5354) );
  NAND2_X1 U5654 ( .A1(n5374), .A2(n5743), .ZN(n5762) );
  NAND2_X1 U5655 ( .A1(n5371), .A2(n5369), .ZN(n5374) );
  AND2_X1 U5656 ( .A1(n5641), .A2(n5660), .ZN(n7005) );
  NAND2_X1 U5657 ( .A1(n5517), .A2(n5184), .ZN(n5603) );
  AND2_X1 U5658 ( .A1(n5600), .A2(n5562), .ZN(n5184) );
  NAND2_X1 U5659 ( .A1(n5605), .A2(n5604), .ZN(n5772) );
  AND2_X1 U5660 ( .A1(n4534), .A2(n6751), .ZN(n5320) );
  AND2_X1 U5661 ( .A1(n6202), .A2(n6201), .ZN(n8232) );
  OAI211_X2 U5662 ( .C1(n7377), .C2(n6700), .A(n6699), .B(n7505), .ZN(n7509)
         );
  AND2_X1 U5663 ( .A1(n8225), .A2(n8881), .ZN(n4908) );
  NAND2_X1 U5664 ( .A1(n4912), .A2(n8225), .ZN(n4906) );
  NAND2_X1 U5665 ( .A1(n8253), .A2(n8252), .ZN(n4912) );
  AND4_X1 U5666 ( .A1(n6360), .A2(n6359), .A3(n6358), .A4(n6357), .ZN(n7685)
         );
  AND3_X1 U5667 ( .A1(n6785), .A2(n6853), .A3(n6793), .ZN(n8324) );
  INV_X1 U5668 ( .A(n8326), .ZN(n8310) );
  INV_X1 U5669 ( .A(n9223), .ZN(n8282) );
  INV_X1 U5670 ( .A(n8316), .ZN(n8332) );
  NAND2_X1 U5671 ( .A1(n6796), .A2(n6795), .ZN(n8329) );
  AND2_X1 U5672 ( .A1(n6578), .A2(n7360), .ZN(n5137) );
  INV_X1 U5673 ( .A(n8213), .ZN(n8896) );
  NOR2_X1 U5674 ( .A1(n10507), .A2(n5001), .ZN(n7166) );
  AND2_X1 U5675 ( .A1(n7164), .A2(n10506), .ZN(n5001) );
  XNOR2_X1 U5676 ( .A(n6280), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7242) );
  NAND2_X1 U5677 ( .A1(n4470), .A2(n5277), .ZN(n6279) );
  OR2_X1 U5678 ( .A1(n7266), .A2(n7267), .ZN(n5006) );
  MUX2_X1 U5679 ( .A(n7169), .B(n8774), .S(n7168), .Z(n8795) );
  OR2_X1 U5680 ( .A1(n8441), .A2(n8440), .ZN(n5104) );
  NAND2_X1 U5681 ( .A1(n5096), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5095) );
  INV_X1 U5682 ( .A(n5099), .ZN(n5096) );
  AND2_X1 U5683 ( .A1(n4690), .A2(n5102), .ZN(n4689) );
  NAND2_X1 U5684 ( .A1(n5088), .A2(n5091), .ZN(n5102) );
  OAI21_X1 U5685 ( .B1(n8472), .B2(n8471), .A(n8470), .ZN(n8482) );
  AND2_X1 U5686 ( .A1(n8797), .A2(n8799), .ZN(n4994) );
  XNOR2_X1 U5687 ( .A(n8801), .B(n8800), .ZN(n4997) );
  OAI21_X1 U5688 ( .B1(n8757), .B2(n8756), .A(n4675), .ZN(n8801) );
  NAND2_X1 U5689 ( .A1(n8754), .A2(n4879), .ZN(n4675) );
  OAI21_X1 U5690 ( .B1(n8778), .B2(n8777), .A(n8776), .ZN(n4996) );
  AND2_X1 U5691 ( .A1(P2_U3893), .A2(n6676), .ZN(n8797) );
  NAND2_X1 U5692 ( .A1(n6781), .A2(n6929), .ZN(n9087) );
  INV_X1 U5693 ( .A(n9090), .ZN(n9029) );
  INV_X1 U5694 ( .A(n7970), .ZN(n9186) );
  XNOR2_X1 U5695 ( .A(n8816), .B(n8815), .ZN(n5173) );
  AND2_X1 U5696 ( .A1(n5169), .A2(n5174), .ZN(n5168) );
  NAND2_X1 U5697 ( .A1(n6883), .A2(n9103), .ZN(n5174) );
  OR2_X1 U5698 ( .A1(n5172), .A2(n5170), .ZN(n5169) );
  NOR2_X1 U5699 ( .A1(n4557), .A2(n4806), .ZN(n4805) );
  NOR2_X1 U5700 ( .A1(n10557), .A2(n9106), .ZN(n4806) );
  NAND2_X1 U5701 ( .A1(n10557), .A2(n10543), .ZN(n9172) );
  INV_X1 U5702 ( .A(n9172), .ZN(n9159) );
  NAND2_X1 U5703 ( .A1(n5270), .A2(n6650), .ZN(n8822) );
  NAND2_X1 U5704 ( .A1(n8831), .A2(n8832), .ZN(n5270) );
  NAND2_X1 U5705 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  NAND2_X1 U5706 ( .A1(n8841), .A2(n9064), .ZN(n4801) );
  INV_X1 U5707 ( .A(n6744), .ZN(n9210) );
  NAND2_X1 U5708 ( .A1(n4883), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U5709 ( .A1(n8857), .A2(n9064), .ZN(n4882) );
  NAND2_X1 U5710 ( .A1(n6498), .A2(n6497), .ZN(n9216) );
  XNOR2_X1 U5711 ( .A(n6293), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7269) );
  NAND2_X1 U5712 ( .A1(n7765), .A2(n5637), .ZN(n4658) );
  AND2_X1 U5713 ( .A1(n9532), .A2(n8172), .ZN(n9350) );
  AND2_X1 U5714 ( .A1(n7070), .A2(n7069), .ZN(n4624) );
  NAND2_X1 U5715 ( .A1(n6919), .A2(n5260), .ZN(n5259) );
  INV_X1 U5716 ( .A(n9900), .ZN(n5260) );
  NAND2_X1 U5717 ( .A1(n9531), .A2(n8159), .ZN(n9532) );
  AND2_X1 U5718 ( .A1(n9534), .A2(n9530), .ZN(n8159) );
  NAND2_X1 U5719 ( .A1(n4631), .A2(n9669), .ZN(n9741) );
  OR2_X1 U5720 ( .A1(n9401), .A2(n5557), .ZN(n5944) );
  NAND2_X1 U5721 ( .A1(n9989), .A2(n9990), .ZN(n4889) );
  NOR2_X1 U5722 ( .A1(n9988), .A2(n9800), .ZN(n4888) );
  NAND2_X1 U5723 ( .A1(n4786), .A2(n4785), .ZN(n4886) );
  AOI21_X1 U5724 ( .B1(n9983), .B2(n9990), .A(n9991), .ZN(n4785) );
  NAND2_X1 U5725 ( .A1(n9986), .A2(n9984), .ZN(n4786) );
  NAND2_X1 U5726 ( .A1(n7999), .A2(n7998), .ZN(n10171) );
  AND2_X1 U5727 ( .A1(n7996), .A2(n10390), .ZN(n7999) );
  OR2_X1 U5728 ( .A1(n7995), .A2(n10168), .ZN(n7996) );
  NAND2_X1 U5729 ( .A1(n5007), .A2(n9999), .ZN(n10172) );
  OAI21_X1 U5730 ( .B1(n10011), .B2(n5974), .A(n5973), .ZN(n10006) );
  OAI21_X1 U5731 ( .B1(n4838), .B2(n7916), .A(n4837), .ZN(n7930) );
  INV_X1 U5732 ( .A(n9403), .ZN(n4837) );
  NAND2_X1 U5733 ( .A1(n4839), .A2(n10377), .ZN(n4838) );
  NAND2_X1 U5734 ( .A1(n7917), .A2(n9689), .ZN(n4839) );
  INV_X1 U5735 ( .A(n5713), .ZN(n5018) );
  INV_X1 U5736 ( .A(n10383), .ZN(n10079) );
  OR2_X1 U5737 ( .A1(n7610), .A2(n7636), .ZN(n10164) );
  OR2_X1 U5738 ( .A1(n7610), .A2(n7611), .ZN(n10383) );
  NAND2_X1 U5739 ( .A1(n10165), .A2(n4790), .ZN(n10255) );
  INV_X1 U5740 ( .A(n4791), .ZN(n4790) );
  OAI21_X1 U5741 ( .B1(n10166), .B2(n10473), .A(n10167), .ZN(n4791) );
  INV_X1 U5742 ( .A(n7914), .ZN(n4851) );
  INV_X1 U5743 ( .A(n5244), .ZN(n6010) );
  NAND2_X1 U5744 ( .A1(n5258), .A2(n5921), .ZN(n7915) );
  NAND2_X1 U5745 ( .A1(n4955), .A2(n4953), .ZN(n5258) );
  AND2_X1 U5746 ( .A1(n10409), .A2(n6916), .ZN(n10405) );
  NAND2_X1 U5747 ( .A1(n5443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5445) );
  NOR2_X2 U5748 ( .A1(n9593), .A2(n9599), .ZN(n4643) );
  NAND2_X1 U5749 ( .A1(n5107), .A2(n9588), .ZN(n4649) );
  NAND2_X1 U5750 ( .A1(n6259), .A2(n6600), .ZN(n4600) );
  NOR2_X1 U5751 ( .A1(n6258), .A2(n6804), .ZN(n4809) );
  INV_X1 U5752 ( .A(n9755), .ZN(n4646) );
  NAND2_X1 U5753 ( .A1(n6270), .A2(n6600), .ZN(n6271) );
  NAND2_X1 U5754 ( .A1(n9619), .A2(n9791), .ZN(n5113) );
  INV_X1 U5755 ( .A(n9621), .ZN(n5114) );
  AND2_X1 U5756 ( .A1(n9613), .A2(n9756), .ZN(n4781) );
  NAND2_X1 U5757 ( .A1(n5181), .A2(n5180), .ZN(n5179) );
  AND2_X1 U5758 ( .A1(n6592), .A2(n6615), .ZN(n5180) );
  NAND2_X1 U5759 ( .A1(n6369), .A2(n4596), .ZN(n5181) );
  INV_X1 U5760 ( .A(n6376), .ZN(n5178) );
  NOR2_X1 U5761 ( .A1(n5188), .A2(n4778), .ZN(n4777) );
  NAND2_X1 U5762 ( .A1(n9625), .A2(n9792), .ZN(n4778) );
  NAND2_X1 U5763 ( .A1(n5121), .A2(n9791), .ZN(n5120) );
  INV_X1 U5764 ( .A(n6634), .ZN(n5032) );
  INV_X1 U5765 ( .A(n4964), .ZN(n4962) );
  NAND2_X1 U5766 ( .A1(n8916), .A2(n6580), .ZN(n4583) );
  NOR2_X1 U5767 ( .A1(n6480), .A2(n5266), .ZN(n4584) );
  NOR2_X1 U5768 ( .A1(n5154), .A2(n6886), .ZN(n4874) );
  NOR2_X1 U5769 ( .A1(n6484), .A2(n4428), .ZN(n5157) );
  NAND2_X1 U5770 ( .A1(n5029), .A2(n5027), .ZN(n6484) );
  INV_X1 U5771 ( .A(n5028), .ZN(n5027) );
  INV_X1 U5772 ( .A(n8905), .ZN(n4825) );
  NOR2_X1 U5773 ( .A1(n6593), .A2(n4820), .ZN(n4819) );
  NAND2_X1 U5774 ( .A1(n4539), .A2(n9042), .ZN(n4820) );
  AND2_X1 U5775 ( .A1(n4651), .A2(n4650), .ZN(n9753) );
  NAND2_X1 U5776 ( .A1(n9751), .A2(n4652), .ZN(n4651) );
  INV_X1 U5777 ( .A(n9597), .ZN(n4652) );
  OR2_X1 U5778 ( .A1(n9661), .A2(n9792), .ZN(n9662) );
  AND2_X1 U5779 ( .A1(n6596), .A2(n4821), .ZN(n6597) );
  NOR2_X1 U5780 ( .A1(n4822), .A2(n8869), .ZN(n4821) );
  NOR2_X1 U5781 ( .A1(n6653), .A2(n4830), .ZN(n4829) );
  OR2_X1 U5782 ( .A1(n6321), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6377) );
  OR2_X1 U5783 ( .A1(n8074), .A2(n8073), .ZN(n5407) );
  INV_X1 U5784 ( .A(n5121), .ZN(n9712) );
  AND2_X1 U5785 ( .A1(n10174), .A2(n9538), .ZN(n6075) );
  NOR2_X1 U5786 ( .A1(n10174), .A2(n9538), .ZN(n9720) );
  INV_X1 U5787 ( .A(n9702), .ZN(n5015) );
  INV_X1 U5788 ( .A(n5191), .ZN(n4653) );
  NOR2_X1 U5789 ( .A1(n5716), .A2(n5715), .ZN(n4892) );
  OR2_X1 U5790 ( .A1(n10225), .A2(n6061), .ZN(n9616) );
  NAND2_X1 U5791 ( .A1(n9473), .A2(n5390), .ZN(n5389) );
  NAND2_X1 U5792 ( .A1(n6119), .A2(n6118), .ZN(n6122) );
  AND2_X1 U5793 ( .A1(n5953), .A2(n5946), .ZN(n5947) );
  AND2_X1 U5794 ( .A1(n4969), .A2(n5853), .ZN(n4966) );
  AOI21_X1 U5795 ( .B1(n4972), .B2(n4971), .A(n4970), .ZN(n4969) );
  INV_X1 U5796 ( .A(n5784), .ZN(n4971) );
  NAND2_X1 U5797 ( .A1(n5785), .A2(n5784), .ZN(n4974) );
  INV_X1 U5798 ( .A(n5826), .ZN(n5356) );
  AOI21_X1 U5799 ( .B1(n5370), .B2(n5372), .A(n4452), .ZN(n5367) );
  INV_X1 U5800 ( .A(n5710), .ZN(n4630) );
  INV_X1 U5801 ( .A(SI_11_), .ZN(n5656) );
  INV_X1 U5802 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5618) );
  INV_X1 U5803 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5328) );
  INV_X1 U5804 ( .A(n6710), .ZN(n4918) );
  AOI21_X1 U5805 ( .B1(n5309), .B2(n4928), .A(n4555), .ZN(n4927) );
  INV_X1 U5806 ( .A(n8322), .ZN(n4928) );
  INV_X1 U5807 ( .A(n5309), .ZN(n4929) );
  AND2_X1 U5808 ( .A1(n6746), .A2(n5315), .ZN(n5314) );
  NAND2_X1 U5809 ( .A1(n5318), .A2(n5316), .ZN(n5315) );
  INV_X1 U5810 ( .A(n8276), .ZN(n5316) );
  INV_X1 U5811 ( .A(n5318), .ZN(n5317) );
  NOR2_X1 U5812 ( .A1(n9177), .A2(n9183), .ZN(n4858) );
  INV_X1 U5813 ( .A(n6578), .ZN(n5136) );
  NOR2_X1 U5814 ( .A1(n6660), .A2(n8794), .ZN(n5067) );
  NOR2_X1 U5815 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  NOR2_X1 U5816 ( .A1(n7574), .A2(n9075), .ZN(n4884) );
  OR2_X1 U5817 ( .A1(n8367), .A2(n8366), .ZN(n8368) );
  NAND2_X1 U5818 ( .A1(n8391), .A2(n8390), .ZN(n4762) );
  INV_X1 U5819 ( .A(n8440), .ZN(n5090) );
  NAND2_X1 U5820 ( .A1(n4752), .A2(n4863), .ZN(n4753) );
  NOR2_X1 U5821 ( .A1(n4990), .A2(n4993), .ZN(n4986) );
  INV_X1 U5822 ( .A(n4988), .ZN(n4987) );
  OAI21_X1 U5823 ( .B1(n8768), .B2(n4990), .A(n4989), .ZN(n4988) );
  INV_X1 U5824 ( .A(n8771), .ZN(n4989) );
  INV_X1 U5825 ( .A(n8768), .ZN(n4982) );
  NAND2_X1 U5826 ( .A1(n4993), .A2(n8768), .ZN(n4980) );
  OR2_X1 U5827 ( .A1(n6532), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8127) );
  AND2_X1 U5828 ( .A1(n6156), .A2(n5077), .ZN(n5076) );
  INV_X1 U5829 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5077) );
  INV_X1 U5830 ( .A(n6197), .ZN(n6157) );
  NOR2_X1 U5831 ( .A1(n6499), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U5832 ( .A1(n5167), .A2(n6825), .ZN(n5164) );
  NOR2_X1 U5833 ( .A1(n6829), .A2(n5166), .ZN(n5165) );
  INV_X1 U5834 ( .A(n6825), .ZN(n5166) );
  INV_X1 U5835 ( .A(n6823), .ZN(n4723) );
  INV_X1 U5836 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8712) );
  NOR2_X1 U5837 ( .A1(n6354), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5064) );
  INV_X1 U5838 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6146) );
  INV_X1 U5839 ( .A(n6685), .ZN(n6786) );
  INV_X1 U5840 ( .A(n5272), .ZN(n5271) );
  OAI21_X1 U5841 ( .B1(n8832), .B2(n5273), .A(n8823), .ZN(n5272) );
  INV_X1 U5842 ( .A(n6650), .ZN(n5273) );
  OR2_X1 U5843 ( .A1(n9192), .A2(n7978), .ZN(n6651) );
  AND2_X1 U5844 ( .A1(n6579), .A2(n8853), .ZN(n6644) );
  NAND2_X1 U5845 ( .A1(n6642), .A2(n5281), .ZN(n5279) );
  NAND2_X1 U5846 ( .A1(n5282), .A2(n6639), .ZN(n5281) );
  INV_X1 U5847 ( .A(n6643), .ZN(n5282) );
  NAND2_X1 U5848 ( .A1(n9210), .A2(n8232), .ZN(n6579) );
  OR2_X1 U5849 ( .A1(n9210), .A2(n8232), .ZN(n6645) );
  INV_X1 U5850 ( .A(n4744), .ZN(n4743) );
  OAI21_X1 U5851 ( .B1(n8916), .B2(n6481), .A(n6637), .ZN(n4744) );
  NAND2_X1 U5852 ( .A1(n5265), .A2(n6633), .ZN(n5264) );
  INV_X1 U5853 ( .A(n6631), .ZN(n5265) );
  INV_X1 U5854 ( .A(n6619), .ZN(n4750) );
  NOR2_X1 U5855 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  INV_X1 U5856 ( .A(n9017), .ZN(n4843) );
  AND2_X1 U5857 ( .A1(n6617), .A2(n9020), .ZN(n6618) );
  NOR2_X2 U5858 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6101) );
  INV_X1 U5859 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6104) );
  INV_X1 U5860 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6103) );
  INV_X1 U5861 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6133) );
  INV_X1 U5862 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U5863 ( .A1(n6377), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U5864 ( .A1(n6206), .A2(n6205), .ZN(n6343) );
  INV_X1 U5865 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6205) );
  INV_X1 U5866 ( .A(n6304), .ZN(n6206) );
  OR2_X1 U5867 ( .A1(n6292), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6304) );
  INV_X1 U5868 ( .A(n5407), .ZN(n5347) );
  NOR2_X1 U5869 ( .A1(n5627), .A2(n5626), .ZN(n4893) );
  NOR2_X1 U5870 ( .A1(n5666), .A2(n5665), .ZN(n5682) );
  NAND2_X1 U5871 ( .A1(n5348), .A2(n5407), .ZN(n9411) );
  NAND2_X1 U5872 ( .A1(n9313), .A2(n5416), .ZN(n5348) );
  NOR2_X1 U5873 ( .A1(n4634), .A2(n10166), .ZN(n4633) );
  OAI21_X1 U5874 ( .B1(n9730), .B2(n9791), .A(n9814), .ZN(n4634) );
  NAND2_X1 U5875 ( .A1(n9730), .A2(n9792), .ZN(n4639) );
  INV_X1 U5876 ( .A(n9735), .ZN(n6085) );
  AND2_X1 U5877 ( .A1(n10166), .A2(n9734), .ZN(n9732) );
  NOR2_X1 U5878 ( .A1(n10016), .A2(n10174), .ZN(n5399) );
  NOR2_X1 U5879 ( .A1(n10005), .A2(n5377), .ZN(n5376) );
  AOI21_X1 U5880 ( .B1(n4653), .B2(n5192), .A(n5188), .ZN(n5187) );
  NAND2_X1 U5881 ( .A1(n10125), .A2(n4653), .ZN(n5189) );
  NAND2_X1 U5882 ( .A1(n5194), .A2(n5195), .ZN(n5193) );
  INV_X1 U5883 ( .A(n6060), .ZN(n5194) );
  NAND2_X1 U5884 ( .A1(n4892), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5753) );
  INV_X1 U5885 ( .A(n4892), .ZN(n5734) );
  OR2_X1 U5886 ( .A1(n8039), .A2(n9831), .ZN(n5236) );
  AND2_X1 U5887 ( .A1(n5236), .A2(n5237), .ZN(n5227) );
  INV_X1 U5888 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5608) );
  OR2_X1 U5889 ( .A1(n5609), .A2(n5608), .ZN(n5627) );
  INV_X1 U5890 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5553) );
  AND2_X1 U5891 ( .A1(n9590), .A2(n9755), .ZN(n7816) );
  AND2_X1 U5892 ( .A1(n5995), .A2(n5983), .ZN(n5993) );
  INV_X1 U5893 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U5894 ( .A1(n4967), .A2(n4969), .ZN(n5854) );
  NAND2_X1 U5895 ( .A1(n5786), .A2(n5784), .ZN(n4968) );
  NAND2_X1 U5896 ( .A1(n5742), .A2(n5741), .ZN(n5743) );
  NAND2_X1 U5897 ( .A1(n5337), .A2(n4466), .ZN(n4977) );
  NAND2_X1 U5898 ( .A1(n5338), .A2(n5690), .ZN(n5337) );
  NOR2_X1 U5899 ( .A1(n5339), .A2(n4522), .ZN(n4975) );
  AND2_X1 U5900 ( .A1(n5674), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5638) );
  AOI21_X1 U5901 ( .B1(n5585), .B2(n5350), .A(n4508), .ZN(n5349) );
  AND2_X1 U5902 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  INV_X1 U5903 ( .A(n6704), .ZN(n5322) );
  NOR2_X1 U5904 ( .A1(n8238), .A2(n5310), .ZN(n5309) );
  INV_X1 U5905 ( .A(n6728), .ZN(n5310) );
  OR2_X1 U5906 ( .A1(n6727), .A2(n8953), .ZN(n6728) );
  NAND2_X1 U5907 ( .A1(n7384), .A2(n6145), .ZN(n6284) );
  INV_X1 U5908 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U5909 ( .A1(n7212), .A2(n6239), .ZN(n6582) );
  OR2_X1 U5910 ( .A1(n6718), .A2(n8291), .ZN(n6719) );
  NAND2_X1 U5911 ( .A1(n7682), .A2(n6710), .ZN(n8286) );
  XNOR2_X1 U5912 ( .A(n6693), .B(n7357), .ZN(n6695) );
  AND2_X1 U5913 ( .A1(n6783), .A2(n6244), .ZN(n6853) );
  NAND2_X1 U5914 ( .A1(n5026), .A2(n5025), .ZN(n5024) );
  INV_X1 U5915 ( .A(n6563), .ZN(n5025) );
  INV_X1 U5916 ( .A(n6564), .ZN(n5026) );
  AOI21_X1 U5917 ( .B1(n6565), .B2(n6563), .A(n6564), .ZN(n6569) );
  AND2_X1 U5918 ( .A1(n6471), .A2(n6470), .ZN(n8204) );
  AND4_X1 U5919 ( .A1(n6278), .A2(n4510), .A3(n6277), .A4(n6276), .ZN(n6809)
         );
  OR2_X1 U5920 ( .A1(n4429), .A2(n7174), .ZN(n6229) );
  NAND2_X1 U5921 ( .A1(n7317), .A2(n7173), .ZN(n4676) );
  AND2_X1 U5922 ( .A1(n4678), .A2(n4677), .ZN(n7214) );
  NAND2_X1 U5923 ( .A1(n7173), .A2(n7174), .ZN(n4677) );
  NOR2_X1 U5924 ( .A1(n7309), .A2(n7182), .ZN(n7217) );
  OAI21_X1 U5925 ( .B1(n7175), .B2(n7162), .A(n7223), .ZN(n10508) );
  INV_X1 U5926 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n6100) );
  NAND2_X1 U5927 ( .A1(n7177), .A2(n5298), .ZN(n5083) );
  INV_X1 U5928 ( .A(n7178), .ZN(n4663) );
  AND2_X1 U5929 ( .A1(n5300), .A2(n4760), .ZN(n7187) );
  AND2_X1 U5930 ( .A1(n4664), .A2(n4663), .ZN(n7228) );
  NOR2_X1 U5931 ( .A1(n7272), .A2(n4847), .ZN(n7234) );
  AND2_X1 U5932 ( .A1(n7233), .A2(n7269), .ZN(n4847) );
  AOI21_X1 U5933 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7229), .A(n7228), .ZN(
        n7268) );
  NAND2_X1 U5934 ( .A1(n4756), .A2(n4754), .ZN(n7556) );
  OR2_X1 U5935 ( .A1(n6343), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U5936 ( .A1(n4765), .A2(n4764), .ZN(n7754) );
  NAND2_X1 U5937 ( .A1(n5082), .A2(n5081), .ZN(n5080) );
  NAND2_X1 U5938 ( .A1(n7755), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U5939 ( .A1(n8346), .A2(n8345), .B1(n8344), .B2(n8343), .ZN(n8363)
         );
  OAI22_X1 U5940 ( .A1(n8363), .A2(n8362), .B1(n8361), .B2(n8360), .ZN(n8385)
         );
  AOI21_X1 U5941 ( .B1(n8399), .B2(n8398), .A(n4562), .ZN(n8418) );
  AOI21_X1 U5942 ( .B1(n8426), .B2(n8425), .A(n4553), .ZN(n8445) );
  NAND2_X1 U5943 ( .A1(n4863), .A2(n8469), .ZN(n8452) );
  AOI21_X1 U5944 ( .B1(n8440), .B2(n5103), .A(n8463), .ZN(n5091) );
  NAND2_X1 U5945 ( .A1(n5088), .A2(n5086), .ZN(n5097) );
  XNOR2_X1 U5946 ( .A(n8754), .B(n4879), .ZN(n8757) );
  AND2_X1 U5947 ( .A1(n6244), .A2(P2_B_REG_SCAN_IN), .ZN(n6854) );
  NAND2_X1 U5948 ( .A1(n6157), .A2(n5076), .ZN(n6522) );
  INV_X1 U5949 ( .A(n4580), .ZN(n6501) );
  OR2_X1 U5950 ( .A1(n8891), .A2(n5154), .ZN(n8851) );
  AOI21_X1 U5951 ( .B1(n8899), .B2(n6534), .A(n6479), .ZN(n8882) );
  NAND2_X1 U5952 ( .A1(n6464), .A2(n6154), .ZN(n6487) );
  NAND2_X1 U5953 ( .A1(n6425), .A2(n4455), .ZN(n6465) );
  INV_X1 U5954 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U5955 ( .A1(n6425), .A2(n5070), .ZN(n6457) );
  NAND2_X1 U5956 ( .A1(n6425), .A2(n6153), .ZN(n6449) );
  INV_X1 U5957 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5072) );
  AND2_X1 U5958 ( .A1(n5419), .A2(n6825), .ZN(n8967) );
  NAND2_X1 U5959 ( .A1(n6151), .A2(n5073), .ZN(n6410) );
  NAND2_X1 U5960 ( .A1(n6151), .A2(n6150), .ZN(n6398) );
  NAND2_X1 U5961 ( .A1(n5062), .A2(n8712), .ZN(n6385) );
  INV_X1 U5962 ( .A(n6221), .ZN(n5062) );
  NAND2_X1 U5963 ( .A1(n5064), .A2(n5063), .ZN(n6221) );
  INV_X1 U5964 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5063) );
  INV_X1 U5965 ( .A(n5064), .ZN(n6356) );
  OR2_X1 U5966 ( .A1(n6337), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6327) );
  AND4_X1 U5967 ( .A1(n6320), .A2(n6319), .A3(n6318), .A4(n6317), .ZN(n7655)
         );
  NOR2_X1 U5968 ( .A1(n7593), .A2(n5151), .ZN(n5150) );
  INV_X1 U5969 ( .A(n6815), .ZN(n5151) );
  NAND2_X1 U5970 ( .A1(n7425), .A2(n7426), .ZN(n5152) );
  NAND2_X1 U5971 ( .A1(n4575), .A2(n6146), .ZN(n6298) );
  INV_X1 U5972 ( .A(n6284), .ZN(n4575) );
  NOR2_X1 U5973 ( .A1(n6610), .A2(n6584), .ZN(n7492) );
  OR2_X1 U5974 ( .A1(n6275), .A2(n6246), .ZN(n6249) );
  NAND2_X1 U5975 ( .A1(n10557), .A2(n9007), .ZN(n5170) );
  NAND2_X1 U5976 ( .A1(n6544), .A2(n6543), .ZN(n6870) );
  NAND2_X1 U5977 ( .A1(n8826), .A2(n9065), .ZN(n4800) );
  NOR2_X1 U5978 ( .A1(n4467), .A2(n5148), .ZN(n5145) );
  INV_X1 U5979 ( .A(n6507), .ZN(n8832) );
  NAND2_X1 U5980 ( .A1(n8858), .A2(n9065), .ZN(n4883) );
  NAND2_X1 U5981 ( .A1(n8850), .A2(n6639), .ZN(n8892) );
  AOI21_X1 U5982 ( .B1(n8917), .B2(n8915), .A(n4831), .ZN(n8906) );
  AND2_X1 U5983 ( .A1(n9238), .A2(n8907), .ZN(n4831) );
  NAND2_X1 U5984 ( .A1(n6448), .A2(n6447), .ZN(n6830) );
  INV_X1 U5985 ( .A(n6827), .ZN(n8940) );
  NAND2_X1 U5986 ( .A1(n5161), .A2(n6825), .ZN(n8937) );
  OR2_X1 U5987 ( .A1(n8962), .A2(n5167), .ZN(n5161) );
  OR2_X1 U5988 ( .A1(n8937), .A2(n8952), .ZN(n8956) );
  INV_X1 U5989 ( .A(n9064), .ZN(n9010) );
  INV_X1 U5990 ( .A(n6826), .ZN(n8952) );
  AND2_X1 U5991 ( .A1(n4736), .A2(n6629), .ZN(n4735) );
  NAND2_X1 U5992 ( .A1(n6628), .A2(n4737), .ZN(n4736) );
  INV_X1 U5993 ( .A(n6628), .ZN(n4738) );
  AND2_X1 U5994 ( .A1(n6626), .A2(n6625), .ZN(n8984) );
  NAND2_X1 U5995 ( .A1(n8989), .A2(n6822), .ZN(n4720) );
  NAND2_X1 U5996 ( .A1(n4749), .A2(n6619), .ZN(n9001) );
  NAND2_X1 U5997 ( .A1(n4840), .A2(n6618), .ZN(n4749) );
  AND2_X1 U5998 ( .A1(n6588), .A2(n6609), .ZN(n7431) );
  OR2_X1 U5999 ( .A1(n6886), .A2(n6685), .ZN(n7336) );
  AND2_X1 U6000 ( .A1(n6793), .A2(n6929), .ZN(n6865) );
  NOR2_X1 U6001 ( .A1(n6789), .A2(n6771), .ZN(n6863) );
  OR2_X1 U6002 ( .A1(n10516), .A2(n6780), .ZN(n10525) );
  AND2_X1 U6003 ( .A1(n6182), .A2(n4930), .ZN(n6185) );
  AND2_X1 U6004 ( .A1(n6136), .A2(n6137), .ZN(n4930) );
  INV_X1 U6005 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6178) );
  INV_X1 U6006 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6113) );
  INV_X1 U6007 ( .A(n6182), .ZN(n6292) );
  NAND2_X1 U6008 ( .A1(n4798), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5609) );
  INV_X1 U6009 ( .A(n5574), .ZN(n4798) );
  NAND2_X1 U6010 ( .A1(n5335), .A2(n5333), .ZN(n5332) );
  INV_X1 U6011 ( .A(n4893), .ZN(n5643) );
  NAND2_X1 U6012 ( .A1(n4527), .A2(n4620), .ZN(n9384) );
  NAND2_X1 U6013 ( .A1(n8029), .A2(n4496), .ZN(n4620) );
  NOR2_X1 U6014 ( .A1(n8090), .A2(n5345), .ZN(n5344) );
  OR2_X1 U6015 ( .A1(n5347), .A2(n5346), .ZN(n5345) );
  INV_X1 U6016 ( .A(n9464), .ZN(n5346) );
  NAND2_X1 U6017 ( .A1(n4610), .A2(n9425), .ZN(n9428) );
  AOI21_X1 U6018 ( .B1(n5056), .B2(n5053), .A(n9426), .ZN(n5052) );
  INV_X1 U6019 ( .A(n5056), .ZN(n5054) );
  OR2_X1 U6020 ( .A1(n5819), .A2(n5818), .ZN(n5833) );
  OR2_X1 U6021 ( .A1(n9377), .A2(n8115), .ZN(n4612) );
  INV_X1 U6022 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5665) );
  INV_X1 U6023 ( .A(n5682), .ZN(n5684) );
  XNOR2_X1 U6024 ( .A(n7119), .B(n8141), .ZN(n7196) );
  NAND2_X1 U6025 ( .A1(n7461), .A2(n7460), .ZN(n9518) );
  INV_X1 U6026 ( .A(n4420), .ZN(n9535) );
  OR2_X1 U6027 ( .A1(n10407), .A2(n7605), .ZN(n7087) );
  INV_X1 U6028 ( .A(n9732), .ZN(n9801) );
  OR2_X1 U6029 ( .A1(n9352), .A2(n5557), .ZN(n6008) );
  AND3_X1 U6030 ( .A1(n5781), .A2(n5780), .A3(n5779), .ZN(n9506) );
  AND4_X1 U6031 ( .A1(n5689), .A2(n5688), .A3(n5687), .A4(n5686), .ZN(n9605)
         );
  AND4_X1 U6032 ( .A1(n5650), .A2(n5649), .A3(n5648), .A4(n5647), .ZN(n8037)
         );
  OR2_X1 U6033 ( .A1(n6081), .A2(n6963), .ZN(n5533) );
  NAND2_X1 U6034 ( .A1(n4438), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U6035 ( .A1(n5552), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5435) );
  OR2_X1 U6036 ( .A1(n7020), .A2(n7019), .ZN(n7022) );
  OR2_X1 U6037 ( .A1(n7044), .A2(n7043), .ZN(n7041) );
  NOR2_X1 U6038 ( .A1(n7391), .A2(n4559), .ZN(n7394) );
  NOR2_X1 U6039 ( .A1(n7394), .A2(n7393), .ZN(n7581) );
  AOI21_X1 U6040 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7582), .A(n7581), .ZN(
        n9929) );
  NOR2_X1 U6041 ( .A1(n9933), .A2(n9932), .ZN(n9941) );
  NAND2_X1 U6042 ( .A1(n7872), .A2(n7871), .ZN(n7886) );
  NAND2_X1 U6043 ( .A1(n7891), .A2(n5380), .ZN(n4640) );
  AND2_X1 U6044 ( .A1(n7890), .A2(n7888), .ZN(n5380) );
  AND2_X1 U6045 ( .A1(n7889), .A2(n4794), .ZN(n4793) );
  NAND2_X1 U6046 ( .A1(n7890), .A2(n4795), .ZN(n4794) );
  NAND2_X1 U6047 ( .A1(n10014), .A2(n5399), .ZN(n10000) );
  INV_X1 U6048 ( .A(n5379), .ZN(n5378) );
  NAND2_X1 U6049 ( .A1(n5376), .A2(n9655), .ZN(n5375) );
  OAI21_X1 U6050 ( .B1(n10005), .B2(n5381), .A(n9647), .ZN(n5379) );
  NAND2_X1 U6051 ( .A1(n10014), .A2(n10180), .ZN(n10013) );
  INV_X1 U6052 ( .A(n5897), .ZN(n5896) );
  NAND2_X1 U6053 ( .A1(n6087), .A2(n4448), .ZN(n10037) );
  NAND2_X1 U6054 ( .A1(n6087), .A2(n5391), .ZN(n7935) );
  NOR2_X1 U6055 ( .A1(n10086), .A2(n5392), .ZN(n10060) );
  NAND2_X1 U6056 ( .A1(n4876), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5819) );
  INV_X1 U6057 ( .A(n9681), .ZN(n4853) );
  NOR2_X1 U6058 ( .A1(n5395), .A2(n8026), .ZN(n5394) );
  INV_X1 U6059 ( .A(n5396), .ZN(n5395) );
  NAND2_X1 U6060 ( .A1(n10368), .A2(n5396), .ZN(n7788) );
  NAND2_X1 U6061 ( .A1(n10368), .A2(n10455), .ZN(n7673) );
  NAND2_X1 U6062 ( .A1(n4797), .A2(n10432), .ZN(n10389) );
  INV_X1 U6063 ( .A(n9568), .ZN(n4845) );
  INV_X1 U6064 ( .A(n7068), .ZN(n7065) );
  AND2_X1 U6065 ( .A1(n7888), .A2(n9648), .ZN(n9694) );
  NAND2_X1 U6066 ( .A1(n5253), .A2(n5246), .ZN(n5245) );
  NAND2_X1 U6067 ( .A1(n5248), .A2(n5250), .ZN(n5247) );
  AOI21_X1 U6068 ( .B1(n4951), .B2(n4949), .A(n5249), .ZN(n4948) );
  INV_X1 U6069 ( .A(n4953), .ZN(n4949) );
  NOR2_X1 U6070 ( .A1(n5922), .A2(n4954), .ZN(n4953) );
  INV_X1 U6071 ( .A(n5904), .ZN(n4954) );
  AOI21_X1 U6072 ( .B1(n4442), .B2(n4440), .A(n4497), .ZN(n4935) );
  NAND2_X1 U6073 ( .A1(n5798), .A2(n4442), .ZN(n4936) );
  NAND2_X1 U6074 ( .A1(n10474), .A2(n9601), .ZN(n4945) );
  INV_X1 U6075 ( .A(n7816), .ZN(n9682) );
  INV_X1 U6076 ( .A(n10390), .ZN(n10475) );
  OR2_X1 U6077 ( .A1(n9791), .A2(n4613), .ZN(n10451) );
  XNOR2_X1 U6078 ( .A(n6542), .B(SI_29_), .ZN(n9298) );
  NAND2_X1 U6079 ( .A1(n5430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U6080 ( .A(n5994), .B(n5993), .ZN(n9304) );
  INV_X1 U6081 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U6082 ( .A1(n6016), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6018) );
  XNOR2_X1 U6083 ( .A(n5828), .B(n5827), .ZN(n7765) );
  NOR2_X1 U6084 ( .A1(n5386), .A2(n5771), .ZN(n5385) );
  NAND2_X1 U6085 ( .A1(n5604), .A2(n5387), .ZN(n5386) );
  INV_X1 U6086 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5387) );
  OAI21_X1 U6087 ( .B1(n5636), .B2(n5339), .A(n5338), .ZN(n5693) );
  NAND2_X1 U6088 ( .A1(n5651), .A2(n5340), .ZN(n4656) );
  INV_X1 U6089 ( .A(n5651), .ZN(n4657) );
  INV_X1 U6090 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5330) );
  INV_X1 U6091 ( .A(n4902), .ZN(n8201) );
  AOI21_X1 U6092 ( .B1(n8299), .B2(n8298), .A(n4461), .ZN(n4902) );
  AND2_X1 U6093 ( .A1(n6494), .A2(n6493), .ZN(n8213) );
  NAND2_X1 U6094 ( .A1(n4901), .A2(n5304), .ZN(n4900) );
  AOI21_X1 U6095 ( .B1(n5306), .B2(n5308), .A(n4507), .ZN(n5304) );
  NAND2_X1 U6096 ( .A1(n4903), .A2(n4461), .ZN(n4901) );
  INV_X1 U6097 ( .A(n8218), .ZN(n4914) );
  OAI21_X1 U6098 ( .B1(n7682), .B2(n4919), .A(n4916), .ZN(n8219) );
  AND2_X1 U6099 ( .A1(n6188), .A2(n6187), .ZN(n8236) );
  NAND2_X1 U6100 ( .A1(n8321), .A2(n6728), .ZN(n8237) );
  AND4_X1 U6101 ( .A1(n6303), .A2(n6302), .A3(n6301), .A4(n6300), .ZN(n7596)
         );
  NAND2_X1 U6102 ( .A1(n5305), .A2(n6735), .ZN(n8260) );
  NAND2_X1 U6103 ( .A1(n8201), .A2(n8202), .ZN(n5305) );
  NAND2_X1 U6104 ( .A1(n8217), .A2(n6719), .ZN(n8268) );
  NOR2_X1 U6105 ( .A1(n7144), .A2(n6692), .ZN(n7151) );
  AND4_X1 U6106 ( .A1(n6342), .A2(n6341), .A3(n6340), .A4(n6339), .ZN(n7656)
         );
  NAND2_X1 U6107 ( .A1(n7509), .A2(n6702), .ZN(n7447) );
  AND2_X1 U6108 ( .A1(n6195), .A2(n6194), .ZN(n8314) );
  INV_X1 U6109 ( .A(n8324), .ZN(n8313) );
  NAND2_X1 U6110 ( .A1(n8323), .A2(n8322), .ZN(n8321) );
  NAND2_X1 U6111 ( .A1(n6409), .A2(n6408), .ZN(n9144) );
  AND2_X1 U6112 ( .A1(n4586), .A2(n4577), .ZN(n5133) );
  NOR2_X1 U6113 ( .A1(n5138), .A2(n5135), .ZN(n4577) );
  INV_X1 U6114 ( .A(n6574), .ZN(n5138) );
  OAI211_X1 U6115 ( .C1(n4586), .C2(n4585), .A(n4835), .B(n4524), .ZN(n4878)
         );
  INV_X1 U6116 ( .A(n5137), .ZN(n4585) );
  AND2_X1 U6117 ( .A1(n6562), .A2(n6169), .ZN(n8808) );
  INV_X1 U6118 ( .A(n7976), .ZN(n8817) );
  NAND2_X1 U6119 ( .A1(n6528), .A2(n6527), .ZN(n8834) );
  INV_X1 U6120 ( .A(n8204), .ZN(n8918) );
  INV_X1 U6121 ( .A(n7656), .ZN(n8336) );
  OR2_X1 U6122 ( .A1(n7170), .A2(P2_U3151), .ZN(n8774) );
  NAND2_X1 U6123 ( .A1(n7305), .A2(n4998), .ZN(n7225) );
  OR2_X1 U6124 ( .A1(n7160), .A2(n4679), .ZN(n4998) );
  NAND2_X1 U6125 ( .A1(n5299), .A2(n5300), .ZN(n10495) );
  NAND2_X1 U6126 ( .A1(n7240), .A2(n5000), .ZN(n7244) );
  OR2_X1 U6127 ( .A1(n7241), .A2(n7242), .ZN(n5000) );
  XNOR2_X1 U6128 ( .A(n7268), .B(n7269), .ZN(n7271) );
  AND2_X1 U6129 ( .A1(n7558), .A2(n7573), .ZN(n7559) );
  INV_X1 U6130 ( .A(n4758), .ZN(n7558) );
  NAND2_X1 U6131 ( .A1(n7621), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7620) );
  XNOR2_X1 U6132 ( .A(n7553), .B(n7573), .ZN(n7619) );
  INV_X1 U6133 ( .A(n5004), .ZN(n7626) );
  OAI22_X1 U6134 ( .A1(n7619), .A2(n7691), .B1(n7573), .B2(n7553), .ZN(n7748)
         );
  XNOR2_X1 U6135 ( .A(n5080), .B(n5079), .ZN(n8341) );
  NAND2_X1 U6136 ( .A1(n5303), .A2(n5301), .ZN(n7757) );
  OAI21_X1 U6137 ( .B1(n8341), .B2(n9170), .A(n5078), .ZN(n8359) );
  NAND2_X1 U6138 ( .A1(n5080), .A2(n5079), .ZN(n5078) );
  XNOR2_X1 U6139 ( .A(n8379), .B(n8383), .ZN(n8380) );
  OAI22_X1 U6140 ( .A1(n8380), .A2(n9158), .B1(n8379), .B2(n8383), .ZN(n8399)
         );
  OAI21_X1 U6141 ( .B1(n8389), .B2(n8391), .A(n8390), .ZN(n8406) );
  XNOR2_X1 U6142 ( .A(n8418), .B(n8420), .ZN(n8421) );
  NAND2_X1 U6143 ( .A1(n5291), .A2(n8431), .ZN(n8411) );
  INV_X1 U6144 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n4864) );
  INV_X1 U6145 ( .A(n8773), .ZN(n8787) );
  NAND2_X1 U6146 ( .A1(n4670), .A2(n4668), .ZN(n4667) );
  NAND2_X1 U6147 ( .A1(n8936), .A2(n6633), .ZN(n8928) );
  NAND2_X1 U6148 ( .A1(n6436), .A2(n6435), .ZN(n8948) );
  OR2_X1 U6149 ( .A1(n7341), .A2(n8995), .ZN(n9090) );
  OAI211_X1 U6150 ( .C1(n6306), .C2(n6907), .A(n6282), .B(n6281), .ZN(n7421)
         );
  INV_X1 U6151 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7384) );
  NOR2_X1 U6152 ( .A1(n7954), .A2(n4705), .ZN(n10526) );
  OAI21_X1 U6153 ( .B1(n6244), .B2(n4751), .A(n4587), .ZN(n7344) );
  NAND2_X1 U6154 ( .A1(n6244), .A2(n9312), .ZN(n4587) );
  NAND2_X1 U6155 ( .A1(n6556), .A2(n6555), .ZN(n9099) );
  INV_X1 U6156 ( .A(n9099), .ZN(n9183) );
  INV_X1 U6157 ( .A(n6870), .ZN(n8129) );
  NAND2_X1 U6158 ( .A1(n6171), .A2(n6170), .ZN(n9198) );
  INV_X1 U6159 ( .A(n8236), .ZN(n9204) );
  NAND2_X1 U6160 ( .A1(n5143), .A2(n5146), .ZN(n8840) );
  NAND2_X1 U6161 ( .A1(n6834), .A2(n4467), .ZN(n5143) );
  AND2_X1 U6162 ( .A1(n6486), .A2(n6485), .ZN(n9223) );
  NAND2_X1 U6163 ( .A1(n6474), .A2(n6473), .ZN(n9226) );
  NAND2_X1 U6164 ( .A1(n6463), .A2(n6462), .ZN(n9232) );
  NAND2_X1 U6165 ( .A1(n8914), .A2(n8916), .ZN(n4742) );
  INV_X1 U6166 ( .A(n6830), .ZN(n9245) );
  NAND2_X1 U6167 ( .A1(n6424), .A2(n6423), .ZN(n9253) );
  NAND2_X1 U6168 ( .A1(n6397), .A2(n6396), .ZN(n9260) );
  AND2_X1 U6169 ( .A1(n8993), .A2(n8992), .ZN(n9264) );
  NAND2_X1 U6170 ( .A1(n6384), .A2(n6383), .ZN(n9266) );
  NAND2_X1 U6171 ( .A1(n9003), .A2(n6621), .ZN(n8988) );
  NAND2_X1 U6172 ( .A1(n4709), .A2(n4708), .ZN(n4711) );
  NAND2_X1 U6173 ( .A1(n5285), .A2(n6611), .ZN(n7599) );
  AND2_X1 U6174 ( .A1(n6158), .A2(n6161), .ZN(n5158) );
  INV_X1 U6175 ( .A(n4746), .ZN(n6159) );
  INV_X1 U6176 ( .A(n6669), .ZN(n6671) );
  NAND2_X1 U6177 ( .A1(n6672), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6673) );
  INV_X1 U6178 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8563) );
  INV_X1 U6179 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7603) );
  INV_X1 U6180 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7476) );
  INV_X1 U6181 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n8654) );
  INV_X1 U6182 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6992) );
  INV_X1 U6183 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6935) );
  INV_X1 U6184 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6932) );
  INV_X1 U6185 ( .A(n7242), .ZN(n7229) );
  NAND2_X1 U6186 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n8579), .ZN(n4869) );
  CLKBUF_X1 U6187 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n4848) );
  NAND2_X1 U6188 ( .A1(n5055), .A2(n4458), .ZN(n8119) );
  OR2_X1 U6189 ( .A1(n9477), .A2(n5058), .ZN(n5055) );
  NAND2_X1 U6190 ( .A1(n5040), .A2(n5041), .ZN(n9337) );
  NAND2_X1 U6191 ( .A1(n9498), .A2(n5042), .ZN(n5040) );
  NAND2_X1 U6192 ( .A1(n5050), .A2(n4488), .ZN(n9362) );
  NAND2_X1 U6193 ( .A1(n5049), .A2(n9533), .ZN(n5048) );
  NAND2_X1 U6194 ( .A1(n5752), .A2(n5751), .ZN(n10220) );
  NAND2_X1 U6195 ( .A1(n5775), .A2(n5774), .ZN(n10215) );
  NAND2_X1 U6196 ( .A1(n7293), .A2(n7292), .ZN(n7461) );
  NAND2_X1 U6197 ( .A1(n8029), .A2(n8028), .ZN(n9441) );
  NAND2_X1 U6198 ( .A1(n4618), .A2(n4616), .ZN(n9455) );
  AOI21_X1 U6199 ( .B1(n4445), .B2(n4617), .A(n4526), .ZN(n4616) );
  NAND2_X1 U6200 ( .A1(n7813), .A2(n5637), .ZN(n5832) );
  NAND2_X1 U6201 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  INV_X1 U6202 ( .A(n5045), .ZN(n4622) );
  INV_X1 U6203 ( .A(n8029), .ZN(n4623) );
  XNOR2_X1 U6204 ( .A(n7196), .B(n7195), .ZN(n7125) );
  NAND2_X1 U6205 ( .A1(n7122), .A2(n4607), .ZN(n7124) );
  INV_X1 U6206 ( .A(n5326), .ZN(n7123) );
  AOI21_X1 U6207 ( .B1(n9498), .B2(n8102), .A(n4464), .ZN(n9502) );
  NAND2_X1 U6208 ( .A1(n7207), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9554) );
  NAND2_X1 U6209 ( .A1(n5384), .A2(n5383), .ZN(n5382) );
  INV_X1 U6210 ( .A(n9534), .ZN(n5383) );
  NAND2_X1 U6211 ( .A1(n9531), .A2(n9530), .ZN(n5384) );
  INV_X1 U6212 ( .A(n9552), .ZN(n9542) );
  OR2_X1 U6213 ( .A1(n7087), .A2(n9787), .ZN(n9552) );
  INV_X1 U6214 ( .A(n9545), .ZN(n9557) );
  NAND2_X1 U6215 ( .A1(n9795), .A2(n9794), .ZN(n9804) );
  NAND2_X1 U6216 ( .A1(n5920), .A2(n5919), .ZN(n9818) );
  NAND2_X1 U6217 ( .A1(n5881), .A2(n5880), .ZN(n9819) );
  OR2_X1 U6218 ( .A1(n5758), .A2(n5757), .ZN(n9825) );
  INV_X1 U6219 ( .A(n9605), .ZN(n9829) );
  INV_X1 U6220 ( .A(n8037), .ZN(n9831) );
  INV_X1 U6221 ( .A(n7526), .ZN(n9834) );
  NAND2_X1 U6222 ( .A1(n4436), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5560) );
  OR2_X2 U6223 ( .A1(n6920), .A2(n10311), .ZN(n9839) );
  NAND2_X1 U6224 ( .A1(n9856), .A2(n9857), .ZN(n9855) );
  NAND2_X1 U6225 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  NAND2_X1 U6226 ( .A1(n6986), .A2(n6987), .ZN(n6994) );
  OR2_X1 U6227 ( .A1(n7016), .A2(n7017), .ZN(n7014) );
  AND2_X1 U6228 ( .A1(n6985), .A2(n8005), .ZN(n9988) );
  NOR2_X1 U6229 ( .A1(n7045), .A2(n4560), .ZN(n6997) );
  NAND2_X1 U6230 ( .A1(n7029), .A2(n7030), .ZN(n7248) );
  NAND2_X1 U6231 ( .A1(n7248), .A2(n4784), .ZN(n7250) );
  OR2_X1 U6232 ( .A1(n7249), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4784) );
  OR2_X1 U6233 ( .A1(n9970), .A2(n9969), .ZN(n9981) );
  INV_X1 U6234 ( .A(n7886), .ZN(n7906) );
  AND2_X1 U6235 ( .A1(n5986), .A2(n5966), .ZN(n10015) );
  AOI21_X1 U6236 ( .B1(n10010), .B2(n10377), .A(n10009), .ZN(n10179) );
  NAND2_X1 U6237 ( .A1(n5016), .A2(n9702), .ZN(n10024) );
  NAND2_X1 U6238 ( .A1(n10125), .A2(n6069), .ZN(n5190) );
  INV_X1 U6239 ( .A(n6067), .ZN(n10112) );
  INV_X1 U6240 ( .A(n10215), .ZN(n10116) );
  INV_X1 U6241 ( .A(n10225), .ZN(n10160) );
  AND2_X1 U6242 ( .A1(n5196), .A2(n9756), .ZN(n7851) );
  NAND2_X1 U6243 ( .A1(n5229), .A2(n5230), .ZN(n10348) );
  INV_X1 U6244 ( .A(n5607), .ZN(n4813) );
  NAND2_X1 U6245 ( .A1(n7702), .A2(n6052), .ZN(n5198) );
  INV_X2 U6246 ( .A(n10421), .ZN(n5481) );
  OAI21_X1 U6247 ( .B1(n10168), .B2(n10473), .A(n10167), .ZN(n10169) );
  NAND2_X1 U6248 ( .A1(n10179), .A2(n5207), .ZN(n10258) );
  AND2_X1 U6249 ( .A1(n10178), .A2(n5208), .ZN(n5207) );
  NAND2_X1 U6250 ( .A1(n10016), .A2(n6090), .ZN(n5208) );
  OR2_X1 U6251 ( .A1(n5798), .A2(n4440), .ZN(n4937) );
  AND2_X1 U6252 ( .A1(n5240), .A2(n5243), .ZN(n10069) );
  NAND2_X1 U6253 ( .A1(n5798), .A2(n5241), .ZN(n5240) );
  NAND2_X1 U6254 ( .A1(n5213), .A2(n5217), .ZN(n10132) );
  NAND2_X1 U6255 ( .A1(n7849), .A2(n5218), .ZN(n5213) );
  AND2_X1 U6256 ( .A1(n5219), .A2(n5222), .ZN(n10147) );
  NAND2_X1 U6257 ( .A1(n7849), .A2(n5723), .ZN(n5219) );
  AND2_X2 U6258 ( .A1(n6096), .A2(n7090), .ZN(n10482) );
  AND2_X1 U6259 ( .A1(n7866), .A2(n6046), .ZN(n10409) );
  AOI21_X1 U6260 ( .B1(n5432), .B2(n4696), .A(n4695), .ZN(n4694) );
  NOR2_X1 U6261 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4695) );
  NOR2_X1 U6262 ( .A1(n4697), .A2(n10312), .ZN(n4696) );
  XNOR2_X1 U6263 ( .A(n6025), .B(n6024), .ZN(n10336) );
  NAND2_X1 U6264 ( .A1(n5948), .A2(n4957), .ZN(n5892) );
  NOR2_X1 U6265 ( .A1(n4551), .A2(n4958), .ZN(n4957) );
  INV_X1 U6266 ( .A(n5946), .ZN(n4958) );
  INV_X1 U6267 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8178) );
  OAI21_X1 U6268 ( .B1(n6016), .B2(n5364), .A(n4516), .ZN(n6013) );
  INV_X1 U6269 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7475) );
  INV_X1 U6270 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7329) );
  INV_X1 U6271 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7095) );
  INV_X1 U6272 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6937) );
  XNOR2_X1 U6273 ( .A(n5261), .B(n5585), .ZN(n6906) );
  NAND2_X1 U6274 ( .A1(n5550), .A2(n5549), .ZN(n5261) );
  INV_X1 U6275 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5210) );
  NOR2_X2 U6276 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7744) );
  NAND2_X1 U6277 ( .A1(n7167), .A2(n4588), .ZN(n6888) );
  NOR2_X1 U6278 ( .A1(n4589), .A2(n6454), .ZN(n4588) );
  OAI21_X1 U6279 ( .B1(n6839), .B2(n8332), .A(n6799), .ZN(n6800) );
  XNOR2_X1 U6280 ( .A(n8189), .B(n8881), .ZN(n8194) );
  NAND2_X1 U6281 ( .A1(n7984), .A2(n4479), .ZN(n7983) );
  INV_X1 U6282 ( .A(n4911), .ZN(n4910) );
  OAI21_X1 U6283 ( .B1(n6744), .B2(n8332), .A(n8258), .ZN(n4911) );
  INV_X1 U6284 ( .A(n5006), .ZN(n7568) );
  OAI211_X1 U6285 ( .C1(n5104), .C2(n5101), .A(n5099), .B(n5100), .ZN(n8460)
         );
  AND2_X1 U6286 ( .A1(n5095), .A2(n4689), .ZN(n8481) );
  AOI21_X1 U6287 ( .B1(n4997), .B2(n10499), .A(n4996), .ZN(n4995) );
  NOR2_X1 U6288 ( .A1(n4447), .A2(n4505), .ZN(n4880) );
  OAI21_X1 U6289 ( .B1(n8783), .B2(n8764), .A(n8763), .ZN(n8780) );
  INV_X1 U6290 ( .A(n4811), .ZN(n4810) );
  OAI21_X1 U6291 ( .B1(n9189), .B2(n9086), .A(n8820), .ZN(n4811) );
  AOI21_X1 U6292 ( .B1(n9208), .B2(n8861), .A(n8981), .ZN(n8862) );
  OAI21_X1 U6293 ( .B1(n5173), .B2(n5171), .A(n5168), .ZN(n9105) );
  OR2_X1 U6294 ( .A1(n5172), .A2(n6883), .ZN(n5171) );
  INV_X1 U6295 ( .A(n4804), .ZN(n4803) );
  OAI21_X1 U6296 ( .B1(n9195), .B2(n9162), .A(n4805), .ZN(n4804) );
  INV_X1 U6297 ( .A(n4833), .ZN(n4832) );
  OAI21_X1 U6298 ( .B1(n9189), .B2(n9280), .A(n9187), .ZN(n4833) );
  NAND2_X1 U6299 ( .A1(n4609), .A2(n4608), .ZN(P1_U3214) );
  AND2_X1 U6300 ( .A1(n8176), .A2(n4556), .ZN(n4608) );
  OAI21_X1 U6301 ( .B1(n8173), .B2(n9350), .A(n9533), .ZN(n4609) );
  OAI21_X1 U6302 ( .B1(n9987), .B2(n4887), .A(n4886), .ZN(n9993) );
  NAND2_X1 U6303 ( .A1(n4889), .A2(n4888), .ZN(n4887) );
  AOI21_X1 U6304 ( .B1(n7992), .B2(n10393), .A(n7991), .ZN(n7993) );
  NAND2_X1 U6305 ( .A1(n4941), .A2(n4940), .ZN(P1_U3266) );
  AOI21_X1 U6306 ( .B1(n10172), .B2(n10162), .A(n10007), .ZN(n4940) );
  NAND2_X1 U6307 ( .A1(n4851), .A2(n10181), .ZN(n4849) );
  NAND2_X1 U6308 ( .A1(n5206), .A2(n5205), .ZN(P1_U3548) );
  NAND2_X1 U6309 ( .A1(n10258), .A2(n10494), .ZN(n5206) );
  AOI22_X1 U6310 ( .A1(n10260), .A2(n10181), .B1(P1_REG1_REG_26__SCAN_IN), 
        .B2(n10492), .ZN(n5205) );
  NAND2_X1 U6311 ( .A1(n4868), .A2(n10181), .ZN(n4867) );
  INV_X1 U6312 ( .A(n7933), .ZN(n4868) );
  NAND2_X1 U6313 ( .A1(n4789), .A2(n4568), .ZN(P1_U3521) );
  NAND2_X1 U6314 ( .A1(n10255), .A2(n10482), .ZN(n4789) );
  INV_X1 U6315 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U6316 ( .A1(n4851), .A2(n6050), .ZN(n4850) );
  NAND2_X1 U6317 ( .A1(n7992), .A2(n6050), .ZN(n6095) );
  AOI21_X1 U6318 ( .B1(n6097), .B2(n10482), .A(n6093), .ZN(n6094) );
  NOR2_X1 U6319 ( .A1(n10482), .A2(n6092), .ZN(n6093) );
  MUX2_X1 U6320 ( .A(n7921), .B(n7923), .S(n10482), .Z(n7922) );
  OR2_X2 U6321 ( .A1(n7068), .A2(n7072), .ZN(n5421) );
  OR2_X1 U6322 ( .A1(n5415), .A2(n4476), .ZN(n4440) );
  NAND2_X1 U6323 ( .A1(n9406), .A2(n9536), .ZN(n5250) );
  INV_X1 U6324 ( .A(n5250), .ZN(n5249) );
  INV_X1 U6325 ( .A(n10506), .ZN(n5298) );
  INV_X1 U6326 ( .A(n9999), .ZN(n5009) );
  AND2_X1 U6327 ( .A1(n5651), .A2(n5635), .ZN(n4441) );
  AND2_X1 U6328 ( .A1(n4938), .A2(n4482), .ZN(n4442) );
  AND2_X1 U6329 ( .A1(n5423), .A2(n5517), .ZN(n5677) );
  NOR2_X1 U6330 ( .A1(n9488), .A2(n5410), .ZN(n4443) );
  INV_X1 U6331 ( .A(n9648), .ZN(n4795) );
  OR3_X1 U6332 ( .A1(n4470), .A2(n4848), .A3(n7159), .ZN(n4444) );
  OAI211_X1 U6333 ( .C1(n6306), .C2(n6893), .A(n6295), .B(n6294), .ZN(n10542)
         );
  INV_X1 U6334 ( .A(n6633), .ZN(n5266) );
  AND2_X1 U6335 ( .A1(n5039), .A2(n5041), .ZN(n4445) );
  NOR2_X1 U6336 ( .A1(n6481), .A2(n6480), .ZN(n4446) );
  AND2_X1 U6337 ( .A1(n8779), .A2(n8786), .ZN(n4447) );
  AOI21_X1 U6338 ( .B1(n5146), .B2(n5145), .A(n4530), .ZN(n5144) );
  AND2_X1 U6339 ( .A1(n10042), .A2(n5391), .ZN(n4448) );
  AND2_X1 U6340 ( .A1(n5944), .A2(n5943), .ZN(n9536) );
  AND2_X1 U6341 ( .A1(n5511), .A2(n5512), .ZN(n4449) );
  AND2_X1 U6342 ( .A1(n5256), .A2(n5247), .ZN(n4450) );
  NOR2_X1 U6343 ( .A1(n9198), .A2(n8841), .ZN(n4451) );
  AND2_X1 U6344 ( .A1(n5760), .A2(SI_16_), .ZN(n4452) );
  NAND3_X1 U6345 ( .A1(n4528), .A2(n4687), .A3(n5097), .ZN(n8754) );
  AND2_X1 U6346 ( .A1(n4762), .A2(n4885), .ZN(n4453) );
  AND2_X1 U6347 ( .A1(n6720), .A2(n6719), .ZN(n4454) );
  INV_X1 U6348 ( .A(n8463), .ZN(n5101) );
  XNOR2_X1 U6349 ( .A(n6018), .B(n6017), .ZN(n9784) );
  NAND2_X1 U6350 ( .A1(n5152), .A2(n6815), .ZN(n7590) );
  AND2_X1 U6351 ( .A1(n5070), .A2(n5069), .ZN(n4455) );
  INV_X1 U6352 ( .A(n10016), .ZN(n10180) );
  NAND2_X1 U6353 ( .A1(n5964), .A2(n5963), .ZN(n10016) );
  NAND2_X2 U6354 ( .A1(n7066), .A2(n9991), .ZN(n9791) );
  AND2_X1 U6355 ( .A1(n8470), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4456) );
  AND2_X1 U6356 ( .A1(n4688), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4457) );
  XNOR2_X1 U6357 ( .A(n6231), .B(n4978), .ZN(n7317) );
  OR2_X1 U6358 ( .A1(n9474), .A2(n9475), .ZN(n4458) );
  OR2_X1 U6359 ( .A1(n10154), .A2(n10220), .ZN(n4459) );
  AND2_X1 U6360 ( .A1(n6291), .A2(n5183), .ZN(n4460) );
  INV_X1 U6361 ( .A(n8883), .ZN(n5156) );
  NAND2_X1 U6362 ( .A1(n4719), .A2(n4718), .ZN(n8962) );
  AND2_X1 U6363 ( .A1(n6732), .A2(n6733), .ZN(n4461) );
  NAND2_X1 U6364 ( .A1(n5189), .A2(n5187), .ZN(n9710) );
  AND2_X1 U6365 ( .A1(n8321), .A2(n5309), .ZN(n4462) );
  NAND2_X1 U6366 ( .A1(n9441), .A2(n8033), .ZN(n4463) );
  NAND2_X1 U6367 ( .A1(n5196), .A2(n5195), .ZN(n7850) );
  NAND2_X1 U6368 ( .A1(n5999), .A2(n5998), .ZN(n9347) );
  NOR2_X1 U6369 ( .A1(n8101), .A2(n9419), .ZN(n4464) );
  NAND2_X1 U6370 ( .A1(n6832), .A2(n8881), .ZN(n4465) );
  NAND2_X1 U6371 ( .A1(n5692), .A2(SI_12_), .ZN(n4466) );
  AND2_X1 U6372 ( .A1(n5149), .A2(n6833), .ZN(n4467) );
  OR2_X1 U6373 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4469) );
  INV_X1 U6374 ( .A(n5239), .ZN(n5235) );
  NAND2_X1 U6375 ( .A1(n7526), .A2(n10455), .ZN(n5239) );
  AND2_X1 U6376 ( .A1(n4751), .A2(n4978), .ZN(n4470) );
  AND3_X1 U6377 ( .A1(n5560), .A2(n5559), .A3(n5558), .ZN(n4471) );
  AOI21_X1 U6378 ( .B1(n9308), .B2(n6472), .A(n5406), .ZN(n6744) );
  XNOR2_X1 U6379 ( .A(n10016), .B(n9816), .ZN(n10012) );
  INV_X1 U6380 ( .A(n10012), .ZN(n5377) );
  XNOR2_X1 U6381 ( .A(n9562), .B(n9561), .ZN(n9688) );
  NAND2_X1 U6382 ( .A1(n9625), .A2(n5190), .ZN(n10092) );
  OR2_X1 U6383 ( .A1(n6081), .A2(n6954), .ZN(n4472) );
  NAND2_X1 U6384 ( .A1(n5798), .A2(n5797), .ZN(n10085) );
  AND2_X1 U6385 ( .A1(n6442), .A2(n8940), .ZN(n4473) );
  NAND2_X1 U6386 ( .A1(n4742), .A2(n6636), .ZN(n8902) );
  AOI21_X1 U6387 ( .B1(n5357), .B2(n5803), .A(n5356), .ZN(n5355) );
  INV_X1 U6388 ( .A(n5355), .ZN(n4970) );
  NAND2_X1 U6389 ( .A1(n5832), .A2(n5831), .ZN(n10197) );
  INV_X1 U6390 ( .A(n10197), .ZN(n5393) );
  NAND2_X1 U6391 ( .A1(n4937), .A2(n4938), .ZN(n10057) );
  AND2_X1 U6392 ( .A1(n6634), .A2(n5264), .ZN(n4474) );
  INV_X1 U6393 ( .A(n6239), .ZN(n6245) );
  AND2_X1 U6394 ( .A1(n5147), .A2(n4465), .ZN(n4475) );
  XNOR2_X1 U6395 ( .A(n6322), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7574) );
  AND2_X1 U6396 ( .A1(n10197), .A2(n9821), .ZN(n4476) );
  INV_X1 U6397 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6161) );
  INV_X1 U6398 ( .A(n7570), .ZN(n7557) );
  XNOR2_X1 U6399 ( .A(n6305), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7570) );
  INV_X1 U6400 ( .A(n8367), .ZN(n8360) );
  XNOR2_X1 U6401 ( .A(n6351), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8367) );
  AND3_X1 U6402 ( .A1(n6576), .A2(n6886), .A3(n6844), .ZN(n4477) );
  AND2_X1 U6403 ( .A1(n6574), .A2(n5136), .ZN(n4478) );
  AND3_X1 U6404 ( .A1(n7979), .A2(n8320), .A3(n7973), .ZN(n4479) );
  AND2_X1 U6405 ( .A1(n5355), .A2(n5353), .ZN(n4480) );
  OR2_X1 U6406 ( .A1(n9155), .A2(n8291), .ZN(n6621) );
  AND2_X1 U6407 ( .A1(n9703), .A2(n9792), .ZN(n4481) );
  OR2_X1 U6408 ( .A1(n10194), .A2(n9820), .ZN(n4482) );
  NOR2_X1 U6409 ( .A1(n7274), .A2(n7494), .ZN(n4483) );
  OR2_X1 U6410 ( .A1(n9076), .A2(n9063), .ZN(n4484) );
  NAND2_X1 U6411 ( .A1(n6140), .A2(n6182), .ZN(n6667) );
  NOR2_X1 U6412 ( .A1(n10206), .A2(n9822), .ZN(n4485) );
  OR2_X1 U6413 ( .A1(n9562), .A2(n9819), .ZN(n4486) );
  AND2_X1 U6414 ( .A1(n10225), .A2(n9826), .ZN(n4487) );
  NOR2_X1 U6415 ( .A1(n9358), .A2(n5048), .ZN(n4488) );
  AND2_X1 U6416 ( .A1(n9260), .A2(n8991), .ZN(n4489) );
  AND2_X1 U6417 ( .A1(n6637), .A2(n6483), .ZN(n4490) );
  OR2_X1 U6418 ( .A1(n6870), .A2(n7976), .ZN(n6845) );
  INV_X1 U6419 ( .A(n6845), .ZN(n4830) );
  AND2_X1 U6420 ( .A1(n5366), .A2(n4630), .ZN(n4491) );
  OR2_X1 U6421 ( .A1(n9245), .A2(n6733), .ZN(n4492) );
  AND2_X1 U6422 ( .A1(n9617), .A2(n9792), .ZN(n4493) );
  AND2_X1 U6423 ( .A1(n4767), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4494) );
  XNOR2_X1 U6424 ( .A(n5691), .B(SI_12_), .ZN(n5690) );
  AND2_X1 U6425 ( .A1(n7069), .A2(n7071), .ZN(n4495) );
  OR2_X1 U6426 ( .A1(n7920), .A2(n9536), .ZN(n9655) );
  INV_X1 U6427 ( .A(n8033), .ZN(n5047) );
  INV_X1 U6428 ( .A(n5724), .ZN(n5725) );
  XNOR2_X1 U6429 ( .A(n5727), .B(SI_14_), .ZN(n5724) );
  AND2_X1 U6430 ( .A1(n5044), .A2(n8048), .ZN(n4496) );
  AND2_X1 U6431 ( .A1(n10194), .A2(n9820), .ZN(n4497) );
  NAND2_X1 U6432 ( .A1(n9497), .A2(n9503), .ZN(n4498) );
  AND2_X1 U6433 ( .A1(n4762), .A2(n4761), .ZN(n4499) );
  AND2_X1 U6434 ( .A1(n9595), .A2(n9594), .ZN(n9751) );
  AND2_X1 U6435 ( .A1(n6603), .A2(n6601), .ZN(n4500) );
  NAND2_X1 U6436 ( .A1(n10206), .A2(n6070), .ZN(n9771) );
  INV_X1 U6437 ( .A(n9771), .ZN(n5188) );
  AND2_X1 U6438 ( .A1(n5130), .A2(n4697), .ZN(n4501) );
  NAND2_X1 U6439 ( .A1(n5740), .A2(SI_15_), .ZN(n4502) );
  NAND2_X1 U6440 ( .A1(n5895), .A2(n5894), .ZN(n10188) );
  INV_X1 U6441 ( .A(n10188), .ZN(n10042) );
  NAND2_X1 U6442 ( .A1(n9638), .A2(n9634), .ZN(n5127) );
  AND2_X1 U6443 ( .A1(n6660), .A2(n8794), .ZN(n4503) );
  OR2_X1 U6444 ( .A1(n7570), .A2(n7440), .ZN(n4504) );
  AND2_X1 U6445 ( .A1(n8775), .A2(n4994), .ZN(n4505) );
  NAND2_X1 U6446 ( .A1(n5619), .A2(n8689), .ZN(n5635) );
  INV_X1 U6447 ( .A(n5635), .ZN(n5340) );
  NOR2_X1 U6448 ( .A1(n10144), .A2(n8083), .ZN(n4506) );
  NOR2_X1 U6449 ( .A1(n6737), .A2(n8918), .ZN(n4507) );
  INV_X1 U6450 ( .A(n6836), .ZN(n5148) );
  NAND2_X1 U6451 ( .A1(n8236), .A2(n8314), .ZN(n6836) );
  AND2_X1 U6452 ( .A1(n5586), .A2(SI_6_), .ZN(n4508) );
  INV_X1 U6453 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5573) );
  AND2_X1 U6454 ( .A1(n8850), .A2(n6637), .ZN(n4509) );
  OR2_X1 U6455 ( .A1(n6074), .A2(n8122), .ZN(n9705) );
  INV_X1 U6456 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8572) );
  INV_X1 U6457 ( .A(n6626), .ZN(n4737) );
  INV_X1 U6458 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6012) );
  NAND2_X1 U6459 ( .A1(n6287), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4510) );
  INV_X1 U6460 ( .A(n5254), .ZN(n5253) );
  OAI21_X1 U6461 ( .B1(n9996), .B2(n5255), .A(n5992), .ZN(n5254) );
  NAND2_X1 U6462 ( .A1(n7412), .A2(n6813), .ZN(n4511) );
  NAND2_X1 U6463 ( .A1(n10176), .A2(n5411), .ZN(n4512) );
  AND2_X1 U6464 ( .A1(n5423), .A2(n5517), .ZN(n4513) );
  NAND2_X1 U6465 ( .A1(n8046), .A2(n9328), .ZN(n4514) );
  AND2_X1 U6466 ( .A1(n4598), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4515) );
  AND2_X1 U6467 ( .A1(n5362), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n4516) );
  AND2_X1 U6468 ( .A1(n5673), .A2(n5659), .ZN(n4517) );
  INV_X1 U6469 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6024) );
  OR2_X1 U6470 ( .A1(n5536), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n4518) );
  NOR2_X1 U6471 ( .A1(n8009), .A2(n8008), .ZN(n9426) );
  AND2_X1 U6472 ( .A1(n6707), .A2(n7595), .ZN(n4519) );
  AND2_X1 U6473 ( .A1(n5031), .A2(n4490), .ZN(n4520) );
  AND2_X1 U6474 ( .A1(n9711), .A2(n9638), .ZN(n4521) );
  NAND2_X1 U6475 ( .A1(n5633), .A2(n4466), .ZN(n4522) );
  NAND2_X1 U6476 ( .A1(n4446), .A2(n4473), .ZN(n4523) );
  NOR2_X1 U6477 ( .A1(n6753), .A2(n8307), .ZN(n4525) );
  AND2_X1 U6478 ( .A1(n6361), .A2(n6612), .ZN(n7593) );
  INV_X1 U6479 ( .A(n7593), .ZN(n5286) );
  AND2_X1 U6480 ( .A1(n8107), .A2(n8106), .ZN(n4526) );
  NAND2_X1 U6481 ( .A1(n9698), .A2(n9726), .ZN(n7890) );
  NAND2_X1 U6482 ( .A1(n10099), .A2(n9624), .ZN(n10123) );
  OR2_X1 U6483 ( .A1(n10220), .A2(n8083), .ZN(n9617) );
  INV_X1 U6484 ( .A(n5370), .ZN(n5369) );
  NAND2_X1 U6485 ( .A1(n5728), .A2(n4502), .ZN(n5370) );
  AND2_X1 U6486 ( .A1(n4619), .A2(n9386), .ZN(n4527) );
  AND2_X1 U6487 ( .A1(n5094), .A2(n5092), .ZN(n4528) );
  AND2_X1 U6488 ( .A1(n5937), .A2(n5936), .ZN(n9406) );
  AND2_X1 U6489 ( .A1(n4698), .A2(n5510), .ZN(n4529) );
  AND2_X1 U6490 ( .A1(n9204), .A2(n8858), .ZN(n4530) );
  AND2_X1 U6491 ( .A1(n4758), .A2(n4757), .ZN(n7560) );
  OR2_X1 U6492 ( .A1(n5220), .A2(n4487), .ZN(n4531) );
  INV_X1 U6493 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6494 ( .A1(n6835), .A2(n4465), .ZN(n4532) );
  OR2_X1 U6495 ( .A1(n7286), .A2(n7285), .ZN(n4533) );
  NOR2_X1 U6496 ( .A1(n8306), .A2(n6753), .ZN(n4534) );
  OR2_X1 U6497 ( .A1(n9622), .A2(n9791), .ZN(n4535) );
  OR2_X1 U6498 ( .A1(n9577), .A2(n9791), .ZN(n4536) );
  NAND2_X1 U6499 ( .A1(n4460), .A2(n6289), .ZN(n8338) );
  INV_X1 U6500 ( .A(n8338), .ZN(n4812) );
  AND2_X1 U6501 ( .A1(n9790), .A2(n4639), .ZN(n4537) );
  AND2_X1 U6502 ( .A1(n9033), .A2(n6817), .ZN(n4538) );
  NAND2_X1 U6503 ( .A1(n6822), .A2(n6823), .ZN(n4539) );
  AND2_X1 U6504 ( .A1(n5400), .A2(n4501), .ZN(n4540) );
  OR2_X1 U6505 ( .A1(n6837), .A2(n6838), .ZN(n4541) );
  INV_X1 U6506 ( .A(n9641), .ZN(n5119) );
  NAND2_X1 U6507 ( .A1(n7183), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4542) );
  AND2_X1 U6508 ( .A1(n4766), .A2(n8344), .ZN(n4543) );
  AND2_X1 U6509 ( .A1(n9276), .A2(n9046), .ZN(n4544) );
  AND2_X1 U6510 ( .A1(n9685), .A2(n9758), .ZN(n4545) );
  INV_X1 U6511 ( .A(n9714), .ZN(n5381) );
  NOR2_X1 U6512 ( .A1(n9192), .A2(n8834), .ZN(n4546) );
  AND2_X1 U6513 ( .A1(n9594), .A2(n9597), .ZN(n10347) );
  INV_X1 U6514 ( .A(n10347), .ZN(n5224) );
  AND2_X1 U6515 ( .A1(n4815), .A2(n4814), .ZN(n4547) );
  OR2_X1 U6516 ( .A1(n8198), .A2(n7685), .ZN(n6615) );
  AND2_X1 U6517 ( .A1(n4598), .A2(n5325), .ZN(n4548) );
  INV_X1 U6518 ( .A(n4973), .ZN(n4972) );
  NAND2_X1 U6519 ( .A1(n5357), .A2(n4974), .ZN(n4973) );
  INV_X1 U6520 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5444) );
  OR2_X1 U6521 ( .A1(n5416), .A2(n5347), .ZN(n4549) );
  INV_X1 U6522 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4978) );
  INV_X1 U6523 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5325) );
  INV_X1 U6524 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U6525 ( .A1(n5146), .A2(n6836), .ZN(n4550) );
  NAND2_X1 U6526 ( .A1(n4710), .A2(n4484), .ZN(n4709) );
  NOR2_X1 U6527 ( .A1(n7756), .A2(n8344), .ZN(n8351) );
  NAND2_X1 U6528 ( .A1(n4621), .A2(n5044), .ZN(n9385) );
  NAND2_X1 U6529 ( .A1(n4923), .A2(n7869), .ZN(n6754) );
  NAND2_X1 U6530 ( .A1(n9463), .A2(n9464), .ZN(n9313) );
  AND2_X1 U6531 ( .A1(n5925), .A2(n5923), .ZN(n4551) );
  NOR2_X1 U6532 ( .A1(n7822), .A2(n5388), .ZN(n7853) );
  NAND2_X1 U6533 ( .A1(n4709), .A2(n6817), .ZN(n9037) );
  OR3_X1 U6534 ( .A1(n7087), .A2(n9735), .A3(n6090), .ZN(n9559) );
  OR2_X1 U6535 ( .A1(n7822), .A2(n10240), .ZN(n4552) );
  INV_X1 U6536 ( .A(n6639), .ZN(n5154) );
  OR2_X1 U6537 ( .A1(n8408), .A2(n8407), .ZN(n4885) );
  OAI21_X1 U6538 ( .B1(n6627), .B2(n4738), .A(n4735), .ZN(n8951) );
  AND2_X1 U6539 ( .A1(n5228), .A2(n5226), .ZN(n7767) );
  NAND2_X1 U6540 ( .A1(n6627), .A2(n6626), .ZN(n8966) );
  NAND2_X1 U6541 ( .A1(n4720), .A2(n6823), .ZN(n8973) );
  NAND2_X1 U6542 ( .A1(n5231), .A2(n5232), .ZN(n7786) );
  AND2_X1 U6543 ( .A1(n8424), .A2(n8423), .ZN(n4553) );
  AND2_X1 U6544 ( .A1(n5103), .A2(n5101), .ZN(n4554) );
  INV_X1 U6545 ( .A(n8226), .ZN(n5312) );
  AND2_X1 U6546 ( .A1(n6729), .A2(n8327), .ZN(n4555) );
  OR2_X1 U6547 ( .A1(n10175), .A2(n9545), .ZN(n4556) );
  NAND2_X1 U6548 ( .A1(n6506), .A2(n6505), .ZN(n8857) );
  INV_X1 U6549 ( .A(n8857), .ZN(n8881) );
  INV_X1 U6550 ( .A(n7317), .ZN(n4679) );
  AND2_X1 U6551 ( .A1(n9192), .A2(n9159), .ZN(n4557) );
  AND2_X1 U6552 ( .A1(n4554), .A2(n4457), .ZN(n4558) );
  AND2_X1 U6553 ( .A1(n7392), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4559) );
  AND2_X1 U6554 ( .A1(n9699), .A2(n9628), .ZN(n6072) );
  INV_X1 U6555 ( .A(n6072), .ZN(n5011) );
  AND2_X1 U6556 ( .A1(n7005), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4560) );
  OR2_X1 U6557 ( .A1(n5772), .A2(n5771), .ZN(n4561) );
  AND2_X1 U6558 ( .A1(n8400), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4562) );
  INV_X1 U6559 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4751) );
  NOR2_X1 U6560 ( .A1(n5101), .A2(n5098), .ZN(n4563) );
  OR2_X1 U6561 ( .A1(n5100), .A2(n5098), .ZN(n4564) );
  OR2_X1 U6562 ( .A1(n7822), .A2(n5389), .ZN(n4565) );
  NAND2_X1 U6563 ( .A1(n6632), .A2(n6631), .ZN(n8936) );
  INV_X1 U6564 ( .A(n8351), .ZN(n5301) );
  AND2_X1 U6565 ( .A1(n5073), .A2(n5072), .ZN(n4566) );
  INV_X1 U6566 ( .A(n5415), .ZN(n5243) );
  NAND2_X1 U6567 ( .A1(n5484), .A2(n5483), .ZN(n7637) );
  AND2_X2 U6568 ( .A1(n6096), .A2(n7606), .ZN(n10494) );
  INV_X1 U6569 ( .A(n10240), .ZN(n5390) );
  AND2_X1 U6570 ( .A1(n6313), .A2(n6350), .ZN(n8344) );
  INV_X1 U6571 ( .A(n8344), .ZN(n5079) );
  NAND2_X2 U6572 ( .A1(n6848), .A2(n6847), .ZN(n9061) );
  INV_X1 U6573 ( .A(n9018), .ZN(n4842) );
  AND2_X1 U6574 ( .A1(n9942), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4567) );
  OR3_X1 U6575 ( .A1(n6887), .A2(n6680), .A3(n6943), .ZN(n7170) );
  INV_X1 U6576 ( .A(n7170), .ZN(n4589) );
  OR2_X1 U6577 ( .A1(n10482), .A2(n4788), .ZN(n4568) );
  INV_X1 U6578 ( .A(n7638), .ZN(n4797) );
  NAND2_X1 U6579 ( .A1(n6852), .A2(n7336), .ZN(n9069) );
  INV_X1 U6580 ( .A(n9069), .ZN(n4725) );
  INV_X1 U6581 ( .A(n4991), .ZN(n4990) );
  INV_X1 U6582 ( .A(n4993), .ZN(n4992) );
  NOR2_X1 U6583 ( .A1(n8488), .A2(n8487), .ZN(n4993) );
  NAND2_X1 U6584 ( .A1(n6053), .A2(n9567), .ZN(n10386) );
  NAND2_X1 U6585 ( .A1(n6245), .A2(n7344), .ZN(n7955) );
  OR2_X1 U6586 ( .A1(n8489), .A2(n4982), .ZN(n4569) );
  NAND2_X1 U6587 ( .A1(n6777), .A2(n6776), .ZN(n8320) );
  INV_X1 U6588 ( .A(n8320), .ZN(n8318) );
  AND2_X1 U6589 ( .A1(n8487), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4570) );
  AND2_X1 U6590 ( .A1(n4991), .A2(n4980), .ZN(n4571) );
  AND2_X1 U6591 ( .A1(n5076), .A2(n5075), .ZN(n4572) );
  INV_X1 U6592 ( .A(n5222), .ZN(n5220) );
  NAND2_X1 U6593 ( .A1(n10230), .A2(n9827), .ZN(n5222) );
  INV_X1 U6594 ( .A(n8767), .ZN(n4879) );
  XNOR2_X1 U6595 ( .A(n6344), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7573) );
  INV_X1 U6596 ( .A(n7573), .ZN(n4757) );
  INV_X1 U6597 ( .A(n7861), .ZN(n5135) );
  INV_X1 U6598 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5098) );
  AND2_X1 U6599 ( .A1(n5814), .A2(n6016), .ZN(n9991) );
  AND2_X1 U6600 ( .A1(n4759), .A2(n5300), .ZN(n4573) );
  INV_X1 U6601 ( .A(n8760), .ZN(n5296) );
  AND2_X1 U6602 ( .A1(n4676), .A2(n4444), .ZN(n4574) );
  INV_X1 U6603 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4922) );
  INV_X1 U6604 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n4783) );
  XNOR2_X1 U6605 ( .A(n4680), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10506) );
  INV_X1 U6606 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n4682) );
  NAND3_X1 U6607 ( .A1(n4579), .A2(n4578), .A3(n4477), .ZN(n4586) );
  OAI21_X1 U6608 ( .B1(n4582), .B2(n4581), .A(n4509), .ZN(n4875) );
  NAND2_X1 U6609 ( .A1(n4590), .A2(n4808), .ZN(n5182) );
  NAND2_X1 U6610 ( .A1(n4591), .A2(n6592), .ZN(n4590) );
  NAND2_X1 U6611 ( .A1(n4592), .A2(n4595), .ZN(n4591) );
  INV_X1 U6612 ( .A(n4593), .ZN(n4592) );
  OAI21_X1 U6613 ( .B1(n6375), .B2(n4594), .A(n9018), .ZN(n4593) );
  NOR2_X1 U6614 ( .A1(n6373), .A2(n6608), .ZN(n4594) );
  NAND3_X1 U6615 ( .A1(n6374), .A2(n6607), .A3(n4596), .ZN(n4595) );
  INV_X1 U6616 ( .A(n6375), .ZN(n4596) );
  NAND2_X1 U6617 ( .A1(n4606), .A2(n4605), .ZN(n5326) );
  INV_X1 U6618 ( .A(n7124), .ZN(n4606) );
  NAND2_X1 U6619 ( .A1(n7121), .A2(n7120), .ZN(n4607) );
  INV_X2 U6620 ( .A(n7205), .ZN(n7072) );
  NAND3_X4 U6621 ( .A1(n4614), .A2(n7205), .A3(n7068), .ZN(n9345) );
  OR2_X2 U6622 ( .A1(n7063), .A2(n4613), .ZN(n7068) );
  INV_X1 U6623 ( .A(n9498), .ZN(n4615) );
  NAND2_X1 U6624 ( .A1(n4615), .A2(n4445), .ZN(n4618) );
  NAND2_X1 U6625 ( .A1(n9455), .A2(n9453), .ZN(n8114) );
  NAND3_X1 U6626 ( .A1(n5044), .A2(n5045), .A3(n8048), .ZN(n4619) );
  NAND2_X2 U6627 ( .A1(n9384), .A2(n8058), .ZN(n9463) );
  NAND2_X1 U6628 ( .A1(n7070), .A2(n4495), .ZN(n7111) );
  NAND2_X1 U6629 ( .A1(n4624), .A2(n8141), .ZN(n7075) );
  NAND2_X1 U6630 ( .A1(n4625), .A2(n5564), .ZN(n5550) );
  NAND3_X1 U6631 ( .A1(n5564), .A2(n4625), .A3(n5585), .ZN(n5017) );
  XNOR2_X1 U6632 ( .A(n5564), .B(n4625), .ZN(n6893) );
  INV_X1 U6633 ( .A(n5711), .ZN(n4626) );
  NAND2_X1 U6634 ( .A1(n4626), .A2(n5366), .ZN(n4629) );
  OR2_X2 U6635 ( .A1(n9789), .A2(n7066), .ZN(n4631) );
  AND2_X2 U6636 ( .A1(n4636), .A2(n4632), .ZN(n9789) );
  NAND2_X1 U6637 ( .A1(n9668), .A2(n9730), .ZN(n4635) );
  NAND2_X1 U6638 ( .A1(n4638), .A2(n4637), .ZN(n4636) );
  NOR2_X1 U6639 ( .A1(n9732), .A2(n9728), .ZN(n4637) );
  OAI21_X1 U6640 ( .B1(n9668), .B2(n9730), .A(n4537), .ZN(n4638) );
  NAND2_X1 U6641 ( .A1(n4640), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U6642 ( .A1(n4643), .A2(n9600), .ZN(n4641) );
  NAND2_X1 U6643 ( .A1(n4649), .A2(n4643), .ZN(n4642) );
  NAND2_X1 U6644 ( .A1(n4647), .A2(n4645), .ZN(n4644) );
  NAND2_X1 U6645 ( .A1(n9753), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U6646 ( .A1(n4649), .A2(n5105), .ZN(n4648) );
  INV_X1 U6647 ( .A(n9599), .ZN(n4650) );
  NAND2_X1 U6648 ( .A1(n5636), .A2(n4655), .ZN(n4654) );
  NAND2_X1 U6649 ( .A1(n4659), .A2(n4777), .ZN(n4817) );
  NAND2_X1 U6650 ( .A1(n9631), .A2(n5111), .ZN(n4659) );
  NAND2_X1 U6651 ( .A1(n4661), .A2(n4660), .ZN(n9631) );
  OAI21_X1 U6652 ( .B1(n9612), .B2(n10124), .A(n4493), .ZN(n4661) );
  NAND2_X2 U6653 ( .A1(n5200), .A2(n5199), .ZN(n5331) );
  NOR2_X1 U6654 ( .A1(n7228), .A2(n4662), .ZN(n7190) );
  NOR2_X1 U6655 ( .A1(n4664), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U6656 ( .A1(n5084), .A2(n5083), .ZN(n4664) );
  NAND2_X1 U6657 ( .A1(n4666), .A2(n10499), .ZN(n8803) );
  XNOR2_X1 U6658 ( .A(n4667), .B(n4673), .ZN(n4666) );
  INV_X1 U6659 ( .A(n4669), .ZN(n4668) );
  INV_X1 U6660 ( .A(n8802), .ZN(n4673) );
  NAND3_X1 U6661 ( .A1(n4679), .A2(n4444), .A3(n7173), .ZN(n4678) );
  XNOR2_X1 U6662 ( .A(n7176), .B(n5298), .ZN(n10497) );
  AND2_X1 U6663 ( .A1(n4681), .A2(n4542), .ZN(n7176) );
  NAND2_X1 U6664 ( .A1(n7214), .A2(n7215), .ZN(n4681) );
  NAND2_X1 U6665 ( .A1(n7552), .A2(n7551), .ZN(n4686) );
  NAND2_X1 U6666 ( .A1(n5085), .A2(n4688), .ZN(n4687) );
  INV_X1 U6667 ( .A(n8480), .ZN(n4688) );
  INV_X1 U6668 ( .A(n5085), .ZN(n4690) );
  OAI211_X1 U6669 ( .C1(n4751), .C2(n4693), .A(n4692), .B(P2_IR_REG_2__SCAN_IN), .ZN(n4870) );
  INV_X1 U6670 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4693) );
  INV_X1 U6671 ( .A(n10322), .ZN(n5433) );
  INV_X1 U6672 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4697) );
  NAND3_X1 U6673 ( .A1(n4513), .A2(n4699), .A3(n5400), .ZN(n5443) );
  NOR2_X1 U6674 ( .A1(n5429), .A2(n5428), .ZN(n4699) );
  AOI21_X2 U6675 ( .B1(n10115), .B2(n5783), .A(n5782), .ZN(n10098) );
  OAI22_X2 U6676 ( .A1(n10022), .A2(n5245), .B1(n5254), .B2(n4450), .ZN(n5244)
         );
  NAND2_X2 U6677 ( .A1(n4955), .A2(n5904), .ZN(n10022) );
  NAND2_X1 U6678 ( .A1(n4771), .A2(n6814), .ZN(n7425) );
  INV_X2 U6679 ( .A(n4704), .ZN(n4855) );
  NAND2_X2 U6680 ( .A1(n6260), .A2(n6600), .ZN(n4704) );
  AND2_X1 U6681 ( .A1(n4855), .A2(n4701), .ZN(n6258) );
  NAND2_X1 U6682 ( .A1(n7348), .A2(n4702), .ZN(n7961) );
  NAND2_X1 U6683 ( .A1(n4703), .A2(n4855), .ZN(n4702) );
  INV_X1 U6684 ( .A(n7957), .ZN(n4703) );
  NAND2_X1 U6685 ( .A1(n4704), .A2(n7957), .ZN(n7348) );
  NOR2_X1 U6686 ( .A1(n7412), .A2(n4704), .ZN(n6585) );
  NOR2_X1 U6687 ( .A1(n4855), .A2(n6599), .ZN(n4705) );
  NAND3_X1 U6688 ( .A1(n4708), .A2(n4709), .A3(n4707), .ZN(n4706) );
  INV_X1 U6689 ( .A(n7654), .ZN(n4710) );
  NAND2_X1 U6690 ( .A1(n4711), .A2(n6819), .ZN(n9023) );
  NAND2_X1 U6691 ( .A1(n4745), .A2(n4712), .ZN(n4713) );
  AND2_X2 U6692 ( .A1(n5277), .A2(n4724), .ZN(n6182) );
  NAND2_X2 U6693 ( .A1(n5285), .A2(n5283), .ZN(n7597) );
  NAND2_X1 U6694 ( .A1(n4731), .A2(n6652), .ZN(n6849) );
  NOR2_X1 U6695 ( .A1(n5414), .A2(n4729), .ZN(n4727) );
  NAND2_X1 U6696 ( .A1(n5414), .A2(n4729), .ZN(n4728) );
  INV_X1 U6697 ( .A(n6652), .ZN(n4729) );
  NAND2_X1 U6698 ( .A1(n4732), .A2(n4733), .ZN(n6632) );
  NAND2_X1 U6699 ( .A1(n4739), .A2(n4740), .ZN(n8891) );
  AND2_X2 U6700 ( .A1(n6182), .A2(n4548), .ZN(n4745) );
  AND3_X2 U6701 ( .A1(n5139), .A2(n5140), .A3(n6136), .ZN(n6140) );
  NAND3_X1 U6702 ( .A1(n5274), .A2(n4748), .A3(n4747), .ZN(n6624) );
  NAND3_X1 U6703 ( .A1(n4840), .A2(n6621), .A3(n6618), .ZN(n4747) );
  NAND3_X1 U6704 ( .A1(n4751), .A2(n4978), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7181) );
  NAND2_X1 U6705 ( .A1(n5288), .A2(n4753), .ZN(n8484) );
  NAND2_X1 U6706 ( .A1(n7234), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7275) );
  NAND2_X1 U6707 ( .A1(n5299), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U6708 ( .A1(n4763), .A2(n4453), .ZN(n8409) );
  NAND3_X1 U6709 ( .A1(n4765), .A2(n4764), .A3(n4543), .ZN(n5303) );
  INV_X1 U6710 ( .A(n7562), .ZN(n4767) );
  NAND2_X1 U6711 ( .A1(n5291), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5290) );
  OAI21_X1 U6712 ( .B1(n5302), .B2(n8351), .A(n8349), .ZN(n8369) );
  OAI22_X2 U6713 ( .A1(n9004), .A2(n6821), .B1(n8291), .B2(n8224), .ZN(n8989)
         );
  AOI21_X1 U6714 ( .B1(n8825), .B2(n6840), .A(n4546), .ZN(n8816) );
  NAND2_X1 U6715 ( .A1(n4812), .A2(n6808), .ZN(n6810) );
  AND2_X1 U6716 ( .A1(n5187), .A2(n6072), .ZN(n5010) );
  NAND2_X2 U6717 ( .A1(n7352), .A2(n7963), .ZN(n6600) );
  INV_X1 U6718 ( .A(n6806), .ZN(n7365) );
  NAND2_X1 U6719 ( .A1(n4769), .A2(n6858), .ZN(n4774) );
  NAND2_X1 U6720 ( .A1(n4770), .A2(n9061), .ZN(n6858) );
  XNOR2_X1 U6721 ( .A(n6846), .B(n5414), .ZN(n4770) );
  INV_X1 U6722 ( .A(n9299), .ZN(n6164) );
  NAND2_X1 U6723 ( .A1(n7363), .A2(n6811), .ZN(n4771) );
  NAND2_X1 U6724 ( .A1(n8816), .A2(n6841), .ZN(n6843) );
  XNOR2_X2 U6725 ( .A(n6162), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9299) );
  NAND2_X1 U6726 ( .A1(n4855), .A2(n6599), .ZN(n7953) );
  NAND2_X1 U6727 ( .A1(n6911), .A2(n6553), .ZN(n6233) );
  INV_X2 U6728 ( .A(n4772), .ZN(n10414) );
  NAND2_X1 U6729 ( .A1(n5459), .A2(n5458), .ZN(n6051) );
  NAND2_X1 U6730 ( .A1(n9674), .A2(n7718), .ZN(n7720) );
  INV_X1 U6731 ( .A(n4872), .ZN(n4871) );
  INV_X1 U6732 ( .A(n7711), .ZN(n9674) );
  NAND2_X1 U6733 ( .A1(n4773), .A2(n9621), .ZN(n10133) );
  OAI21_X1 U6734 ( .B1(n7818), .B2(n5019), .A(n4866), .ZN(n4773) );
  INV_X1 U6735 ( .A(n6804), .ZN(n7350) );
  NAND2_X1 U6736 ( .A1(n4774), .A2(n6869), .ZN(n6871) );
  NAND2_X1 U6737 ( .A1(n4775), .A2(n5401), .ZN(n6884) );
  NAND2_X1 U6738 ( .A1(n4890), .A2(n6858), .ZN(n4775) );
  NAND2_X1 U6739 ( .A1(n8339), .A2(n5142), .ZN(n5141) );
  INV_X4 U6740 ( .A(n4429), .ZN(n6535) );
  NAND2_X1 U6741 ( .A1(n4870), .A2(n4869), .ZN(n6253) );
  XNOR2_X1 U6743 ( .A(n7080), .B(n8141), .ZN(n7081) );
  NAND2_X1 U6744 ( .A1(n7198), .A2(n5458), .ZN(n7079) );
  NAND2_X1 U6745 ( .A1(n7288), .A2(n7287), .ZN(n5035) );
  AND3_X2 U6746 ( .A1(n6232), .A2(n6233), .A3(n6234), .ZN(n7963) );
  NAND2_X1 U6747 ( .A1(n6831), .A2(n8866), .ZN(n6834) );
  NAND2_X1 U6748 ( .A1(n7591), .A2(n6816), .ZN(n7654) );
  MUX2_X2 U6749 ( .A(n6368), .B(n6367), .S(n6886), .Z(n6375) );
  OAI21_X1 U6750 ( .B1(n9615), .B2(n9609), .A(n4545), .ZN(n9611) );
  NAND2_X1 U6751 ( .A1(n8388), .A2(n4779), .ZN(n8372) );
  NAND2_X1 U6752 ( .A1(n8371), .A2(n8370), .ZN(n8388) );
  XNOR2_X1 U6753 ( .A(n4780), .B(n8753), .ZN(P2_U3199) );
  NAND2_X1 U6754 ( .A1(n4873), .A2(n4871), .ZN(n4780) );
  NOR2_X1 U6755 ( .A1(n8372), .A2(n9026), .ZN(n8389) );
  NAND2_X1 U6756 ( .A1(n4915), .A2(n4913), .ZN(n8217) );
  NAND2_X1 U6757 ( .A1(n8266), .A2(n6723), .ZN(n8180) );
  INV_X1 U6758 ( .A(n6419), .ZN(n6108) );
  INV_X1 U6759 ( .A(n6421), .ZN(n6110) );
  INV_X1 U6760 ( .A(n9578), .ZN(n5109) );
  NOR2_X1 U6761 ( .A1(n6565), .A2(n5024), .ZN(n6566) );
  NAND2_X1 U6762 ( .A1(n6097), .A2(n10494), .ZN(n6098) );
  OAI21_X1 U6763 ( .B1(n9615), .B2(n9614), .A(n4781), .ZN(n9618) );
  NAND2_X1 U6764 ( .A1(n5189), .A2(n5010), .ZN(n10071) );
  NAND2_X1 U6765 ( .A1(n5185), .A2(n9594), .ZN(n7768) );
  NAND2_X1 U6766 ( .A1(n7819), .A2(n9589), .ZN(n4787) );
  NAND2_X1 U6767 ( .A1(n10414), .A2(n10253), .ZN(n7715) );
  OAI21_X2 U6768 ( .B1(n7898), .B2(n4792), .A(n7897), .ZN(n7909) );
  INV_X1 U6769 ( .A(n10389), .ZN(n4796) );
  NAND2_X1 U6770 ( .A1(n4891), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5965) );
  AOI21_X1 U6771 ( .B1(n4802), .B2(n9061), .A(n4799), .ZN(n9190) );
  XNOR2_X1 U6772 ( .A(n8825), .B(n8824), .ZN(n4802) );
  NAND2_X1 U6773 ( .A1(n4807), .A2(n4803), .ZN(P2_U3486) );
  OR2_X1 U6774 ( .A1(n9190), .A2(n6883), .ZN(n4807) );
  NAND2_X2 U6775 ( .A1(n6676), .A2(n6677), .ZN(n6244) );
  INV_X1 U6776 ( .A(n6573), .ZN(n5132) );
  OAI21_X1 U6777 ( .B1(n6531), .B2(n8824), .A(n6530), .ZN(n6565) );
  NAND2_X1 U6778 ( .A1(n9188), .A2(n4832), .ZN(P2_U3455) );
  NAND2_X1 U6779 ( .A1(n8821), .A2(n4810), .ZN(P2_U3205) );
  NAND2_X1 U6780 ( .A1(n7244), .A2(n7243), .ZN(n7264) );
  BUF_X4 U6781 ( .A(n6677), .Z(n8770) );
  NAND2_X1 U6782 ( .A1(n7166), .A2(n7165), .ZN(n7240) );
  NAND2_X1 U6783 ( .A1(n7306), .A2(n7319), .ZN(n7305) );
  NAND2_X1 U6784 ( .A1(n4979), .A2(n4992), .ZN(n8769) );
  OAI21_X1 U6785 ( .B1(n8496), .B2(n8781), .A(n8495), .ZN(n4872) );
  NAND2_X1 U6786 ( .A1(n4511), .A2(n6812), .ZN(n6814) );
  AOI21_X2 U6787 ( .B1(n6912), .B2(n5637), .A(n4813), .ZN(n9370) );
  AND2_X1 U6788 ( .A1(n6057), .A2(n9583), .ZN(n9581) );
  NAND2_X1 U6789 ( .A1(n4817), .A2(n4535), .ZN(n4894) );
  INV_X1 U6790 ( .A(n6856), .ZN(n6857) );
  NAND2_X1 U6791 ( .A1(n5129), .A2(n5130), .ZN(n5432) );
  NAND2_X1 U6792 ( .A1(n7767), .A2(n9681), .ZN(n4946) );
  NAND2_X1 U6793 ( .A1(n4936), .A2(n4935), .ZN(n7934) );
  NAND2_X1 U6794 ( .A1(n7840), .A2(n7839), .ZN(n4943) );
  NAND3_X1 U6795 ( .A1(n8930), .A2(n4825), .A3(n8940), .ZN(n4824) );
  OAI21_X1 U6796 ( .B1(n6849), .B2(n4830), .A(n4857), .ZN(n4856) );
  AND2_X1 U6797 ( .A1(n6812), .A2(n7414), .ZN(n6811) );
  AND2_X1 U6798 ( .A1(n6290), .A2(n6288), .ZN(n5183) );
  AOI21_X1 U6799 ( .B1(n5173), .B2(n9061), .A(n5172), .ZN(n9184) );
  NAND2_X1 U6800 ( .A1(n5068), .A2(n4503), .ZN(n4834) );
  NAND2_X1 U6801 ( .A1(n8186), .A2(n8188), .ZN(n8253) );
  NAND2_X1 U6802 ( .A1(n6108), .A2(n6107), .ZN(n6421) );
  NAND2_X1 U6803 ( .A1(n6110), .A2(n6109), .ZN(n6445) );
  NAND2_X1 U6804 ( .A1(n8275), .A2(n8276), .ZN(n4896) );
  NAND2_X1 U6805 ( .A1(n4926), .A2(n4924), .ZN(n8245) );
  AOI21_X2 U6806 ( .B1(n7544), .B2(n6708), .A(n4519), .ZN(n7684) );
  NAND2_X1 U6807 ( .A1(n4920), .A2(n4836), .ZN(n6758) );
  NAND3_X1 U6808 ( .A1(n6944), .A2(n6681), .A3(n6680), .ZN(n4836) );
  NAND2_X2 U6809 ( .A1(n6058), .A2(n9677), .ZN(n10339) );
  OAI21_X1 U6810 ( .B1(n6069), .B2(n5192), .A(n10093), .ZN(n5191) );
  NAND2_X1 U6811 ( .A1(n7659), .A2(n4841), .ZN(n4840) );
  NAND2_X1 U6812 ( .A1(n4875), .A2(n4874), .ZN(n5153) );
  INV_X1 U6813 ( .A(n7768), .ZN(n4854) );
  AOI21_X1 U6814 ( .B1(n8471), .B2(n8470), .A(n4570), .ZN(n5288) );
  NAND2_X1 U6815 ( .A1(n8369), .A2(n8368), .ZN(n8371) );
  NAND2_X1 U6816 ( .A1(n7913), .A2(n4849), .ZN(P1_U3551) );
  NAND2_X1 U6817 ( .A1(n7902), .A2(n4850), .ZN(P1_U3519) );
  NAND2_X1 U6818 ( .A1(n4852), .A2(n8762), .ZN(n8486) );
  NAND2_X1 U6819 ( .A1(n4865), .A2(n4864), .ZN(n4852) );
  NAND2_X1 U6820 ( .A1(n6807), .A2(n6806), .ZN(n7363) );
  NAND2_X1 U6821 ( .A1(n8906), .A2(n5420), .ZN(n8866) );
  NAND2_X2 U6822 ( .A1(n4860), .A2(n5594), .ZN(n5617) );
  NAND2_X1 U6823 ( .A1(n5592), .A2(n5591), .ZN(n4860) );
  NAND2_X1 U6824 ( .A1(n4976), .A2(n4861), .ZN(n5711) );
  NAND2_X1 U6825 ( .A1(n5634), .A2(n4975), .ZN(n4976) );
  NAND4_X1 U6826 ( .A1(n4862), .A2(n5131), .A3(n5134), .A4(n6679), .ZN(
        P2_U3296) );
  NAND2_X1 U6827 ( .A1(n4878), .A2(n7861), .ZN(n4862) );
  NAND2_X4 U6828 ( .A1(n7635), .A2(n7067), .ZN(n8165) );
  INV_X1 U6829 ( .A(n5335), .ZN(n5334) );
  NAND2_X1 U6830 ( .A1(n5017), .A2(n5349), .ZN(n5592) );
  INV_X1 U6831 ( .A(n9350), .ZN(n5050) );
  NAND2_X1 U6832 ( .A1(n8485), .A2(n8761), .ZN(n4865) );
  NOR2_X1 U6833 ( .A1(n7233), .A2(n7269), .ZN(n7272) );
  AND2_X1 U6834 ( .A1(n6063), .A2(n5193), .ZN(n4866) );
  NAND2_X1 U6835 ( .A1(n6051), .A2(n9745), .ZN(n7711) );
  NAND2_X1 U6836 ( .A1(n7925), .A2(n4867), .ZN(P1_U3547) );
  INV_X1 U6837 ( .A(n10054), .ZN(n5200) );
  NAND2_X1 U6838 ( .A1(n8486), .A2(n8763), .ZN(n4873) );
  NAND2_X1 U6839 ( .A1(n5682), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5700) );
  INV_X1 U6840 ( .A(n5127), .ZN(n5126) );
  NAND2_X1 U6841 ( .A1(n4893), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U6842 ( .A1(n5182), .A2(n4539), .ZN(n5020) );
  NOR2_X1 U6843 ( .A1(n5122), .A2(n5119), .ZN(n5118) );
  NOR2_X2 U6844 ( .A1(n5753), .A2(n9414), .ZN(n4876) );
  NAND2_X1 U6845 ( .A1(n4877), .A2(n4963), .ZN(n4961) );
  NAND2_X1 U6846 ( .A1(n4894), .A2(n9641), .ZN(n4877) );
  NAND2_X1 U6847 ( .A1(n5280), .A2(n5278), .ZN(n6646) );
  NAND2_X1 U6848 ( .A1(n6159), .A2(n5158), .ZN(n9292) );
  NAND2_X1 U6849 ( .A1(n6649), .A2(n6648), .ZN(n8831) );
  NAND2_X1 U6850 ( .A1(n8441), .A2(n5103), .ZN(n5088) );
  NAND3_X1 U6851 ( .A1(n4995), .A2(n8780), .A3(n4880), .ZN(P2_U3200) );
  NAND2_X2 U6852 ( .A1(n6353), .A2(n6352), .ZN(n8198) );
  NAND2_X1 U6853 ( .A1(n6834), .A2(n6833), .ZN(n5147) );
  XNOR2_X2 U6854 ( .A(n5504), .B(n5503), .ZN(n9852) );
  NAND2_X1 U6855 ( .A1(n5872), .A2(n5871), .ZN(n5897) );
  AOI211_X2 U6856 ( .C1(n9791), .C2(n9659), .A(n9652), .B(n9660), .ZN(n9658)
         );
  NOR2_X2 U6857 ( .A1(n5914), .A2(n9432), .ZN(n4891) );
  NAND2_X1 U6858 ( .A1(n10071), .A2(n9699), .ZN(n10054) );
  NAND2_X1 U6859 ( .A1(n9743), .A2(n5186), .ZN(n5185) );
  NAND2_X1 U6860 ( .A1(n5133), .A2(n5132), .ZN(n5131) );
  NOR2_X1 U6861 ( .A1(n6105), .A2(n6139), .ZN(n5140) );
  OAI21_X1 U6862 ( .B1(n9580), .B2(n5108), .A(n4547), .ZN(n5107) );
  NAND2_X1 U6863 ( .A1(n7748), .A2(n7747), .ZN(n5082) );
  NAND3_X1 U6864 ( .A1(n4895), .A2(n5110), .A3(n9576), .ZN(n5108) );
  OAI21_X1 U6865 ( .B1(n9651), .B2(n5116), .A(n9662), .ZN(n5115) );
  INV_X1 U6866 ( .A(n6106), .ZN(n5139) );
  NAND2_X1 U6867 ( .A1(n6646), .A2(n6645), .ZN(n8845) );
  NAND2_X1 U6868 ( .A1(n5269), .A2(n5267), .ZN(n8814) );
  INV_X1 U6869 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U6870 ( .A1(n4898), .A2(n8572), .ZN(n6672) );
  INV_X1 U6871 ( .A(n4899), .ZN(n8209) );
  INV_X1 U6872 ( .A(n8189), .ZN(n4909) );
  NAND2_X1 U6873 ( .A1(n4905), .A2(n4910), .ZN(P2_U3169) );
  NAND3_X1 U6874 ( .A1(n4907), .A2(n4906), .A3(n8320), .ZN(n4905) );
  NAND2_X1 U6875 ( .A1(n4909), .A2(n4908), .ZN(n4907) );
  NAND2_X1 U6876 ( .A1(n7682), .A2(n4916), .ZN(n4915) );
  NAND2_X1 U6877 ( .A1(n6681), .A2(n6680), .ZN(n4923) );
  NAND2_X1 U6878 ( .A1(n8323), .A2(n4927), .ZN(n4926) );
  OAI21_X2 U6879 ( .B1(n5617), .B2(n5616), .A(n5615), .ZN(n5634) );
  OAI21_X2 U6880 ( .B1(n7817), .B2(n7816), .A(n4944), .ZN(n7840) );
  OR2_X1 U6881 ( .A1(n10036), .A2(n4950), .ZN(n4947) );
  NAND2_X1 U6882 ( .A1(n4947), .A2(n4948), .ZN(n10011) );
  MUX2_X1 U6883 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6142), .Z(n5471) );
  MUX2_X1 U6884 ( .A(n6992), .B(n5655), .S(n6142), .Z(n5657) );
  MUX2_X1 U6885 ( .A(n6935), .B(n6937), .S(n6142), .Z(n5652) );
  MUX2_X1 U6886 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6142), .Z(n5593) );
  MUX2_X1 U6887 ( .A(n6932), .B(n5618), .S(n4956), .Z(n5619) );
  MUX2_X1 U6888 ( .A(n6914), .B(n5595), .S(n4956), .Z(n5597) );
  MUX2_X1 U6889 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n4956), .Z(n5727) );
  MUX2_X1 U6890 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4956), .Z(n5709) );
  MUX2_X1 U6891 ( .A(n8654), .B(n7329), .S(n4956), .Z(n5759) );
  MUX2_X1 U6892 ( .A(n7476), .B(n7475), .S(n4956), .Z(n5764) );
  MUX2_X1 U6893 ( .A(n8563), .B(n8717), .S(n4956), .Z(n5805) );
  MUX2_X1 U6894 ( .A(n7603), .B(n5787), .S(n4956), .Z(n5800) );
  MUX2_X1 U6895 ( .A(n7831), .B(n5830), .S(n4956), .Z(n5855) );
  MUX2_X1 U6896 ( .A(n5842), .B(n7834), .S(n4956), .Z(n5858) );
  MUX2_X1 U6897 ( .A(n5888), .B(n5893), .S(n4956), .Z(n5890) );
  MUX2_X1 U6898 ( .A(n7837), .B(n8178), .S(n4956), .Z(n5866) );
  MUX2_X1 U6899 ( .A(n8135), .B(n10329), .S(n4956), .Z(n5932) );
  MUX2_X1 U6900 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n4956), .Z(n5907) );
  MUX2_X1 U6901 ( .A(n5958), .B(n10326), .S(n4956), .Z(n5960) );
  MUX2_X1 U6902 ( .A(n5979), .B(n10325), .S(n4956), .Z(n5981) );
  MUX2_X1 U6903 ( .A(n5997), .B(n8006), .S(n4956), .Z(n6117) );
  MUX2_X1 U6904 ( .A(n6120), .B(n10323), .S(n4956), .Z(n6121) );
  NAND2_X1 U6905 ( .A1(n5120), .A2(n9640), .ZN(n4964) );
  NAND2_X1 U6906 ( .A1(n4964), .A2(n9641), .ZN(n4963) );
  NAND2_X1 U6907 ( .A1(n4959), .A2(n5117), .ZN(n5125) );
  NAND2_X1 U6908 ( .A1(n4961), .A2(n4960), .ZN(n4959) );
  NAND2_X1 U6909 ( .A1(n4962), .A2(n5127), .ZN(n4960) );
  AND2_X1 U6910 ( .A1(n4976), .A2(n4977), .ZN(n5708) );
  OR2_X1 U6911 ( .A1(n8490), .A2(n8489), .ZN(n4979) );
  OR2_X1 U6912 ( .A1(n8490), .A2(n4569), .ZN(n4981) );
  NAND2_X1 U6913 ( .A1(n8489), .A2(n4986), .ZN(n4984) );
  NAND2_X1 U6914 ( .A1(n8490), .A2(n4986), .ZN(n4985) );
  NAND2_X1 U6915 ( .A1(n8766), .A2(n8767), .ZN(n4991) );
  OAI211_X1 U6916 ( .C1(n10177), .C2(n10249), .A(n5008), .B(n5007), .ZN(n10257) );
  INV_X1 U6917 ( .A(n5201), .ZN(n10023) );
  OR2_X1 U6918 ( .A1(n6073), .A2(n4521), .ZN(n5013) );
  NAND3_X1 U6920 ( .A1(n10148), .A2(n9756), .A3(n9613), .ZN(n5019) );
  NAND2_X1 U6921 ( .A1(n5034), .A2(n4473), .ZN(n6482) );
  NAND2_X1 U6922 ( .A1(n5034), .A2(n5030), .ZN(n5029) );
  OAI211_X2 U6923 ( .C1(n5334), .C2(n7293), .A(n5332), .B(n7523), .ZN(n7536)
         );
  NAND2_X1 U6924 ( .A1(n5326), .A2(n7197), .ZN(n7288) );
  INV_X1 U6925 ( .A(n5429), .ZN(n5036) );
  NAND4_X1 U6926 ( .A1(n5423), .A2(n5517), .A3(n5037), .A4(n5036), .ZN(n5038)
         );
  NAND4_X1 U6927 ( .A1(n6659), .A2(n6660), .A3(n8794), .A4(n6658), .ZN(n5065)
         );
  NAND2_X1 U6928 ( .A1(n6151), .A2(n4566), .ZN(n6426) );
  NAND2_X1 U6929 ( .A1(n6157), .A2(n4572), .ZN(n6532) );
  NAND2_X1 U6930 ( .A1(n6157), .A2(n6156), .ZN(n6190) );
  NAND2_X1 U6931 ( .A1(n10497), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5084) );
  AOI21_X1 U6932 ( .B1(n4558), .B2(n8440), .A(n5093), .ZN(n5092) );
  NAND2_X1 U6933 ( .A1(n8441), .A2(n4558), .ZN(n5094) );
  NAND2_X1 U6934 ( .A1(n5104), .A2(n4554), .ZN(n5099) );
  OR2_X1 U6935 ( .A1(n5103), .A2(n5101), .ZN(n5100) );
  AOI21_X1 U6936 ( .B1(n5115), .B2(n9695), .A(n9665), .ZN(n9668) );
  NAND2_X1 U6937 ( .A1(n9657), .A2(n9658), .ZN(n5116) );
  NAND2_X1 U6938 ( .A1(n9635), .A2(n5126), .ZN(n5122) );
  NOR2_X1 U6939 ( .A1(n5118), .A2(n4481), .ZN(n5117) );
  NAND2_X1 U6940 ( .A1(n5123), .A2(n9642), .ZN(n9656) );
  NAND2_X1 U6941 ( .A1(n5125), .A2(n5124), .ZN(n5123) );
  INV_X1 U6942 ( .A(n9643), .ZN(n5124) );
  NAND2_X2 U6943 ( .A1(n9570), .A2(n9567), .ZN(n10374) );
  AND2_X4 U6944 ( .A1(n5433), .A2(n10318), .ZN(n5508) );
  NAND3_X1 U6945 ( .A1(n6573), .A2(n7861), .A3(n5137), .ZN(n5134) );
  INV_X1 U6946 ( .A(n7357), .ZN(n5142) );
  NAND2_X1 U6947 ( .A1(n5152), .A2(n5150), .ZN(n7591) );
  XNOR2_X2 U6948 ( .A(n5159), .B(n6160), .ZN(n6165) );
  NAND2_X1 U6949 ( .A1(n8962), .A2(n5165), .ZN(n5160) );
  INV_X1 U6950 ( .A(n5419), .ZN(n5167) );
  AND2_X1 U6951 ( .A1(n8834), .A2(n9064), .ZN(n5176) );
  OR2_X1 U6952 ( .A1(n6592), .A2(n5178), .ZN(n5177) );
  XNOR2_X1 U6953 ( .A(n5198), .B(n9673), .ZN(n7634) );
  OAI21_X1 U6954 ( .B1(n5201), .B2(n9689), .A(n5202), .ZN(n5204) );
  XNOR2_X1 U6955 ( .A(n5204), .B(n5377), .ZN(n10010) );
  INV_X1 U6956 ( .A(n5204), .ZN(n10008) );
  XNOR2_X2 U6957 ( .A(n5209), .B(n5431), .ZN(n5434) );
  NOR2_X1 U6958 ( .A1(n10310), .A2(n10312), .ZN(n5209) );
  XNOR2_X1 U6959 ( .A(n5447), .B(n5210), .ZN(n10337) );
  AND2_X1 U6960 ( .A1(n6889), .A2(SI_0_), .ZN(n5447) );
  OAI21_X1 U6961 ( .B1(n7849), .B2(n5216), .A(n5214), .ZN(n10131) );
  NAND2_X1 U6962 ( .A1(n5224), .A2(n5230), .ZN(n5225) );
  NAND2_X1 U6963 ( .A1(n5225), .A2(n5236), .ZN(n5228) );
  NAND3_X1 U6964 ( .A1(n5232), .A2(n5231), .A3(n5237), .ZN(n5229) );
  NAND3_X1 U6965 ( .A1(n5232), .A2(n5231), .A3(n5227), .ZN(n5226) );
  INV_X1 U6966 ( .A(n5233), .ZN(n5231) );
  NAND2_X1 U6967 ( .A1(n5234), .A2(n7648), .ZN(n5232) );
  AOI21_X1 U6968 ( .B1(n7648), .B2(n9578), .A(n5235), .ZN(n7676) );
  OR2_X1 U6969 ( .A1(n10245), .A2(n9833), .ZN(n5238) );
  OAI211_X2 U6970 ( .C1(n6906), .C2(n5587), .A(n5551), .B(n5259), .ZN(n9527)
         );
  NAND2_X1 U6971 ( .A1(n6632), .A2(n4474), .ZN(n5262) );
  NAND2_X1 U6972 ( .A1(n8831), .A2(n5271), .ZN(n5269) );
  NAND2_X1 U6973 ( .A1(n8891), .A2(n6642), .ZN(n5280) );
  NAND3_X1 U6974 ( .A1(n6140), .A2(n5325), .A3(n6182), .ZN(n5287) );
  INV_X1 U6975 ( .A(n5287), .ZN(n6670) );
  AND2_X1 U6976 ( .A1(n6858), .A2(n6857), .ZN(n8126) );
  INV_X1 U6977 ( .A(n8484), .ZN(n8483) );
  NAND2_X1 U6978 ( .A1(n5290), .A2(n8431), .ZN(n8429) );
  NAND3_X1 U6979 ( .A1(n5294), .A2(n8782), .A3(n5293), .ZN(n8784) );
  NAND3_X1 U6980 ( .A1(n8485), .A2(P2_REG2_REG_17__SCAN_IN), .A3(n8761), .ZN(
        n8762) );
  NAND2_X1 U6981 ( .A1(n5294), .A2(n5293), .ZN(n8783) );
  NAND2_X1 U6982 ( .A1(n7185), .A2(n10506), .ZN(n5299) );
  INV_X1 U6983 ( .A(n7185), .ZN(n5297) );
  OAI21_X1 U6984 ( .B1(n8275), .B2(n5317), .A(n5314), .ZN(n8225) );
  NAND2_X1 U6985 ( .A1(n5313), .A2(n5311), .ZN(n6748) );
  NAND2_X1 U6986 ( .A1(n8275), .A2(n5314), .ZN(n5313) );
  NAND2_X1 U6987 ( .A1(n8228), .A2(n6751), .ZN(n8305) );
  AOI21_X2 U6988 ( .B1(n8228), .B2(n5320), .A(n4525), .ZN(n7984) );
  NAND2_X1 U6989 ( .A1(n8217), .A2(n4454), .ZN(n8266) );
  NAND3_X1 U6990 ( .A1(n5324), .A2(n6702), .A3(n7509), .ZN(n5323) );
  NOR2_X1 U6991 ( .A1(n7446), .A2(n6704), .ZN(n7482) );
  AND2_X1 U6992 ( .A1(n5322), .A2(n7481), .ZN(n5321) );
  NAND2_X4 U6993 ( .A1(n5329), .A2(n5327), .ZN(n6889) );
  NAND2_X1 U6994 ( .A1(n7744), .A2(n5446), .ZN(n5329) );
  NAND2_X1 U6995 ( .A1(n5331), .A2(n9711), .ZN(n7938) );
  INV_X1 U6996 ( .A(n7460), .ZN(n5336) );
  OAI21_X1 U6997 ( .B1(n4549), .B2(n8090), .A(n8089), .ZN(n5342) );
  NAND2_X2 U6998 ( .A1(n5343), .A2(n5341), .ZN(n9498) );
  OAI21_X1 U6999 ( .B1(n5804), .B2(n5803), .A(n5802), .ZN(n5828) );
  INV_X1 U7000 ( .A(n5359), .ZN(n6043) );
  OAI21_X1 U7001 ( .B1(n6016), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7002 ( .A1(n5726), .A2(n5725), .ZN(n5371) );
  NAND2_X1 U7003 ( .A1(n5371), .A2(n5728), .ZN(n5744) );
  AOI21_X1 U7004 ( .B1(n10008), .B2(n10012), .A(n9714), .ZN(n9997) );
  NAND3_X1 U7005 ( .A1(n9532), .A2(n9533), .A3(n5382), .ZN(n9544) );
  NAND2_X1 U7006 ( .A1(n5605), .A2(n5385), .ZN(n5811) );
  NAND2_X1 U7007 ( .A1(n7853), .A2(n10160), .ZN(n10154) );
  AND2_X2 U7008 ( .A1(n10368), .A2(n5394), .ZN(n10351) );
  NAND2_X1 U7009 ( .A1(n9804), .A2(n9803), .ZN(n9811) );
  NAND2_X1 U7010 ( .A1(n10171), .A2(n10170), .ZN(n10256) );
  XNOR2_X1 U7011 ( .A(n6688), .B(n7963), .ZN(n6689) );
  OR2_X1 U7012 ( .A1(n6701), .A2(n8338), .ZN(n6702) );
  XNOR2_X1 U7013 ( .A(n7915), .B(n9689), .ZN(n7933) );
  INV_X1 U7014 ( .A(n7412), .ZN(n7415) );
  OAI21_X1 U7015 ( .B1(n9801), .B2(n9800), .A(n9799), .ZN(n9802) );
  XNOR2_X1 U7016 ( .A(n6015), .B(n6014), .ZN(n7063) );
  INV_X1 U7017 ( .A(n5811), .ZN(n5813) );
  BUF_X4 U7018 ( .A(n7198), .Z(n8137) );
  NAND2_X1 U7019 ( .A1(n6689), .A2(n7352), .ZN(n6691) );
  NAND2_X1 U7020 ( .A1(n7899), .A2(n7906), .ZN(n7994) );
  XNOR2_X1 U7021 ( .A(n5482), .B(n5481), .ZN(n7703) );
  INV_X1 U7022 ( .A(n6859), .ZN(n8131) );
  INV_X1 U7023 ( .A(n6165), .ZN(n9296) );
  XNOR2_X1 U7024 ( .A(n5477), .B(n5476), .ZN(n6899) );
  XNOR2_X1 U7025 ( .A(n5471), .B(n5489), .ZN(n5477) );
  OR2_X1 U7026 ( .A1(n10557), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5401) );
  AND2_X1 U7027 ( .A1(n6929), .A2(n6754), .ZN(n6942) );
  INV_X1 U7028 ( .A(n6942), .ZN(n6946) );
  INV_X1 U7029 ( .A(n10557), .ZN(n6883) );
  INV_X2 U7030 ( .A(n10550), .ZN(n10548) );
  OR2_X1 U7031 ( .A1(n10494), .A2(n6005), .ZN(n5402) );
  INV_X2 U7032 ( .A(n7610), .ZN(n10162) );
  INV_X1 U7033 ( .A(n10306), .ZN(n6050) );
  NAND2_X1 U7034 ( .A1(n6810), .A2(n7489), .ZN(n5404) );
  AOI21_X1 U7035 ( .B1(n6086), .B2(n10377), .A(n9356), .ZN(n7986) );
  OR2_X1 U7036 ( .A1(n8129), .A2(n9172), .ZN(n5405) );
  AND2_X1 U7037 ( .A1(n6554), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5406) );
  NOR2_X1 U7038 ( .A1(n8099), .A2(n9499), .ZN(n5409) );
  AND2_X1 U7039 ( .A1(n9326), .A2(n8047), .ZN(n5410) );
  OR2_X1 U7040 ( .A1(n10175), .A2(n10473), .ZN(n5411) );
  OR2_X1 U7041 ( .A1(n8129), .A2(n9289), .ZN(n5412) );
  OR2_X1 U7042 ( .A1(n10254), .A2(n9806), .ZN(n10473) );
  INV_X1 U7043 ( .A(n10473), .ZN(n6090) );
  AND4_X1 U7044 ( .A1(n8856), .A2(n6597), .A3(n8846), .A4(n8883), .ZN(n5413)
         );
  AND3_X2 U7045 ( .A1(n5480), .A2(n5479), .A3(n5478), .ZN(n10421) );
  AND2_X1 U7046 ( .A1(n6845), .A2(n6844), .ZN(n5414) );
  AND2_X1 U7047 ( .A1(n10206), .A2(n9822), .ZN(n5415) );
  AND2_X1 U7048 ( .A1(n8072), .A2(n9314), .ZN(n5416) );
  OR2_X1 U7049 ( .A1(n6830), .A2(n8943), .ZN(n5417) );
  NOR2_X2 U7050 ( .A1(n4459), .A2(n10215), .ZN(n10105) );
  AND2_X1 U7051 ( .A1(n7990), .A2(n6091), .ZN(n5418) );
  NAND2_X1 U7052 ( .A1(n9144), .A2(n8976), .ZN(n5419) );
  AND2_X1 U7053 ( .A1(n8892), .A2(n8905), .ZN(n5420) );
  OR2_X1 U7054 ( .A1(n5582), .A2(n9852), .ZN(n5422) );
  AND2_X1 U7055 ( .A1(n7183), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7184) );
  OR2_X1 U7056 ( .A1(n9316), .A2(n9315), .ZN(n8072) );
  INV_X1 U7057 ( .A(n5706), .ZN(n5707) );
  INV_X1 U7058 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5626) );
  INV_X1 U7059 ( .A(n8943), .ZN(n6733) );
  INV_X1 U7060 ( .A(n9198), .ZN(n6837) );
  INV_X1 U7061 ( .A(n6426), .ZN(n6152) );
  INV_X1 U7062 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6107) );
  INV_X1 U7063 ( .A(n5875), .ZN(n5872) );
  NAND2_X1 U7064 ( .A1(n9347), .A2(n6090), .ZN(n6091) );
  NAND2_X1 U7065 ( .A1(n5994), .A2(n5993), .ZN(n5996) );
  AND2_X1 U7066 ( .A1(n5926), .A2(n5923), .ZN(n5949) );
  INV_X1 U7067 ( .A(SI_19_), .ZN(n8513) );
  INV_X1 U7068 ( .A(n5759), .ZN(n5760) );
  INV_X1 U7069 ( .A(SI_9_), .ZN(n8689) );
  INV_X1 U7070 ( .A(n8975), .ZN(n6722) );
  AND2_X1 U7071 ( .A1(n8290), .A2(n6711), .ZN(n6712) );
  INV_X1 U7072 ( .A(n9024), .ZN(n8291) );
  OR2_X1 U7073 ( .A1(n6709), .A2(n7655), .ZN(n6710) );
  NAND2_X1 U7074 ( .A1(n6603), .A2(n6581), .ZN(n6806) );
  INV_X1 U7075 ( .A(n6185), .ZN(n6183) );
  OR2_X1 U7076 ( .A1(n5557), .A2(n7805), .ZN(n5559) );
  INV_X1 U7077 ( .A(n10117), .ZN(n10380) );
  OR2_X1 U7078 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  AND2_X1 U7079 ( .A1(n5929), .A2(n5928), .ZN(n5953) );
  INV_X1 U7080 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7081 ( .A1(n5764), .A2(n5763), .ZN(n5784) );
  NAND2_X1 U7082 ( .A1(n5657), .A2(n5656), .ZN(n5673) );
  NAND2_X1 U7083 ( .A1(n5597), .A2(n5596), .ZN(n5615) );
  NAND2_X1 U7084 ( .A1(n6721), .A2(n6722), .ZN(n6723) );
  INV_X1 U7085 ( .A(n8834), .ZN(n7978) );
  INV_X1 U7086 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8738) );
  INV_X1 U7087 ( .A(n6575), .ZN(n6660) );
  OR2_X1 U7088 ( .A1(n7172), .A2(n9302), .ZN(n7318) );
  NAND2_X1 U7089 ( .A1(n7953), .A2(n6600), .ZN(n7346) );
  INV_X1 U7090 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6216) );
  NAND2_X1 U7091 ( .A1(n4437), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5510) );
  INV_X1 U7092 ( .A(n8005), .ZN(n7112) );
  AND2_X1 U7093 ( .A1(n6077), .A2(n9798), .ZN(n10152) );
  AND2_X1 U7094 ( .A1(n5635), .A2(n5621), .ZN(n5633) );
  XNOR2_X1 U7095 ( .A(n6734), .B(n8907), .ZN(n8202) );
  AOI21_X1 U7096 ( .B1(n6690), .B2(n7212), .A(n6599), .ZN(n7146) );
  INV_X1 U7097 ( .A(n7838), .ZN(n6780) );
  INV_X1 U7098 ( .A(n8778), .ZN(n10513) );
  NOR2_X1 U7099 ( .A1(n7318), .A2(n8788), .ZN(n10499) );
  OR2_X1 U7100 ( .A1(n10537), .A2(n7360), .ZN(n8995) );
  INV_X1 U7101 ( .A(n10537), .ZN(n10543) );
  AND3_X1 U7102 ( .A1(n6879), .A2(n6878), .A3(n6877), .ZN(n7333) );
  AND2_X1 U7103 ( .A1(n6648), .A2(n6647), .ZN(n8846) );
  AND2_X1 U7104 ( .A1(n8978), .A2(n8977), .ZN(n9258) );
  OR2_X1 U7105 ( .A1(n4435), .A2(n6780), .ZN(n10537) );
  INV_X1 U7106 ( .A(n9289), .ZN(n9277) );
  NAND2_X1 U7107 ( .A1(n9069), .A2(n10525), .ZN(n10544) );
  XNOR2_X1 U7108 ( .A(n6673), .B(n8573), .ZN(n6680) );
  XNOR2_X1 U7109 ( .A(n6405), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8448) );
  INV_X1 U7110 ( .A(n9559), .ZN(n9533) );
  INV_X1 U7111 ( .A(n9802), .ZN(n9803) );
  INV_X1 U7112 ( .A(n9960), .ZN(n9984) );
  AND2_X1 U7113 ( .A1(n6923), .A2(n6922), .ZN(n6985) );
  AND2_X1 U7114 ( .A1(n7059), .A2(n9784), .ZN(n10390) );
  INV_X1 U7115 ( .A(n10082), .ZN(n10392) );
  INV_X1 U7116 ( .A(n10152), .ZN(n10377) );
  OR2_X1 U7117 ( .A1(n7061), .A2(n7060), .ZN(n10117) );
  INV_X1 U7118 ( .A(n9671), .ZN(n10149) );
  NAND2_X1 U7119 ( .A1(n10410), .A2(n10451), .ZN(n10480) );
  AND2_X1 U7120 ( .A1(n6047), .A2(n7608), .ZN(n6096) );
  AND2_X1 U7121 ( .A1(n6049), .A2(n6048), .ZN(n7606) );
  AND2_X1 U7122 ( .A1(n5696), .A2(n5712), .ZN(n7392) );
  INV_X1 U7123 ( .A(n6800), .ZN(n6801) );
  INV_X1 U7124 ( .A(n8329), .ZN(n8294) );
  INV_X1 U7125 ( .A(n8232), .ZN(n8871) );
  INV_X1 U7126 ( .A(n7685), .ZN(n9066) );
  INV_X1 U7127 ( .A(n10499), .ZN(n8781) );
  OR2_X1 U7128 ( .A1(n8981), .A2(n7361), .ZN(n9086) );
  NAND2_X1 U7129 ( .A1(n10557), .A2(n10544), .ZN(n9162) );
  AND3_X2 U7130 ( .A1(n6882), .A2(n7333), .A3(n6881), .ZN(n10557) );
  OR2_X1 U7131 ( .A1(n10550), .A2(n9119), .ZN(n9280) );
  OR2_X1 U7132 ( .A1(n10550), .A2(n10537), .ZN(n9289) );
  AND2_X1 U7133 ( .A1(n6867), .A2(n6866), .ZN(n10550) );
  AND2_X1 U7134 ( .A1(n6787), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6929) );
  INV_X1 U7135 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8549) );
  INV_X1 U7136 ( .A(n7574), .ZN(n7755) );
  INV_X1 U7137 ( .A(n9603), .ZN(n10474) );
  AND2_X1 U7138 ( .A1(n7062), .A2(n10117), .ZN(n9545) );
  INV_X1 U7139 ( .A(n7892), .ZN(n9815) );
  INV_X1 U7140 ( .A(n9990), .ZN(n9939) );
  OR2_X1 U7141 ( .A1(n7609), .A2(n9991), .ZN(n10082) );
  NAND2_X1 U7142 ( .A1(n10494), .A2(n10480), .ZN(n10243) );
  INV_X1 U7143 ( .A(n10494), .ZN(n10492) );
  XNOR2_X1 U7144 ( .A(n7887), .B(n7890), .ZN(n7914) );
  NAND2_X1 U7145 ( .A1(n10482), .A2(n10480), .ZN(n10306) );
  INV_X1 U7146 ( .A(n10482), .ZN(n10481) );
  INV_X1 U7147 ( .A(n10405), .ZN(n10406) );
  INV_X1 U7148 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8717) );
  INV_X1 U7149 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6891) );
  INV_X1 U7150 ( .A(n10315), .ZN(n10332) );
  INV_X1 U7151 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10562) );
  INV_X2 U7152 ( .A(n8774), .ZN(P2_U3893) );
  INV_X1 U7153 ( .A(n9839), .ZN(P1_U3973) );
  OAI211_X1 U7154 ( .C1(n6099), .C2(n10243), .A(n6098), .B(n5402), .ZN(
        P1_U3550) );
  NAND2_X1 U7155 ( .A1(n6095), .A2(n6094), .ZN(P1_U3518) );
  NOR2_X1 U7156 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5426) );
  NOR2_X1 U7157 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5425) );
  NOR2_X1 U7158 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5424) );
  NAND4_X1 U7159 ( .A1(n5426), .A2(n5425), .A3(n5424), .A4(n6017), .ZN(n5429)
         );
  NAND4_X1 U7160 ( .A1(n8556), .A2(n5749), .A3(n6012), .A4(n5427), .ZN(n5428)
         );
  NAND2_X1 U7161 ( .A1(n5509), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5438) );
  NAND2_X1 U7162 ( .A1(n5508), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7163 ( .A1(n5572), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5436) );
  NAND4_X1 U7164 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n7077)
         );
  INV_X1 U7165 ( .A(n7077), .ZN(n5459) );
  OAI21_X1 U7166 ( .B1(n5439), .B2(n10312), .A(P1_IR_REG_28__SCAN_IN), .ZN(
        n5441) );
  NAND2_X1 U7167 ( .A1(n5441), .A2(n5440), .ZN(n5442) );
  NAND2_X1 U7168 ( .A1(n5432), .A2(n5442), .ZN(n6084) );
  XNOR2_X2 U7169 ( .A(n5445), .B(n5444), .ZN(n6924) );
  INV_X1 U7170 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U7171 ( .A1(n5447), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5450) );
  AND2_X1 U7172 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7173 ( .A1(n5450), .A2(n6242), .ZN(n5493) );
  INV_X1 U7174 ( .A(SI_1_), .ZN(n5472) );
  XNOR2_X1 U7175 ( .A(n5493), .B(n5472), .ZN(n5452) );
  MUX2_X1 U7176 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6142), .Z(n5451) );
  NOR2_X1 U7177 ( .A1(n4431), .A2(n6911), .ZN(n5453) );
  NAND2_X1 U7178 ( .A1(n5582), .A2(n5453), .ZN(n5457) );
  INV_X1 U7179 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U7180 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5454) );
  NAND2_X1 U7181 ( .A1(n4438), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U7182 ( .A1(n4436), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5462) );
  NAND2_X1 U7183 ( .A1(n5508), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U7184 ( .A1(n5572), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5460) );
  NAND4_X2 U7185 ( .A1(n5463), .A2(n5462), .A3(n5461), .A4(n5460), .ZN(n9840)
         );
  MUX2_X1 U7186 ( .A(P1_IR_REG_0__SCAN_IN), .B(n10337), .S(n4432), .Z(n7141)
         );
  NAND2_X1 U7187 ( .A1(n9840), .A2(n7141), .ZN(n7713) );
  NAND2_X1 U7188 ( .A1(n7712), .A2(n7713), .ZN(n5466) );
  CLKBUF_X1 U7189 ( .A(n7077), .Z(n5464) );
  OR2_X1 U7190 ( .A1(n5464), .A2(n5458), .ZN(n5465) );
  NAND2_X1 U7191 ( .A1(n5466), .A2(n5465), .ZN(n7696) );
  NAND2_X1 U7192 ( .A1(n4439), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7193 ( .A1(n5572), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U7194 ( .A1(n4436), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U7195 ( .A1(n5508), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5467) );
  NAND4_X2 U7196 ( .A1(n5470), .A2(n5469), .A3(n5468), .A4(n5467), .ZN(n5482)
         );
  INV_X1 U7197 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6896) );
  OR2_X1 U7198 ( .A1(n7876), .A2(n6896), .ZN(n5480) );
  INV_X1 U7199 ( .A(SI_2_), .ZN(n5489) );
  INV_X1 U7200 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U7201 ( .A1(n6889), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5473) );
  OAI211_X1 U7202 ( .C1(n6889), .C2(n6910), .A(n5473), .B(n5472), .ZN(n5490)
         );
  NAND2_X1 U7203 ( .A1(n5493), .A2(n5490), .ZN(n5475) );
  NAND2_X1 U7204 ( .A1(n6142), .A2(n6895), .ZN(n5474) );
  OAI211_X1 U7205 ( .C1(n6142), .C2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .B(
        n5474), .ZN(n5498) );
  NAND2_X1 U7206 ( .A1(n5475), .A2(n5498), .ZN(n5476) );
  INV_X1 U7207 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5500) );
  OR2_X1 U7208 ( .A1(n5582), .A2(n7106), .ZN(n5478) );
  INV_X1 U7209 ( .A(n7703), .ZN(n9675) );
  NAND2_X1 U7210 ( .A1(n7696), .A2(n9675), .ZN(n5484) );
  OR2_X1 U7211 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  INV_X2 U7212 ( .A(n5572), .ZN(n5557) );
  OR2_X1 U7213 ( .A1(n5557), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5487) );
  INV_X1 U7214 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6954) );
  NAND2_X1 U7215 ( .A1(n4438), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5486) );
  INV_X1 U7216 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5485) );
  INV_X1 U7217 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6894) );
  OR2_X1 U7218 ( .A1(n7876), .A2(n6894), .ZN(n5507) );
  INV_X1 U7219 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6898) );
  NAND2_X1 U7220 ( .A1(n6889), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5488) );
  OAI211_X1 U7221 ( .C1(n6889), .C2(n6898), .A(n5489), .B(n5488), .ZN(n5491)
         );
  INV_X1 U7222 ( .A(n5491), .ZN(n5497) );
  NAND2_X1 U7223 ( .A1(n5493), .A2(n5492), .ZN(n5496) );
  NAND2_X1 U7224 ( .A1(n6142), .A2(n6896), .ZN(n5494) );
  OAI211_X1 U7225 ( .C1(n6142), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5494), .B(
        SI_2_), .ZN(n5495) );
  MUX2_X1 U7226 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6889), .Z(n5521) );
  INV_X1 U7227 ( .A(SI_3_), .ZN(n5499) );
  XNOR2_X1 U7228 ( .A(n5521), .B(n5499), .ZN(n5519) );
  XNOR2_X1 U7229 ( .A(n5519), .B(n5520), .ZN(n6909) );
  OR2_X1 U7230 ( .A1(n5587), .A2(n6909), .ZN(n5505) );
  NAND2_X1 U7231 ( .A1(n5501), .A2(n5500), .ZN(n5502) );
  NAND2_X1 U7232 ( .A1(n5502), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5504) );
  INV_X1 U7233 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5503) );
  AND2_X1 U7234 ( .A1(n5505), .A2(n5422), .ZN(n5506) );
  NAND2_X1 U7235 ( .A1(n5508), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5512) );
  INV_X1 U7236 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6978) );
  OAI21_X1 U7237 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5554), .ZN(n10379) );
  OR2_X1 U7238 ( .A1(n5557), .A2(n10379), .ZN(n5511) );
  AND2_X1 U7239 ( .A1(n5513), .A2(n5601), .ZN(n5514) );
  NOR2_X1 U7240 ( .A1(n5514), .A2(n10312), .ZN(n5515) );
  MUX2_X1 U7241 ( .A(n10312), .B(n5515), .S(P1_IR_REG_4__SCAN_IN), .Z(n5516)
         );
  INV_X1 U7242 ( .A(n5516), .ZN(n5518) );
  INV_X1 U7243 ( .A(n5517), .ZN(n5536) );
  NAND2_X1 U7244 ( .A1(n5518), .A2(n5536), .ZN(n9870) );
  INV_X1 U7245 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8686) );
  INV_X1 U7246 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6890) );
  MUX2_X1 U7247 ( .A(n8686), .B(n6890), .S(n6142), .Z(n5542) );
  NAND2_X1 U7248 ( .A1(n5520), .A2(n5519), .ZN(n5523) );
  NAND2_X1 U7249 ( .A1(n5521), .A2(SI_3_), .ZN(n5522) );
  NAND2_X1 U7250 ( .A1(n5523), .A2(n5522), .ZN(n5541) );
  XNOR2_X1 U7251 ( .A(n5541), .B(n5540), .ZN(n6907) );
  OR2_X1 U7252 ( .A1(n5587), .A2(n6907), .ZN(n5525) );
  OR2_X1 U7253 ( .A1(n7876), .A2(n6890), .ZN(n5524) );
  OAI211_X1 U7254 ( .C1(n4432), .C2(n9870), .A(n5525), .B(n5524), .ZN(n7298)
         );
  NAND2_X1 U7255 ( .A1(n7291), .A2(n7298), .ZN(n9568) );
  INV_X1 U7256 ( .A(n7298), .ZN(n10432) );
  NAND2_X1 U7257 ( .A1(n9837), .A2(n10432), .ZN(n6054) );
  NAND2_X1 U7258 ( .A1(n9568), .A2(n6054), .ZN(n9672) );
  NAND3_X1 U7259 ( .A1(n7637), .A2(n10386), .A3(n9672), .ZN(n5528) );
  NOR2_X1 U7260 ( .A1(n9838), .A2(n7203), .ZN(n10385) );
  NOR2_X1 U7261 ( .A1(n9837), .A2(n7298), .ZN(n5526) );
  AOI21_X1 U7262 ( .B1(n9672), .B2(n10385), .A(n5526), .ZN(n5527) );
  NAND2_X1 U7263 ( .A1(n5528), .A2(n5527), .ZN(n7803) );
  NAND2_X1 U7264 ( .A1(n4436), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5535) );
  INV_X1 U7265 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6981) );
  OR2_X1 U7266 ( .A1(n5625), .A2(n6981), .ZN(n5534) );
  INV_X1 U7267 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6963) );
  NOR2_X2 U7268 ( .A1(n5554), .A2(n5553), .ZN(n5529) );
  INV_X1 U7269 ( .A(n5529), .ZN(n5556) );
  INV_X1 U7270 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7271 ( .A1(n5556), .A2(n5530), .ZN(n5531) );
  NAND2_X1 U7272 ( .A1(n5574), .A2(n5531), .ZN(n10360) );
  OR2_X1 U7273 ( .A1(n5557), .A2(n10360), .ZN(n5532) );
  INV_X1 U7274 ( .A(n7538), .ZN(n9835) );
  NAND2_X1 U7275 ( .A1(n4518), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5538) );
  INV_X1 U7276 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7277 ( .A1(n5538), .A2(n5537), .ZN(n5583) );
  OR2_X1 U7278 ( .A1(n5538), .A2(n5537), .ZN(n5539) );
  NAND2_X1 U7279 ( .A1(n5583), .A2(n5539), .ZN(n9900) );
  NAND2_X1 U7280 ( .A1(n5541), .A2(n5540), .ZN(n5545) );
  INV_X1 U7281 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7282 ( .A1(n5543), .A2(SI_4_), .ZN(n5544) );
  INV_X1 U7283 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5546) );
  MUX2_X1 U7284 ( .A(n5546), .B(n6891), .S(n6142), .Z(n5547) );
  XNOR2_X1 U7285 ( .A(n5547), .B(SI_5_), .ZN(n5564) );
  INV_X1 U7286 ( .A(n5547), .ZN(n5548) );
  NAND2_X1 U7287 ( .A1(n5548), .A2(SI_5_), .ZN(n5549) );
  XNOR2_X1 U7288 ( .A(n5586), .B(n8588), .ZN(n5585) );
  INV_X1 U7289 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6897) );
  OR2_X1 U7290 ( .A1(n7876), .A2(n6897), .ZN(n5551) );
  INV_X1 U7291 ( .A(n9527), .ZN(n10445) );
  NAND2_X1 U7292 ( .A1(n7538), .A2(n9527), .ZN(n9577) );
  NAND2_X1 U7293 ( .A1(n7643), .A2(n9577), .ZN(n10356) );
  NAND2_X1 U7294 ( .A1(n5554), .A2(n5553), .ZN(n5555) );
  NAND2_X1 U7295 ( .A1(n5556), .A2(n5555), .ZN(n7805) );
  NAND2_X1 U7296 ( .A1(n4439), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5558) );
  INV_X1 U7297 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6958) );
  OR2_X1 U7298 ( .A1(n6081), .A2(n6958), .ZN(n5561) );
  OR2_X1 U7299 ( .A1(n5517), .A2(n10312), .ZN(n5563) );
  INV_X1 U7300 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5562) );
  XNOR2_X1 U7301 ( .A(n5563), .B(n5562), .ZN(n9886) );
  OR2_X1 U7302 ( .A1(n7876), .A2(n6891), .ZN(n5565) );
  OAI211_X1 U7303 ( .C1(n5582), .C2(n9886), .A(n5566), .B(n5565), .ZN(n7808)
         );
  NAND2_X1 U7304 ( .A1(n7463), .A2(n7808), .ZN(n9571) );
  NAND2_X1 U7305 ( .A1(n9836), .A2(n10439), .ZN(n9746) );
  AND2_X1 U7306 ( .A1(n10356), .A2(n7798), .ZN(n5567) );
  NAND2_X1 U7307 ( .A1(n7803), .A2(n5567), .ZN(n5570) );
  NOR2_X1 U7308 ( .A1(n9836), .A2(n7808), .ZN(n10364) );
  NOR2_X1 U7309 ( .A1(n9835), .A2(n9527), .ZN(n5568) );
  AOI21_X1 U7310 ( .B1(n10356), .B2(n10364), .A(n5568), .ZN(n5569) );
  NAND2_X1 U7311 ( .A1(n5570), .A2(n5569), .ZN(n7648) );
  NAND2_X1 U7312 ( .A1(n4438), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5581) );
  INV_X1 U7313 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5571) );
  OR2_X1 U7314 ( .A1(n6081), .A2(n5571), .ZN(n5580) );
  NAND2_X1 U7315 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  NAND2_X1 U7316 ( .A1(n5609), .A2(n5575), .ZN(n7649) );
  OR2_X1 U7317 ( .A1(n5557), .A2(n7649), .ZN(n5579) );
  INV_X1 U7318 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5577) );
  OR2_X1 U7319 ( .A1(n5576), .A2(n5577), .ZN(n5578) );
  NAND2_X1 U7320 ( .A1(n5583), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5584) );
  XNOR2_X1 U7321 ( .A(n5584), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9916) );
  AOI22_X1 U7322 ( .A1(n5815), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6919), .B2(
        n9916), .ZN(n5589) );
  XNOR2_X1 U7323 ( .A(n5592), .B(n5590), .ZN(n6900) );
  INV_X2 U7324 ( .A(n5587), .ZN(n5637) );
  NAND2_X1 U7325 ( .A1(n6900), .A2(n5637), .ZN(n5588) );
  NAND2_X1 U7326 ( .A1(n7526), .A2(n7528), .ZN(n7666) );
  NAND2_X1 U7327 ( .A1(n9834), .A2(n10455), .ZN(n6057) );
  NAND2_X1 U7328 ( .A1(n7666), .A2(n6057), .ZN(n9578) );
  NAND2_X1 U7329 ( .A1(n5593), .A2(SI_7_), .ZN(n5594) );
  INV_X1 U7330 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6914) );
  INV_X1 U7331 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5595) );
  INV_X1 U7332 ( .A(SI_8_), .ZN(n5596) );
  INV_X1 U7333 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7334 ( .A1(n5598), .A2(SI_8_), .ZN(n5599) );
  NOR2_X1 U7335 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5600) );
  NAND2_X1 U7336 ( .A1(n5603), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5602) );
  MUX2_X1 U7337 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5602), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5606) );
  AND2_X1 U7338 ( .A1(n5606), .A2(n5772), .ZN(n7000) );
  AOI22_X1 U7339 ( .A1(n5815), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6919), .B2(
        n7000), .ZN(n5607) );
  NAND2_X1 U7340 ( .A1(n4439), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7341 ( .A1(n5609), .A2(n5608), .ZN(n5610) );
  NAND2_X1 U7342 ( .A1(n5627), .A2(n5610), .ZN(n9369) );
  OR2_X1 U7343 ( .A1(n5557), .A2(n9369), .ZN(n5613) );
  NAND2_X1 U7344 ( .A1(n5508), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7345 ( .A1(n4436), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5611) );
  NAND4_X1 U7346 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n9833)
         );
  NAND2_X1 U7347 ( .A1(n9370), .A2(n9833), .ZN(n9583) );
  INV_X1 U7348 ( .A(n9833), .ZN(n8015) );
  NAND2_X1 U7349 ( .A1(n10245), .A2(n8015), .ZN(n9584) );
  INV_X1 U7350 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7351 ( .A1(n5620), .A2(SI_9_), .ZN(n5621) );
  XNOR2_X1 U7352 ( .A(n5634), .B(n5633), .ZN(n6930) );
  NAND2_X1 U7353 ( .A1(n6930), .A2(n5637), .ZN(n5624) );
  NAND2_X1 U7354 ( .A1(n5772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5622) );
  XNOR2_X1 U7355 ( .A(n5622), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7025) );
  AOI22_X1 U7356 ( .A1(n5815), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6919), .B2(
        n7025), .ZN(n5623) );
  NAND2_X1 U7357 ( .A1(n4436), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5632) );
  INV_X1 U7358 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7792) );
  OR2_X1 U7359 ( .A1(n5625), .A2(n7792), .ZN(n5631) );
  INV_X1 U7360 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n7003) );
  OR2_X1 U7361 ( .A1(n6081), .A2(n7003), .ZN(n5630) );
  NAND2_X1 U7362 ( .A1(n5627), .A2(n5626), .ZN(n5628) );
  NAND2_X1 U7363 ( .A1(n5643), .A2(n5628), .ZN(n9446) );
  OR2_X1 U7364 ( .A1(n5557), .A2(n9446), .ZN(n5629) );
  NAND2_X1 U7365 ( .A1(n8026), .A2(n7668), .ZN(n9596) );
  NAND2_X1 U7366 ( .A1(n9591), .A2(n9596), .ZN(n7787) );
  INV_X1 U7367 ( .A(n8026), .ZN(n10462) );
  OR2_X1 U7368 ( .A1(n5772), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U7369 ( .A1(n5638), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5641) );
  INV_X1 U7370 ( .A(n5638), .ZN(n5640) );
  INV_X1 U7371 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5639) );
  NAND2_X1 U7372 ( .A1(n5640), .A2(n5639), .ZN(n5660) );
  AOI22_X1 U7373 ( .A1(n5815), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6919), .B2(
        n7005), .ZN(n5642) );
  NAND2_X1 U7374 ( .A1(n4437), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5650) );
  INV_X1 U7375 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U7376 ( .A1(n5643), .A2(n8722), .ZN(n5644) );
  NAND2_X1 U7377 ( .A1(n5666), .A2(n5644), .ZN(n10343) );
  OR2_X1 U7378 ( .A1(n5557), .A2(n10343), .ZN(n5649) );
  INV_X1 U7379 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5645) );
  OR2_X1 U7380 ( .A1(n5625), .A2(n5645), .ZN(n5648) );
  INV_X1 U7381 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5646) );
  OR2_X1 U7382 ( .A1(n6081), .A2(n5646), .ZN(n5647) );
  INV_X1 U7383 ( .A(n5652), .ZN(n5653) );
  NAND2_X1 U7384 ( .A1(n5653), .A2(SI_10_), .ZN(n5654) );
  INV_X1 U7385 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7386 ( .A1(n5658), .A2(SI_11_), .ZN(n5659) );
  NAND2_X1 U7387 ( .A1(n6947), .A2(n5637), .ZN(n5663) );
  NAND2_X1 U7388 ( .A1(n5660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5661) );
  XNOR2_X1 U7389 ( .A(n5661), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7033) );
  AOI22_X1 U7390 ( .A1(n5815), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6919), .B2(
        n7033), .ZN(n5662) );
  NAND2_X1 U7391 ( .A1(n4439), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5672) );
  INV_X1 U7392 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5664) );
  OR2_X1 U7393 ( .A1(n5576), .A2(n5664), .ZN(n5671) );
  NAND2_X1 U7394 ( .A1(n5666), .A2(n5665), .ZN(n5667) );
  NAND2_X1 U7395 ( .A1(n5684), .A2(n5667), .ZN(n9492) );
  OR2_X1 U7396 ( .A1(n5557), .A2(n9492), .ZN(n5670) );
  INV_X1 U7397 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5668) );
  OR2_X1 U7398 ( .A1(n6081), .A2(n5668), .ZN(n5669) );
  OR2_X2 U7399 ( .A1(n9603), .A2(n9601), .ZN(n9589) );
  NAND2_X1 U7400 ( .A1(n9603), .A2(n9601), .ZN(n9595) );
  NAND2_X1 U7401 ( .A1(n9589), .A2(n9595), .ZN(n9681) );
  MUX2_X1 U7402 ( .A(n8549), .B(n7095), .S(n4956), .Z(n5691) );
  XNOR2_X1 U7403 ( .A(n5693), .B(n5690), .ZN(n7093) );
  INV_X1 U7404 ( .A(n5674), .ZN(n5675) );
  AOI21_X1 U7405 ( .B1(n5675), .B2(n5770), .A(n10312), .ZN(n5676) );
  MUX2_X1 U7406 ( .A(n10312), .B(n5676), .S(P1_IR_REG_12__SCAN_IN), .Z(n5678)
         );
  OR2_X1 U7407 ( .A1(n5678), .A2(n5677), .ZN(n7252) );
  INV_X1 U7408 ( .A(n7252), .ZN(n7249) );
  AOI22_X1 U7409 ( .A1(n5815), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6919), .B2(
        n7249), .ZN(n5679) );
  NAND2_X1 U7410 ( .A1(n4437), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5689) );
  INV_X1 U7411 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10241) );
  OR2_X1 U7412 ( .A1(n6081), .A2(n10241), .ZN(n5688) );
  INV_X1 U7413 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5681) );
  OR2_X1 U7414 ( .A1(n5625), .A2(n5681), .ZN(n5687) );
  INV_X1 U7415 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5683) );
  NAND2_X1 U7416 ( .A1(n5684), .A2(n5683), .ZN(n5685) );
  NAND2_X1 U7417 ( .A1(n5700), .A2(n5685), .ZN(n9392) );
  OR2_X1 U7418 ( .A1(n5557), .A2(n9392), .ZN(n5686) );
  NAND2_X1 U7419 ( .A1(n10240), .A2(n9605), .ZN(n9755) );
  INV_X1 U7420 ( .A(n5691), .ZN(n5692) );
  XNOR2_X1 U7421 ( .A(n5708), .B(n5706), .ZN(n7096) );
  NAND2_X1 U7422 ( .A1(n7096), .A2(n5637), .ZN(n5698) );
  INV_X1 U7423 ( .A(n5677), .ZN(n5695) );
  NAND2_X1 U7424 ( .A1(n5695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5694) );
  MUX2_X1 U7425 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5694), .S(
        P1_IR_REG_13__SCAN_IN), .Z(n5696) );
  OR2_X1 U7426 ( .A1(n5695), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5712) );
  AOI22_X1 U7427 ( .A1(n5815), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6919), .B2(
        n7392), .ZN(n5697) );
  NAND2_X1 U7428 ( .A1(n4438), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5705) );
  INV_X1 U7429 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10300) );
  OR2_X1 U7430 ( .A1(n5576), .A2(n10300), .ZN(n5704) );
  INV_X1 U7431 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5699) );
  OR2_X2 U7432 ( .A1(n5700), .A2(n5699), .ZN(n5716) );
  NAND2_X1 U7433 ( .A1(n5700), .A2(n5699), .ZN(n5701) );
  NAND2_X1 U7434 ( .A1(n5716), .A2(n5701), .ZN(n9468) );
  OR2_X1 U7435 ( .A1(n5557), .A2(n9468), .ZN(n5703) );
  INV_X1 U7436 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10236) );
  OR2_X1 U7437 ( .A1(n6081), .A2(n10236), .ZN(n5702) );
  NAND2_X1 U7438 ( .A1(n10235), .A2(n8062), .ZN(n9756) );
  NAND2_X1 U7439 ( .A1(n9758), .A2(n9756), .ZN(n7839) );
  INV_X1 U7440 ( .A(n10235), .ZN(n9473) );
  NAND2_X1 U7441 ( .A1(n5709), .A2(SI_13_), .ZN(n5710) );
  NAND2_X1 U7442 ( .A1(n5712), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5748) );
  XNOR2_X1 U7443 ( .A(n5748), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7582) );
  AOI22_X1 U7444 ( .A1(n5815), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6919), .B2(
        n7582), .ZN(n5713) );
  NAND2_X1 U7445 ( .A1(n5508), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5722) );
  INV_X1 U7446 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5714) );
  OR2_X1 U7447 ( .A1(n5625), .A2(n5714), .ZN(n5721) );
  INV_X1 U7448 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7449 ( .A1(n5716), .A2(n5715), .ZN(n5717) );
  NAND2_X1 U7450 ( .A1(n5734), .A2(n5717), .ZN(n9321) );
  OR2_X1 U7451 ( .A1(n5557), .A2(n9321), .ZN(n5720) );
  INV_X1 U7452 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5718) );
  OR2_X1 U7453 ( .A1(n5576), .A2(n5718), .ZN(n5719) );
  NAND2_X1 U7454 ( .A1(n8066), .A2(n8064), .ZN(n5723) );
  INV_X1 U7455 ( .A(n8064), .ZN(n9827) );
  NAND2_X1 U7456 ( .A1(n5727), .A2(SI_14_), .ZN(n5728) );
  MUX2_X1 U7457 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4956), .Z(n5740) );
  XNOR2_X1 U7458 ( .A(n5740), .B(SI_15_), .ZN(n5729) );
  XNOR2_X1 U7459 ( .A(n5744), .B(n5729), .ZN(n7301) );
  NAND2_X1 U7460 ( .A1(n7301), .A2(n5637), .ZN(n5733) );
  INV_X1 U7461 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U7462 ( .A1(n5748), .A2(n8724), .ZN(n5730) );
  NAND2_X1 U7463 ( .A1(n5730), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5731) );
  XNOR2_X1 U7464 ( .A(n5731), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7583) );
  AOI22_X1 U7465 ( .A1(n5815), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6919), .B2(
        n7583), .ZN(n5732) );
  INV_X1 U7466 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U7467 ( .A1(n5734), .A2(n9553), .ZN(n5735) );
  NAND2_X1 U7468 ( .A1(n5753), .A2(n5735), .ZN(n10156) );
  OR2_X1 U7469 ( .A1(n5557), .A2(n10156), .ZN(n5739) );
  INV_X1 U7470 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10295) );
  OR2_X1 U7471 ( .A1(n5576), .A2(n10295), .ZN(n5738) );
  NAND2_X1 U7472 ( .A1(n5508), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7473 ( .A1(n4439), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5736) );
  NAND4_X1 U7474 ( .A1(n5739), .A2(n5738), .A3(n5737), .A4(n5736), .ZN(n9826)
         );
  INV_X1 U7475 ( .A(n9826), .ZN(n6061) );
  INV_X1 U7476 ( .A(n5740), .ZN(n5742) );
  INV_X1 U7477 ( .A(SI_15_), .ZN(n5741) );
  XNOR2_X1 U7478 ( .A(n5759), .B(SI_16_), .ZN(n5745) );
  XNOR2_X1 U7479 ( .A(n5762), .B(n5745), .ZN(n7327) );
  NAND2_X1 U7480 ( .A1(n7327), .A2(n5637), .ZN(n5752) );
  OR2_X1 U7481 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5746) );
  NAND2_X1 U7482 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5746), .ZN(n5747) );
  NAND2_X1 U7483 ( .A1(n5748), .A2(n5747), .ZN(n5750) );
  XNOR2_X1 U7484 ( .A(n5750), .B(n5749), .ZN(n9942) );
  AOI22_X1 U7485 ( .A1(n5815), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6919), .B2(
        n9942), .ZN(n5751) );
  INV_X1 U7486 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U7487 ( .A1(n5753), .A2(n9414), .ZN(n5754) );
  NAND2_X1 U7488 ( .A1(n5777), .A2(n5754), .ZN(n10140) );
  NAND2_X1 U7489 ( .A1(n4436), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5755) );
  OAI21_X1 U7490 ( .B1(n10140), .B2(n5557), .A(n5755), .ZN(n5758) );
  INV_X1 U7491 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10221) );
  INV_X1 U7492 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5756) );
  OAI22_X1 U7493 ( .A1(n6081), .A2(n10221), .B1(n5625), .B2(n5756), .ZN(n5757)
         );
  NAND2_X1 U7494 ( .A1(n10220), .A2(n8083), .ZN(n9619) );
  NAND2_X1 U7495 ( .A1(n9617), .A2(n9619), .ZN(n10135) );
  INV_X1 U7496 ( .A(n10220), .ZN(n10144) );
  INV_X1 U7497 ( .A(SI_17_), .ZN(n5763) );
  INV_X1 U7498 ( .A(n5764), .ZN(n5765) );
  NAND2_X1 U7499 ( .A1(n5765), .A2(SI_17_), .ZN(n5766) );
  XNOR2_X1 U7500 ( .A(n5786), .B(n5785), .ZN(n7474) );
  NAND2_X1 U7501 ( .A1(n7474), .A2(n5637), .ZN(n5775) );
  NOR2_X1 U7502 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5768) );
  NOR2_X1 U7503 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5767) );
  NAND4_X1 U7504 ( .A1(n5769), .A2(n5770), .A3(n5768), .A4(n5767), .ZN(n5771)
         );
  NAND2_X1 U7505 ( .A1(n4561), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5773) );
  XNOR2_X1 U7506 ( .A(n5773), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9943) );
  AOI22_X1 U7507 ( .A1(n5815), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6919), .B2(
        n9943), .ZN(n5774) );
  INV_X1 U7508 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7509 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  NAND2_X1 U7510 ( .A1(n5819), .A2(n5778), .ZN(n10118) );
  OR2_X1 U7511 ( .A1(n10118), .A2(n5557), .ZN(n5781) );
  AOI22_X1 U7512 ( .A1(n5508), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n4439), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n5780) );
  NAND2_X1 U7513 ( .A1(n4437), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7514 ( .A1(n10116), .A2(n9506), .ZN(n5783) );
  NOR2_X1 U7515 ( .A1(n10116), .A2(n9506), .ZN(n5782) );
  INV_X1 U7516 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U7517 ( .A(n5804), .B(n5799), .ZN(n7499) );
  NAND2_X1 U7518 ( .A1(n7499), .A2(n5637), .ZN(n5790) );
  NAND2_X1 U7519 ( .A1(n5811), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5788) );
  XNOR2_X1 U7520 ( .A(n5788), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U7521 ( .A1(n5815), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6919), .B2(
        n9979), .ZN(n5789) );
  XNOR2_X1 U7522 ( .A(n5819), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U7523 ( .A1(n10109), .A2(n6083), .ZN(n5795) );
  INV_X1 U7524 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10211) );
  NAND2_X1 U7525 ( .A1(n4436), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7526 ( .A1(n4438), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5791) );
  OAI211_X1 U7527 ( .C1(n6081), .C2(n10211), .A(n5792), .B(n5791), .ZN(n5793)
         );
  INV_X1 U7528 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U7529 ( .A1(n5795), .A2(n5794), .ZN(n9823) );
  NAND2_X1 U7530 ( .A1(n6067), .A2(n9823), .ZN(n5796) );
  INV_X1 U7531 ( .A(n9823), .ZN(n6066) );
  NAND2_X1 U7532 ( .A1(n10112), .A2(n6066), .ZN(n5797) );
  INV_X1 U7533 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U7534 ( .A1(n5801), .A2(SI_18_), .ZN(n5802) );
  INV_X1 U7535 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U7536 ( .A1(n5806), .A2(SI_19_), .ZN(n5807) );
  AND2_X1 U7537 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5810) );
  NAND2_X1 U7538 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5808) );
  AOI22_X1 U7539 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(n10312), .B1(n5808), .B2(
        P1_IR_REG_31__SCAN_IN), .ZN(n5809) );
  AOI22_X1 U7540 ( .A1(n5815), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9991), .B2(
        n6919), .ZN(n5816) );
  INV_X1 U7541 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9507) );
  INV_X1 U7542 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5817) );
  OAI21_X1 U7543 ( .B1(n5819), .B2(n9507), .A(n5817), .ZN(n5820) );
  NAND2_X1 U7544 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5818) );
  NAND2_X1 U7545 ( .A1(n5820), .A2(n5833), .ZN(n10088) );
  OR2_X1 U7546 ( .A1(n10088), .A2(n5557), .ZN(n5825) );
  INV_X1 U7547 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U7548 ( .A1(n4437), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7549 ( .A1(n4438), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5821) );
  OAI211_X1 U7550 ( .C1(n6081), .C2(n10207), .A(n5822), .B(n5821), .ZN(n5823)
         );
  INV_X1 U7551 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U7552 ( .A1(n5825), .A2(n5824), .ZN(n9822) );
  INV_X1 U7553 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7831) );
  INV_X1 U7554 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U7555 ( .A(n5855), .B(SI_20_), .ZN(n5829) );
  OR2_X1 U7556 ( .A1(n7876), .A2(n5830), .ZN(n5831) );
  INV_X1 U7557 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9458) );
  OR2_X2 U7558 ( .A1(n5833), .A2(n9458), .ZN(n5875) );
  NAND2_X1 U7559 ( .A1(n5833), .A2(n9458), .ZN(n5834) );
  NAND2_X1 U7560 ( .A1(n5875), .A2(n5834), .ZN(n10077) );
  INV_X1 U7561 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10275) );
  NAND2_X1 U7562 ( .A1(n5508), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7563 ( .A1(n4439), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5835) );
  OAI211_X1 U7564 ( .C1(n10275), .C2(n5576), .A(n5836), .B(n5835), .ZN(n5837)
         );
  INV_X1 U7565 ( .A(n5837), .ZN(n5838) );
  OAI21_X1 U7566 ( .B1(n10077), .B2(n5557), .A(n5838), .ZN(n9821) );
  INV_X1 U7567 ( .A(n9821), .ZN(n6071) );
  NAND2_X1 U7568 ( .A1(n5393), .A2(n6071), .ZN(n5839) );
  INV_X1 U7569 ( .A(SI_20_), .ZN(n5852) );
  OAI21_X1 U7570 ( .B1(n5854), .B2(n5852), .A(n5855), .ZN(n5841) );
  NAND2_X1 U7571 ( .A1(n5854), .A2(n5852), .ZN(n5840) );
  NAND2_X1 U7572 ( .A1(n5841), .A2(n5840), .ZN(n5844) );
  INV_X1 U7573 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5842) );
  INV_X1 U7574 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7834) );
  XNOR2_X1 U7575 ( .A(n5858), .B(SI_21_), .ZN(n5843) );
  NAND2_X1 U7576 ( .A1(n7832), .A2(n5637), .ZN(n5846) );
  OR2_X1 U7577 ( .A1(n7876), .A2(n7834), .ZN(n5845) );
  XNOR2_X1 U7578 ( .A(n5875), .B(P1_REG3_REG_21__SCAN_IN), .ZN(n10062) );
  NAND2_X1 U7579 ( .A1(n10062), .A2(n6083), .ZN(n5851) );
  INV_X1 U7580 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10195) );
  NAND2_X1 U7581 ( .A1(n4438), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U7582 ( .A1(n4436), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5847) );
  OAI211_X1 U7583 ( .C1(n10195), .C2(n6081), .A(n5848), .B(n5847), .ZN(n5849)
         );
  INV_X1 U7584 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7585 ( .A1(n5851), .A2(n5850), .ZN(n9820) );
  INV_X1 U7586 ( .A(SI_21_), .ZN(n5856) );
  AOI22_X1 U7587 ( .A1(n5852), .A2(n5855), .B1(n5858), .B2(n5856), .ZN(n5853)
         );
  INV_X1 U7588 ( .A(n5855), .ZN(n5860) );
  NAND2_X1 U7589 ( .A1(n5860), .A2(SI_20_), .ZN(n5857) );
  NAND2_X1 U7590 ( .A1(n5857), .A2(n5856), .ZN(n5862) );
  INV_X1 U7591 ( .A(n5858), .ZN(n5861) );
  AND2_X1 U7592 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5859) );
  AOI22_X1 U7593 ( .A1(n5862), .A2(n5861), .B1(n5860), .B2(n5859), .ZN(n5863)
         );
  NAND2_X1 U7594 ( .A1(n5864), .A2(n5863), .ZN(n5884) );
  INV_X1 U7595 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7837) );
  INV_X1 U7596 ( .A(SI_22_), .ZN(n5865) );
  NAND2_X1 U7597 ( .A1(n5866), .A2(n5865), .ZN(n5946) );
  INV_X1 U7598 ( .A(n5866), .ZN(n5867) );
  NAND2_X1 U7599 ( .A1(n5867), .A2(SI_22_), .ZN(n5868) );
  NAND2_X1 U7600 ( .A1(n5946), .A2(n5868), .ZN(n5885) );
  XNOR2_X1 U7601 ( .A(n5884), .B(n5885), .ZN(n7836) );
  NAND2_X1 U7602 ( .A1(n7836), .A2(n5637), .ZN(n5870) );
  OR2_X1 U7603 ( .A1(n4426), .A2(n8178), .ZN(n5869) );
  AND2_X1 U7604 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_21__SCAN_IN), 
        .ZN(n5871) );
  INV_X1 U7605 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5874) );
  INV_X1 U7606 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5873) );
  OAI21_X1 U7607 ( .B1(n5875), .B2(n5874), .A(n5873), .ZN(n5876) );
  AND2_X1 U7608 ( .A1(n5897), .A2(n5876), .ZN(n9479) );
  NAND2_X1 U7609 ( .A1(n9479), .A2(n6083), .ZN(n5881) );
  INV_X1 U7610 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U7611 ( .A1(n4437), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7612 ( .A1(n4439), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5877) );
  OAI211_X1 U7613 ( .C1(n6081), .C2(n7944), .A(n5878), .B(n5877), .ZN(n5879)
         );
  INV_X1 U7614 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U7615 ( .A1(n7934), .A2(n4486), .ZN(n5883) );
  NAND2_X1 U7616 ( .A1(n9562), .A2(n9819), .ZN(n5882) );
  NAND2_X1 U7617 ( .A1(n5883), .A2(n5882), .ZN(n10036) );
  INV_X1 U7618 ( .A(n5884), .ZN(n5887) );
  INV_X1 U7619 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5888) );
  INV_X1 U7620 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5893) );
  INV_X1 U7621 ( .A(SI_23_), .ZN(n5889) );
  NAND2_X1 U7622 ( .A1(n5890), .A2(n5889), .ZN(n5925) );
  INV_X1 U7623 ( .A(n5890), .ZN(n5891) );
  NAND2_X1 U7624 ( .A1(n5891), .A2(SI_23_), .ZN(n5923) );
  NAND2_X1 U7625 ( .A1(n7865), .A2(n5637), .ZN(n5895) );
  OR2_X1 U7626 ( .A1(n4426), .A2(n5893), .ZN(n5894) );
  INV_X1 U7627 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U7628 ( .A1(n5897), .A2(n8716), .ZN(n5898) );
  NAND2_X1 U7629 ( .A1(n5914), .A2(n5898), .ZN(n10039) );
  OR2_X1 U7630 ( .A1(n10039), .A2(n5557), .ZN(n5903) );
  INV_X1 U7631 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10189) );
  NAND2_X1 U7632 ( .A1(n4438), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7633 ( .A1(n4436), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5899) );
  OAI211_X1 U7634 ( .C1(n6081), .C2(n10189), .A(n5900), .B(n5899), .ZN(n5901)
         );
  INV_X1 U7635 ( .A(n5901), .ZN(n5902) );
  NOR2_X1 U7636 ( .A1(n10042), .A2(n9431), .ZN(n5905) );
  NAND2_X1 U7637 ( .A1(n10042), .A2(n9431), .ZN(n5904) );
  NAND2_X1 U7638 ( .A1(n5907), .A2(SI_24_), .ZN(n5926) );
  INV_X1 U7639 ( .A(n5907), .ZN(n5909) );
  INV_X1 U7640 ( .A(SI_24_), .ZN(n5908) );
  NAND2_X1 U7641 ( .A1(n5909), .A2(n5908), .ZN(n5928) );
  AND2_X1 U7642 ( .A1(n5926), .A2(n5928), .ZN(n5910) );
  NAND2_X1 U7643 ( .A1(n9308), .A2(n5637), .ZN(n5913) );
  INV_X1 U7644 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10333) );
  OR2_X1 U7645 ( .A1(n7876), .A2(n10333), .ZN(n5912) );
  INV_X1 U7646 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9432) );
  NAND2_X1 U7647 ( .A1(n5914), .A2(n9432), .ZN(n5915) );
  AND2_X1 U7648 ( .A1(n5938), .A2(n5915), .ZN(n10030) );
  NAND2_X1 U7649 ( .A1(n10030), .A2(n6083), .ZN(n5920) );
  INV_X1 U7650 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U7651 ( .A1(n4439), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U7652 ( .A1(n4437), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5916) );
  OAI211_X1 U7653 ( .C1(n6081), .C2(n10184), .A(n5917), .B(n5916), .ZN(n5918)
         );
  INV_X1 U7654 ( .A(n5918), .ZN(n5919) );
  NOR2_X1 U7655 ( .A1(n6074), .A2(n9818), .ZN(n5922) );
  NAND2_X1 U7656 ( .A1(n6074), .A2(n9818), .ZN(n5921) );
  INV_X1 U7657 ( .A(n5925), .ZN(n5927) );
  NAND2_X1 U7658 ( .A1(n5927), .A2(n5926), .ZN(n5929) );
  INV_X1 U7659 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8135) );
  INV_X1 U7660 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10329) );
  INV_X1 U7661 ( .A(SI_25_), .ZN(n5931) );
  NAND2_X1 U7662 ( .A1(n5932), .A2(n5931), .ZN(n5956) );
  INV_X1 U7663 ( .A(n5932), .ZN(n5933) );
  NAND2_X1 U7664 ( .A1(n5933), .A2(SI_25_), .ZN(n5934) );
  NAND2_X1 U7665 ( .A1(n8133), .A2(n5637), .ZN(n5937) );
  OR2_X1 U7666 ( .A1(n7876), .A2(n10329), .ZN(n5936) );
  INV_X1 U7667 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9400) );
  NAND2_X1 U7668 ( .A1(n5938), .A2(n9400), .ZN(n5939) );
  NAND2_X1 U7669 ( .A1(n5965), .A2(n5939), .ZN(n9401) );
  INV_X1 U7670 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U7671 ( .A1(n4436), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7672 ( .A1(n5508), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5940) );
  OAI211_X1 U7673 ( .C1(n5625), .C2(n7926), .A(n5941), .B(n5940), .ZN(n5942)
         );
  INV_X1 U7674 ( .A(n5942), .ZN(n5943) );
  NOR2_X1 U7675 ( .A1(n9406), .A2(n9536), .ZN(n5945) );
  INV_X1 U7676 ( .A(n9536), .ZN(n9817) );
  NAND2_X1 U7677 ( .A1(n5948), .A2(n5947), .ZN(n5955) );
  INV_X1 U7678 ( .A(n5949), .ZN(n5952) );
  INV_X1 U7679 ( .A(n5950), .ZN(n5951) );
  AOI21_X1 U7680 ( .B1(n5953), .B2(n5952), .A(n5951), .ZN(n5954) );
  NAND2_X1 U7681 ( .A1(n5955), .A2(n5954), .ZN(n5957) );
  INV_X1 U7682 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5958) );
  INV_X1 U7683 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10326) );
  INV_X1 U7684 ( .A(SI_26_), .ZN(n5959) );
  NAND2_X1 U7685 ( .A1(n5960), .A2(n5959), .ZN(n5977) );
  INV_X1 U7686 ( .A(n5960), .ZN(n5961) );
  NAND2_X1 U7687 ( .A1(n5961), .A2(SI_26_), .ZN(n5962) );
  NAND2_X1 U7688 ( .A1(n7868), .A2(n5637), .ZN(n5964) );
  OR2_X1 U7689 ( .A1(n7876), .A2(n10326), .ZN(n5963) );
  INV_X1 U7690 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9539) );
  NAND2_X1 U7691 ( .A1(n5965), .A2(n9539), .ZN(n5966) );
  NAND2_X1 U7692 ( .A1(n10015), .A2(n6083), .ZN(n5972) );
  INV_X1 U7693 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7694 ( .A1(n4437), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7695 ( .A1(n5508), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5967) );
  OAI211_X1 U7696 ( .C1(n5625), .C2(n5969), .A(n5968), .B(n5967), .ZN(n5970)
         );
  INV_X1 U7697 ( .A(n5970), .ZN(n5971) );
  NOR2_X1 U7698 ( .A1(n10016), .A2(n9816), .ZN(n5974) );
  NAND2_X1 U7699 ( .A1(n10016), .A2(n9816), .ZN(n5973) );
  NAND2_X1 U7700 ( .A1(n5976), .A2(n5975), .ZN(n5978) );
  INV_X1 U7701 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5979) );
  INV_X1 U7702 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10325) );
  INV_X1 U7703 ( .A(SI_27_), .ZN(n5980) );
  NAND2_X1 U7704 ( .A1(n5981), .A2(n5980), .ZN(n5995) );
  INV_X1 U7705 ( .A(n5981), .ZN(n5982) );
  NAND2_X1 U7706 ( .A1(n5982), .A2(SI_27_), .ZN(n5983) );
  NAND2_X1 U7707 ( .A1(n9304), .A2(n5637), .ZN(n5985) );
  OR2_X1 U7708 ( .A1(n7876), .A2(n10325), .ZN(n5984) );
  INV_X1 U7709 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8723) );
  OR2_X2 U7710 ( .A1(n5986), .A2(n8723), .ZN(n6001) );
  NAND2_X1 U7711 ( .A1(n5986), .A2(n8723), .ZN(n5987) );
  INV_X1 U7712 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7713 ( .A1(n4436), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U7714 ( .A1(n5508), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5988) );
  OAI211_X1 U7715 ( .C1(n5625), .C2(n5990), .A(n5989), .B(n5988), .ZN(n5991)
         );
  NAND2_X1 U7716 ( .A1(n10175), .A2(n9538), .ZN(n5992) );
  INV_X1 U7717 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5997) );
  INV_X1 U7718 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8006) );
  XNOR2_X1 U7719 ( .A(n6117), .B(SI_28_), .ZN(n6114) );
  NAND2_X1 U7720 ( .A1(n8004), .A2(n5637), .ZN(n5999) );
  OR2_X1 U7721 ( .A1(n4426), .A2(n8006), .ZN(n5998) );
  INV_X1 U7722 ( .A(n6001), .ZN(n6000) );
  NAND2_X1 U7723 ( .A1(n6000), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n6078) );
  INV_X1 U7724 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U7725 ( .A1(n6001), .A2(n9351), .ZN(n6002) );
  INV_X1 U7726 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7727 ( .A1(n4438), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7728 ( .A1(n4437), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6003) );
  OAI211_X1 U7729 ( .C1(n6005), .C2(n6081), .A(n6004), .B(n6003), .ZN(n6006)
         );
  INV_X1 U7730 ( .A(n6006), .ZN(n6007) );
  AND2_X2 U7731 ( .A1(n6008), .A2(n6007), .ZN(n7892) );
  NAND2_X1 U7732 ( .A1(n9347), .A2(n7892), .ZN(n9648) );
  INV_X1 U7733 ( .A(n9694), .ZN(n6009) );
  NAND2_X1 U7734 ( .A1(n6010), .A2(n9694), .ZN(n6011) );
  NAND2_X1 U7735 ( .A1(n10390), .A2(n9991), .ZN(n7060) );
  NAND2_X1 U7736 ( .A1(n10331), .A2(P1_B_REG_SCAN_IN), .ZN(n6026) );
  INV_X1 U7737 ( .A(n6022), .ZN(n6023) );
  NAND2_X1 U7738 ( .A1(n6023), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6025) );
  MUX2_X1 U7739 ( .A(P1_B_REG_SCAN_IN), .B(n6026), .S(n10336), .Z(n6031) );
  INV_X1 U7740 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6028) );
  INV_X1 U7741 ( .A(n10328), .ZN(n6030) );
  INV_X1 U7742 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U7743 ( .A1(n7056), .A2(n6918), .ZN(n6041) );
  NAND2_X1 U7744 ( .A1(n10328), .A2(n10331), .ZN(n7057) );
  NOR4_X1 U7745 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n8731) );
  NOR2_X1 U7746 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6034) );
  NOR4_X1 U7747 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6033) );
  NOR4_X1 U7748 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6032) );
  AND4_X1 U7749 ( .A1(n8731), .A2(n6034), .A3(n6033), .A4(n6032), .ZN(n6040)
         );
  NOR4_X1 U7750 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6038) );
  NOR4_X1 U7751 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6037) );
  NOR4_X1 U7752 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n6036) );
  NOR4_X1 U7753 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6035) );
  AND4_X1 U7754 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n6039)
         );
  NAND2_X1 U7755 ( .A1(n6040), .A2(n6039), .ZN(n7053) );
  AOI22_X1 U7756 ( .A1(n6041), .A2(n7057), .B1(n7056), .B2(n7053), .ZN(n6042)
         );
  AND2_X1 U7757 ( .A1(n7060), .A2(n6042), .ZN(n6047) );
  NAND2_X1 U7758 ( .A1(n6043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6045) );
  INV_X1 U7759 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6044) );
  AND2_X1 U7760 ( .A1(n7205), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6046) );
  INV_X1 U7761 ( .A(n7066), .ZN(n9796) );
  INV_X1 U7762 ( .A(n7063), .ZN(n6076) );
  NAND2_X1 U7763 ( .A1(n9735), .A2(n9787), .ZN(n7204) );
  INV_X1 U7764 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U7765 ( .A1(n7056), .A2(n10408), .ZN(n6049) );
  NAND2_X1 U7766 ( .A1(n10328), .A2(n10336), .ZN(n6048) );
  INV_X1 U7767 ( .A(n7606), .ZN(n7090) );
  NOR2_X1 U7768 ( .A1(n7066), .A2(n9991), .ZN(n7064) );
  NAND2_X1 U7769 ( .A1(n9735), .A2(n9806), .ZN(n7612) );
  OAI211_X1 U7770 ( .C1(n7064), .C2(n9806), .A(n7612), .B(n10254), .ZN(n10410)
         );
  INV_X2 U7771 ( .A(n7141), .ZN(n10253) );
  NOR2_X1 U7772 ( .A1(n9840), .A2(n10253), .ZN(n7718) );
  NAND2_X1 U7773 ( .A1(n7720), .A2(n6051), .ZN(n7704) );
  OR2_X1 U7774 ( .A1(n5482), .A2(n10421), .ZN(n6052) );
  NAND2_X1 U7775 ( .A1(n9584), .A2(n7666), .ZN(n9582) );
  NAND2_X1 U7776 ( .A1(n9582), .A2(n9583), .ZN(n7780) );
  NAND2_X1 U7777 ( .A1(n7780), .A2(n9596), .ZN(n6055) );
  NAND2_X1 U7778 ( .A1(n6055), .A2(n9591), .ZN(n9677) );
  AND2_X1 U7779 ( .A1(n9677), .A2(n9577), .ZN(n6056) );
  NAND2_X1 U7780 ( .A1(n9678), .A2(n7643), .ZN(n6058) );
  INV_X1 U7781 ( .A(n9590), .ZN(n6059) );
  NOR2_X1 U7782 ( .A1(n7839), .A2(n6059), .ZN(n6060) );
  INV_X1 U7783 ( .A(n9756), .ZN(n9609) );
  NAND2_X1 U7784 ( .A1(n10230), .A2(n8064), .ZN(n9613) );
  NAND2_X1 U7785 ( .A1(n10225), .A2(n6061), .ZN(n9621) );
  NAND2_X1 U7786 ( .A1(n9616), .A2(n9621), .ZN(n9671) );
  INV_X1 U7787 ( .A(n10148), .ZN(n6062) );
  NOR2_X1 U7788 ( .A1(n9671), .A2(n6062), .ZN(n6063) );
  INV_X1 U7789 ( .A(n10135), .ZN(n6064) );
  NAND2_X1 U7790 ( .A1(n10215), .A2(n9506), .ZN(n9624) );
  INV_X1 U7791 ( .A(n9619), .ZN(n10124) );
  NOR2_X1 U7792 ( .A1(n10123), .A2(n10124), .ZN(n6065) );
  OR2_X1 U7793 ( .A1(n6067), .A2(n6066), .ZN(n9768) );
  NAND2_X1 U7794 ( .A1(n6067), .A2(n6066), .ZN(n9625) );
  INV_X1 U7795 ( .A(n10099), .ZN(n6068) );
  INV_X1 U7796 ( .A(n9822), .ZN(n6070) );
  NAND2_X1 U7797 ( .A1(n10197), .A2(n6071), .ZN(n9628) );
  INV_X1 U7798 ( .A(n9820), .ZN(n7939) );
  XNOR2_X1 U7799 ( .A(n10194), .B(n7939), .ZN(n10058) );
  NAND2_X1 U7800 ( .A1(n10194), .A2(n7939), .ZN(n9636) );
  NAND2_X1 U7801 ( .A1(n9636), .A2(n9628), .ZN(n9633) );
  OR2_X1 U7802 ( .A1(n10194), .A2(n7939), .ZN(n9700) );
  NAND2_X1 U7803 ( .A1(n9633), .A2(n9700), .ZN(n9711) );
  INV_X1 U7804 ( .A(n9819), .ZN(n9561) );
  OR2_X1 U7805 ( .A1(n10188), .A2(n9431), .ZN(n9641) );
  OR2_X1 U7806 ( .A1(n9562), .A2(n9561), .ZN(n10045) );
  NAND2_X1 U7807 ( .A1(n10047), .A2(n10045), .ZN(n6073) );
  INV_X1 U7808 ( .A(n9818), .ZN(n8122) );
  NAND2_X1 U7809 ( .A1(n6074), .A2(n8122), .ZN(n9713) );
  NAND2_X1 U7810 ( .A1(n9705), .A2(n9713), .ZN(n10025) );
  NAND2_X1 U7811 ( .A1(n7920), .A2(n9536), .ZN(n9653) );
  INV_X1 U7812 ( .A(n9655), .ZN(n9645) );
  INV_X1 U7813 ( .A(n9816), .ZN(n9654) );
  AND2_X1 U7814 ( .A1(n10016), .A2(n9654), .ZN(n9714) );
  INV_X1 U7815 ( .A(n9996), .ZN(n10005) );
  INV_X1 U7816 ( .A(n6075), .ZN(n9647) );
  XNOR2_X1 U7817 ( .A(n7891), .B(n9694), .ZN(n6086) );
  OR2_X1 U7818 ( .A1(n7066), .A2(n9800), .ZN(n6077) );
  NAND2_X1 U7819 ( .A1(n6076), .A2(n4613), .ZN(n9798) );
  INV_X1 U7820 ( .A(n6078), .ZN(n7904) );
  INV_X1 U7821 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7912) );
  NAND2_X1 U7822 ( .A1(n4439), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7823 ( .A1(n4436), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6079) );
  OAI211_X1 U7824 ( .C1(n6081), .C2(n7912), .A(n6080), .B(n6079), .ZN(n6082)
         );
  AOI21_X1 U7825 ( .B1(n7904), .B2(n6083), .A(n6082), .ZN(n7885) );
  INV_X1 U7826 ( .A(n9551), .ZN(n9537) );
  OAI22_X1 U7827 ( .A1(n7885), .A2(n9537), .B1(n9538), .B2(n9535), .ZN(n9356)
         );
  NOR2_X2 U7828 ( .A1(n7715), .A2(n5481), .ZN(n7699) );
  NAND2_X1 U7829 ( .A1(n7699), .A2(n10426), .ZN(n7638) );
  INV_X1 U7830 ( .A(n8039), .ZN(n10469) );
  AND2_X2 U7831 ( .A1(n10351), .A2(n10469), .ZN(n10349) );
  NAND2_X1 U7832 ( .A1(n10105), .A2(n10112), .ZN(n10106) );
  NOR2_X2 U7833 ( .A1(n10106), .A2(n10206), .ZN(n6087) );
  INV_X1 U7834 ( .A(n6087), .ZN(n10086) );
  INV_X1 U7835 ( .A(n10194), .ZN(n10059) );
  INV_X1 U7836 ( .A(n9562), .ZN(n8118) );
  OR2_X2 U7837 ( .A1(n10037), .A2(n6074), .ZN(n10028) );
  NOR2_X4 U7838 ( .A1(n10028), .A2(n7920), .ZN(n10014) );
  NAND2_X1 U7839 ( .A1(n10000), .A2(n9347), .ZN(n6088) );
  NAND2_X1 U7840 ( .A1(n6088), .A2(n10390), .ZN(n6089) );
  INV_X1 U7841 ( .A(n9347), .ZN(n9353) );
  OR2_X1 U7842 ( .A1(n6089), .A2(n7899), .ZN(n7990) );
  NAND2_X1 U7843 ( .A1(n7986), .A2(n5418), .ZN(n6097) );
  INV_X1 U7844 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6092) );
  INV_X1 U7845 ( .A(n7992), .ZN(n6099) );
  NOR2_X2 U7846 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n6379) );
  NAND4_X1 U7847 ( .A1(n8661), .A2(n6104), .A3(n6103), .A4(n6404), .ZN(n6105)
         );
  NAND2_X1 U7848 ( .A1(n6182), .A2(n6137), .ZN(n6419) );
  OAI21_X2 U7849 ( .B1(n6445), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7850 ( .A1(n6112), .A2(n6113), .ZN(n6111) );
  NAND2_X1 U7851 ( .A1(n7829), .A2(n6772), .ZN(n10516) );
  INV_X1 U7852 ( .A(n10516), .ZN(n7360) );
  NAND2_X1 U7853 ( .A1(n6115), .A2(n6114), .ZN(n6119) );
  INV_X1 U7854 ( .A(SI_28_), .ZN(n6116) );
  NAND2_X1 U7855 ( .A1(n6117), .A2(n6116), .ZN(n6118) );
  INV_X1 U7856 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6120) );
  INV_X1 U7857 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10323) );
  INV_X1 U7858 ( .A(SI_29_), .ZN(n8701) );
  INV_X1 U7859 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10320) );
  INV_X1 U7860 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n6124) );
  MUX2_X1 U7861 ( .A(n10320), .B(n6124), .S(n4431), .Z(n6126) );
  INV_X1 U7862 ( .A(SI_30_), .ZN(n6125) );
  NAND2_X1 U7863 ( .A1(n6126), .A2(n6125), .ZN(n6129) );
  INV_X1 U7864 ( .A(n6126), .ZN(n6127) );
  NAND2_X1 U7865 ( .A1(n6127), .A2(SI_30_), .ZN(n6128) );
  NAND2_X1 U7866 ( .A1(n6129), .A2(n6128), .ZN(n6551) );
  MUX2_X1 U7867 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4431), .Z(n6130) );
  INV_X1 U7868 ( .A(SI_31_), .ZN(n8548) );
  XNOR2_X1 U7869 ( .A(n6130), .B(n8548), .ZN(n6131) );
  NOR2_X1 U7870 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n6135) );
  NOR2_X1 U7871 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n6134) );
  NAND4_X1 U7872 ( .A1(n8578), .A2(n8573), .A3(n8572), .A4(n6138), .ZN(n6139)
         );
  NAND2_X1 U7873 ( .A1(n9291), .A2(n6553), .ZN(n6144) );
  AND2_X4 U7874 ( .A1(n6244), .A2(n4956), .ZN(n6554) );
  NAND2_X1 U7875 ( .A1(n6554), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6143) );
  INV_X1 U7876 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6153) );
  INV_X1 U7877 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6154) );
  INV_X1 U7878 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6155) );
  INV_X1 U7879 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6156) );
  INV_X1 U7880 ( .A(n8127), .ZN(n6163) );
  INV_X1 U7881 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7882 ( .A1(n6163), .A2(n6534), .ZN(n6562) );
  INV_X1 U7883 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U7884 ( .A1(n6545), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6167) );
  INV_X1 U7885 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9098) );
  OR2_X1 U7886 ( .A1(n4430), .A2(n9098), .ZN(n6166) );
  OAI211_X1 U7887 ( .C1(n8811), .C2(n6428), .A(n6167), .B(n6166), .ZN(n6168)
         );
  INV_X1 U7888 ( .A(n6168), .ZN(n6169) );
  NOR2_X1 U7889 ( .A1(n6575), .A2(n6685), .ZN(n6574) );
  NAND2_X1 U7890 ( .A1(n7868), .A2(n6472), .ZN(n6171) );
  NAND2_X1 U7891 ( .A1(n6554), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7892 ( .A1(n6190), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7893 ( .A1(n6522), .A2(n6172), .ZN(n8837) );
  NAND2_X1 U7894 ( .A1(n8837), .A2(n6534), .ZN(n6177) );
  INV_X1 U7895 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U7896 ( .A1(n6545), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7897 ( .A1(n6535), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7898 ( .C1(n8836), .C2(n6453), .A(n6174), .B(n6173), .ZN(n6175)
         );
  INV_X1 U7899 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U7900 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  NAND2_X1 U7901 ( .A1(n6183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7902 ( .A(n6184), .B(P2_IR_REG_31__SCAN_IN), .S(n8578), .Z(n6186)
         );
  NAND2_X1 U7903 ( .A1(n6185), .A2(n8578), .ZN(n6662) );
  NAND2_X1 U7904 ( .A1(n6186), .A2(n6662), .ZN(n7838) );
  NAND2_X2 U7905 ( .A1(n4434), .A2(n6780), .ZN(n6886) );
  NOR3_X1 U7906 ( .A1(n9198), .A2(n6838), .A3(n6886), .ZN(n6513) );
  NAND2_X1 U7907 ( .A1(n8133), .A2(n6472), .ZN(n6188) );
  NAND2_X1 U7908 ( .A1(n6554), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7909 ( .A1(n6197), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7910 ( .A1(n6190), .A2(n6189), .ZN(n8843) );
  NAND2_X1 U7911 ( .A1(n8843), .A2(n6534), .ZN(n6195) );
  INV_X1 U7912 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U7913 ( .A1(n6535), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6192) );
  INV_X1 U7914 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9203) );
  OR2_X1 U7915 ( .A1(n6489), .A2(n9203), .ZN(n6191) );
  OAI211_X1 U7916 ( .C1(n8847), .C2(n6453), .A(n6192), .B(n6191), .ZN(n6193)
         );
  INV_X1 U7917 ( .A(n6193), .ZN(n6194) );
  INV_X1 U7918 ( .A(n6648), .ZN(n6204) );
  NAND2_X1 U7919 ( .A1(n6501), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6196) );
  NAND2_X1 U7920 ( .A1(n6197), .A2(n6196), .ZN(n8860) );
  NAND2_X1 U7921 ( .A1(n8860), .A2(n6534), .ZN(n6202) );
  INV_X1 U7922 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U7923 ( .A1(n6545), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6199) );
  INV_X1 U7924 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9113) );
  OR2_X1 U7925 ( .A1(n4429), .A2(n9113), .ZN(n6198) );
  OAI211_X1 U7926 ( .C1(n6453), .C2(n8713), .A(n6199), .B(n6198), .ZN(n6200)
         );
  INV_X1 U7927 ( .A(n6200), .ZN(n6201) );
  INV_X1 U7928 ( .A(n6645), .ZN(n6203) );
  NAND2_X1 U7929 ( .A1(n9204), .A2(n8314), .ZN(n6647) );
  NAND2_X1 U7930 ( .A1(n6647), .A2(n4428), .ZN(n6512) );
  NOR4_X1 U7931 ( .A1(n6513), .A2(n6204), .A3(n6203), .A4(n6512), .ZN(n6519)
         );
  NAND2_X1 U7932 ( .A1(n7093), .A2(n6472), .ZN(n6210) );
  OAI21_X1 U7933 ( .B1(P2_IR_REG_10__SCAN_IN), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7934 ( .A1(n6312), .A2(n6207), .ZN(n6217) );
  OAI21_X1 U7935 ( .B1(n6217), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6208) );
  AOI22_X1 U7936 ( .A1(n8408), .A2(n4776), .B1(n6554), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6209) );
  NAND2_X1 U7937 ( .A1(n6535), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6215) );
  INV_X1 U7938 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9271) );
  OR2_X1 U7939 ( .A1(n6489), .A2(n9271), .ZN(n6214) );
  NAND2_X1 U7940 ( .A1(n6221), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6211) );
  AND2_X1 U7941 ( .A1(n6385), .A2(n6211), .ZN(n9012) );
  OR2_X1 U7942 ( .A1(n4768), .A2(n9012), .ZN(n6213) );
  INV_X1 U7943 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8407) );
  OR2_X1 U7944 ( .A1(n6453), .A2(n8407), .ZN(n6212) );
  NAND4_X1 U7945 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n9024)
         );
  INV_X1 U7946 ( .A(n6621), .ZN(n6226) );
  NAND2_X1 U7947 ( .A1(n6947), .A2(n6472), .ZN(n6219) );
  XNOR2_X1 U7948 ( .A(n6217), .B(n6216), .ZN(n8383) );
  AOI22_X1 U7949 ( .A1(n6554), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n8383), .B2(
        n4776), .ZN(n6218) );
  NAND2_X2 U7950 ( .A1(n6219), .A2(n6218), .ZN(n9276) );
  NAND2_X1 U7951 ( .A1(n6535), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6225) );
  INV_X1 U7952 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9275) );
  OR2_X1 U7953 ( .A1(n6489), .A2(n9275), .ZN(n6224) );
  NAND2_X1 U7954 ( .A1(n6356), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6220) );
  AND2_X1 U7955 ( .A1(n6221), .A2(n6220), .ZN(n9027) );
  OR2_X1 U7956 ( .A1(n4768), .A2(n9027), .ZN(n6223) );
  INV_X1 U7957 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n9026) );
  OR2_X1 U7958 ( .A1(n6453), .A2(n9026), .ZN(n6222) );
  NAND4_X1 U7959 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n9046)
         );
  INV_X1 U7960 ( .A(n9046), .ZN(n9009) );
  NAND2_X1 U7961 ( .A1(n9276), .A2(n9009), .ZN(n6619) );
  NAND2_X1 U7962 ( .A1(n9155), .A2(n8291), .ZN(n6370) );
  OAI21_X1 U7963 ( .B1(n6226), .B2(n6619), .A(n6370), .ZN(n6376) );
  INV_X1 U7964 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7962) );
  OR2_X1 U7965 ( .A1(n6428), .A2(n7962), .ZN(n6230) );
  INV_X1 U7966 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U7967 ( .A1(n6287), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6228) );
  INV_X1 U7968 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U7969 ( .A1(n6554), .A2(n6910), .ZN(n6234) );
  NAND2_X1 U7970 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6231) );
  NAND2_X1 U7971 ( .A1(n6454), .A2(n7317), .ZN(n6232) );
  OR2_X1 U7972 ( .A1(n6428), .A2(n7179), .ZN(n6238) );
  INV_X1 U7973 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7159) );
  OR2_X1 U7974 ( .A1(n4430), .A2(n7159), .ZN(n6237) );
  NAND2_X1 U7975 ( .A1(n6287), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6236) );
  INV_X1 U7976 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7340) );
  OR2_X1 U7977 ( .A1(n6275), .A2(n7340), .ZN(n6235) );
  NAND4_X1 U7978 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n6239)
         );
  NAND2_X1 U7979 ( .A1(n4431), .A2(SI_0_), .ZN(n6241) );
  INV_X1 U7980 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7981 ( .A1(n6241), .A2(n6240), .ZN(n6243) );
  AND2_X1 U7982 ( .A1(n6243), .A2(n6242), .ZN(n9312) );
  INV_X1 U7983 ( .A(n7955), .ZN(n6599) );
  INV_X1 U7984 ( .A(n7344), .ZN(n7212) );
  OAI22_X1 U7985 ( .A1(n6599), .A2(n4435), .B1(n6780), .B2(n6582), .ZN(n6259)
         );
  NAND2_X1 U7986 ( .A1(n6535), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6250) );
  INV_X1 U7987 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6246) );
  INV_X1 U7988 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6247) );
  OR2_X1 U7989 ( .A1(n6428), .A2(n6247), .ZN(n6248) );
  NAND2_X1 U7990 ( .A1(n6554), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6256) );
  INV_X1 U7991 ( .A(n6899), .ZN(n6251) );
  NAND2_X1 U7992 ( .A1(n6553), .A2(n6251), .ZN(n6255) );
  NAND2_X1 U7993 ( .A1(n6454), .A2(n7175), .ZN(n6254) );
  INV_X1 U7994 ( .A(n6270), .ZN(n6269) );
  INV_X1 U7995 ( .A(n6260), .ZN(n6268) );
  NAND2_X1 U7996 ( .A1(n6535), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6265) );
  OR2_X1 U7997 ( .A1(n6275), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6264) );
  INV_X1 U7998 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10496) );
  INV_X1 U7999 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6261) );
  OR2_X1 U8000 ( .A1(n6489), .A2(n6261), .ZN(n6262) );
  NAND2_X1 U8001 ( .A1(n6554), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U8002 ( .A1(n6454), .A2(n10506), .ZN(n6266) );
  OAI211_X1 U8003 ( .C1(n6306), .C2(n6909), .A(n6267), .B(n6266), .ZN(n7369)
         );
  NAND2_X1 U8004 ( .A1(n7375), .A2(n7369), .ZN(n6603) );
  NAND2_X1 U8005 ( .A1(n7958), .A2(n5142), .ZN(n6601) );
  INV_X1 U8006 ( .A(n7369), .ZN(n10533) );
  OAI211_X1 U8007 ( .C1(n7958), .C2(n5142), .A(n6271), .B(n6581), .ZN(n6272)
         );
  MUX2_X1 U8008 ( .A(n6273), .B(n6272), .S(n4428), .Z(n6283) );
  NAND2_X1 U8009 ( .A1(n6535), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U8010 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6274) );
  AND2_X1 U8011 ( .A1(n6284), .A2(n6274), .ZN(n7419) );
  OR2_X1 U8012 ( .A1(n6275), .A2(n7419), .ZN(n6277) );
  INV_X1 U8013 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7418) );
  OR2_X1 U8014 ( .A1(n6453), .A2(n7418), .ZN(n6276) );
  NAND2_X1 U8015 ( .A1(n6554), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6282) );
  NAND2_X1 U8016 ( .A1(n6279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6280) );
  NAND2_X1 U8017 ( .A1(n6454), .A2(n7242), .ZN(n6281) );
  NAND2_X1 U8018 ( .A1(n6809), .A2(n7421), .ZN(n6605) );
  INV_X1 U8019 ( .A(n6809), .ZN(n7367) );
  INV_X1 U8020 ( .A(n7421), .ZN(n10538) );
  NAND2_X1 U8021 ( .A1(n7367), .A2(n10538), .ZN(n6296) );
  NAND2_X1 U8022 ( .A1(n6605), .A2(n6296), .ZN(n7412) );
  NAND2_X1 U8023 ( .A1(n6283), .A2(n7415), .ZN(n6372) );
  INV_X1 U8024 ( .A(n6603), .ZN(n6297) );
  NAND2_X1 U8025 ( .A1(n6284), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6285) );
  AND2_X1 U8026 ( .A1(n6298), .A2(n6285), .ZN(n7495) );
  OR2_X1 U8027 ( .A1(n6275), .A2(n7495), .ZN(n6291) );
  INV_X1 U8028 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7270) );
  OR2_X1 U8029 ( .A1(n4430), .A2(n7270), .ZN(n6290) );
  INV_X1 U8030 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7494) );
  OR2_X1 U8031 ( .A1(n6453), .A2(n7494), .ZN(n6289) );
  NAND2_X1 U8032 ( .A1(n6287), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U8033 ( .A1(n6554), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U8034 ( .A1(n6292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U8035 ( .A1(n6454), .A2(n7269), .ZN(n6294) );
  INV_X1 U8036 ( .A(n10542), .ZN(n6808) );
  NAND2_X1 U8037 ( .A1(n8338), .A2(n6808), .ZN(n6583) );
  OAI211_X1 U8038 ( .C1(n6372), .C2(n6297), .A(n6583), .B(n6296), .ZN(n6309)
         );
  NAND2_X1 U8039 ( .A1(n6535), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6303) );
  INV_X1 U8040 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7433) );
  OR2_X1 U8041 ( .A1(n6489), .A2(n7433), .ZN(n6302) );
  NAND2_X1 U8042 ( .A1(n6298), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6299) );
  AND2_X1 U8043 ( .A1(n6335), .A2(n6299), .ZN(n7456) );
  OR2_X1 U8044 ( .A1(n6275), .A2(n7456), .ZN(n6301) );
  INV_X1 U8045 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7440) );
  OR2_X1 U8046 ( .A1(n6453), .A2(n7440), .ZN(n6300) );
  NAND2_X1 U8047 ( .A1(n6304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6305) );
  AOI22_X1 U8048 ( .A1(n6554), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7570), .B2(
        n6454), .ZN(n6308) );
  OR2_X1 U8049 ( .A1(n6906), .A2(n6306), .ZN(n6307) );
  NAND2_X1 U8050 ( .A1(n6308), .A2(n6307), .ZN(n7453) );
  NAND2_X1 U8051 ( .A1(n7596), .A2(n7453), .ZN(n6588) );
  NOR2_X1 U8052 ( .A1(n8338), .A2(n6808), .ZN(n6610) );
  INV_X1 U8053 ( .A(n6610), .ZN(n7430) );
  NAND3_X1 U8054 ( .A1(n6309), .A2(n6588), .A3(n7430), .ZN(n6349) );
  NAND2_X1 U8055 ( .A1(n6930), .A2(n6472), .ZN(n6315) );
  INV_X1 U8056 ( .A(n6312), .ZN(n6310) );
  NAND2_X1 U8057 ( .A1(n6310), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6313) );
  INV_X1 U8058 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U8059 ( .A1(n6312), .A2(n6311), .ZN(n6350) );
  AOI22_X1 U8060 ( .A1(n6554), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n8344), .B2(
        n4776), .ZN(n6314) );
  NAND2_X1 U8061 ( .A1(n6315), .A2(n6314), .ZN(n7681) );
  NAND2_X1 U8062 ( .A1(n6557), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6320) );
  INV_X1 U8063 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9287) );
  OR2_X1 U8064 ( .A1(n6489), .A2(n9287), .ZN(n6319) );
  INV_X1 U8065 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9170) );
  OR2_X1 U8066 ( .A1(n4430), .A2(n9170), .ZN(n6318) );
  NAND2_X1 U8067 ( .A1(n6327), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6316) );
  AND2_X1 U8068 ( .A1(n6354), .A2(n6316), .ZN(n9057) );
  OR2_X1 U8069 ( .A1(n4768), .A2(n9057), .ZN(n6317) );
  INV_X1 U8070 ( .A(n9034), .ZN(n6333) );
  NAND2_X1 U8071 ( .A1(n6912), .A2(n6472), .ZN(n6324) );
  NAND2_X1 U8072 ( .A1(n6321), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6322) );
  AOI22_X1 U8073 ( .A1(n6554), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7574), .B2(
        n4776), .ZN(n6323) );
  NAND2_X1 U8074 ( .A1(n6535), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6331) );
  INV_X1 U8075 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6325) );
  OR2_X1 U8076 ( .A1(n6489), .A2(n6325), .ZN(n6330) );
  NAND2_X1 U8077 ( .A1(n6337), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6326) );
  AND2_X1 U8078 ( .A1(n6327), .A2(n6326), .ZN(n9077) );
  OR2_X1 U8079 ( .A1(n6275), .A2(n9077), .ZN(n6329) );
  INV_X1 U8080 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9075) );
  OR2_X1 U8081 ( .A1(n6453), .A2(n9075), .ZN(n6328) );
  INV_X1 U8082 ( .A(n9032), .ZN(n6332) );
  NOR3_X1 U8083 ( .A1(n6333), .A2(n6332), .A3(n6886), .ZN(n6347) );
  NAND2_X1 U8084 ( .A1(n7681), .A2(n7655), .ZN(n6614) );
  NAND2_X1 U8085 ( .A1(n9076), .A2(n7595), .ZN(n6613) );
  AND2_X1 U8086 ( .A1(n6613), .A2(n6886), .ZN(n6334) );
  AND2_X1 U8087 ( .A1(n6334), .A2(n6614), .ZN(n6364) );
  NAND2_X1 U8088 ( .A1(n6545), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6342) );
  INV_X1 U8089 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7691) );
  OR2_X1 U8090 ( .A1(n4430), .A2(n7691), .ZN(n6341) );
  NAND2_X1 U8091 ( .A1(n6335), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6336) );
  AND2_X1 U8092 ( .A1(n6337), .A2(n6336), .ZN(n9088) );
  OR2_X1 U8093 ( .A1(n6275), .A2(n9088), .ZN(n6340) );
  INV_X1 U8094 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6338) );
  OR2_X1 U8095 ( .A1(n6453), .A2(n6338), .ZN(n6339) );
  NAND2_X1 U8096 ( .A1(n6900), .A2(n6472), .ZN(n6346) );
  NAND2_X1 U8097 ( .A1(n6343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  AOI22_X1 U8098 ( .A1(n6554), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7573), .B2(
        n6454), .ZN(n6345) );
  NAND2_X1 U8099 ( .A1(n6346), .A2(n6345), .ZN(n7692) );
  NAND2_X1 U8100 ( .A1(n7656), .A2(n7692), .ZN(n6361) );
  INV_X1 U8101 ( .A(n7692), .ZN(n9089) );
  NAND2_X1 U8102 ( .A1(n9089), .A2(n8336), .ZN(n6612) );
  OAI21_X1 U8103 ( .B1(n6347), .B2(n6364), .A(n7593), .ZN(n6373) );
  INV_X1 U8104 ( .A(n6373), .ZN(n6348) );
  INV_X1 U8105 ( .A(n7453), .ZN(n7441) );
  NAND2_X1 U8106 ( .A1(n8337), .A2(n7441), .ZN(n6609) );
  NAND3_X1 U8107 ( .A1(n6349), .A2(n6348), .A3(n6609), .ZN(n6369) );
  NAND2_X1 U8108 ( .A1(n6934), .A2(n6472), .ZN(n6353) );
  NAND2_X1 U8109 ( .A1(n6350), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6351) );
  AOI22_X1 U8110 ( .A1(n8367), .A2(n4776), .B1(n6554), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8111 ( .A1(n6545), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6360) );
  INV_X1 U8112 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9165) );
  OR2_X1 U8113 ( .A1(n4430), .A2(n9165), .ZN(n6359) );
  NAND2_X1 U8114 ( .A1(n6354), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6355) );
  AND2_X1 U8115 ( .A1(n6356), .A2(n6355), .ZN(n9036) );
  OR2_X1 U8116 ( .A1(n4768), .A2(n9036), .ZN(n6358) );
  INV_X1 U8117 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8366) );
  OR2_X1 U8118 ( .A1(n6453), .A2(n8366), .ZN(n6357) );
  NAND2_X1 U8119 ( .A1(n8198), .A2(n7685), .ZN(n9018) );
  NAND2_X1 U8120 ( .A1(n6613), .A2(n6361), .ZN(n6362) );
  NAND3_X1 U8121 ( .A1(n9034), .A2(n9032), .A3(n6362), .ZN(n6363) );
  NAND3_X1 U8122 ( .A1(n9018), .A2(n6614), .A3(n6363), .ZN(n6368) );
  INV_X1 U8123 ( .A(n6364), .ZN(n6366) );
  AND2_X1 U8124 ( .A1(n9032), .A2(n6612), .ZN(n6365) );
  OAI211_X1 U8125 ( .C1(n6366), .C2(n6365), .A(n6615), .B(n9034), .ZN(n6367)
         );
  INV_X1 U8126 ( .A(n6581), .ZN(n6371) );
  OAI211_X1 U8127 ( .C1(n6372), .C2(n6371), .A(n6605), .B(n7430), .ZN(n6374)
         );
  AND2_X1 U8128 ( .A1(n6583), .A2(n6609), .ZN(n6607) );
  INV_X1 U8129 ( .A(n6588), .ZN(n6608) );
  NAND2_X1 U8130 ( .A1(n7096), .A2(n6472), .ZN(n6384) );
  INV_X1 U8131 ( .A(n6377), .ZN(n6381) );
  NOR2_X1 U8132 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n6378) );
  AND2_X1 U8133 ( .A1(n6379), .A2(n6378), .ZN(n6380) );
  NAND2_X1 U8134 ( .A1(n6381), .A2(n6380), .ZN(n6392) );
  NAND2_X1 U8135 ( .A1(n6392), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6382) );
  XNOR2_X1 U8136 ( .A(n6382), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8424) );
  AOI22_X1 U8137 ( .A1(n8424), .A2(n4776), .B1(n6554), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6383) );
  NAND2_X1 U8138 ( .A1(n6535), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6390) );
  INV_X1 U8139 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9265) );
  OR2_X1 U8140 ( .A1(n6489), .A2(n9265), .ZN(n6389) );
  NAND2_X1 U8141 ( .A1(n6385), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6386) );
  AND2_X1 U8142 ( .A1(n6398), .A2(n6386), .ZN(n8994) );
  OR2_X1 U8143 ( .A1(n4768), .A2(n8994), .ZN(n6388) );
  INV_X1 U8144 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8410) );
  OR2_X1 U8145 ( .A1(n6453), .A2(n8410), .ZN(n6387) );
  NAND4_X1 U8146 ( .A1(n6390), .A2(n6389), .A3(n6388), .A4(n6387), .ZN(n8975)
         );
  OR2_X1 U8147 ( .A1(n9266), .A2(n8975), .ZN(n6822) );
  NAND2_X1 U8148 ( .A1(n9266), .A2(n8975), .ZN(n6823) );
  NAND2_X1 U8149 ( .A1(n9266), .A2(n6722), .ZN(n6622) );
  OR2_X1 U8150 ( .A1(n9266), .A2(n6722), .ZN(n6623) );
  MUX2_X1 U8151 ( .A(n6622), .B(n6623), .S(n4428), .Z(n6391) );
  NAND2_X1 U8152 ( .A1(n7132), .A2(n6472), .ZN(n6397) );
  INV_X1 U8153 ( .A(n6392), .ZN(n6394) );
  INV_X1 U8154 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6393) );
  NAND2_X1 U8155 ( .A1(n6394), .A2(n6393), .ZN(n6395) );
  NAND2_X1 U8156 ( .A1(n6395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6405) );
  AOI22_X1 U8157 ( .A1(n8448), .A2(n4776), .B1(n6554), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6396) );
  NAND2_X1 U8158 ( .A1(n6398), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U8159 ( .A1(n6410), .A2(n6399), .ZN(n8979) );
  NAND2_X1 U8160 ( .A1(n6534), .A2(n8979), .ZN(n6403) );
  INV_X1 U8161 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9259) );
  OR2_X1 U8162 ( .A1(n6489), .A2(n9259), .ZN(n6402) );
  INV_X1 U8163 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9148) );
  OR2_X1 U8164 ( .A1(n4430), .A2(n9148), .ZN(n6401) );
  INV_X1 U8165 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8985) );
  OR2_X1 U8166 ( .A1(n6453), .A2(n8985), .ZN(n6400) );
  NAND4_X1 U8167 ( .A1(n6403), .A2(n6402), .A3(n6401), .A4(n6400), .ZN(n8991)
         );
  INV_X1 U8168 ( .A(n8991), .ZN(n6724) );
  OR2_X1 U8169 ( .A1(n9260), .A2(n6724), .ZN(n6626) );
  NAND2_X1 U8170 ( .A1(n9260), .A2(n6724), .ZN(n6625) );
  NAND2_X1 U8171 ( .A1(n7301), .A2(n6472), .ZN(n6409) );
  NAND2_X1 U8172 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  NAND2_X1 U8173 ( .A1(n6406), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6407) );
  XNOR2_X1 U8174 ( .A(n6407), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8463) );
  AOI22_X1 U8175 ( .A1(n8463), .A2(n4776), .B1(n6554), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6408) );
  NAND2_X1 U8176 ( .A1(n6410), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6411) );
  NAND2_X1 U8177 ( .A1(n6426), .A2(n6411), .ZN(n8968) );
  NAND2_X1 U8178 ( .A1(n8968), .A2(n6534), .ZN(n6415) );
  NAND2_X1 U8179 ( .A1(n6545), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8180 ( .A1(n6535), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6413) );
  NAND2_X1 U8181 ( .A1(n6557), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6412) );
  NAND4_X1 U8182 ( .A1(n6415), .A2(n6414), .A3(n6413), .A4(n6412), .ZN(n8976)
         );
  OR2_X1 U8183 ( .A1(n9144), .A2(n8976), .ZN(n6825) );
  INV_X1 U8184 ( .A(n6625), .ZN(n6416) );
  MUX2_X1 U8185 ( .A(n6416), .B(n4737), .S(n4428), .Z(n6417) );
  AOI211_X1 U8186 ( .C1(n6418), .C2(n8984), .A(n8967), .B(n6417), .ZN(n6444)
         );
  NAND2_X1 U8187 ( .A1(n7327), .A2(n6472), .ZN(n6424) );
  NAND2_X1 U8188 ( .A1(n6419), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6420) );
  MUX2_X1 U8189 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6420), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6422) );
  AND2_X1 U8190 ( .A1(n6422), .A2(n6421), .ZN(n8479) );
  AOI22_X1 U8191 ( .A1(n6554), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n8479), .B2(
        n4776), .ZN(n6423) );
  INV_X1 U8192 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9252) );
  INV_X1 U8193 ( .A(n6425), .ZN(n6437) );
  NAND2_X1 U8194 ( .A1(n6426), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8195 ( .A1(n6437), .A2(n6427), .ZN(n8959) );
  NAND2_X1 U8196 ( .A1(n8959), .A2(n6534), .ZN(n6432) );
  INV_X1 U8197 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9141) );
  OR2_X1 U8198 ( .A1(n4430), .A2(n9141), .ZN(n6430) );
  INV_X1 U8199 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8958) );
  OR2_X1 U8200 ( .A1(n6453), .A2(n8958), .ZN(n6429) );
  AND2_X1 U8201 ( .A1(n6430), .A2(n6429), .ZN(n6431) );
  OAI211_X1 U8202 ( .C1(n6489), .C2(n9252), .A(n6432), .B(n6431), .ZN(n8964)
         );
  INV_X1 U8203 ( .A(n8964), .ZN(n8327) );
  NAND2_X1 U8204 ( .A1(n9253), .A2(n8327), .ZN(n6630) );
  NAND2_X1 U8205 ( .A1(n6631), .A2(n6630), .ZN(n6826) );
  INV_X1 U8206 ( .A(n8976), .ZN(n8953) );
  NAND2_X1 U8207 ( .A1(n9144), .A2(n8953), .ZN(n6628) );
  OR2_X1 U8208 ( .A1(n9144), .A2(n8953), .ZN(n6629) );
  MUX2_X1 U8209 ( .A(n6628), .B(n6629), .S(n6886), .Z(n6433) );
  NAND2_X1 U8210 ( .A1(n8952), .A2(n6433), .ZN(n6443) );
  NAND2_X1 U8211 ( .A1(n7474), .A2(n6472), .ZN(n6436) );
  NAND2_X1 U8212 ( .A1(n6421), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6434) );
  XNOR2_X1 U8213 ( .A(n6434), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8767) );
  AOI22_X1 U8214 ( .A1(n6554), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n8767), .B2(
        n4776), .ZN(n6435) );
  NAND2_X1 U8215 ( .A1(n6437), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8216 ( .A1(n6449), .A2(n6438), .ZN(n8947) );
  NAND2_X1 U8217 ( .A1(n8947), .A2(n6534), .ZN(n6441) );
  AOI22_X1 U8218 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n6535), .B1(n6545), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U8219 ( .A1(n6557), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8220 ( .A1(n8948), .A2(n8954), .ZN(n6633) );
  NAND2_X1 U8221 ( .A1(n8927), .A2(n6633), .ZN(n6827) );
  MUX2_X1 U8222 ( .A(n6630), .B(n6631), .S(n4428), .Z(n6442) );
  NAND2_X1 U8223 ( .A1(n7499), .A2(n6472), .ZN(n6448) );
  NAND2_X1 U8224 ( .A1(n6445), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U8225 ( .A(n6446), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8786) );
  AOI22_X1 U8226 ( .A1(n6554), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n8786), .B2(
        n4776), .ZN(n6447) );
  INV_X1 U8227 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U8228 ( .A1(n6449), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8229 ( .A1(n6457), .A2(n6450), .ZN(n8931) );
  NAND2_X1 U8230 ( .A1(n8931), .A2(n6534), .ZN(n6452) );
  AOI22_X1 U8231 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n6535), .B1(n6545), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6451) );
  OAI211_X1 U8232 ( .C1(n6453), .C2(n8758), .A(n6452), .B(n6451), .ZN(n8943)
         );
  NAND2_X1 U8233 ( .A1(n6830), .A2(n6733), .ZN(n6635) );
  NAND2_X1 U8234 ( .A1(n7765), .A2(n6472), .ZN(n6456) );
  AOI22_X1 U8235 ( .A1(n6554), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6772), .B2(
        n4776), .ZN(n6455) );
  NAND2_X1 U8236 ( .A1(n6457), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U8237 ( .A1(n6465), .A2(n6458), .ZN(n8921) );
  INV_X1 U8238 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U8239 ( .A1(n6557), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U8240 ( .A1(n6545), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6459) );
  OAI211_X1 U8241 ( .C1(n4430), .C2(n9132), .A(n6460), .B(n6459), .ZN(n6461)
         );
  AOI21_X1 U8242 ( .B1(n8921), .B2(n6534), .A(n6461), .ZN(n8926) );
  OR2_X1 U8243 ( .A1(n9238), .A2(n8926), .ZN(n6483) );
  NAND2_X1 U8244 ( .A1(n9238), .A2(n8926), .ZN(n6636) );
  NAND2_X1 U8245 ( .A1(n6483), .A2(n6636), .ZN(n8915) );
  INV_X1 U8246 ( .A(n8915), .ZN(n8916) );
  OR2_X1 U8247 ( .A1(n6830), .A2(n6733), .ZN(n6580) );
  NAND2_X1 U8248 ( .A1(n7813), .A2(n6472), .ZN(n6463) );
  NAND2_X1 U8249 ( .A1(n6554), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6462) );
  INV_X1 U8250 ( .A(n6464), .ZN(n6475) );
  NAND2_X1 U8251 ( .A1(n6465), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8252 ( .A1(n6475), .A2(n6466), .ZN(n8911) );
  NAND2_X1 U8253 ( .A1(n8911), .A2(n6534), .ZN(n6471) );
  INV_X1 U8254 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8910) );
  NAND2_X1 U8255 ( .A1(n6545), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8256 ( .A1(n6535), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6467) );
  OAI211_X1 U8257 ( .C1(n8910), .C2(n6453), .A(n6468), .B(n6467), .ZN(n6469)
         );
  INV_X1 U8258 ( .A(n6469), .ZN(n6470) );
  NAND2_X1 U8259 ( .A1(n9232), .A2(n8204), .ZN(n6638) );
  NAND2_X1 U8260 ( .A1(n7832), .A2(n6472), .ZN(n6474) );
  NAND2_X1 U8261 ( .A1(n6554), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8262 ( .A1(n6475), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8263 ( .A1(n6487), .A2(n6476), .ZN(n8899) );
  INV_X1 U8264 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8898) );
  NAND2_X1 U8265 ( .A1(n6545), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8266 ( .A1(n6535), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6477) );
  OAI211_X1 U8267 ( .C1(n8898), .C2(n6453), .A(n6478), .B(n6477), .ZN(n6479)
         );
  NAND2_X1 U8268 ( .A1(n9226), .A2(n8882), .ZN(n6639) );
  AND2_X1 U8269 ( .A1(n6580), .A2(n8927), .ZN(n6634) );
  INV_X1 U8270 ( .A(n6636), .ZN(n6481) );
  INV_X1 U8271 ( .A(n6635), .ZN(n6480) );
  NAND2_X1 U8272 ( .A1(n7836), .A2(n6553), .ZN(n6486) );
  NAND2_X1 U8273 ( .A1(n6554), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6485) );
  NAND2_X1 U8274 ( .A1(n6487), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U8275 ( .A1(n6499), .A2(n6488), .ZN(n8886) );
  NAND2_X1 U8276 ( .A1(n8886), .A2(n6534), .ZN(n6494) );
  INV_X1 U8277 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U8278 ( .A1(n6557), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6491) );
  INV_X1 U8279 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9221) );
  OR2_X1 U8280 ( .A1(n6489), .A2(n9221), .ZN(n6490) );
  OAI211_X1 U8281 ( .C1(n4430), .C2(n9124), .A(n6491), .B(n6490), .ZN(n6492)
         );
  INV_X1 U8282 ( .A(n6492), .ZN(n6493) );
  XNOR2_X1 U8283 ( .A(n9223), .B(n8213), .ZN(n8883) );
  INV_X1 U8284 ( .A(n8852), .ZN(n6495) );
  AND2_X1 U8285 ( .A1(n8282), .A2(n8213), .ZN(n6643) );
  MUX2_X1 U8286 ( .A(n6495), .B(n6643), .S(n4428), .Z(n6496) );
  NAND2_X1 U8287 ( .A1(n7865), .A2(n6553), .ZN(n6498) );
  NAND2_X1 U8288 ( .A1(n6554), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U8289 ( .A1(n6499), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6500) );
  NAND2_X1 U8290 ( .A1(n6501), .A2(n6500), .ZN(n8874) );
  NAND2_X1 U8291 ( .A1(n8874), .A2(n6534), .ZN(n6506) );
  INV_X1 U8292 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U8293 ( .A1(n6545), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8294 ( .A1(n6557), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6502) );
  OAI211_X1 U8295 ( .C1(n4430), .C2(n9116), .A(n6503), .B(n6502), .ZN(n6504)
         );
  INV_X1 U8296 ( .A(n6504), .ZN(n6505) );
  OR2_X1 U8297 ( .A1(n9216), .A2(n8881), .ZN(n6640) );
  INV_X1 U8298 ( .A(n6640), .ZN(n8854) );
  NAND2_X1 U8299 ( .A1(n9216), .A2(n8881), .ZN(n8853) );
  OAI21_X1 U8300 ( .B1(n6511), .B2(n8854), .A(n6644), .ZN(n6518) );
  INV_X1 U8301 ( .A(n6644), .ZN(n6510) );
  NAND3_X1 U8302 ( .A1(n6645), .A2(n6886), .A3(n6648), .ZN(n6508) );
  OAI21_X1 U8303 ( .B1(n6511), .B2(n6510), .A(n6509), .ZN(n6517) );
  OAI21_X1 U8304 ( .B1(n4428), .B2(n6647), .A(n6512), .ZN(n6515) );
  NOR3_X1 U8305 ( .A1(n6837), .A2(n4428), .A3(n8841), .ZN(n6514) );
  AOI211_X1 U8306 ( .C1(n8832), .C2(n6515), .A(n6514), .B(n6513), .ZN(n6516)
         );
  AOI22_X1 U8307 ( .A1(n6519), .A2(n6518), .B1(n6517), .B2(n6516), .ZN(n6531)
         );
  NAND2_X1 U8308 ( .A1(n9304), .A2(n6472), .ZN(n6521) );
  NAND2_X1 U8309 ( .A1(n6554), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6520) );
  NAND2_X1 U8310 ( .A1(n6522), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6523) );
  NAND2_X1 U8311 ( .A1(n6532), .A2(n6523), .ZN(n8828) );
  NAND2_X1 U8312 ( .A1(n8828), .A2(n6534), .ZN(n6528) );
  INV_X1 U8313 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U8314 ( .A1(n6545), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6525) );
  INV_X1 U8315 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9106) );
  OR2_X1 U8316 ( .A1(n4429), .A2(n9106), .ZN(n6524) );
  OAI211_X1 U8317 ( .C1(n8827), .C2(n6453), .A(n6525), .B(n6524), .ZN(n6526)
         );
  INV_X1 U8318 ( .A(n6526), .ZN(n6527) );
  INV_X1 U8319 ( .A(n8823), .ZN(n8824) );
  NAND2_X1 U8320 ( .A1(n9192), .A2(n7978), .ZN(n6529) );
  MUX2_X1 U8321 ( .A(n6651), .B(n6529), .S(n4428), .Z(n6530) );
  NAND2_X1 U8322 ( .A1(n6532), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6533) );
  INV_X1 U8323 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U8324 ( .A1(n6535), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8325 ( .A1(n6545), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6536) );
  OAI211_X1 U8326 ( .C1(n8818), .C2(n6453), .A(n6537), .B(n6536), .ZN(n6538)
         );
  INV_X1 U8327 ( .A(n6538), .ZN(n6539) );
  NAND2_X1 U8328 ( .A1(n8004), .A2(n6553), .ZN(n6541) );
  NAND2_X1 U8329 ( .A1(n6554), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6540) );
  MUX2_X1 U8330 ( .A(n7968), .B(n7970), .S(n6886), .Z(n6563) );
  NAND2_X1 U8331 ( .A1(n9298), .A2(n6553), .ZN(n6544) );
  NAND2_X1 U8332 ( .A1(n6554), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6543) );
  INV_X1 U8333 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8651) );
  NAND2_X1 U8334 ( .A1(n6545), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8335 ( .A1(n6557), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6546) );
  OAI211_X1 U8336 ( .C1(n4430), .C2(n8651), .A(n6547), .B(n6546), .ZN(n6548)
         );
  INV_X1 U8337 ( .A(n6548), .ZN(n6549) );
  NAND2_X1 U8338 ( .A1(n6870), .A2(n4428), .ZN(n6550) );
  AOI22_X1 U8339 ( .A1(n6845), .A2(n6550), .B1(n4428), .B2(n8817), .ZN(n6564)
         );
  NAND2_X1 U8340 ( .A1(n9295), .A2(n6553), .ZN(n6556) );
  NAND2_X1 U8341 ( .A1(n6554), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6555) );
  INV_X1 U8342 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9102) );
  NAND2_X1 U8343 ( .A1(n6545), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U8344 ( .A1(n6557), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6558) );
  OAI211_X1 U8345 ( .C1(n4430), .C2(n9102), .A(n6559), .B(n6558), .ZN(n6560)
         );
  INV_X1 U8346 ( .A(n6560), .ZN(n6561) );
  NAND2_X1 U8347 ( .A1(n6562), .A2(n6561), .ZN(n8334) );
  INV_X1 U8348 ( .A(n8334), .ZN(n6567) );
  NAND2_X1 U8349 ( .A1(n9099), .A2(n6567), .ZN(n6576) );
  NAND2_X1 U8350 ( .A1(n6870), .A2(n7976), .ZN(n6844) );
  NOR2_X1 U8351 ( .A1(n9099), .A2(n6567), .ZN(n6653) );
  NOR3_X1 U8352 ( .A1(n6566), .A2(n4830), .A3(n6653), .ZN(n6572) );
  OAI21_X1 U8353 ( .B1(n6567), .B2(n6886), .A(n9099), .ZN(n6568) );
  OAI21_X1 U8354 ( .B1(n4428), .B2(n8334), .A(n6568), .ZN(n6571) );
  NAND4_X1 U8355 ( .A1(n6569), .A2(n7970), .A3(n4428), .A4(n6576), .ZN(n6570)
         );
  OAI21_X1 U8356 ( .B1(n6572), .B2(n6571), .A(n6570), .ZN(n6573) );
  AND2_X1 U8357 ( .A1(n6576), .A2(n6844), .ZN(n6577) );
  NAND2_X1 U8358 ( .A1(n6578), .A2(n6577), .ZN(n6655) );
  NAND2_X1 U8359 ( .A1(n6640), .A2(n8853), .ZN(n8869) );
  NAND2_X1 U8360 ( .A1(n6637), .A2(n6638), .ZN(n8905) );
  INV_X1 U8361 ( .A(n8967), .ZN(n8963) );
  INV_X1 U8362 ( .A(n8984), .ZN(n6593) );
  NAND2_X1 U8363 ( .A1(n6615), .A2(n9018), .ZN(n9039) );
  INV_X1 U8364 ( .A(n9039), .ZN(n9042) );
  NOR2_X1 U8365 ( .A1(n6804), .A2(n4435), .ZN(n6587) );
  NAND2_X1 U8366 ( .A1(n7955), .A2(n6582), .ZN(n7337) );
  NOR2_X1 U8367 ( .A1(n6806), .A2(n7337), .ZN(n6586) );
  INV_X1 U8368 ( .A(n6583), .ZN(n6584) );
  NAND4_X1 U8369 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n7492), .ZN(n6589)
         );
  INV_X1 U8370 ( .A(n7431), .ZN(n7426) );
  OR3_X1 U8371 ( .A1(n6589), .A2(n5286), .A3(n7426), .ZN(n6590) );
  NAND2_X1 U8372 ( .A1(n9034), .A2(n6614), .ZN(n9033) );
  NAND2_X1 U8373 ( .A1(n9032), .A2(n6613), .ZN(n7660) );
  NOR3_X1 U8374 ( .A1(n6590), .A2(n9033), .A3(n7660), .ZN(n6591) );
  NAND2_X1 U8375 ( .A1(n8963), .A2(n6594), .ZN(n6595) );
  NOR2_X1 U8376 ( .A1(n6826), .A2(n6595), .ZN(n6596) );
  AND4_X1 U8377 ( .A1(n8815), .A2(n5413), .A3(n8832), .A4(n8823), .ZN(n6598)
         );
  INV_X1 U8378 ( .A(n7829), .ZN(n6658) );
  NAND3_X1 U8379 ( .A1(n6657), .A2(n6658), .A3(n6772), .ZN(n6656) );
  NAND2_X1 U8380 ( .A1(n7346), .A2(n7350), .ZN(n6602) );
  NAND2_X1 U8381 ( .A1(n6602), .A2(n6601), .ZN(n7362) );
  NAND2_X1 U8382 ( .A1(n7362), .A2(n7365), .ZN(n6604) );
  NAND2_X1 U8383 ( .A1(n6604), .A2(n6603), .ZN(n7411) );
  NAND2_X1 U8384 ( .A1(n7411), .A2(n7415), .ZN(n6606) );
  AOI21_X1 U8385 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(n6611) );
  AND2_X1 U8386 ( .A1(n6614), .A2(n6613), .ZN(n9017) );
  INV_X1 U8387 ( .A(n6614), .ZN(n6616) );
  OAI211_X1 U8388 ( .C1(n6616), .C2(n9032), .A(n6615), .B(n9034), .ZN(n9016)
         );
  NAND2_X1 U8389 ( .A1(n9016), .A2(n9018), .ZN(n6617) );
  INV_X1 U8390 ( .A(n9005), .ZN(n6620) );
  NAND2_X1 U8391 ( .A1(n6624), .A2(n6623), .ZN(n8983) );
  NAND2_X1 U8392 ( .A1(n8983), .A2(n6625), .ZN(n6627) );
  OAI211_X1 U8393 ( .C1(n6643), .C2(n8850), .A(n6640), .B(n8852), .ZN(n6641)
         );
  INV_X1 U8394 ( .A(n6641), .ZN(n6642) );
  NAND2_X1 U8395 ( .A1(n8845), .A2(n6647), .ZN(n6649) );
  OR2_X1 U8396 ( .A1(n9198), .A2(n6838), .ZN(n6650) );
  OR2_X1 U8397 ( .A1(n9186), .A2(n7968), .ZN(n6652) );
  NAND2_X1 U8398 ( .A1(n4435), .A2(n6658), .ZN(n6848) );
  AOI21_X1 U8399 ( .B1(n6653), .B2(n9177), .A(n6848), .ZN(n6654) );
  INV_X1 U8400 ( .A(n6657), .ZN(n6659) );
  NAND2_X1 U8401 ( .A1(n6662), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6661) );
  MUX2_X1 U8402 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6661), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n6664) );
  INV_X1 U8403 ( .A(n6662), .ZN(n6663) );
  NAND2_X1 U8404 ( .A1(n6663), .A2(n6138), .ZN(n6665) );
  NAND2_X1 U8405 ( .A1(n6664), .A2(n6665), .ZN(n6885) );
  NOR2_X1 U8406 ( .A1(n6885), .A2(P2_U3151), .ZN(n7861) );
  INV_X1 U8407 ( .A(n7336), .ZN(n6675) );
  INV_X1 U8408 ( .A(n6682), .ZN(n9310) );
  NAND2_X1 U8409 ( .A1(n6667), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6668) );
  MUX2_X1 U8410 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6668), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6669) );
  NAND2_X1 U8411 ( .A1(n9310), .A2(n7869), .ZN(n6887) );
  NAND2_X1 U8412 ( .A1(n6675), .A2(n6929), .ZN(n6794) );
  INV_X1 U8413 ( .A(n6794), .ZN(n6785) );
  INV_X1 U8414 ( .A(n6676), .ZN(n7168) );
  NAND3_X1 U8415 ( .A1(n6785), .A2(n7168), .A3(n8770), .ZN(n6678) );
  OAI211_X1 U8416 ( .C1(n6780), .C2(n5135), .A(n6678), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6679) );
  XNOR2_X1 U8417 ( .A(n6682), .B(P2_B_REG_SCAN_IN), .ZN(n6681) );
  INV_X1 U8418 ( .A(n7869), .ZN(n6755) );
  NAND2_X1 U8419 ( .A1(n6682), .A2(n6755), .ZN(n6944) );
  NOR2_X1 U8420 ( .A1(n4435), .A2(n7829), .ZN(n6683) );
  NAND2_X1 U8421 ( .A1(n6758), .A2(n6683), .ZN(n6687) );
  NAND2_X1 U8422 ( .A1(n4434), .A2(n7829), .ZN(n6850) );
  AND2_X1 U8423 ( .A1(n6685), .A2(n6850), .ZN(n6686) );
  INV_X2 U8424 ( .A(n6688), .ZN(n6690) );
  INV_X2 U8425 ( .A(n6690), .ZN(n6693) );
  XNOR2_X1 U8426 ( .A(n9192), .B(n7967), .ZN(n7977) );
  NOR2_X1 U8427 ( .A1(n7977), .A2(n7978), .ZN(n7972) );
  AOI21_X1 U8428 ( .B1(n7978), .B2(n7977), .A(n7972), .ZN(n6779) );
  XNOR2_X1 U8429 ( .A(n8948), .B(n7967), .ZN(n6730) );
  INV_X1 U8430 ( .A(n6730), .ZN(n6731) );
  INV_X1 U8431 ( .A(n8954), .ZN(n8335) );
  XNOR2_X1 U8432 ( .A(n7967), .B(n7692), .ZN(n6705) );
  INV_X1 U8433 ( .A(n6705), .ZN(n6706) );
  OAI21_X1 U8434 ( .B1(n6689), .B2(n7352), .A(n6691), .ZN(n7145) );
  NOR2_X1 U8435 ( .A1(n7145), .A2(n7146), .ZN(n7144) );
  INV_X1 U8436 ( .A(n6691), .ZN(n6692) );
  XNOR2_X1 U8437 ( .A(n6695), .B(n8339), .ZN(n7152) );
  NOR2_X1 U8438 ( .A1(n7151), .A2(n7152), .ZN(n7377) );
  XNOR2_X1 U8439 ( .A(n6693), .B(n7369), .ZN(n7376) );
  INV_X1 U8440 ( .A(n7376), .ZN(n6697) );
  XNOR2_X1 U8441 ( .A(n6693), .B(n7421), .ZN(n6698) );
  NAND2_X1 U8442 ( .A1(n6698), .A2(n6809), .ZN(n7506) );
  INV_X1 U8443 ( .A(n6695), .ZN(n6696) );
  NAND2_X1 U8444 ( .A1(n6696), .A2(n7958), .ZN(n7378) );
  OAI211_X1 U8445 ( .C1(n6697), .C2(n6694), .A(n7506), .B(n7378), .ZN(n6700)
         );
  NOR2_X1 U8446 ( .A1(n7376), .A2(n7375), .ZN(n7399) );
  NOR2_X1 U8447 ( .A1(n6698), .A2(n6809), .ZN(n7402) );
  OAI21_X1 U8448 ( .B1(n7399), .B2(n7402), .A(n7506), .ZN(n6699) );
  XNOR2_X1 U8449 ( .A(n6693), .B(n6808), .ZN(n6701) );
  XNOR2_X1 U8450 ( .A(n6701), .B(n4812), .ZN(n7505) );
  XNOR2_X1 U8451 ( .A(n7967), .B(n7441), .ZN(n6703) );
  XNOR2_X1 U8452 ( .A(n6703), .B(n8337), .ZN(n7448) );
  AND2_X1 U8453 ( .A1(n6703), .A2(n8337), .ZN(n6704) );
  XNOR2_X1 U8454 ( .A(n6705), .B(n8336), .ZN(n7481) );
  OAI21_X1 U8455 ( .B1(n6706), .B2(n8336), .A(n7480), .ZN(n7544) );
  XOR2_X1 U8456 ( .A(n7967), .B(n9076), .Z(n7542) );
  NAND2_X1 U8457 ( .A1(n7542), .A2(n9063), .ZN(n6708) );
  INV_X1 U8458 ( .A(n7542), .ZN(n6707) );
  XNOR2_X1 U8459 ( .A(n7681), .B(n7967), .ZN(n6709) );
  INV_X1 U8460 ( .A(n7655), .ZN(n9047) );
  XNOR2_X1 U8461 ( .A(n6709), .B(n9047), .ZN(n7683) );
  XNOR2_X1 U8462 ( .A(n9020), .B(n7967), .ZN(n8290) );
  XOR2_X1 U8463 ( .A(n7967), .B(n8198), .Z(n8287) );
  NOR3_X1 U8464 ( .A1(n8198), .A2(n7685), .A3(n6690), .ZN(n6713) );
  AOI211_X1 U8465 ( .C1(n6690), .C2(n9046), .A(n6713), .B(n9022), .ZN(n6716)
         );
  INV_X1 U8466 ( .A(n8198), .ZN(n9285) );
  NOR3_X1 U8467 ( .A1(n9285), .A2(n7685), .A3(n7967), .ZN(n6714) );
  AOI211_X1 U8468 ( .C1(n9046), .C2(n7967), .A(n6714), .B(n9020), .ZN(n6715)
         );
  XNOR2_X1 U8469 ( .A(n9155), .B(n7967), .ZN(n6718) );
  XNOR2_X1 U8470 ( .A(n6718), .B(n9024), .ZN(n8218) );
  XNOR2_X1 U8471 ( .A(n9266), .B(n7967), .ZN(n6721) );
  XNOR2_X1 U8472 ( .A(n6721), .B(n6722), .ZN(n8269) );
  INV_X1 U8473 ( .A(n8269), .ZN(n6720) );
  XNOR2_X1 U8474 ( .A(n9260), .B(n7967), .ZN(n6725) );
  XNOR2_X1 U8475 ( .A(n6725), .B(n8991), .ZN(n8179) );
  AND2_X1 U8476 ( .A1(n6725), .A2(n6724), .ZN(n6726) );
  AOI21_X2 U8477 ( .B1(n8180), .B2(n8179), .A(n6726), .ZN(n8323) );
  XNOR2_X1 U8478 ( .A(n9144), .B(n7967), .ZN(n6727) );
  XNOR2_X1 U8479 ( .A(n6727), .B(n8976), .ZN(n8322) );
  XNOR2_X1 U8480 ( .A(n9253), .B(n7967), .ZN(n6729) );
  XNOR2_X1 U8481 ( .A(n6729), .B(n8327), .ZN(n8238) );
  XNOR2_X1 U8482 ( .A(n6730), .B(n8335), .ZN(n8244) );
  XNOR2_X1 U8483 ( .A(n6830), .B(n7967), .ZN(n6732) );
  XNOR2_X1 U8484 ( .A(n6732), .B(n8943), .ZN(n8298) );
  XNOR2_X1 U8485 ( .A(n9238), .B(n7967), .ZN(n6734) );
  INV_X1 U8486 ( .A(n8926), .ZN(n8907) );
  NAND2_X1 U8487 ( .A1(n6734), .A2(n8926), .ZN(n6735) );
  XOR2_X1 U8488 ( .A(n7967), .B(n9232), .Z(n6737) );
  INV_X1 U8489 ( .A(n6737), .ZN(n6736) );
  XNOR2_X1 U8490 ( .A(n6736), .B(n8918), .ZN(n8259) );
  XNOR2_X1 U8491 ( .A(n9226), .B(n7967), .ZN(n6739) );
  XNOR2_X1 U8492 ( .A(n6739), .B(n8882), .ZN(n8210) );
  INV_X1 U8493 ( .A(n8210), .ZN(n6738) );
  NAND2_X1 U8494 ( .A1(n8209), .A2(n6738), .ZN(n6741) );
  NAND2_X1 U8495 ( .A1(n6739), .A2(n8882), .ZN(n6740) );
  XNOR2_X1 U8496 ( .A(n9223), .B(n7967), .ZN(n6742) );
  NAND2_X1 U8497 ( .A1(n6742), .A2(n8896), .ZN(n8276) );
  INV_X1 U8498 ( .A(n6742), .ZN(n6743) );
  NAND2_X1 U8499 ( .A1(n6743), .A2(n8213), .ZN(n8277) );
  XNOR2_X1 U8500 ( .A(n9216), .B(n6690), .ZN(n8187) );
  NOR2_X1 U8501 ( .A1(n8187), .A2(n8857), .ZN(n6747) );
  XNOR2_X1 U8502 ( .A(n6744), .B(n6690), .ZN(n6745) );
  NAND2_X1 U8503 ( .A1(n6745), .A2(n8232), .ZN(n8226) );
  OAI21_X1 U8504 ( .B1(n6745), .B2(n8232), .A(n8226), .ZN(n8252) );
  AOI21_X1 U8505 ( .B1(n8187), .B2(n8857), .A(n8252), .ZN(n6746) );
  XNOR2_X1 U8506 ( .A(n8236), .B(n7967), .ZN(n6749) );
  XNOR2_X1 U8507 ( .A(n6749), .B(n8314), .ZN(n8227) );
  NAND2_X1 U8508 ( .A1(n6748), .A2(n8227), .ZN(n8228) );
  INV_X1 U8509 ( .A(n6749), .ZN(n6750) );
  NAND2_X1 U8510 ( .A1(n6750), .A2(n8314), .ZN(n6751) );
  XNOR2_X1 U8511 ( .A(n6837), .B(n7967), .ZN(n6752) );
  NOR2_X1 U8512 ( .A1(n6752), .A2(n8841), .ZN(n8306) );
  NAND2_X1 U8513 ( .A1(n6752), .A2(n8841), .ZN(n8307) );
  OAI21_X1 U8514 ( .B1(n8305), .B2(n8306), .A(n8307), .ZN(n6778) );
  INV_X1 U8515 ( .A(n6779), .ZN(n6753) );
  OR2_X1 U8516 ( .A1(n6754), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6757) );
  NAND2_X1 U8517 ( .A1(n6680), .A2(n6755), .ZN(n6756) );
  NAND2_X1 U8518 ( .A1(n6757), .A2(n6756), .ZN(n6880) );
  INV_X1 U8519 ( .A(n6880), .ZN(n7330) );
  NAND2_X1 U8520 ( .A1(n7330), .A2(n6758), .ZN(n6879) );
  NOR2_X1 U8521 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n6762) );
  NOR4_X1 U8522 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6761) );
  NOR4_X1 U8523 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6760) );
  NOR4_X1 U8524 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6759) );
  NAND4_X1 U8525 ( .A1(n6762), .A2(n6761), .A3(n6760), .A4(n6759), .ZN(n6768)
         );
  NOR4_X1 U8526 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6766) );
  NOR4_X1 U8527 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6765) );
  NOR4_X1 U8528 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6764) );
  NOR4_X1 U8529 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6763) );
  NAND4_X1 U8530 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6767)
         );
  NOR2_X1 U8531 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  OR2_X1 U8532 ( .A1(n6754), .A2(n6769), .ZN(n6876) );
  INV_X1 U8533 ( .A(n6876), .ZN(n6770) );
  INV_X1 U8534 ( .A(n6929), .ZN(n6771) );
  NAND2_X1 U8535 ( .A1(n6772), .A2(n6780), .ZN(n6847) );
  OR3_X1 U8536 ( .A1(n4435), .A2(n7829), .A3(n6847), .ZN(n6861) );
  NAND3_X1 U8537 ( .A1(n10537), .A2(n6861), .A3(n6886), .ZN(n6788) );
  INV_X1 U8538 ( .A(n6788), .ZN(n6773) );
  NAND2_X1 U8539 ( .A1(n6863), .A2(n6773), .ZN(n6777) );
  NAND2_X1 U8540 ( .A1(n6880), .A2(n6876), .ZN(n6774) );
  INV_X1 U8541 ( .A(n6861), .ZN(n6775) );
  NAND2_X1 U8542 ( .A1(n6865), .A2(n6775), .ZN(n6776) );
  OAI211_X1 U8543 ( .C1(n6779), .C2(n6778), .A(n7984), .B(n8320), .ZN(n6802)
         );
  INV_X1 U8544 ( .A(n9192), .ZN(n6839) );
  INV_X1 U8545 ( .A(n8995), .ZN(n8980) );
  NAND2_X1 U8546 ( .A1(n6863), .A2(n8980), .ZN(n6782) );
  OR2_X1 U8547 ( .A1(n10525), .A2(n4435), .ZN(n6872) );
  INV_X1 U8548 ( .A(n6872), .ZN(n6781) );
  INV_X1 U8549 ( .A(n8770), .ZN(n8788) );
  NAND2_X1 U8550 ( .A1(n8788), .A2(n7168), .ZN(n6783) );
  INV_X1 U8551 ( .A(n6853), .ZN(n6784) );
  NAND3_X1 U8552 ( .A1(n6785), .A2(n6793), .A3(n6784), .ZN(n8326) );
  OR2_X1 U8553 ( .A1(n6886), .A2(n6786), .ZN(n6877) );
  AND2_X1 U8554 ( .A1(n6877), .A2(n6787), .ZN(n6791) );
  NAND2_X1 U8555 ( .A1(n6788), .A2(n8995), .ZN(n6864) );
  NAND2_X1 U8556 ( .A1(n6789), .A2(n6864), .ZN(n6790) );
  OAI211_X1 U8557 ( .C1(n6793), .C2(n6861), .A(n6791), .B(n6790), .ZN(n6792)
         );
  NAND2_X1 U8558 ( .A1(n6792), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6796) );
  OR2_X1 U8559 ( .A1(n6794), .A2(n6793), .ZN(n6795) );
  AOI22_X1 U8560 ( .A1(n8828), .A2(n8329), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6797) );
  OAI21_X1 U8561 ( .B1(n6838), .B2(n8313), .A(n6797), .ZN(n6798) );
  AOI21_X1 U8562 ( .B1(n8826), .B2(n8310), .A(n6798), .ZN(n6799) );
  NAND2_X1 U8563 ( .A1(n6802), .A2(n6801), .ZN(P2_U3154) );
  NOR2_X1 U8564 ( .A1(n9232), .A2(n8918), .ZN(n8893) );
  INV_X1 U8565 ( .A(n8882), .ZN(n8908) );
  NOR2_X1 U8566 ( .A1(n9226), .A2(n8908), .ZN(n8877) );
  AOI21_X1 U8567 ( .B1(n8893), .B2(n8892), .A(n8877), .ZN(n8865) );
  NAND2_X1 U8568 ( .A1(n9223), .A2(n8213), .ZN(n8867) );
  AND2_X1 U8569 ( .A1(n8865), .A2(n8867), .ZN(n6831) );
  NAND2_X1 U8570 ( .A1(n6239), .A2(n7344), .ZN(n7957) );
  NAND2_X1 U8571 ( .A1(n7352), .A2(n6803), .ZN(n7349) );
  NAND2_X1 U8572 ( .A1(n7348), .A2(n7349), .ZN(n6805) );
  NAND2_X1 U8573 ( .A1(n6805), .A2(n6804), .ZN(n7347) );
  NAND2_X1 U8574 ( .A1(n7347), .A2(n7364), .ZN(n6807) );
  NAND2_X1 U8575 ( .A1(n7375), .A2(n10533), .ZN(n7414) );
  NAND2_X1 U8576 ( .A1(n6809), .A2(n10538), .ZN(n7489) );
  NAND2_X1 U8577 ( .A1(n8338), .A2(n10542), .ZN(n6813) );
  NAND2_X1 U8578 ( .A1(n8337), .A2(n7453), .ZN(n6815) );
  NAND2_X1 U8579 ( .A1(n7656), .A2(n9089), .ZN(n6816) );
  NAND2_X1 U8580 ( .A1(n9076), .A2(n9063), .ZN(n6817) );
  NOR2_X1 U8581 ( .A1(n7681), .A2(n9047), .ZN(n9038) );
  NOR2_X1 U8582 ( .A1(n8198), .A2(n9066), .ZN(n6818) );
  AOI21_X1 U8583 ( .B1(n9039), .B2(n9038), .A(n6818), .ZN(n6819) );
  OR2_X1 U8584 ( .A1(n9276), .A2(n9046), .ZN(n6820) );
  NOR2_X1 U8585 ( .A1(n9155), .A2(n9024), .ZN(n6821) );
  INV_X1 U8586 ( .A(n9155), .ZN(n8224) );
  OR2_X1 U8587 ( .A1(n9260), .A2(n8991), .ZN(n6824) );
  NAND2_X1 U8588 ( .A1(n6827), .A2(n6826), .ZN(n6829) );
  AND2_X1 U8589 ( .A1(n9253), .A2(n8964), .ZN(n8938) );
  AOI22_X1 U8590 ( .A1(n6827), .A2(n8938), .B1(n8948), .B2(n8335), .ZN(n6828)
         );
  AOI22_X1 U8591 ( .A1(n9216), .A2(n8857), .B1(n8282), .B2(n8896), .ZN(n6833)
         );
  INV_X1 U8592 ( .A(n9216), .ZN(n6832) );
  NAND2_X1 U8593 ( .A1(n6744), .A2(n8232), .ZN(n6835) );
  NAND2_X1 U8594 ( .A1(n9192), .A2(n8834), .ZN(n6840) );
  NAND2_X1 U8595 ( .A1(n7970), .A2(n7968), .ZN(n6841) );
  NAND2_X1 U8596 ( .A1(n9186), .A2(n8826), .ZN(n6842) );
  NAND2_X1 U8597 ( .A1(n6843), .A2(n6842), .ZN(n6846) );
  NAND2_X1 U8598 ( .A1(n6850), .A2(n7838), .ZN(n6851) );
  NAND2_X1 U8599 ( .A1(n6851), .A2(n8794), .ZN(n6873) );
  INV_X1 U8600 ( .A(n6873), .ZN(n6852) );
  NOR2_X1 U8601 ( .A1(n9008), .A2(n6854), .ZN(n8806) );
  AOI22_X1 U8602 ( .A1(n9064), .A2(n8826), .B1(n8334), .B2(n8806), .ZN(n6855)
         );
  INV_X1 U8603 ( .A(n10525), .ZN(n9169) );
  NAND2_X1 U8604 ( .A1(n8131), .A2(n9169), .ZN(n6860) );
  NAND2_X1 U8605 ( .A1(n7336), .A2(n6861), .ZN(n6862) );
  NAND2_X1 U8606 ( .A1(n6863), .A2(n6862), .ZN(n6867) );
  NAND2_X1 U8607 ( .A1(n6865), .A2(n6864), .ZN(n6866) );
  INV_X1 U8608 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8609 ( .A1(n10550), .A2(n6868), .ZN(n6869) );
  NAND2_X1 U8610 ( .A1(n6871), .A2(n5412), .ZN(P2_U3456) );
  AND2_X1 U8611 ( .A1(n6872), .A2(n6758), .ZN(n6875) );
  OR2_X1 U8612 ( .A1(n6873), .A2(n7829), .ZN(n6874) );
  NAND2_X1 U8613 ( .A1(n6874), .A2(n6886), .ZN(n7332) );
  OR2_X1 U8614 ( .A1(n6875), .A2(n7332), .ZN(n6882) );
  AND2_X1 U8615 ( .A1(n6929), .A2(n6876), .ZN(n6878) );
  NAND2_X1 U8616 ( .A1(n7332), .A2(n6880), .ZN(n6881) );
  NAND2_X1 U8617 ( .A1(n6884), .A2(n5405), .ZN(P2_U3488) );
  NAND2_X1 U8618 ( .A1(n7866), .A2(n7072), .ZN(n6920) );
  INV_X1 U8619 ( .A(n6885), .ZN(n6943) );
  OR2_X1 U8620 ( .A1(n6886), .A2(n6943), .ZN(n7167) );
  NAND2_X1 U8621 ( .A1(n6888), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  XNOR2_X1 U8622 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8623 ( .A1(n4431), .A2(P1_U3086), .ZN(n10315) );
  AND2_X1 U8624 ( .A1(n4956), .A2(P1_U3086), .ZN(n7864) );
  OAI222_X1 U8625 ( .A1(n10332), .A2(n6890), .B1(n10335), .B2(n6907), .C1(
        P1_U3086), .C2(n9870), .ZN(P1_U3351) );
  OAI222_X1 U8626 ( .A1(n10332), .A2(n6891), .B1(n10335), .B2(n6893), .C1(
        n10311), .C2(n9886), .ZN(P1_U3350) );
  NOR2_X1 U8627 ( .A1(n4431), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9309) );
  AOI22_X1 U8628 ( .A1(n7269), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n9309), .ZN(n6892) );
  OAI21_X1 U8629 ( .B1(n6893), .B2(n9307), .A(n6892), .ZN(P2_U3290) );
  INV_X2 U8630 ( .A(n7864), .ZN(n10335) );
  OAI222_X1 U8631 ( .A1(P1_U3086), .A2(n9852), .B1(n10335), .B2(n6909), .C1(
        n6894), .C2(n10332), .ZN(P1_U3352) );
  OAI222_X1 U8632 ( .A1(n10332), .A2(n6897), .B1(n10335), .B2(n6906), .C1(
        P1_U3086), .C2(n9900), .ZN(P1_U3349) );
  INV_X1 U8633 ( .A(n9309), .ZN(n8134) );
  OAI222_X1 U8634 ( .A1(P2_U3151), .A2(n7183), .B1(n9307), .B2(n6899), .C1(
        n6898), .C2(n8134), .ZN(P2_U3293) );
  INV_X1 U8635 ( .A(n6900), .ZN(n6905) );
  AOI22_X1 U8636 ( .A1(n9916), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10315), .ZN(n6901) );
  OAI21_X1 U8637 ( .B1(n6905), .B2(n10335), .A(n6901), .ZN(P1_U3348) );
  INV_X1 U8638 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U8639 ( .A1(n7330), .A2(n6929), .ZN(n6902) );
  OAI21_X1 U8640 ( .B1(n6929), .B2(n6903), .A(n6902), .ZN(P2_U3377) );
  INV_X1 U8641 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6904) );
  OAI222_X1 U8642 ( .A1(n4757), .A2(P2_U3151), .B1(n9307), .B2(n6905), .C1(
        n6904), .C2(n8134), .ZN(P2_U3288) );
  OAI222_X1 U8643 ( .A1(n7557), .A2(P2_U3151), .B1(n9307), .B2(n6906), .C1(
        n4783), .C2(n8134), .ZN(P2_U3289) );
  OAI222_X1 U8644 ( .A1(n7229), .A2(P2_U3151), .B1(n9307), .B2(n6907), .C1(
        n8686), .C2(n8134), .ZN(P2_U3291) );
  INV_X1 U8645 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6908) );
  OAI222_X1 U8646 ( .A1(n5298), .A2(P2_U3151), .B1(n9307), .B2(n6909), .C1(
        n6908), .C2(n8134), .ZN(P2_U3292) );
  INV_X1 U8647 ( .A(n6912), .ZN(n6915) );
  AOI22_X1 U8648 ( .A1(n7000), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10315), .ZN(n6913) );
  OAI21_X1 U8649 ( .B1(n6915), .B2(n10335), .A(n6913), .ZN(P1_U3347) );
  OAI222_X1 U8650 ( .A1(n7755), .A2(P2_U3151), .B1(n9307), .B2(n6915), .C1(
        n6914), .C2(n8134), .ZN(P2_U3287) );
  INV_X1 U8651 ( .A(n7056), .ZN(n6916) );
  NAND2_X1 U8652 ( .A1(n10405), .A2(n7057), .ZN(n6917) );
  OAI21_X1 U8653 ( .B1(n10405), .B2(n6918), .A(n6917), .ZN(P1_U3440) );
  AOI21_X1 U8654 ( .B1(n7866), .B2(n9735), .A(n6919), .ZN(n6922) );
  INV_X1 U8655 ( .A(n6922), .ZN(n6921) );
  AND2_X1 U8656 ( .A1(n6920), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8657 ( .A1(n6921), .A2(n6923), .ZN(n9994) );
  INV_X1 U8658 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6928) );
  INV_X1 U8659 ( .A(n6924), .ZN(n9807) );
  INV_X1 U8660 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7615) );
  AOI21_X1 U8661 ( .B1(n9807), .B2(n7615), .A(n8005), .ZN(n7115) );
  OAI21_X1 U8662 ( .B1(n9807), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7115), .ZN(
        n6925) );
  XNOR2_X1 U8663 ( .A(n6925), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6926) );
  AOI22_X1 U8664 ( .A1(n6985), .A2(n6926), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10311), .ZN(n6927) );
  OAI21_X1 U8665 ( .B1(n9994), .B2(n6928), .A(n6927), .ZN(P1_U3243) );
  INV_X1 U8666 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n8698) );
  NOR2_X1 U8667 ( .A1(n6942), .A2(n8698), .ZN(P2_U3259) );
  INV_X1 U8668 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n8541) );
  NOR2_X1 U8669 ( .A1(n6942), .A2(n8541), .ZN(P2_U3248) );
  INV_X1 U8670 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n8666) );
  NOR2_X1 U8671 ( .A1(n6942), .A2(n8666), .ZN(P2_U3260) );
  INV_X1 U8672 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n8508) );
  NOR2_X1 U8673 ( .A1(n6942), .A2(n8508), .ZN(P2_U3244) );
  INV_X1 U8674 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n8564) );
  NOR2_X1 U8675 ( .A1(n6942), .A2(n8564), .ZN(P2_U3235) );
  INV_X1 U8676 ( .A(n6930), .ZN(n6933) );
  AOI22_X1 U8677 ( .A1(n7025), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10315), .ZN(n6931) );
  OAI21_X1 U8678 ( .B1(n6933), .B2(n10335), .A(n6931), .ZN(P1_U3346) );
  OAI222_X1 U8679 ( .A1(P2_U3151), .A2(n5079), .B1(n9307), .B2(n6933), .C1(
        n6932), .C2(n8134), .ZN(P2_U3286) );
  INV_X1 U8680 ( .A(n6934), .ZN(n6936) );
  OAI222_X1 U8681 ( .A1(P2_U3151), .A2(n8360), .B1(n9307), .B2(n6936), .C1(
        n6935), .C2(n8134), .ZN(P2_U3285) );
  INV_X1 U8682 ( .A(n7005), .ZN(n7049) );
  OAI222_X1 U8683 ( .A1(n10332), .A2(n6937), .B1(n10335), .B2(n6936), .C1(
        n7049), .C2(n10311), .ZN(P1_U3345) );
  INV_X1 U8684 ( .A(n9994), .ZN(n9965) );
  NOR2_X1 U8685 ( .A1(n9965), .A2(P1_U3973), .ZN(P1_U3085) );
  AND2_X1 U8686 ( .A1(n6946), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8687 ( .A1(n6946), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8688 ( .A1(n6946), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8689 ( .A1(n6946), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8690 ( .A1(n6946), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8691 ( .A1(n6946), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8692 ( .A1(n6946), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8693 ( .A1(n6946), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8694 ( .A1(n6946), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8695 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8663) );
  NAND2_X1 U8696 ( .A1(n5508), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8697 ( .A1(n4438), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U8698 ( .A1(n4437), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6938) );
  NAND3_X1 U8699 ( .A1(n6940), .A2(n6939), .A3(n6938), .ZN(n9734) );
  NAND2_X1 U8700 ( .A1(P1_U3973), .A2(n9734), .ZN(n6941) );
  OAI21_X1 U8701 ( .B1(P1_U3973), .B2(n8663), .A(n6941), .ZN(P1_U3585) );
  NOR3_X1 U8702 ( .A1(n6944), .A2(n6943), .A3(P2_U3151), .ZN(n6945) );
  AOI21_X1 U8703 ( .B1(n6946), .B2(n4922), .A(n6945), .ZN(P2_U3376) );
  AND2_X1 U8704 ( .A1(n6946), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8705 ( .A1(n6946), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8706 ( .A1(n6946), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8707 ( .A1(n6946), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8708 ( .A1(n6946), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8709 ( .A1(n6946), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8710 ( .A1(n6946), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8711 ( .A1(n6946), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8712 ( .A1(n6946), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8713 ( .A1(n6946), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8714 ( .A1(n6946), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8715 ( .A1(n6946), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8716 ( .A1(n6946), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8717 ( .A1(n6946), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8718 ( .A1(n6946), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8719 ( .A1(n6946), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  INV_X1 U8720 ( .A(n6947), .ZN(n6991) );
  AOI22_X1 U8721 ( .A1(n7033), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10315), .ZN(n6948) );
  OAI21_X1 U8722 ( .B1(n6991), .B2(n10335), .A(n6948), .ZN(P1_U3344) );
  INV_X1 U8723 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6949) );
  MUX2_X1 U8724 ( .A(n6949), .B(P1_REG1_REG_2__SCAN_IN), .S(n7106), .Z(n7100)
         );
  INV_X1 U8725 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6950) );
  MUX2_X1 U8726 ( .A(n6950), .B(P1_REG1_REG_1__SCAN_IN), .S(n6972), .Z(n9842)
         );
  AND2_X1 U8727 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9843) );
  NAND2_X1 U8728 ( .A1(n9842), .A2(n9843), .ZN(n9841) );
  OR2_X1 U8729 ( .A1(n6972), .A2(n6950), .ZN(n6951) );
  NAND2_X1 U8730 ( .A1(n9841), .A2(n6951), .ZN(n7101) );
  NAND2_X1 U8731 ( .A1(n7100), .A2(n7101), .ZN(n6953) );
  INV_X1 U8732 ( .A(n7106), .ZN(n6974) );
  NAND2_X1 U8733 ( .A1(n6974), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6952) );
  NAND2_X1 U8734 ( .A1(n6953), .A2(n6952), .ZN(n9858) );
  MUX2_X1 U8735 ( .A(n6954), .B(P1_REG1_REG_3__SCAN_IN), .S(n9852), .Z(n9859)
         );
  NAND2_X1 U8736 ( .A1(n9858), .A2(n9859), .ZN(n9873) );
  OR2_X1 U8737 ( .A1(n9852), .A2(n6954), .ZN(n9872) );
  NAND2_X1 U8738 ( .A1(n9873), .A2(n9872), .ZN(n6957) );
  INV_X1 U8739 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6955) );
  MUX2_X1 U8740 ( .A(n6955), .B(P1_REG1_REG_4__SCAN_IN), .S(n9870), .Z(n6956)
         );
  NAND2_X1 U8741 ( .A1(n6957), .A2(n6956), .ZN(n9889) );
  OR2_X1 U8742 ( .A1(n9870), .A2(n6955), .ZN(n9888) );
  NAND2_X1 U8743 ( .A1(n9889), .A2(n9888), .ZN(n6960) );
  MUX2_X1 U8744 ( .A(n6958), .B(P1_REG1_REG_5__SCAN_IN), .S(n9886), .Z(n6959)
         );
  NAND2_X1 U8745 ( .A1(n6960), .A2(n6959), .ZN(n9903) );
  INV_X1 U8746 ( .A(n9886), .ZN(n9882) );
  NAND2_X1 U8747 ( .A1(n9882), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9902) );
  NAND2_X1 U8748 ( .A1(n9903), .A2(n9902), .ZN(n6962) );
  MUX2_X1 U8749 ( .A(n6963), .B(P1_REG1_REG_6__SCAN_IN), .S(n9900), .Z(n6961)
         );
  NAND2_X1 U8750 ( .A1(n6962), .A2(n6961), .ZN(n9910) );
  OR2_X1 U8751 ( .A1(n9900), .A2(n6963), .ZN(n9909) );
  NAND2_X1 U8752 ( .A1(n9910), .A2(n9909), .ZN(n6965) );
  MUX2_X1 U8753 ( .A(n5571), .B(P1_REG1_REG_7__SCAN_IN), .S(n9916), .Z(n9908)
         );
  INV_X1 U8754 ( .A(n9908), .ZN(n6964) );
  NAND2_X1 U8755 ( .A1(n6965), .A2(n6964), .ZN(n9912) );
  NAND2_X1 U8756 ( .A1(n9916), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8757 ( .A1(n9912), .A2(n6966), .ZN(n6999) );
  INV_X1 U8758 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6967) );
  XNOR2_X1 U8759 ( .A(n7000), .B(n6967), .ZN(n6998) );
  XNOR2_X1 U8760 ( .A(n6999), .B(n6998), .ZN(n6990) );
  INV_X1 U8761 ( .A(n6985), .ZN(n9985) );
  NOR2_X2 U8762 ( .A1(n9985), .A2(n9807), .ZN(n9990) );
  INV_X1 U8763 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6968) );
  NAND2_X1 U8764 ( .A1(n10311), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9368) );
  OAI21_X1 U8765 ( .B1(n9994), .B2(n6968), .A(n9368), .ZN(n6969) );
  AOI21_X1 U8766 ( .B1(n7000), .B2(n9988), .A(n6969), .ZN(n6989) );
  INV_X1 U8767 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6970) );
  XNOR2_X1 U8768 ( .A(n7000), .B(n6970), .ZN(n6987) );
  INV_X1 U8769 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6971) );
  MUX2_X1 U8770 ( .A(n6971), .B(P1_REG2_REG_1__SCAN_IN), .S(n6972), .Z(n9847)
         );
  AND2_X1 U8771 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9846) );
  NAND2_X1 U8772 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  INV_X1 U8773 ( .A(n6972), .ZN(n9844) );
  NAND2_X1 U8774 ( .A1(n9844), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6973) );
  NAND2_X1 U8775 ( .A1(n9845), .A2(n6973), .ZN(n7103) );
  XNOR2_X1 U8776 ( .A(n7106), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7104) );
  NAND2_X1 U8777 ( .A1(n7103), .A2(n7104), .ZN(n7102) );
  NAND2_X1 U8778 ( .A1(n6974), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6975) );
  NAND2_X1 U8779 ( .A1(n7102), .A2(n6975), .ZN(n9856) );
  XNOR2_X1 U8780 ( .A(n9852), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9857) );
  INV_X1 U8781 ( .A(n9852), .ZN(n6976) );
  NAND2_X1 U8782 ( .A1(n6976), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8783 ( .A1(n9855), .A2(n6977), .ZN(n9868) );
  MUX2_X1 U8784 ( .A(n6978), .B(P1_REG2_REG_4__SCAN_IN), .S(n9870), .Z(n9869)
         );
  NAND2_X1 U8785 ( .A1(n9868), .A2(n9869), .ZN(n9867) );
  OR2_X1 U8786 ( .A1(n9870), .A2(n6978), .ZN(n6979) );
  NAND2_X1 U8787 ( .A1(n9867), .A2(n6979), .ZN(n9884) );
  XNOR2_X1 U8788 ( .A(n9886), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9885) );
  NAND2_X1 U8789 ( .A1(n9884), .A2(n9885), .ZN(n9883) );
  NAND2_X1 U8790 ( .A1(n9882), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8791 ( .A1(n9883), .A2(n6980), .ZN(n9898) );
  XNOR2_X1 U8792 ( .A(n9900), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9899) );
  OR2_X1 U8793 ( .A1(n9900), .A2(n6981), .ZN(n6982) );
  NAND2_X1 U8794 ( .A1(n9897), .A2(n6982), .ZN(n9918) );
  INV_X1 U8795 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8539) );
  MUX2_X1 U8796 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n8539), .S(n9916), .Z(n9919)
         );
  NAND2_X1 U8797 ( .A1(n9918), .A2(n9919), .ZN(n9917) );
  NAND2_X1 U8798 ( .A1(n9916), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6983) );
  NAND2_X1 U8799 ( .A1(n9917), .A2(n6983), .ZN(n6986) );
  NOR2_X1 U8800 ( .A1(n8005), .A2(n6924), .ZN(n6984) );
  NAND2_X1 U8801 ( .A1(n6985), .A2(n6984), .ZN(n9960) );
  OAI211_X1 U8802 ( .C1(n6987), .C2(n6986), .A(n9984), .B(n6994), .ZN(n6988)
         );
  OAI211_X1 U8803 ( .C1(n6990), .C2(n9939), .A(n6989), .B(n6988), .ZN(P1_U3251) );
  INV_X1 U8804 ( .A(n8383), .ZN(n8370) );
  OAI222_X1 U8805 ( .A1(n8134), .A2(n6992), .B1(n9307), .B2(n6991), .C1(
        P2_U3151), .C2(n8370), .ZN(P2_U3284) );
  NAND2_X1 U8806 ( .A1(n7000), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8807 ( .A1(n6994), .A2(n6993), .ZN(n7016) );
  XNOR2_X1 U8808 ( .A(n7025), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7017) );
  OR2_X1 U8809 ( .A1(n7025), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6995) );
  NAND2_X1 U8810 ( .A1(n7014), .A2(n6995), .ZN(n7046) );
  XNOR2_X1 U8811 ( .A(n7005), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U8812 ( .A1(n7046), .A2(n7047), .ZN(n7045) );
  XNOR2_X1 U8813 ( .A(n7033), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n6996) );
  AOI211_X1 U8814 ( .C1(n6997), .C2(n6996), .A(n9960), .B(n7028), .ZN(n7013)
         );
  NAND2_X1 U8815 ( .A1(n6999), .A2(n6998), .ZN(n7002) );
  NAND2_X1 U8816 ( .A1(n7000), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8817 ( .A1(n7002), .A2(n7001), .ZN(n7020) );
  MUX2_X1 U8818 ( .A(n7003), .B(P1_REG1_REG_9__SCAN_IN), .S(n7025), .Z(n7019)
         );
  OR2_X1 U8819 ( .A1(n7025), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8820 ( .A1(n7022), .A2(n7004), .ZN(n7044) );
  MUX2_X1 U8821 ( .A(n5646), .B(P1_REG1_REG_10__SCAN_IN), .S(n7005), .Z(n7043)
         );
  NAND2_X1 U8822 ( .A1(n7005), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7007) );
  MUX2_X1 U8823 ( .A(n5668), .B(P1_REG1_REG_11__SCAN_IN), .S(n7033), .Z(n7006)
         );
  AOI21_X1 U8824 ( .B1(n7041), .B2(n7007), .A(n7006), .ZN(n7032) );
  AND3_X1 U8825 ( .A1(n7041), .A2(n7007), .A3(n7006), .ZN(n7008) );
  NOR3_X1 U8826 ( .A1(n9939), .A2(n7032), .A3(n7008), .ZN(n7012) );
  INV_X1 U8827 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7010) );
  NAND2_X1 U8828 ( .A1(n9988), .A2(n7033), .ZN(n7009) );
  NAND2_X1 U8829 ( .A1(n10311), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9491) );
  OAI211_X1 U8830 ( .C1(n9994), .C2(n7010), .A(n7009), .B(n9491), .ZN(n7011)
         );
  OR3_X1 U8831 ( .A1(n7013), .A2(n7012), .A3(n7011), .ZN(P1_U3254) );
  INV_X1 U8832 ( .A(n7014), .ZN(n7015) );
  AOI21_X1 U8833 ( .B1(n7017), .B2(n7016), .A(n7015), .ZN(n7027) );
  INV_X1 U8834 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n7018) );
  NAND2_X1 U8835 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9448) );
  OAI21_X1 U8836 ( .B1(n9994), .B2(n7018), .A(n9448), .ZN(n7024) );
  NAND2_X1 U8837 ( .A1(n7020), .A2(n7019), .ZN(n7021) );
  AOI21_X1 U8838 ( .B1(n7022), .B2(n7021), .A(n9939), .ZN(n7023) );
  AOI211_X1 U8839 ( .C1(n9988), .C2(n7025), .A(n7024), .B(n7023), .ZN(n7026)
         );
  OAI21_X1 U8840 ( .B1(n7027), .B2(n9960), .A(n7026), .ZN(P1_U3252) );
  XNOR2_X1 U8841 ( .A(n7252), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n7030) );
  AOI21_X1 U8842 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n7033), .A(n7028), .ZN(
        n7029) );
  OAI21_X1 U8843 ( .B1(n7030), .B2(n7029), .A(n7248), .ZN(n7031) );
  NAND2_X1 U8844 ( .A1(n7031), .A2(n9984), .ZN(n7040) );
  XNOR2_X1 U8845 ( .A(n7252), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7035) );
  AOI21_X1 U8846 ( .B1(n7033), .B2(P1_REG1_REG_11__SCAN_IN), .A(n7032), .ZN(
        n7034) );
  NAND2_X1 U8847 ( .A1(n7034), .A2(n7035), .ZN(n7255) );
  OAI21_X1 U8848 ( .B1(n7035), .B2(n7034), .A(n7255), .ZN(n7038) );
  INV_X1 U8849 ( .A(n9988), .ZN(n9975) );
  NAND2_X1 U8850 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9391) );
  NAND2_X1 U8851 ( .A1(n9965), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n7036) );
  OAI211_X1 U8852 ( .C1(n9975), .C2(n7252), .A(n9391), .B(n7036), .ZN(n7037)
         );
  AOI21_X1 U8853 ( .B1(n7038), .B2(n9990), .A(n7037), .ZN(n7039) );
  NAND2_X1 U8854 ( .A1(n7040), .A2(n7039), .ZN(P1_U3255) );
  INV_X1 U8855 ( .A(n7041), .ZN(n7042) );
  AOI211_X1 U8856 ( .C1(n7044), .C2(n7043), .A(n7042), .B(n9939), .ZN(n7052)
         );
  AOI211_X1 U8857 ( .C1(n7047), .C2(n7046), .A(n9960), .B(n7045), .ZN(n7051)
         );
  NAND2_X1 U8858 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U8859 ( .A1(n9965), .A2(P1_ADDR_REG_10__SCAN_IN), .ZN(n7048) );
  OAI211_X1 U8860 ( .C1(n9975), .C2(n7049), .A(n9332), .B(n7048), .ZN(n7050)
         );
  OR3_X1 U8861 ( .A1(n7052), .A2(n7051), .A3(n7050), .ZN(P1_U3253) );
  NAND2_X1 U8862 ( .A1(n10409), .A2(n7606), .ZN(n10407) );
  INV_X1 U8863 ( .A(n7053), .ZN(n7054) );
  NAND2_X1 U8864 ( .A1(n7054), .A2(P1_D_REG_1__SCAN_IN), .ZN(n7055) );
  NAND2_X1 U8865 ( .A1(n7056), .A2(n7055), .ZN(n7058) );
  NAND2_X1 U8866 ( .A1(n7058), .A2(n7057), .ZN(n7605) );
  NAND2_X1 U8867 ( .A1(n7059), .A2(n4613), .ZN(n7611) );
  OR2_X1 U8868 ( .A1(n7087), .A2(n7611), .ZN(n7062) );
  INV_X1 U8869 ( .A(n10409), .ZN(n7061) );
  NAND2_X1 U8870 ( .A1(n7065), .A2(n9991), .ZN(n7635) );
  NAND2_X1 U8871 ( .A1(n7198), .A2(n7141), .ZN(n7070) );
  NAND2_X1 U8872 ( .A1(n9840), .A2(n8108), .ZN(n7069) );
  NAND2_X1 U8873 ( .A1(n7072), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U8874 ( .A1(n9342), .A2(n9840), .ZN(n7074) );
  AOI22_X1 U8875 ( .A1(n8108), .A2(n7141), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n7072), .ZN(n7073) );
  NAND2_X1 U8876 ( .A1(n7074), .A2(n7073), .ZN(n7110) );
  NAND2_X1 U8877 ( .A1(n7111), .A2(n7110), .ZN(n7076) );
  NAND2_X1 U8878 ( .A1(n7076), .A2(n7075), .ZN(n7121) );
  NAND2_X1 U8879 ( .A1(n5464), .A2(n8108), .ZN(n7078) );
  NAND2_X1 U8880 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  AOI22_X1 U8881 ( .A1(n9342), .A2(n5464), .B1(n5458), .B2(n4427), .ZN(n7082)
         );
  NAND2_X1 U8882 ( .A1(n7081), .A2(n7082), .ZN(n7120) );
  INV_X1 U8883 ( .A(n7081), .ZN(n7084) );
  INV_X1 U8884 ( .A(n7082), .ZN(n7083) );
  NAND2_X1 U8885 ( .A1(n7084), .A2(n7083), .ZN(n7122) );
  NAND2_X1 U8886 ( .A1(n7120), .A2(n7122), .ZN(n7085) );
  XNOR2_X1 U8887 ( .A(n7121), .B(n7085), .ZN(n7086) );
  NAND2_X1 U8888 ( .A1(n7086), .A2(n9533), .ZN(n7092) );
  NAND2_X1 U8889 ( .A1(n4420), .A2(n9840), .ZN(n7089) );
  NAND2_X1 U8890 ( .A1(n9551), .A2(n5482), .ZN(n7088) );
  NAND2_X1 U8891 ( .A1(n7089), .A2(n7088), .ZN(n7722) );
  NOR2_X1 U8892 ( .A1(n9784), .A2(P1_U3086), .ZN(n7814) );
  OAI22_X1 U8893 ( .A1(n10473), .A2(n7814), .B1(n7090), .B2(n7605), .ZN(n7206)
         );
  NAND2_X1 U8894 ( .A1(n7608), .A2(n7206), .ZN(n7138) );
  AOI22_X1 U8895 ( .A1(n9542), .A2(n7722), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n7138), .ZN(n7091) );
  OAI211_X1 U8896 ( .C1(n10414), .C2(n9545), .A(n7092), .B(n7091), .ZN(
        P1_U3222) );
  INV_X1 U8897 ( .A(n8408), .ZN(n8400) );
  INV_X1 U8898 ( .A(n7093), .ZN(n7094) );
  OAI222_X1 U8899 ( .A1(P2_U3151), .A2(n8400), .B1(n9307), .B2(n7094), .C1(
        n8549), .C2(n8134), .ZN(P2_U3283) );
  OAI222_X1 U8900 ( .A1(n10332), .A2(n7095), .B1(n10335), .B2(n7094), .C1(
        n7252), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8901 ( .A(n8424), .ZN(n8420) );
  INV_X1 U8902 ( .A(n7096), .ZN(n7098) );
  INV_X1 U8903 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7097) );
  OAI222_X1 U8904 ( .A1(n8420), .A2(P2_U3151), .B1(n9307), .B2(n7098), .C1(
        n7097), .C2(n8134), .ZN(P2_U3282) );
  INV_X1 U8905 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7099) );
  INV_X1 U8906 ( .A(n7392), .ZN(n7388) );
  OAI222_X1 U8907 ( .A1(n10332), .A2(n7099), .B1(n10335), .B2(n7098), .C1(
        n10311), .C2(n7388), .ZN(P1_U3342) );
  XOR2_X1 U8908 ( .A(n7101), .B(n7100), .Z(n7109) );
  INV_X1 U8909 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U8910 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n10311), .ZN(n8699) );
  OAI21_X1 U8911 ( .B1(n9994), .B2(n8605), .A(n8699), .ZN(n7108) );
  OAI211_X1 U8912 ( .C1(n7104), .C2(n7103), .A(n9984), .B(n7102), .ZN(n7105)
         );
  OAI21_X1 U8913 ( .B1(n9975), .B2(n7106), .A(n7105), .ZN(n7107) );
  AOI211_X1 U8914 ( .C1(n9990), .C2(n7109), .A(n7108), .B(n7107), .ZN(n7116)
         );
  XNOR2_X1 U8915 ( .A(n7111), .B(n7110), .ZN(n7143) );
  MUX2_X1 U8916 ( .A(n9846), .B(n7143), .S(n6924), .Z(n7113) );
  NAND2_X1 U8917 ( .A1(n7113), .A2(n7112), .ZN(n7114) );
  OAI211_X1 U8918 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n7115), .A(n7114), .B(
        P1_U3973), .ZN(n9878) );
  NAND2_X1 U8919 ( .A1(n7116), .A2(n9878), .ZN(P1_U3245) );
  NAND2_X1 U8920 ( .A1(n7198), .A2(n5481), .ZN(n7118) );
  NAND2_X1 U8921 ( .A1(n5482), .A2(n8108), .ZN(n7117) );
  NAND2_X1 U8922 ( .A1(n7118), .A2(n7117), .ZN(n7119) );
  AOI22_X1 U8923 ( .A1(n9342), .A2(n5482), .B1(n5481), .B2(n4427), .ZN(n7195)
         );
  AOI21_X1 U8924 ( .B1(n7125), .B2(n7124), .A(n7123), .ZN(n7128) );
  OAI22_X1 U8925 ( .A1(n7201), .A2(n9537), .B1(n9535), .B2(n5459), .ZN(n7705)
         );
  AOI22_X1 U8926 ( .A1(n9542), .A2(n7705), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n7138), .ZN(n7127) );
  NAND2_X1 U8927 ( .A1(n9557), .A2(n5481), .ZN(n7126) );
  OAI211_X1 U8928 ( .C1(n7128), .C2(n9559), .A(n7127), .B(n7126), .ZN(P1_U3237) );
  INV_X1 U8929 ( .A(n7337), .ZN(n7131) );
  NAND2_X1 U8930 ( .A1(n8294), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7155) );
  NAND2_X1 U8931 ( .A1(n7155), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7130) );
  AOI22_X1 U8932 ( .A1(n8316), .A2(n7344), .B1(n8310), .B2(n8340), .ZN(n7129)
         );
  OAI211_X1 U8933 ( .C1(n7131), .C2(n8318), .A(n7130), .B(n7129), .ZN(P2_U3172) );
  INV_X1 U8934 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7133) );
  INV_X1 U8935 ( .A(n7132), .ZN(n7135) );
  INV_X1 U8936 ( .A(n7582), .ZN(n7390) );
  OAI222_X1 U8937 ( .A1(n10332), .A2(n7133), .B1(n10335), .B2(n7135), .C1(
        P1_U3086), .C2(n7390), .ZN(P1_U3341) );
  INV_X1 U8938 ( .A(n8448), .ZN(n8442) );
  INV_X1 U8939 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7134) );
  OAI222_X1 U8940 ( .A1(n8442), .A2(P2_U3151), .B1(n9307), .B2(n7135), .C1(
        n7134), .C2(n8134), .ZN(P2_U3281) );
  INV_X1 U8941 ( .A(n9431), .ZN(n7136) );
  NAND2_X1 U8942 ( .A1(n7136), .A2(P1_U3973), .ZN(n7137) );
  OAI21_X1 U8943 ( .B1(P1_U3973), .B2(n5888), .A(n7137), .ZN(P1_U3577) );
  NAND2_X1 U8944 ( .A1(n9522), .A2(n5464), .ZN(n10251) );
  INV_X1 U8945 ( .A(n7138), .ZN(n7139) );
  INV_X1 U8946 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7614) );
  OAI22_X1 U8947 ( .A1(n9552), .A2(n10251), .B1(n7139), .B2(n7614), .ZN(n7140)
         );
  AOI21_X1 U8948 ( .B1(n7141), .B2(n9557), .A(n7140), .ZN(n7142) );
  OAI21_X1 U8949 ( .B1(n9559), .B2(n7143), .A(n7142), .ZN(P1_U3232) );
  AOI21_X1 U8950 ( .B1(n7146), .B2(n7145), .A(n7144), .ZN(n7150) );
  AOI22_X1 U8951 ( .A1(n8310), .A2(n8339), .B1(n8324), .B2(n6239), .ZN(n7147)
         );
  OAI21_X1 U8952 ( .B1(n8332), .B2(n6803), .A(n7147), .ZN(n7148) );
  AOI21_X1 U8953 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7155), .A(n7148), .ZN(
        n7149) );
  OAI21_X1 U8954 ( .B1(n7150), .B2(n8318), .A(n7149), .ZN(P2_U3162) );
  AOI21_X1 U8955 ( .B1(n7152), .B2(n7151), .A(n7377), .ZN(n7157) );
  AOI22_X1 U8956 ( .A1(n8310), .A2(n6694), .B1(n8324), .B2(n8340), .ZN(n7153)
         );
  OAI21_X1 U8957 ( .B1(n8332), .B2(n7357), .A(n7153), .ZN(n7154) );
  AOI21_X1 U8958 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7155), .A(n7154), .ZN(
        n7156) );
  OAI21_X1 U8959 ( .B1(n7157), .B2(n8318), .A(n7156), .ZN(P2_U3177) );
  MUX2_X1 U8960 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8770), .Z(n7163) );
  INV_X1 U8961 ( .A(n7163), .ZN(n7164) );
  MUX2_X1 U8962 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8770), .Z(n7161) );
  INV_X1 U8963 ( .A(n7161), .ZN(n7162) );
  INV_X1 U8964 ( .A(n7158), .ZN(n7160) );
  INV_X1 U8965 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7179) );
  MUX2_X1 U8966 ( .A(n7179), .B(n7159), .S(n8770), .Z(n7320) );
  NAND2_X1 U8967 ( .A1(n7320), .A2(n4848), .ZN(n7319) );
  XNOR2_X1 U8968 ( .A(n7161), .B(n7175), .ZN(n7224) );
  NAND2_X1 U8969 ( .A1(n7225), .A2(n7224), .ZN(n7223) );
  XOR2_X1 U8970 ( .A(n10506), .B(n7163), .Z(n10509) );
  NOR2_X1 U8971 ( .A1(n10508), .A2(n10509), .ZN(n10507) );
  MUX2_X1 U8972 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8770), .Z(n7239) );
  XNOR2_X1 U8973 ( .A(n7239), .B(n7242), .ZN(n7165) );
  OAI211_X1 U8974 ( .C1(n7166), .C2(n7165), .A(n7240), .B(n8797), .ZN(n7194)
         );
  NAND2_X1 U8975 ( .A1(n7167), .A2(n7170), .ZN(n7172) );
  NAND2_X1 U8976 ( .A1(n8788), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9306) );
  OR2_X1 U8977 ( .A1(n7172), .A2(n9306), .ZN(n7169) );
  INV_X1 U8978 ( .A(n8795), .ZN(n10505) );
  INV_X1 U8979 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7171) );
  NAND2_X1 U8980 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7406) );
  OAI21_X1 U8981 ( .B1(n8778), .B2(n7171), .A(n7406), .ZN(n7192) );
  OR2_X1 U8982 ( .A1(n6676), .A2(P2_U3151), .ZN(n9302) );
  INV_X1 U8983 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10554) );
  MUX2_X1 U8984 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10554), .S(n7242), .Z(n7178)
         );
  NAND2_X1 U8985 ( .A1(n4470), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7173) );
  INV_X1 U8986 ( .A(n7176), .ZN(n7177) );
  NOR2_X1 U8987 ( .A1(n7179), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7180) );
  INV_X1 U8988 ( .A(n7181), .ZN(n7182) );
  NOR2_X1 U8989 ( .A1(n7217), .A2(n7218), .ZN(n7216) );
  NOR2_X1 U8990 ( .A1(n7216), .A2(n7184), .ZN(n7185) );
  NAND2_X1 U8991 ( .A1(n7229), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7230) );
  OAI21_X1 U8992 ( .B1(n7229), .B2(P2_REG2_REG_4__SCAN_IN), .A(n7230), .ZN(
        n7186) );
  AOI21_X1 U8993 ( .B1(n7187), .B2(n7186), .A(n7232), .ZN(n7189) );
  INV_X1 U8994 ( .A(n7318), .ZN(n7188) );
  NAND2_X1 U8995 ( .A1(n7188), .A2(n8788), .ZN(n10503) );
  OAI22_X1 U8996 ( .A1(n8781), .A2(n7190), .B1(n7189), .B2(n10503), .ZN(n7191)
         );
  AOI211_X1 U8997 ( .C1(n7242), .C2(n10505), .A(n7192), .B(n7191), .ZN(n7193)
         );
  NAND2_X1 U8998 ( .A1(n7194), .A2(n7193), .ZN(P2_U3186) );
  NAND2_X1 U8999 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  NAND2_X1 U9000 ( .A1(n8137), .A2(n7203), .ZN(n7199) );
  OAI21_X1 U9001 ( .B1(n7201), .B2(n5421), .A(n7199), .ZN(n7200) );
  XNOR2_X1 U9002 ( .A(n7200), .B(n8141), .ZN(n7284) );
  OAI22_X1 U9003 ( .A1(n7201), .A2(n8165), .B1(n10426), .B2(n5421), .ZN(n7285)
         );
  XNOR2_X1 U9004 ( .A(n7284), .B(n7285), .ZN(n7287) );
  XOR2_X1 U9005 ( .A(n7288), .B(n7287), .Z(n7210) );
  INV_X1 U9006 ( .A(n5482), .ZN(n7202) );
  OAI22_X1 U9007 ( .A1(n7202), .A2(n9535), .B1(n9537), .B2(n7291), .ZN(n7633)
         );
  AOI22_X1 U9008 ( .A1(n9557), .A2(n7203), .B1(n9542), .B2(n7633), .ZN(n7209)
         );
  NAND4_X1 U9009 ( .A1(n7206), .A2(n7866), .A3(n7205), .A4(n7204), .ZN(n7207)
         );
  MUX2_X1 U9010 ( .A(n9554), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n7208) );
  OAI211_X1 U9011 ( .C1(n7210), .C2(n9559), .A(n7209), .B(n7208), .ZN(P1_U3218) );
  INV_X1 U9012 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8502) );
  OAI21_X1 U9013 ( .B1(n10544), .B2(n9061), .A(n7337), .ZN(n7211) );
  OR2_X1 U9014 ( .A1(n7352), .A2(n9008), .ZN(n7338) );
  OAI211_X1 U9015 ( .C1(n10537), .C2(n7212), .A(n7211), .B(n7338), .ZN(n9176)
         );
  NAND2_X1 U9016 ( .A1(n10548), .A2(n9176), .ZN(n7213) );
  OAI21_X1 U9017 ( .B1(n10548), .B2(n8502), .A(n7213), .ZN(P2_U3390) );
  NOR2_X1 U9018 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6246), .ZN(n7222) );
  XOR2_X1 U9019 ( .A(n7215), .B(n7214), .Z(n7220) );
  AOI21_X1 U9020 ( .B1(n7218), .B2(n7217), .A(n7216), .ZN(n7219) );
  OAI22_X1 U9021 ( .A1(n8781), .A2(n7220), .B1(n7219), .B2(n10503), .ZN(n7221)
         );
  AOI211_X1 U9022 ( .C1(n10513), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n7222), .B(
        n7221), .ZN(n7227) );
  OAI211_X1 U9023 ( .C1(n7225), .C2(n7224), .A(n7223), .B(n8797), .ZN(n7226)
         );
  OAI211_X1 U9024 ( .C1(n8795), .C2(n7183), .A(n7227), .B(n7226), .ZN(P2_U3184) );
  XNOR2_X1 U9025 ( .A(n7271), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7247) );
  INV_X1 U9026 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n7237) );
  INV_X1 U9027 ( .A(n7230), .ZN(n7231) );
  OAI21_X1 U9028 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7234), .A(n7275), .ZN(
        n7235) );
  INV_X1 U9029 ( .A(n10503), .ZN(n8763) );
  NAND2_X1 U9030 ( .A1(n7235), .A2(n8763), .ZN(n7236) );
  NAND2_X1 U9031 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7501) );
  OAI211_X1 U9032 ( .C1(n8778), .C2(n7237), .A(n7236), .B(n7501), .ZN(n7238)
         );
  AOI21_X1 U9033 ( .B1(n7269), .B2(n10505), .A(n7238), .ZN(n7246) );
  INV_X1 U9034 ( .A(n7239), .ZN(n7241) );
  MUX2_X1 U9035 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8770), .Z(n7263) );
  XNOR2_X1 U9036 ( .A(n7263), .B(n7269), .ZN(n7243) );
  OAI211_X1 U9037 ( .C1(n7244), .C2(n7243), .A(n7264), .B(n8797), .ZN(n7245)
         );
  OAI211_X1 U9038 ( .C1(n7247), .C2(n8781), .A(n7246), .B(n7245), .ZN(P2_U3187) );
  XNOR2_X1 U9039 ( .A(n7392), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n7251) );
  NOR2_X1 U9040 ( .A1(n7250), .A2(n7251), .ZN(n7391) );
  AOI211_X1 U9041 ( .C1(n7251), .C2(n7250), .A(n9960), .B(n7391), .ZN(n7262)
         );
  XOR2_X1 U9042 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7392), .Z(n7253) );
  NAND2_X1 U9043 ( .A1(n7252), .A2(n10241), .ZN(n7254) );
  NAND3_X1 U9044 ( .A1(n7255), .A2(n7253), .A3(n7254), .ZN(n7387) );
  INV_X1 U9045 ( .A(n7387), .ZN(n7257) );
  AOI21_X1 U9046 ( .B1(n7255), .B2(n7254), .A(n7253), .ZN(n7256) );
  NOR3_X1 U9047 ( .A1(n7257), .A2(n7256), .A3(n9939), .ZN(n7261) );
  INV_X1 U9048 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7259) );
  NAND2_X1 U9049 ( .A1(n9988), .A2(n7392), .ZN(n7258) );
  NAND2_X1 U9050 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9467) );
  OAI211_X1 U9051 ( .C1(n9994), .C2(n7259), .A(n7258), .B(n9467), .ZN(n7260)
         );
  OR3_X1 U9052 ( .A1(n7262), .A2(n7261), .A3(n7260), .ZN(P1_U3256) );
  MUX2_X1 U9053 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8770), .Z(n7567) );
  XOR2_X1 U9054 ( .A(n7570), .B(n7567), .Z(n7267) );
  INV_X1 U9055 ( .A(n7263), .ZN(n7265) );
  OAI21_X1 U9056 ( .B1(n7269), .B2(n7265), .A(n7264), .ZN(n7266) );
  AOI21_X1 U9057 ( .B1(n7267), .B2(n7266), .A(n7568), .ZN(n7283) );
  INV_X1 U9058 ( .A(n8797), .ZN(n10510) );
  XNOR2_X1 U9059 ( .A(n7570), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n7551) );
  XNOR2_X1 U9060 ( .A(n7552), .B(n7551), .ZN(n7281) );
  NOR2_X1 U9061 ( .A1(n8795), .A2(n7557), .ZN(n7280) );
  INV_X1 U9062 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7278) );
  INV_X1 U9063 ( .A(n7272), .ZN(n7273) );
  XNOR2_X1 U9064 ( .A(n7570), .B(n7440), .ZN(n7274) );
  AND3_X1 U9065 ( .A1(n7275), .A2(n7274), .A3(n7273), .ZN(n7276) );
  OAI21_X1 U9066 ( .B1(n7556), .B2(n7276), .A(n8763), .ZN(n7277) );
  NAND2_X1 U9067 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7450) );
  OAI211_X1 U9068 ( .C1(n8778), .C2(n7278), .A(n7277), .B(n7450), .ZN(n7279)
         );
  AOI211_X1 U9069 ( .C1(n10499), .C2(n7281), .A(n7280), .B(n7279), .ZN(n7282)
         );
  OAI21_X1 U9070 ( .B1(n7283), .B2(n10510), .A(n7282), .ZN(P2_U3188) );
  INV_X1 U9071 ( .A(n7284), .ZN(n7286) );
  NAND2_X1 U9072 ( .A1(n8137), .A2(n7298), .ZN(n7289) );
  OAI21_X1 U9073 ( .B1(n7291), .B2(n5421), .A(n7289), .ZN(n7290) );
  XNOR2_X1 U9074 ( .A(n7290), .B(n8141), .ZN(n7457) );
  OAI22_X1 U9075 ( .A1(n7291), .A2(n8165), .B1(n10432), .B2(n5421), .ZN(n7458)
         );
  XNOR2_X1 U9076 ( .A(n7457), .B(n7458), .ZN(n7292) );
  OAI211_X1 U9077 ( .C1(n7293), .C2(n7292), .A(n7461), .B(n9533), .ZN(n7300)
         );
  NAND2_X1 U9078 ( .A1(n9838), .A2(n4420), .ZN(n7295) );
  NAND2_X1 U9079 ( .A1(n9836), .A2(n9522), .ZN(n7294) );
  AND2_X1 U9080 ( .A1(n7295), .A2(n7294), .ZN(n10375) );
  NAND2_X1 U9081 ( .A1(n10311), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9863) );
  OR2_X1 U9082 ( .A1(n9554), .A2(n10379), .ZN(n7296) );
  OAI211_X1 U9083 ( .C1(n9552), .C2(n10375), .A(n9863), .B(n7296), .ZN(n7297)
         );
  AOI21_X1 U9084 ( .B1(n7298), .B2(n9557), .A(n7297), .ZN(n7299) );
  NAND2_X1 U9085 ( .A1(n7300), .A2(n7299), .ZN(P1_U3230) );
  INV_X1 U9086 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7302) );
  INV_X1 U9087 ( .A(n7301), .ZN(n7304) );
  INV_X1 U9088 ( .A(n7583), .ZN(n9928) );
  OAI222_X1 U9089 ( .A1(n10332), .A2(n7302), .B1(n10335), .B2(n7304), .C1(
        n10311), .C2(n9928), .ZN(P1_U3340) );
  INV_X1 U9090 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7303) );
  OAI222_X1 U9091 ( .A1(n5101), .A2(P2_U3151), .B1(n9307), .B2(n7304), .C1(
        n7303), .C2(n8134), .ZN(P2_U3280) );
  XNOR2_X1 U9092 ( .A(n4574), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n7308) );
  OAI211_X1 U9093 ( .C1(n7306), .C2(n7319), .A(n7305), .B(n8797), .ZN(n7307)
         );
  OAI21_X1 U9094 ( .B1(n8781), .B2(n7308), .A(n7307), .ZN(n7315) );
  AOI21_X1 U9095 ( .B1(n7962), .B2(n7310), .A(n7309), .ZN(n7311) );
  NOR2_X1 U9096 ( .A1(n10503), .A2(n7311), .ZN(n7314) );
  OAI22_X1 U9097 ( .A1(n8778), .A2(n10562), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7312), .ZN(n7313) );
  NOR3_X1 U9098 ( .A1(n7315), .A2(n7314), .A3(n7313), .ZN(n7316) );
  OAI21_X1 U9099 ( .B1(n7317), .B2(n8795), .A(n7316), .ZN(P2_U3183) );
  INV_X1 U9100 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7325) );
  NAND2_X1 U9101 ( .A1(n10505), .A2(n4848), .ZN(n7324) );
  NAND2_X1 U9102 ( .A1(n7318), .A2(n10510), .ZN(n7322) );
  OAI21_X1 U9103 ( .B1(n4848), .B2(n7320), .A(n7319), .ZN(n7321) );
  AOI22_X1 U9104 ( .A1(n7322), .A2(n7321), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n7323) );
  OAI211_X1 U9105 ( .C1(n8778), .C2(n7325), .A(n7324), .B(n7323), .ZN(P2_U3182) );
  NAND2_X1 U9106 ( .A1(n8857), .A2(P2_U3893), .ZN(n7326) );
  OAI21_X1 U9107 ( .B1(P2_U3893), .B2(n5893), .A(n7326), .ZN(P2_U3514) );
  INV_X1 U9108 ( .A(n8479), .ZN(n8487) );
  INV_X1 U9109 ( .A(n7327), .ZN(n7328) );
  OAI222_X1 U9110 ( .A1(P2_U3151), .A2(n8487), .B1(n9307), .B2(n7328), .C1(
        n8654), .C2(n8134), .ZN(P2_U3279) );
  INV_X1 U9111 ( .A(n9942), .ZN(n9945) );
  OAI222_X1 U9112 ( .A1(n10332), .A2(n7329), .B1(n10311), .B2(n9945), .C1(
        n7328), .C2(n10335), .ZN(P1_U3339) );
  OR2_X1 U9113 ( .A1(n7332), .A2(n7330), .ZN(n7335) );
  INV_X1 U9114 ( .A(n6758), .ZN(n7331) );
  NAND2_X1 U9115 ( .A1(n7332), .A2(n7331), .ZN(n7334) );
  NAND3_X1 U9116 ( .A1(n7335), .A2(n7334), .A3(n7333), .ZN(n7341) );
  NAND3_X1 U9117 ( .A1(n7337), .A2(n7336), .A3(n10537), .ZN(n7339) );
  OAI211_X1 U9118 ( .C1(n9087), .C2(n7340), .A(n7339), .B(n7338), .ZN(n7342)
         );
  MUX2_X1 U9119 ( .A(n7342), .B(P2_REG2_REG_0__SCAN_IN), .S(n8981), .Z(n7343)
         );
  AOI21_X1 U9120 ( .B1(n9029), .B2(n7344), .A(n7343), .ZN(n7345) );
  INV_X1 U9121 ( .A(n7345), .ZN(P2_U3233) );
  XNOR2_X1 U9122 ( .A(n7346), .B(n7350), .ZN(n10519) );
  NAND2_X1 U9123 ( .A1(n10519), .A2(n4725), .ZN(n7356) );
  NAND3_X1 U9124 ( .A1(n7350), .A2(n7349), .A3(n7348), .ZN(n7351) );
  NAND2_X1 U9125 ( .A1(n7347), .A2(n7351), .ZN(n7354) );
  OAI22_X1 U9126 ( .A1(n9010), .A2(n7352), .B1(n7375), .B2(n9008), .ZN(n7353)
         );
  AOI21_X1 U9127 ( .B1(n7354), .B2(n9061), .A(n7353), .ZN(n7355) );
  AND2_X1 U9128 ( .A1(n7356), .A2(n7355), .ZN(n10523) );
  NOR2_X1 U9129 ( .A1(n7357), .A2(n10537), .ZN(n10517) );
  AOI21_X1 U9130 ( .B1(n10519), .B2(n9169), .A(n10517), .ZN(n7358) );
  AND2_X1 U9131 ( .A1(n10523), .A2(n7358), .ZN(n10530) );
  MUX2_X1 U9132 ( .A(n10530), .B(n4682), .S(n6883), .Z(n7359) );
  INV_X1 U9133 ( .A(n7359), .ZN(P2_U3461) );
  NAND2_X1 U9134 ( .A1(n7360), .A2(n4435), .ZN(n7956) );
  AND2_X1 U9135 ( .A1(n9069), .A2(n7956), .ZN(n7361) );
  XNOR2_X1 U9136 ( .A(n7365), .B(n7362), .ZN(n10535) );
  INV_X1 U9137 ( .A(n10535), .ZN(n7372) );
  NAND3_X1 U9138 ( .A1(n7347), .A2(n7365), .A3(n7364), .ZN(n7366) );
  NAND2_X1 U9139 ( .A1(n7363), .A2(n7366), .ZN(n7368) );
  AOI222_X1 U9140 ( .A1(n9061), .A2(n7368), .B1(n7367), .B2(n9065), .C1(n8339), 
        .C2(n9064), .ZN(n10532) );
  INV_X2 U9141 ( .A(n8981), .ZN(n9091) );
  MUX2_X1 U9142 ( .A(n10496), .B(n10532), .S(n9091), .Z(n7371) );
  AOI22_X1 U9143 ( .A1(n9029), .A2(n7369), .B1(n10518), .B2(n7384), .ZN(n7370)
         );
  OAI211_X1 U9144 ( .C1(n9086), .C2(n7372), .A(n7371), .B(n7370), .ZN(P2_U3230) );
  NAND2_X1 U9145 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10500) );
  OAI21_X1 U9146 ( .B1(n8313), .B2(n7958), .A(n10500), .ZN(n7373) );
  AOI21_X1 U9147 ( .B1(n8310), .B2(n7367), .A(n7373), .ZN(n7374) );
  OAI21_X1 U9148 ( .B1(n10533), .B2(n8332), .A(n7374), .ZN(n7383) );
  XNOR2_X1 U9149 ( .A(n7376), .B(n7375), .ZN(n7381) );
  INV_X1 U9150 ( .A(n7377), .ZN(n7379) );
  NAND2_X1 U9151 ( .A1(n7379), .A2(n7378), .ZN(n7380) );
  NOR2_X1 U9152 ( .A1(n7380), .A2(n7381), .ZN(n7400) );
  AOI211_X1 U9153 ( .C1(n7381), .C2(n7380), .A(n8318), .B(n7400), .ZN(n7382)
         );
  AOI211_X1 U9154 ( .C1(n7384), .C2(n8329), .A(n7383), .B(n7382), .ZN(n7385)
         );
  INV_X1 U9155 ( .A(n7385), .ZN(P2_U3158) );
  INV_X1 U9156 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7386) );
  XNOR2_X1 U9157 ( .A(n7582), .B(n7386), .ZN(n7579) );
  OAI21_X1 U9158 ( .B1(n7388), .B2(n10236), .A(n7387), .ZN(n7580) );
  XOR2_X1 U9159 ( .A(n7579), .B(n7580), .Z(n7397) );
  NAND2_X1 U9160 ( .A1(n10311), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9320) );
  NAND2_X1 U9161 ( .A1(n9965), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n7389) );
  OAI211_X1 U9162 ( .C1(n9975), .C2(n7390), .A(n9320), .B(n7389), .ZN(n7396)
         );
  XNOR2_X1 U9163 ( .A(n7582), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n7393) );
  AOI211_X1 U9164 ( .C1(n7394), .C2(n7393), .A(n9960), .B(n7581), .ZN(n7395)
         );
  AOI211_X1 U9165 ( .C1(n9990), .C2(n7397), .A(n7396), .B(n7395), .ZN(n7398)
         );
  INV_X1 U9166 ( .A(n7398), .ZN(P1_U3257) );
  NOR2_X1 U9167 ( .A1(n7400), .A2(n7399), .ZN(n7404) );
  INV_X1 U9168 ( .A(n7506), .ZN(n7401) );
  NOR2_X1 U9169 ( .A1(n7402), .A2(n7401), .ZN(n7403) );
  NAND2_X1 U9170 ( .A1(n7404), .A2(n7403), .ZN(n7508) );
  OAI21_X1 U9171 ( .B1(n7404), .B2(n7403), .A(n7508), .ZN(n7405) );
  NAND2_X1 U9172 ( .A1(n7405), .A2(n8320), .ZN(n7410) );
  NAND2_X1 U9173 ( .A1(n8324), .A2(n6694), .ZN(n7407) );
  OAI211_X1 U9174 ( .C1(n4812), .C2(n8326), .A(n7407), .B(n7406), .ZN(n7408)
         );
  AOI21_X1 U9175 ( .B1(n7421), .B2(n8316), .A(n7408), .ZN(n7409) );
  OAI211_X1 U9176 ( .C1(n7419), .C2(n8294), .A(n7410), .B(n7409), .ZN(P2_U3170) );
  XNOR2_X1 U9177 ( .A(n7411), .B(n7415), .ZN(n10540) );
  INV_X1 U9178 ( .A(n10540), .ZN(n7424) );
  NAND2_X1 U9179 ( .A1(n7363), .A2(n7414), .ZN(n7413) );
  NAND2_X1 U9180 ( .A1(n7413), .A2(n7412), .ZN(n7490) );
  NAND3_X1 U9181 ( .A1(n7363), .A2(n7415), .A3(n7414), .ZN(n7416) );
  NAND2_X1 U9182 ( .A1(n7490), .A2(n7416), .ZN(n7417) );
  AOI222_X1 U9183 ( .A1(n9061), .A2(n7417), .B1(n6694), .B2(n9064), .C1(n8338), 
        .C2(n9065), .ZN(n10536) );
  MUX2_X1 U9184 ( .A(n7418), .B(n10536), .S(n9091), .Z(n7423) );
  INV_X1 U9185 ( .A(n7419), .ZN(n7420) );
  AOI22_X1 U9186 ( .A1(n9029), .A2(n7421), .B1(n10518), .B2(n7420), .ZN(n7422)
         );
  OAI211_X1 U9187 ( .C1(n9086), .C2(n7424), .A(n7423), .B(n7422), .ZN(P2_U3229) );
  INV_X1 U9188 ( .A(n7425), .ZN(n7427) );
  XNOR2_X1 U9189 ( .A(n7427), .B(n7426), .ZN(n7428) );
  AOI222_X1 U9190 ( .A1(n9061), .A2(n7428), .B1(n8336), .B2(n9065), .C1(n8338), 
        .C2(n9064), .ZN(n7439) );
  NAND2_X1 U9191 ( .A1(n7429), .A2(n7492), .ZN(n7488) );
  NAND2_X1 U9192 ( .A1(n7488), .A2(n7430), .ZN(n7432) );
  XNOR2_X1 U9193 ( .A(n7432), .B(n7431), .ZN(n7443) );
  INV_X1 U9194 ( .A(n10544), .ZN(n9119) );
  INV_X1 U9195 ( .A(n9280), .ZN(n7600) );
  OAI22_X1 U9196 ( .A1(n7441), .A2(n9289), .B1(n10548), .B2(n7433), .ZN(n7434)
         );
  AOI21_X1 U9197 ( .B1(n7443), .B2(n7600), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9198 ( .B1(n7439), .B2(n10550), .A(n7435), .ZN(P2_U3408) );
  INV_X1 U9199 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7436) );
  MUX2_X1 U9200 ( .A(n7436), .B(n7439), .S(n10557), .Z(n7438) );
  INV_X1 U9201 ( .A(n9162), .ZN(n7693) );
  AOI22_X1 U9202 ( .A1(n7443), .A2(n7693), .B1(n9159), .B2(n7453), .ZN(n7437)
         );
  NAND2_X1 U9203 ( .A1(n7438), .A2(n7437), .ZN(P2_U3465) );
  MUX2_X1 U9204 ( .A(n7440), .B(n7439), .S(n9091), .Z(n7445) );
  INV_X1 U9205 ( .A(n9086), .ZN(n9080) );
  OAI22_X1 U9206 ( .A1(n9090), .A2(n7441), .B1(n7456), .B2(n9087), .ZN(n7442)
         );
  AOI21_X1 U9207 ( .B1(n7443), .B2(n9080), .A(n7442), .ZN(n7444) );
  NAND2_X1 U9208 ( .A1(n7445), .A2(n7444), .ZN(P2_U3227) );
  AOI211_X1 U9209 ( .C1(n7448), .C2(n7447), .A(n8318), .B(n7446), .ZN(n7449)
         );
  INV_X1 U9210 ( .A(n7449), .ZN(n7455) );
  NAND2_X1 U9211 ( .A1(n8324), .A2(n8338), .ZN(n7451) );
  OAI211_X1 U9212 ( .C1(n7656), .C2(n8326), .A(n7451), .B(n7450), .ZN(n7452)
         );
  AOI21_X1 U9213 ( .B1(n7453), .B2(n8316), .A(n7452), .ZN(n7454) );
  OAI211_X1 U9214 ( .C1(n7456), .C2(n8294), .A(n7455), .B(n7454), .ZN(P2_U3179) );
  OAI22_X1 U9215 ( .A1(n7463), .A2(n8165), .B1(n10439), .B2(n5421), .ZN(n7519)
         );
  INV_X1 U9216 ( .A(n7519), .ZN(n7466) );
  INV_X1 U9217 ( .A(n7457), .ZN(n7459) );
  NAND2_X1 U9218 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  NAND2_X1 U9219 ( .A1(n8137), .A2(n7808), .ZN(n7462) );
  OAI21_X1 U9220 ( .B1(n7463), .B2(n5421), .A(n7462), .ZN(n7464) );
  XNOR2_X1 U9221 ( .A(n7464), .B(n9345), .ZN(n9519) );
  INV_X1 U9222 ( .A(n9519), .ZN(n7521) );
  XNOR2_X1 U9223 ( .A(n9518), .B(n7521), .ZN(n7465) );
  NAND2_X1 U9224 ( .A1(n7465), .A2(n7466), .ZN(n9517) );
  OAI21_X1 U9225 ( .B1(n7466), .B2(n7465), .A(n9517), .ZN(n7467) );
  NAND2_X1 U9226 ( .A1(n7467), .A2(n9533), .ZN(n7473) );
  NAND2_X1 U9227 ( .A1(n9837), .A2(n4420), .ZN(n7469) );
  NAND2_X1 U9228 ( .A1(n9835), .A2(n9522), .ZN(n7468) );
  NAND2_X1 U9229 ( .A1(n7469), .A2(n7468), .ZN(n7800) );
  NAND2_X1 U9230 ( .A1(n10311), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9879) );
  OAI21_X1 U9231 ( .B1(n9554), .B2(n7805), .A(n9879), .ZN(n7471) );
  NOR2_X1 U9232 ( .A1(n9545), .A2(n10439), .ZN(n7470) );
  AOI211_X1 U9233 ( .C1(n9542), .C2(n7800), .A(n7471), .B(n7470), .ZN(n7472)
         );
  NAND2_X1 U9234 ( .A1(n7473), .A2(n7472), .ZN(P1_U3227) );
  INV_X1 U9235 ( .A(n7474), .ZN(n7477) );
  INV_X1 U9236 ( .A(n9943), .ZN(n9966) );
  OAI222_X1 U9237 ( .A1(n10332), .A2(n7475), .B1(n10335), .B2(n7477), .C1(
        n10311), .C2(n9966), .ZN(P1_U3338) );
  OAI222_X1 U9238 ( .A1(n4879), .A2(P2_U3151), .B1(n9307), .B2(n7477), .C1(
        n7476), .C2(n8134), .ZN(P2_U3278) );
  NAND2_X1 U9239 ( .A1(n9839), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7478) );
  OAI21_X1 U9240 ( .B1(n7885), .B2(n9839), .A(n7478), .ZN(P1_U3583) );
  NAND2_X1 U9241 ( .A1(n9839), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7479) );
  OAI21_X1 U9242 ( .B1(n9538), .B2(n9839), .A(n7479), .ZN(P1_U3581) );
  OAI21_X1 U9243 ( .B1(n7482), .B2(n7481), .A(n7480), .ZN(n7483) );
  NAND2_X1 U9244 ( .A1(n7483), .A2(n8320), .ZN(n7487) );
  AND2_X1 U9245 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7622) );
  AOI21_X1 U9246 ( .B1(n8324), .B2(n8337), .A(n7622), .ZN(n7484) );
  OAI21_X1 U9247 ( .B1(n7595), .B2(n8326), .A(n7484), .ZN(n7485) );
  AOI21_X1 U9248 ( .B1(n7692), .B2(n8316), .A(n7485), .ZN(n7486) );
  OAI211_X1 U9249 ( .C1(n9088), .C2(n8294), .A(n7487), .B(n7486), .ZN(P2_U3153) );
  OAI21_X1 U9250 ( .B1(n7429), .B2(n7492), .A(n7488), .ZN(n10545) );
  INV_X1 U9251 ( .A(n10545), .ZN(n7498) );
  NAND2_X1 U9252 ( .A1(n7490), .A2(n7489), .ZN(n7491) );
  XOR2_X1 U9253 ( .A(n7492), .B(n7491), .Z(n7493) );
  AOI222_X1 U9254 ( .A1(n9061), .A2(n7493), .B1(n7367), .B2(n9064), .C1(n8337), 
        .C2(n9065), .ZN(n10547) );
  MUX2_X1 U9255 ( .A(n7494), .B(n10547), .S(n9091), .Z(n7497) );
  INV_X1 U9256 ( .A(n7495), .ZN(n7513) );
  AOI22_X1 U9257 ( .A1(n9029), .A2(n10542), .B1(n10518), .B2(n7513), .ZN(n7496) );
  OAI211_X1 U9258 ( .C1(n7498), .C2(n9086), .A(n7497), .B(n7496), .ZN(P2_U3228) );
  INV_X1 U9259 ( .A(n7499), .ZN(n7604) );
  AOI22_X1 U9260 ( .A1(n9979), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10315), .ZN(n7500) );
  OAI21_X1 U9261 ( .B1(n7604), .B2(n10335), .A(n7500), .ZN(P1_U3337) );
  NAND2_X1 U9262 ( .A1(n8316), .A2(n10542), .ZN(n7504) );
  INV_X1 U9263 ( .A(n7501), .ZN(n7502) );
  AOI21_X1 U9264 ( .B1(n8324), .B2(n7367), .A(n7502), .ZN(n7503) );
  OAI211_X1 U9265 ( .C1(n7596), .C2(n8326), .A(n7504), .B(n7503), .ZN(n7512)
         );
  INV_X1 U9266 ( .A(n7505), .ZN(n7507) );
  NAND3_X1 U9267 ( .A1(n7508), .A2(n7507), .A3(n7506), .ZN(n7510) );
  AOI21_X1 U9268 ( .B1(n7510), .B2(n7509), .A(n8318), .ZN(n7511) );
  AOI211_X1 U9269 ( .C1(n7513), .C2(n8329), .A(n7512), .B(n7511), .ZN(n7514)
         );
  INV_X1 U9270 ( .A(n7514), .ZN(P2_U3167) );
  AND2_X1 U9271 ( .A1(n9519), .A2(n7519), .ZN(n7517) );
  NAND2_X1 U9272 ( .A1(n8137), .A2(n9527), .ZN(n7515) );
  OAI21_X1 U9273 ( .B1(n7538), .B2(n5421), .A(n7515), .ZN(n7516) );
  XNOR2_X1 U9274 ( .A(n7516), .B(n9345), .ZN(n7518) );
  OAI22_X1 U9275 ( .A1(n7538), .A2(n8165), .B1(n10445), .B2(n5421), .ZN(n9513)
         );
  AND2_X1 U9276 ( .A1(n7518), .A2(n9513), .ZN(n9514) );
  OR2_X1 U9277 ( .A1(n7517), .A2(n9514), .ZN(n7524) );
  OAI21_X1 U9278 ( .B1(n9519), .B2(n7519), .A(n9513), .ZN(n7522) );
  INV_X1 U9279 ( .A(n7518), .ZN(n9516) );
  NOR2_X1 U9280 ( .A1(n7519), .A2(n9513), .ZN(n7520) );
  AOI22_X1 U9281 ( .A1(n7522), .A2(n9516), .B1(n7521), .B2(n7520), .ZN(n7523)
         );
  NAND2_X1 U9282 ( .A1(n8137), .A2(n7528), .ZN(n7525) );
  OAI21_X1 U9283 ( .B1(n7526), .B2(n5421), .A(n7525), .ZN(n7527) );
  XNOR2_X1 U9284 ( .A(n7527), .B(n8141), .ZN(n7530) );
  AND2_X1 U9285 ( .A1(n7528), .A2(n4427), .ZN(n7529) );
  AOI21_X1 U9286 ( .B1(n9834), .B2(n9342), .A(n7529), .ZN(n7531) );
  NAND2_X1 U9287 ( .A1(n7530), .A2(n7531), .ZN(n8020) );
  INV_X1 U9288 ( .A(n7530), .ZN(n7533) );
  INV_X1 U9289 ( .A(n7531), .ZN(n7532) );
  NAND2_X1 U9290 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  AND2_X1 U9291 ( .A1(n8020), .A2(n7534), .ZN(n7535) );
  NOR2_X1 U9292 ( .A1(n7536), .A2(n7535), .ZN(n7537) );
  OAI21_X1 U9293 ( .B1(n9364), .B2(n7537), .A(n9533), .ZN(n7541) );
  OAI22_X1 U9294 ( .A1(n7538), .A2(n9535), .B1(n9537), .B2(n8015), .ZN(n7646)
         );
  NAND2_X1 U9295 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9913) );
  OAI21_X1 U9296 ( .B1(n9554), .B2(n7649), .A(n9913), .ZN(n7539) );
  AOI21_X1 U9297 ( .B1(n9542), .B2(n7646), .A(n7539), .ZN(n7540) );
  OAI211_X1 U9298 ( .C1(n10455), .C2(n9545), .A(n7541), .B(n7540), .ZN(
        P1_U3213) );
  XNOR2_X1 U9299 ( .A(n7542), .B(n9063), .ZN(n7543) );
  XNOR2_X1 U9300 ( .A(n7544), .B(n7543), .ZN(n7550) );
  NAND2_X1 U9301 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7554) );
  INV_X1 U9302 ( .A(n7554), .ZN(n7546) );
  NOR2_X1 U9303 ( .A1(n8326), .A2(n7655), .ZN(n7545) );
  AOI211_X1 U9304 ( .C1(n8324), .C2(n8336), .A(n7546), .B(n7545), .ZN(n7547)
         );
  OAI21_X1 U9305 ( .B1(n9077), .B2(n8294), .A(n7547), .ZN(n7548) );
  AOI21_X1 U9306 ( .B1(n9076), .B2(n8316), .A(n7548), .ZN(n7549) );
  OAI21_X1 U9307 ( .B1(n7550), .B2(n8318), .A(n7549), .ZN(P2_U3161) );
  XNOR2_X1 U9308 ( .A(n7574), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7747) );
  XOR2_X1 U9309 ( .A(n7748), .B(n7747), .Z(n7578) );
  INV_X1 U9310 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7555) );
  OAI21_X1 U9311 ( .B1(n8778), .B2(n7555), .A(n7554), .ZN(n7566) );
  INV_X1 U9312 ( .A(n7560), .ZN(n7561) );
  XNOR2_X1 U9313 ( .A(n7574), .B(n9075), .ZN(n7562) );
  INV_X1 U9314 ( .A(n7754), .ZN(n7564) );
  NAND3_X1 U9315 ( .A1(n7620), .A2(n7562), .A3(n7561), .ZN(n7563) );
  AOI21_X1 U9316 ( .B1(n7564), .B2(n7563), .A(n10503), .ZN(n7565) );
  AOI211_X1 U9317 ( .C1(n10505), .C2(n7574), .A(n7566), .B(n7565), .ZN(n7577)
         );
  MUX2_X1 U9318 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8770), .Z(n7571) );
  INV_X1 U9319 ( .A(n7571), .ZN(n7572) );
  INV_X1 U9320 ( .A(n7567), .ZN(n7569) );
  XOR2_X1 U9321 ( .A(n7573), .B(n7571), .Z(n7625) );
  MUX2_X1 U9322 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8770), .Z(n7749) );
  XOR2_X1 U9323 ( .A(n7574), .B(n7749), .Z(n7750) );
  XNOR2_X1 U9324 ( .A(n7751), .B(n7750), .ZN(n7575) );
  NAND2_X1 U9325 ( .A1(n7575), .A2(n8797), .ZN(n7576) );
  OAI211_X1 U9326 ( .C1(n7578), .C2(n8781), .A(n7577), .B(n7576), .ZN(P2_U3190) );
  AOI22_X1 U9327 ( .A1(n7580), .A2(n7579), .B1(n7582), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n9923) );
  XOR2_X1 U9328 ( .A(n7583), .B(n9923), .Z(n9924) );
  INV_X1 U9329 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10226) );
  XNOR2_X1 U9330 ( .A(n9924), .B(n10226), .ZN(n7589) );
  XNOR2_X1 U9331 ( .A(n9929), .B(n7583), .ZN(n7584) );
  NAND2_X1 U9332 ( .A1(n7584), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n9927) );
  OAI211_X1 U9333 ( .C1(n7584), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9927), .B(
        n9984), .ZN(n7588) );
  NOR2_X1 U9334 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9553), .ZN(n7586) );
  NOR2_X1 U9335 ( .A1(n9975), .A2(n9928), .ZN(n7585) );
  AOI211_X1 U9336 ( .C1(n9965), .C2(P1_ADDR_REG_15__SCAN_IN), .A(n7586), .B(
        n7585), .ZN(n7587) );
  OAI211_X1 U9337 ( .C1(n7589), .C2(n9939), .A(n7588), .B(n7587), .ZN(P1_U3258) );
  INV_X1 U9338 ( .A(n9061), .ZN(n9007) );
  INV_X1 U9339 ( .A(n7591), .ZN(n7592) );
  AOI21_X1 U9340 ( .B1(n7593), .B2(n7590), .A(n7592), .ZN(n7594) );
  OAI222_X1 U9341 ( .A1(n9010), .A2(n7596), .B1(n9008), .B2(n7595), .C1(n9007), 
        .C2(n7594), .ZN(n9092) );
  INV_X1 U9342 ( .A(n9092), .ZN(n7690) );
  AOI22_X1 U9343 ( .A1(n9277), .A2(n7692), .B1(P2_REG0_REG_7__SCAN_IN), .B2(
        n10550), .ZN(n7602) );
  INV_X1 U9344 ( .A(n7597), .ZN(n7598) );
  AOI21_X1 U9345 ( .B1(n7599), .B2(n5286), .A(n7598), .ZN(n9095) );
  NAND2_X1 U9346 ( .A1(n9095), .A2(n7600), .ZN(n7601) );
  OAI211_X1 U9347 ( .C1(n7690), .C2(n10550), .A(n7602), .B(n7601), .ZN(
        P2_U3411) );
  INV_X1 U9348 ( .A(n8786), .ZN(n8799) );
  OAI222_X1 U9349 ( .A1(P2_U3151), .A2(n8799), .B1(n9307), .B2(n7604), .C1(
        n7603), .C2(n8134), .ZN(P2_U3277) );
  NOR2_X1 U9350 ( .A1(n7606), .A2(n7605), .ZN(n7607) );
  NAND2_X1 U9351 ( .A1(n7608), .A2(n7607), .ZN(n7609) );
  NAND2_X1 U9352 ( .A1(n10392), .A2(n10390), .ZN(n7776) );
  AND2_X2 U9353 ( .A1(n7609), .A2(n10117), .ZN(n7610) );
  AOI21_X1 U9354 ( .B1(n7776), .B2(n10383), .A(n10253), .ZN(n7618) );
  XNOR2_X1 U9355 ( .A(n9840), .B(n10253), .ZN(n10250) );
  NAND3_X1 U9356 ( .A1(n10250), .A2(n10254), .A3(n7612), .ZN(n7613) );
  AOI21_X1 U9357 ( .B1(n10251), .B2(n7613), .A(n7610), .ZN(n7617) );
  OAI22_X1 U9358 ( .A1(n10162), .A2(n7615), .B1(n7614), .B2(n10117), .ZN(n7616) );
  OR3_X1 U9359 ( .A1(n7618), .A2(n7617), .A3(n7616), .ZN(P1_U3293) );
  XNOR2_X1 U9360 ( .A(n7619), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7632) );
  OAI21_X1 U9361 ( .B1(P2_REG2_REG_7__SCAN_IN), .B2(n7621), .A(n7620), .ZN(
        n7630) );
  AOI21_X1 U9362 ( .B1(n10513), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7622), .ZN(
        n7623) );
  OAI21_X1 U9363 ( .B1(n4757), .B2(n8795), .A(n7623), .ZN(n7629) );
  AOI21_X1 U9364 ( .B1(n7626), .B2(n7625), .A(n7624), .ZN(n7627) );
  NOR2_X1 U9365 ( .A1(n7627), .A2(n10510), .ZN(n7628) );
  AOI211_X1 U9366 ( .C1(n8763), .C2(n7630), .A(n7629), .B(n7628), .ZN(n7631)
         );
  OAI21_X1 U9367 ( .B1(n7632), .B2(n8781), .A(n7631), .ZN(P2_U3189) );
  AOI21_X1 U9368 ( .B1(n7634), .B2(n10377), .A(n7633), .ZN(n10427) );
  AND2_X1 U9369 ( .A1(n10410), .A2(n7635), .ZN(n7636) );
  XNOR2_X1 U9370 ( .A(n7637), .B(n10386), .ZN(n10430) );
  OAI211_X1 U9371 ( .C1(n7699), .C2(n10426), .A(n10390), .B(n7638), .ZN(n10425) );
  OAI22_X1 U9372 ( .A1(n10082), .A2(n10425), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10117), .ZN(n7639) );
  AOI21_X1 U9373 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n7610), .A(n7639), .ZN(
        n7640) );
  OAI21_X1 U9374 ( .B1(n10426), .B2(n10383), .A(n7640), .ZN(n7641) );
  AOI21_X1 U9375 ( .B1(n10393), .B2(n10430), .A(n7641), .ZN(n7642) );
  OAI21_X1 U9376 ( .B1(n7610), .B2(n10427), .A(n7642), .ZN(P1_U3290) );
  INV_X1 U9377 ( .A(n9574), .ZN(n9572) );
  INV_X1 U9378 ( .A(n9577), .ZN(n7644) );
  AOI21_X1 U9379 ( .B1(n7645), .B2(n9572), .A(n7644), .ZN(n7667) );
  XNOR2_X1 U9380 ( .A(n7667), .B(n9578), .ZN(n7647) );
  AOI21_X1 U9381 ( .B1(n7647), .B2(n10377), .A(n7646), .ZN(n10456) );
  MUX2_X1 U9382 ( .A(n8539), .B(n10456), .S(n10162), .Z(n7653) );
  XNOR2_X1 U9383 ( .A(n7648), .B(n9578), .ZN(n10459) );
  OAI22_X1 U9384 ( .A1(n10383), .A2(n10455), .B1(n10117), .B2(n7649), .ZN(
        n7651) );
  OAI211_X1 U9385 ( .C1(n10368), .C2(n10455), .A(n10390), .B(n7673), .ZN(
        n10453) );
  NOR2_X1 U9386 ( .A1(n10453), .A2(n10082), .ZN(n7650) );
  AOI211_X1 U9387 ( .C1(n10393), .C2(n10459), .A(n7651), .B(n7650), .ZN(n7652)
         );
  NAND2_X1 U9388 ( .A1(n7653), .A2(n7652), .ZN(P1_U3286) );
  XNOR2_X1 U9389 ( .A(n7654), .B(n7660), .ZN(n7658) );
  OAI22_X1 U9390 ( .A1(n9010), .A2(n7656), .B1(n7655), .B2(n9008), .ZN(n7657)
         );
  AOI21_X1 U9391 ( .B1(n7658), .B2(n9061), .A(n7657), .ZN(n9074) );
  INV_X1 U9392 ( .A(n7660), .ZN(n7661) );
  OR2_X1 U9393 ( .A1(n7659), .A2(n7661), .ZN(n9082) );
  NAND2_X1 U9394 ( .A1(n7659), .A2(n7661), .ZN(n9081) );
  NAND3_X1 U9395 ( .A1(n9082), .A2(n9081), .A3(n10544), .ZN(n7663) );
  NAND2_X1 U9396 ( .A1(n9076), .A2(n10543), .ZN(n7662) );
  AND2_X1 U9397 ( .A1(n7663), .A2(n7662), .ZN(n7664) );
  AND2_X1 U9398 ( .A1(n9074), .A2(n7664), .ZN(n9173) );
  NAND2_X1 U9399 ( .A1(n10550), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7665) );
  OAI21_X1 U9400 ( .B1(n9173), .B2(n10550), .A(n7665), .ZN(P2_U3414) );
  OAI21_X1 U9401 ( .B1(n7667), .B2(n9578), .A(n7666), .ZN(n7783) );
  XNOR2_X1 U9402 ( .A(n7783), .B(n7782), .ZN(n7671) );
  NAND2_X1 U9403 ( .A1(n9834), .A2(n4420), .ZN(n7670) );
  INV_X1 U9404 ( .A(n7668), .ZN(n9832) );
  NAND2_X1 U9405 ( .A1(n9832), .A2(n9551), .ZN(n7669) );
  NAND2_X1 U9406 ( .A1(n7670), .A2(n7669), .ZN(n9373) );
  AOI21_X1 U9407 ( .B1(n7671), .B2(n10377), .A(n9373), .ZN(n10247) );
  INV_X1 U9408 ( .A(n7788), .ZN(n7672) );
  AOI211_X1 U9409 ( .C1(n10245), .C2(n7673), .A(n10475), .B(n7672), .ZN(n10244) );
  INV_X1 U9410 ( .A(n9369), .ZN(n7674) );
  AOI22_X1 U9411 ( .A1(n7610), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7674), .B2(
        n10380), .ZN(n7675) );
  OAI21_X1 U9412 ( .B1(n10383), .B2(n9370), .A(n7675), .ZN(n7678) );
  XOR2_X1 U9413 ( .A(n7782), .B(n7676), .Z(n10248) );
  NOR2_X1 U9414 ( .A1(n10248), .A2(n10164), .ZN(n7677) );
  AOI211_X1 U9415 ( .C1(n10244), .C2(n10392), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI21_X1 U9416 ( .B1(n10247), .B2(n7610), .A(n7679), .ZN(P1_U3285) );
  NAND2_X1 U9417 ( .A1(n8774), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7680) );
  OAI21_X1 U9418 ( .B1(n8808), .B2(n8774), .A(n7680), .ZN(P2_U3522) );
  INV_X1 U9419 ( .A(n7681), .ZN(n9290) );
  OAI211_X1 U9420 ( .C1(n7684), .C2(n7683), .A(n7682), .B(n8320), .ZN(n7689)
         );
  NAND2_X1 U9421 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7753) );
  OAI21_X1 U9422 ( .B1(n8326), .B2(n7685), .A(n7753), .ZN(n7687) );
  NOR2_X1 U9423 ( .A1(n8294), .A2(n9057), .ZN(n7686) );
  AOI211_X1 U9424 ( .C1(n8324), .C2(n9063), .A(n7687), .B(n7686), .ZN(n7688)
         );
  OAI211_X1 U9425 ( .C1(n9290), .C2(n8332), .A(n7689), .B(n7688), .ZN(P2_U3171) );
  MUX2_X1 U9426 ( .A(n7691), .B(n7690), .S(n10557), .Z(n7695) );
  AOI22_X1 U9427 ( .A1(n9095), .A2(n7693), .B1(n9159), .B2(n7692), .ZN(n7694)
         );
  NAND2_X1 U9428 ( .A1(n7695), .A2(n7694), .ZN(P2_U3466) );
  XNOR2_X1 U9429 ( .A(n9675), .B(n7696), .ZN(n10423) );
  INV_X1 U9430 ( .A(n10423), .ZN(n7710) );
  NAND2_X1 U9431 ( .A1(n7715), .A2(n5481), .ZN(n7697) );
  NAND2_X1 U9432 ( .A1(n7697), .A2(n10390), .ZN(n7698) );
  OR2_X1 U9433 ( .A1(n7699), .A2(n7698), .ZN(n10419) );
  NAND2_X1 U9434 ( .A1(n7610), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7701) );
  NAND2_X1 U9435 ( .A1(n10380), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7700) );
  OAI211_X1 U9436 ( .C1(n10419), .C2(n10082), .A(n7701), .B(n7700), .ZN(n7708)
         );
  OAI21_X1 U9437 ( .B1(n7704), .B2(n7703), .A(n7702), .ZN(n7706) );
  AOI21_X1 U9438 ( .B1(n7706), .B2(n10377), .A(n7705), .ZN(n10420) );
  NOR2_X1 U9439 ( .A1(n10420), .A2(n7610), .ZN(n7707) );
  AOI211_X1 U9440 ( .C1(n10079), .C2(n5481), .A(n7708), .B(n7707), .ZN(n7709)
         );
  OAI21_X1 U9441 ( .B1(n10164), .B2(n7710), .A(n7709), .ZN(P1_U3291) );
  CLKBUF_X1 U9442 ( .A(n7711), .Z(n7712) );
  INV_X1 U9443 ( .A(n7713), .ZN(n7714) );
  XNOR2_X1 U9444 ( .A(n7712), .B(n7714), .ZN(n10411) );
  OAI211_X1 U9445 ( .C1(n10253), .C2(n10414), .A(n10390), .B(n7715), .ZN(
        n10412) );
  INV_X1 U9446 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7716) );
  OAI22_X1 U9447 ( .A1(n10082), .A2(n10412), .B1(n7716), .B2(n10117), .ZN(
        n7717) );
  AOI21_X1 U9448 ( .B1(n10079), .B2(n5458), .A(n7717), .ZN(n7725) );
  INV_X1 U9449 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U9450 ( .A1(n7719), .A2(n7712), .ZN(n7721) );
  NAND2_X1 U9451 ( .A1(n7721), .A2(n7720), .ZN(n7723) );
  AOI21_X1 U9452 ( .B1(n7723), .B2(n10377), .A(n7722), .ZN(n10413) );
  MUX2_X1 U9453 ( .A(n10413), .B(n6971), .S(n7610), .Z(n7724) );
  OAI211_X1 U9454 ( .C1(n10411), .C2(n10164), .A(n7725), .B(n7724), .ZN(
        P1_U3292) );
  INV_X1 U9455 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10564) );
  NOR2_X1 U9456 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7726) );
  AOI21_X1 U9457 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7726), .ZN(n10569) );
  NOR2_X1 U9458 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7727) );
  AOI21_X1 U9459 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7727), .ZN(n10572) );
  NOR2_X1 U9460 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7728) );
  AOI21_X1 U9461 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7728), .ZN(n10575) );
  NOR2_X1 U9462 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7729) );
  AOI21_X1 U9463 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7729), .ZN(n10578) );
  NOR2_X1 U9464 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7730) );
  AOI21_X1 U9465 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n7730), .ZN(n10581) );
  NOR2_X1 U9466 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7731) );
  AOI21_X1 U9467 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7731), .ZN(n10589) );
  NOR2_X1 U9468 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7732) );
  AOI21_X1 U9469 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7732), .ZN(n10592) );
  NOR2_X1 U9470 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7733) );
  AOI21_X1 U9471 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7733), .ZN(n10601) );
  NOR2_X1 U9472 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7734) );
  AOI21_X1 U9473 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7734), .ZN(n10607) );
  NOR2_X1 U9474 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7735) );
  AOI21_X1 U9475 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7735), .ZN(n10604) );
  NOR2_X1 U9476 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7736) );
  AOI21_X1 U9477 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7736), .ZN(n10595) );
  NOR2_X1 U9478 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7737) );
  AOI21_X1 U9479 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7737), .ZN(n10598) );
  AND2_X1 U9480 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7738) );
  NOR2_X1 U9481 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7738), .ZN(n10559) );
  INV_X1 U9482 ( .A(n10559), .ZN(n10560) );
  NAND3_X1 U9483 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10561) );
  NAND2_X1 U9484 ( .A1(n10562), .A2(n10561), .ZN(n10558) );
  NAND2_X1 U9485 ( .A1(n10560), .A2(n10558), .ZN(n10610) );
  NAND2_X1 U9486 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7739) );
  OAI21_X1 U9487 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7739), .ZN(n10609) );
  NOR2_X1 U9488 ( .A1(n10610), .A2(n10609), .ZN(n10608) );
  AOI21_X1 U9489 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10608), .ZN(n10613) );
  NAND2_X1 U9490 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7740) );
  OAI21_X1 U9491 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7740), .ZN(n10612) );
  NOR2_X1 U9492 ( .A1(n10613), .A2(n10612), .ZN(n10611) );
  AOI21_X1 U9493 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10611), .ZN(n10616) );
  NOR2_X1 U9494 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7741) );
  AOI21_X1 U9495 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7741), .ZN(n10615) );
  NAND2_X1 U9496 ( .A1(n10616), .A2(n10615), .ZN(n10614) );
  OAI21_X1 U9497 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10614), .ZN(n10597) );
  NAND2_X1 U9498 ( .A1(n10598), .A2(n10597), .ZN(n10596) );
  OAI21_X1 U9499 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10596), .ZN(n10594) );
  NAND2_X1 U9500 ( .A1(n10595), .A2(n10594), .ZN(n10593) );
  OAI21_X1 U9501 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10593), .ZN(n10603) );
  NAND2_X1 U9502 ( .A1(n10604), .A2(n10603), .ZN(n10602) );
  OAI21_X1 U9503 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10602), .ZN(n10606) );
  NAND2_X1 U9504 ( .A1(n10607), .A2(n10606), .ZN(n10605) );
  OAI21_X1 U9505 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10605), .ZN(n10600) );
  NAND2_X1 U9506 ( .A1(n10601), .A2(n10600), .ZN(n10599) );
  OAI21_X1 U9507 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10599), .ZN(n10591) );
  NAND2_X1 U9508 ( .A1(n10592), .A2(n10591), .ZN(n10590) );
  OAI21_X1 U9509 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10590), .ZN(n10588) );
  NAND2_X1 U9510 ( .A1(n10589), .A2(n10588), .ZN(n10587) );
  OAI21_X1 U9511 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10587), .ZN(n10585) );
  NAND2_X1 U9512 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8704) );
  OAI211_X1 U9513 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10585), .B(n8704), .ZN(n10584) );
  OAI21_X1 U9514 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10584), .ZN(n10580) );
  NAND2_X1 U9515 ( .A1(n10581), .A2(n10580), .ZN(n10579) );
  OAI21_X1 U9516 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10579), .ZN(n10577) );
  NAND2_X1 U9517 ( .A1(n10578), .A2(n10577), .ZN(n10576) );
  OAI21_X1 U9518 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10576), .ZN(n10574) );
  NAND2_X1 U9519 ( .A1(n10575), .A2(n10574), .ZN(n10573) );
  OAI21_X1 U9520 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10573), .ZN(n10571) );
  NAND2_X1 U9521 ( .A1(n10572), .A2(n10571), .ZN(n10570) );
  OAI21_X1 U9522 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10570), .ZN(n10568) );
  NAND2_X1 U9523 ( .A1(n10569), .A2(n10568), .ZN(n10567) );
  OAI21_X1 U9524 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10567), .ZN(n10565) );
  NOR2_X1 U9525 ( .A1(n10564), .A2(n10565), .ZN(n7742) );
  NAND2_X1 U9526 ( .A1(n10564), .A2(n10565), .ZN(n10563) );
  OAI21_X1 U9527 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7742), .A(n10563), .ZN(
        n7746) );
  NOR2_X1 U9528 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  XNOR2_X1 U9529 ( .A(n7746), .B(n7745), .ZN(ADD_1068_U4) );
  XNOR2_X1 U9530 ( .A(n8341), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n7764) );
  OAI22_X1 U9531 ( .A1(n7751), .A2(n7750), .B1(n7749), .B2(n7755), .ZN(n8346)
         );
  MUX2_X1 U9532 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8770), .Z(n8342) );
  XNOR2_X1 U9533 ( .A(n8342), .B(n8344), .ZN(n8345) );
  XNOR2_X1 U9534 ( .A(n8346), .B(n8345), .ZN(n7762) );
  NAND2_X1 U9535 ( .A1(n10513), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7752) );
  OAI211_X1 U9536 ( .C1(n8795), .C2(n5079), .A(n7753), .B(n7752), .ZN(n7761)
         );
  INV_X1 U9537 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7758) );
  AOI21_X1 U9538 ( .B1(n7758), .B2(n7757), .A(n8350), .ZN(n7759) );
  NOR2_X1 U9539 ( .A1(n7759), .A2(n10503), .ZN(n7760) );
  AOI211_X1 U9540 ( .C1(n8797), .C2(n7762), .A(n7761), .B(n7760), .ZN(n7763)
         );
  OAI21_X1 U9541 ( .B1(n7764), .B2(n8781), .A(n7763), .ZN(P2_U3191) );
  INV_X1 U9542 ( .A(n7765), .ZN(n7766) );
  OAI222_X1 U9543 ( .A1(n8794), .A2(P2_U3151), .B1(n9307), .B2(n7766), .C1(
        n8563), .C2(n8134), .ZN(P2_U3276) );
  OAI222_X1 U9544 ( .A1(n10332), .A2(n8717), .B1(n10335), .B2(n7766), .C1(
        n9800), .C2(n10311), .ZN(P1_U3336) );
  XNOR2_X1 U9545 ( .A(n7767), .B(n9681), .ZN(n10479) );
  INV_X1 U9546 ( .A(n10479), .ZN(n7779) );
  XNOR2_X1 U9547 ( .A(n7768), .B(n9681), .ZN(n7772) );
  NAND2_X1 U9548 ( .A1(n9829), .A2(n9522), .ZN(n7770) );
  NAND2_X1 U9549 ( .A1(n9831), .A2(n4420), .ZN(n7769) );
  NAND2_X1 U9550 ( .A1(n7770), .A2(n7769), .ZN(n9494) );
  INV_X1 U9551 ( .A(n9494), .ZN(n7771) );
  OAI21_X1 U9552 ( .B1(n7772), .B2(n10152), .A(n7771), .ZN(n10477) );
  OAI21_X1 U9553 ( .B1(n10349), .B2(n10474), .A(n7822), .ZN(n10476) );
  INV_X1 U9554 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7773) );
  OAI22_X1 U9555 ( .A1(n10162), .A2(n7773), .B1(n9492), .B2(n10117), .ZN(n7774) );
  AOI21_X1 U9556 ( .B1(n10079), .B2(n9603), .A(n7774), .ZN(n7775) );
  OAI21_X1 U9557 ( .B1(n10476), .B2(n7776), .A(n7775), .ZN(n7777) );
  AOI21_X1 U9558 ( .B1(n10477), .B2(n10162), .A(n7777), .ZN(n7778) );
  OAI21_X1 U9559 ( .B1(n7779), .B2(n10164), .A(n7778), .ZN(P1_U3282) );
  INV_X1 U9560 ( .A(n7780), .ZN(n7781) );
  AOI21_X1 U9561 ( .B1(n7783), .B2(n7782), .A(n7781), .ZN(n7784) );
  XOR2_X1 U9562 ( .A(n7787), .B(n7784), .Z(n7785) );
  NAND2_X1 U9563 ( .A1(n4420), .A2(n9833), .ZN(n9444) );
  OAI21_X1 U9564 ( .B1(n7785), .B2(n10152), .A(n9444), .ZN(n10463) );
  INV_X1 U9565 ( .A(n10463), .ZN(n7797) );
  XNOR2_X1 U9566 ( .A(n7786), .B(n7787), .ZN(n10465) );
  NAND2_X1 U9567 ( .A1(n7788), .A2(n8026), .ZN(n7789) );
  NAND2_X1 U9568 ( .A1(n7789), .A2(n10390), .ZN(n7790) );
  OR2_X1 U9569 ( .A1(n7790), .A2(n10351), .ZN(n7791) );
  NAND2_X1 U9570 ( .A1(n9831), .A2(n9551), .ZN(n9445) );
  AND2_X1 U9571 ( .A1(n7791), .A2(n9445), .ZN(n10461) );
  OAI22_X1 U9572 ( .A1(n10162), .A2(n7792), .B1(n9446), .B2(n10117), .ZN(n7793) );
  AOI21_X1 U9573 ( .B1(n10079), .B2(n8026), .A(n7793), .ZN(n7794) );
  OAI21_X1 U9574 ( .B1(n10461), .B2(n10082), .A(n7794), .ZN(n7795) );
  AOI21_X1 U9575 ( .B1(n10465), .B2(n10393), .A(n7795), .ZN(n7796) );
  OAI21_X1 U9576 ( .B1(n7797), .B2(n7610), .A(n7796), .ZN(P1_U3284) );
  XOR2_X1 U9577 ( .A(n7799), .B(n7798), .Z(n7802) );
  INV_X1 U9578 ( .A(n7800), .ZN(n7801) );
  OAI21_X1 U9579 ( .B1(n7802), .B2(n10152), .A(n7801), .ZN(n10440) );
  INV_X1 U9580 ( .A(n10440), .ZN(n7812) );
  XNOR2_X1 U9581 ( .A(n7803), .B(n7798), .ZN(n10442) );
  AOI21_X1 U9582 ( .B1(n10389), .B2(n7808), .A(n10475), .ZN(n7804) );
  NAND2_X1 U9583 ( .A1(n7804), .A2(n10367), .ZN(n10438) );
  INV_X1 U9584 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7806) );
  OAI22_X1 U9585 ( .A1(n10162), .A2(n7806), .B1(n7805), .B2(n10117), .ZN(n7807) );
  AOI21_X1 U9586 ( .B1(n10079), .B2(n7808), .A(n7807), .ZN(n7809) );
  OAI21_X1 U9587 ( .B1(n10082), .B2(n10438), .A(n7809), .ZN(n7810) );
  AOI21_X1 U9588 ( .B1(n10393), .B2(n10442), .A(n7810), .ZN(n7811) );
  OAI21_X1 U9589 ( .B1(n7812), .B2(n7610), .A(n7811), .ZN(P1_U3288) );
  INV_X1 U9590 ( .A(n7813), .ZN(n7830) );
  AOI21_X1 U9591 ( .B1(n10315), .B2(P2_DATAO_REG_20__SCAN_IN), .A(n7814), .ZN(
        n7815) );
  OAI21_X1 U9592 ( .B1(n7830), .B2(n10335), .A(n7815), .ZN(P1_U3335) );
  XNOR2_X1 U9593 ( .A(n7817), .B(n9682), .ZN(n10307) );
  NAND3_X1 U9594 ( .A1(n7819), .A2(n9682), .A3(n9589), .ZN(n7820) );
  NAND3_X1 U9595 ( .A1(n7818), .A2(n10377), .A3(n7820), .ZN(n7821) );
  INV_X1 U9596 ( .A(n9601), .ZN(n9830) );
  INV_X1 U9597 ( .A(n8062), .ZN(n9828) );
  AOI22_X1 U9598 ( .A1(n4420), .A2(n9830), .B1(n9828), .B2(n9522), .ZN(n9390)
         );
  NAND2_X1 U9599 ( .A1(n7821), .A2(n9390), .ZN(n10238) );
  AOI21_X1 U9600 ( .B1(n7822), .B2(n10240), .A(n10475), .ZN(n7823) );
  AND2_X1 U9601 ( .A1(n7823), .A2(n4552), .ZN(n10239) );
  NAND2_X1 U9602 ( .A1(n10239), .A2(n10392), .ZN(n7826) );
  INV_X1 U9603 ( .A(n9392), .ZN(n7824) );
  AOI22_X1 U9604 ( .A1(n7610), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7824), .B2(
        n10380), .ZN(n7825) );
  OAI211_X1 U9605 ( .C1(n5390), .C2(n10383), .A(n7826), .B(n7825), .ZN(n7827)
         );
  AOI21_X1 U9606 ( .B1(n10238), .B2(n10162), .A(n7827), .ZN(n7828) );
  OAI21_X1 U9607 ( .B1(n10307), .B2(n10164), .A(n7828), .ZN(P1_U3281) );
  OAI222_X1 U9608 ( .A1(n8134), .A2(n7831), .B1(n9307), .B2(n7830), .C1(
        P2_U3151), .C2(n7829), .ZN(P2_U3275) );
  INV_X1 U9609 ( .A(n7832), .ZN(n7835) );
  AOI22_X1 U9610 ( .A1(n4435), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9309), .ZN(n7833) );
  OAI21_X1 U9611 ( .B1(n7835), .B2(n9307), .A(n7833), .ZN(P2_U3274) );
  OAI222_X1 U9612 ( .A1(n10311), .A2(n7063), .B1(n10335), .B2(n7835), .C1(
        n7834), .C2(n10332), .ZN(P1_U3334) );
  INV_X1 U9613 ( .A(n7836), .ZN(n8177) );
  OAI222_X1 U9614 ( .A1(P2_U3151), .A2(n7838), .B1(n9307), .B2(n8177), .C1(
        n7837), .C2(n8134), .ZN(P2_U3273) );
  INV_X1 U9615 ( .A(n7839), .ZN(n9684) );
  XNOR2_X1 U9616 ( .A(n7840), .B(n9684), .ZN(n10302) );
  NAND2_X1 U9617 ( .A1(n7818), .A2(n9590), .ZN(n7841) );
  XNOR2_X1 U9618 ( .A(n7841), .B(n9684), .ZN(n7842) );
  AOI22_X1 U9619 ( .A1(n4420), .A2(n9829), .B1(n9827), .B2(n9522), .ZN(n9466)
         );
  OAI21_X1 U9620 ( .B1(n7842), .B2(n10152), .A(n9466), .ZN(n10233) );
  AOI21_X1 U9621 ( .B1(n4552), .B2(n10235), .A(n10475), .ZN(n7843) );
  AND2_X1 U9622 ( .A1(n4565), .A2(n7843), .ZN(n10234) );
  NAND2_X1 U9623 ( .A1(n10234), .A2(n10392), .ZN(n7846) );
  INV_X1 U9624 ( .A(n9468), .ZN(n7844) );
  AOI22_X1 U9625 ( .A1(n7610), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7844), .B2(
        n10380), .ZN(n7845) );
  OAI211_X1 U9626 ( .C1(n9473), .C2(n10383), .A(n7846), .B(n7845), .ZN(n7847)
         );
  AOI21_X1 U9627 ( .B1(n10233), .B2(n10162), .A(n7847), .ZN(n7848) );
  OAI21_X1 U9628 ( .B1(n10302), .B2(n10164), .A(n7848), .ZN(P1_U3280) );
  XOR2_X1 U9629 ( .A(n9685), .B(n7849), .Z(n10232) );
  OAI211_X1 U9630 ( .C1(n9685), .C2(n7851), .A(n7850), .B(n10377), .ZN(n7852)
         );
  AOI22_X1 U9631 ( .A1(n9828), .A2(n4420), .B1(n9522), .B2(n9826), .ZN(n9319)
         );
  NAND2_X1 U9632 ( .A1(n7852), .A2(n9319), .ZN(n10228) );
  NAND2_X1 U9633 ( .A1(n4565), .A2(n10230), .ZN(n7854) );
  NAND2_X1 U9634 ( .A1(n7854), .A2(n10390), .ZN(n7855) );
  NOR2_X1 U9635 ( .A1(n7853), .A2(n7855), .ZN(n10229) );
  NAND2_X1 U9636 ( .A1(n10229), .A2(n10392), .ZN(n7858) );
  INV_X1 U9637 ( .A(n9321), .ZN(n7856) );
  AOI22_X1 U9638 ( .A1(n7610), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7856), .B2(
        n10380), .ZN(n7857) );
  OAI211_X1 U9639 ( .C1(n8066), .C2(n10383), .A(n7858), .B(n7857), .ZN(n7859)
         );
  AOI21_X1 U9640 ( .B1(n10228), .B2(n10162), .A(n7859), .ZN(n7860) );
  OAI21_X1 U9641 ( .B1(n10232), .B2(n10164), .A(n7860), .ZN(P1_U3279) );
  INV_X1 U9642 ( .A(n7865), .ZN(n7863) );
  AOI21_X1 U9643 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9309), .A(n7861), .ZN(
        n7862) );
  OAI21_X1 U9644 ( .B1(n7863), .B2(n9307), .A(n7862), .ZN(P2_U3272) );
  NAND2_X1 U9645 ( .A1(n7865), .A2(n7864), .ZN(n7867) );
  OR2_X1 U9646 ( .A1(n7866), .A2(n10311), .ZN(n9797) );
  OAI211_X1 U9647 ( .C1(n5893), .C2(n10332), .A(n7867), .B(n9797), .ZN(
        P1_U3332) );
  INV_X1 U9648 ( .A(n7868), .ZN(n10327) );
  AOI22_X1 U9649 ( .A1(n7869), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9309), .ZN(n7870) );
  OAI21_X1 U9650 ( .B1(n10327), .B2(n9307), .A(n7870), .ZN(P2_U3269) );
  NAND2_X1 U9651 ( .A1(n9298), .A2(n5637), .ZN(n7872) );
  OR2_X1 U9652 ( .A1(n4426), .A2(n10323), .ZN(n7871) );
  NAND2_X1 U9653 ( .A1(n9295), .A2(n5637), .ZN(n7874) );
  OR2_X1 U9654 ( .A1(n7876), .A2(n10320), .ZN(n7873) );
  NOR2_X2 U9655 ( .A1(n7994), .A2(n9730), .ZN(n7997) );
  NAND2_X1 U9656 ( .A1(n9291), .A2(n5637), .ZN(n7878) );
  INV_X1 U9657 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7875) );
  OR2_X1 U9658 ( .A1(n4426), .A2(n7875), .ZN(n7877) );
  XNOR2_X1 U9659 ( .A(n7997), .B(n9666), .ZN(n7879) );
  NAND2_X1 U9660 ( .A1(n7879), .A2(n10390), .ZN(n10165) );
  NAND2_X1 U9661 ( .A1(n9807), .A2(P1_B_REG_SCAN_IN), .ZN(n7880) );
  AND2_X1 U9662 ( .A1(n9522), .A2(n7880), .ZN(n7896) );
  NAND2_X1 U9663 ( .A1(n7896), .A2(n9734), .ZN(n10167) );
  NOR2_X1 U9664 ( .A1(n7610), .A2(n10167), .ZN(n8001) );
  NOR2_X1 U9665 ( .A1(n10166), .A2(n10383), .ZN(n7881) );
  AOI211_X1 U9666 ( .C1(n7610), .C2(P1_REG2_REG_31__SCAN_IN), .A(n8001), .B(
        n7881), .ZN(n7882) );
  OAI21_X1 U9667 ( .B1(n10082), .B2(n10165), .A(n7882), .ZN(P1_U3263) );
  NAND2_X1 U9668 ( .A1(n9347), .A2(n9815), .ZN(n7883) );
  NAND2_X1 U9669 ( .A1(n7884), .A2(n7883), .ZN(n7887) );
  NAND2_X1 U9670 ( .A1(n7886), .A2(n7885), .ZN(n9726) );
  INV_X1 U9671 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n7901) );
  INV_X1 U9672 ( .A(n7890), .ZN(n9695) );
  AOI21_X1 U9673 ( .B1(n9695), .B2(n9660), .A(n10152), .ZN(n7889) );
  NOR3_X1 U9674 ( .A1(n7891), .A2(n4795), .A3(n7890), .ZN(n7898) );
  INV_X1 U9675 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7895) );
  NAND2_X1 U9676 ( .A1(n5508), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n7894) );
  NAND2_X1 U9677 ( .A1(n4436), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7893) );
  OAI211_X1 U9678 ( .C1(n5625), .C2(n7895), .A(n7894), .B(n7893), .ZN(n9814)
         );
  AOI22_X1 U9679 ( .A1(n9815), .A2(n4420), .B1(n7896), .B2(n9814), .ZN(n7897)
         );
  OAI211_X1 U9680 ( .C1(n7899), .C2(n7906), .A(n10390), .B(n7994), .ZN(n7903)
         );
  OAI21_X1 U9681 ( .B1(n7906), .B2(n10473), .A(n7903), .ZN(n7900) );
  NOR2_X1 U9682 ( .A1(n7909), .A2(n7900), .ZN(n7911) );
  MUX2_X1 U9683 ( .A(n7901), .B(n7911), .S(n10482), .Z(n7902) );
  NOR2_X1 U9684 ( .A1(n7903), .A2(n10082), .ZN(n7908) );
  AOI22_X1 U9685 ( .A1(n7904), .A2(n10380), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n7610), .ZN(n7905) );
  OAI21_X1 U9686 ( .B1(n7906), .B2(n10383), .A(n7905), .ZN(n7907) );
  AOI211_X1 U9687 ( .C1(n7909), .C2(n10162), .A(n7908), .B(n7907), .ZN(n7910)
         );
  OAI21_X1 U9688 ( .B1(n7914), .B2(n10164), .A(n7910), .ZN(P1_U3356) );
  MUX2_X1 U9689 ( .A(n7912), .B(n7911), .S(n10494), .Z(n7913) );
  INV_X1 U9690 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n7921) );
  AOI211_X1 U9691 ( .C1(n7920), .C2(n10028), .A(n10475), .B(n10014), .ZN(n7929) );
  NAND2_X1 U9692 ( .A1(n9816), .A2(n9551), .ZN(n7919) );
  NAND2_X1 U9693 ( .A1(n9818), .A2(n4420), .ZN(n7918) );
  NAND2_X1 U9694 ( .A1(n7919), .A2(n7918), .ZN(n9403) );
  OAI21_X1 U9695 ( .B1(n7933), .B2(n10306), .A(n7922), .ZN(P1_U3515) );
  INV_X1 U9696 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n7924) );
  MUX2_X1 U9697 ( .A(n7924), .B(n7923), .S(n10494), .Z(n7925) );
  NOR2_X1 U9698 ( .A1(n9406), .A2(n10383), .ZN(n7928) );
  OAI22_X1 U9699 ( .A1(n9401), .A2(n10117), .B1(n7926), .B2(n10162), .ZN(n7927) );
  AOI211_X1 U9700 ( .C1(n7929), .C2(n10392), .A(n7928), .B(n7927), .ZN(n7932)
         );
  NAND2_X1 U9701 ( .A1(n7930), .A2(n10162), .ZN(n7931) );
  OAI211_X1 U9702 ( .C1(n7933), .C2(n10164), .A(n7932), .B(n7931), .ZN(
        P1_U3268) );
  XNOR2_X1 U9703 ( .A(n7934), .B(n9688), .ZN(n7952) );
  INV_X1 U9704 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n7941) );
  INV_X1 U9705 ( .A(n10060), .ZN(n7937) );
  INV_X1 U9706 ( .A(n7935), .ZN(n7936) );
  AOI211_X1 U9707 ( .C1(n9562), .C2(n7937), .A(n10475), .B(n7936), .ZN(n7946)
         );
  AOI211_X1 U9708 ( .C1(n9688), .C2(n7938), .A(n10152), .B(n10044), .ZN(n7940)
         );
  OAI22_X1 U9709 ( .A1(n9431), .A2(n9537), .B1(n7939), .B2(n9535), .ZN(n9478)
         );
  OR2_X1 U9710 ( .A1(n7940), .A2(n9478), .ZN(n7950) );
  AOI211_X1 U9711 ( .C1(n6090), .C2(n9562), .A(n7946), .B(n7950), .ZN(n7943)
         );
  MUX2_X1 U9712 ( .A(n7941), .B(n7943), .S(n10482), .Z(n7942) );
  OAI21_X1 U9713 ( .B1(n7952), .B2(n10306), .A(n7942), .ZN(P1_U3512) );
  MUX2_X1 U9714 ( .A(n7944), .B(n7943), .S(n10494), .Z(n7945) );
  OAI21_X1 U9715 ( .B1(n7952), .B2(n10243), .A(n7945), .ZN(P1_U3544) );
  NAND2_X1 U9716 ( .A1(n7946), .A2(n10392), .ZN(n7948) );
  AOI22_X1 U9717 ( .A1(n7610), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9479), .B2(
        n10380), .ZN(n7947) );
  OAI211_X1 U9718 ( .C1(n8118), .C2(n10383), .A(n7948), .B(n7947), .ZN(n7949)
         );
  AOI21_X1 U9719 ( .B1(n7950), .B2(n10162), .A(n7949), .ZN(n7951) );
  OAI21_X1 U9720 ( .B1(n7952), .B2(n10164), .A(n7951), .ZN(P1_U3271) );
  INV_X1 U9721 ( .A(n7953), .ZN(n7954) );
  NOR2_X1 U9722 ( .A1(n8981), .A2(n7956), .ZN(n10520) );
  INV_X1 U9723 ( .A(n10520), .ZN(n7966) );
  OAI22_X1 U9724 ( .A1(n9010), .A2(n6245), .B1(n7958), .B2(n9008), .ZN(n7960)
         );
  NOR2_X1 U9725 ( .A1(n10526), .A2(n9069), .ZN(n7959) );
  AOI211_X1 U9726 ( .C1(n9061), .C2(n7961), .A(n7960), .B(n7959), .ZN(n10524)
         );
  MUX2_X1 U9727 ( .A(n7962), .B(n10524), .S(n9091), .Z(n7965) );
  AOI22_X1 U9728 ( .A1(n9029), .A2(n7963), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10518), .ZN(n7964) );
  OAI211_X1 U9729 ( .C1(n10526), .C2(n7966), .A(n7965), .B(n7964), .ZN(
        P2_U3232) );
  XNOR2_X1 U9730 ( .A(n7968), .B(n7967), .ZN(n7969) );
  XNOR2_X1 U9731 ( .A(n7970), .B(n7969), .ZN(n7979) );
  INV_X1 U9732 ( .A(n7979), .ZN(n7971) );
  NAND2_X1 U9733 ( .A1(n7971), .A2(n8320), .ZN(n7985) );
  INV_X1 U9734 ( .A(n7972), .ZN(n7973) );
  AOI22_X1 U9735 ( .A1(n8819), .A2(n8329), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7975) );
  NAND2_X1 U9736 ( .A1(n8834), .A2(n8324), .ZN(n7974) );
  OAI211_X1 U9737 ( .C1(n7976), .C2(n8326), .A(n7975), .B(n7974), .ZN(n7981)
         );
  NOR4_X1 U9738 ( .A1(n7979), .A2(n7978), .A3(n7977), .A4(n8318), .ZN(n7980)
         );
  AOI211_X1 U9739 ( .C1(n9186), .C2(n8316), .A(n7981), .B(n7980), .ZN(n7982)
         );
  OAI211_X1 U9740 ( .C1(n7985), .C2(n7984), .A(n7983), .B(n7982), .ZN(P2_U3160) );
  INV_X1 U9741 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7987) );
  OAI22_X1 U9742 ( .A1(n9352), .A2(n10117), .B1(n7987), .B2(n10162), .ZN(n7988) );
  AOI21_X1 U9743 ( .B1(n9347), .B2(n10079), .A(n7988), .ZN(n7989) );
  OAI21_X1 U9744 ( .B1(n7990), .B2(n10082), .A(n7989), .ZN(n7991) );
  OAI21_X1 U9745 ( .B1(n7986), .B2(n7610), .A(n7993), .ZN(P1_U3265) );
  INV_X1 U9746 ( .A(n7994), .ZN(n7995) );
  INV_X1 U9747 ( .A(n7997), .ZN(n7998) );
  AND2_X1 U9748 ( .A1(n7610), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8000) );
  NOR2_X1 U9749 ( .A1(n8001), .A2(n8000), .ZN(n8003) );
  NAND2_X1 U9750 ( .A1(n9730), .A2(n10079), .ZN(n8002) );
  OAI211_X1 U9751 ( .C1(n10171), .C2(n10082), .A(n8003), .B(n8002), .ZN(
        P1_U3264) );
  INV_X1 U9752 ( .A(n8004), .ZN(n9303) );
  OAI222_X1 U9753 ( .A1(n10332), .A2(n8006), .B1(n10311), .B2(n8005), .C1(
        n10335), .C2(n9303), .ZN(P1_U3327) );
  OAI22_X1 U9754 ( .A1(n10042), .A2(n8163), .B1(n9431), .B2(n5421), .ZN(n8007)
         );
  XNOR2_X1 U9755 ( .A(n8007), .B(n9345), .ZN(n8009) );
  OAI22_X1 U9756 ( .A1(n10042), .A2(n5421), .B1(n9431), .B2(n8165), .ZN(n8008)
         );
  AOI21_X1 U9757 ( .B1(n8009), .B2(n8008), .A(n9426), .ZN(n8120) );
  NAND2_X1 U9758 ( .A1(n10194), .A2(n8137), .ZN(n8011) );
  NAND2_X1 U9759 ( .A1(n9820), .A2(n8108), .ZN(n8010) );
  NAND2_X1 U9760 ( .A1(n8011), .A2(n8010), .ZN(n8012) );
  XNOR2_X1 U9761 ( .A(n8012), .B(n9345), .ZN(n9377) );
  NAND2_X1 U9762 ( .A1(n10194), .A2(n4427), .ZN(n8014) );
  NAND2_X1 U9763 ( .A1(n9820), .A2(n9342), .ZN(n8013) );
  NAND2_X1 U9764 ( .A1(n8014), .A2(n8013), .ZN(n8115) );
  OAI22_X1 U9765 ( .A1(n8163), .A2(n9370), .B1(n8015), .B2(n5421), .ZN(n8016)
         );
  XNOR2_X1 U9766 ( .A(n8016), .B(n9345), .ZN(n9365) );
  OR2_X1 U9767 ( .A1(n9370), .A2(n5421), .ZN(n8018) );
  NAND2_X1 U9768 ( .A1(n9342), .A2(n9833), .ZN(n8017) );
  NAND2_X1 U9769 ( .A1(n8018), .A2(n8017), .ZN(n9366) );
  NAND2_X1 U9770 ( .A1(n9365), .A2(n9366), .ZN(n8019) );
  NAND2_X1 U9771 ( .A1(n9364), .A2(n8019), .ZN(n8029) );
  INV_X1 U9772 ( .A(n9365), .ZN(n9440) );
  NAND2_X1 U9773 ( .A1(n8020), .A2(n9366), .ZN(n8022) );
  INV_X1 U9774 ( .A(n8020), .ZN(n9363) );
  INV_X1 U9775 ( .A(n9366), .ZN(n8021) );
  AOI22_X1 U9776 ( .A1(n9440), .A2(n8022), .B1(n9363), .B2(n8021), .ZN(n8027)
         );
  NAND2_X1 U9777 ( .A1(n8026), .A2(n8137), .ZN(n8024) );
  NAND2_X1 U9778 ( .A1(n9832), .A2(n4427), .ZN(n8023) );
  NAND2_X1 U9779 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  XNOR2_X1 U9780 ( .A(n8025), .B(n9345), .ZN(n8030) );
  AOI22_X1 U9781 ( .A1(n8026), .A2(n4427), .B1(n9342), .B2(n9832), .ZN(n8031)
         );
  XNOR2_X1 U9782 ( .A(n8030), .B(n8031), .ZN(n9442) );
  AND2_X1 U9783 ( .A1(n8027), .A2(n9442), .ZN(n8028) );
  INV_X1 U9784 ( .A(n8030), .ZN(n8032) );
  OR2_X1 U9785 ( .A1(n8032), .A2(n8031), .ZN(n8033) );
  NAND2_X1 U9786 ( .A1(n8039), .A2(n8137), .ZN(n8035) );
  NAND2_X1 U9787 ( .A1(n9831), .A2(n4427), .ZN(n8034) );
  NAND2_X1 U9788 ( .A1(n8035), .A2(n8034), .ZN(n8036) );
  XNOR2_X1 U9789 ( .A(n8036), .B(n8141), .ZN(n8046) );
  NOR2_X1 U9790 ( .A1(n8037), .A2(n8165), .ZN(n8038) );
  AOI21_X1 U9791 ( .B1(n8039), .B2(n4427), .A(n8038), .ZN(n9328) );
  NAND2_X1 U9792 ( .A1(n9603), .A2(n8137), .ZN(n8041) );
  NAND2_X1 U9793 ( .A1(n9830), .A2(n4427), .ZN(n8040) );
  NAND2_X1 U9794 ( .A1(n8041), .A2(n8040), .ZN(n8042) );
  XNOR2_X1 U9795 ( .A(n8042), .B(n8141), .ZN(n8045) );
  NOR2_X1 U9796 ( .A1(n9601), .A2(n8165), .ZN(n8043) );
  AOI21_X1 U9797 ( .B1(n9603), .B2(n4427), .A(n8043), .ZN(n8044) );
  NAND2_X1 U9798 ( .A1(n8045), .A2(n8044), .ZN(n8048) );
  OAI21_X1 U9799 ( .B1(n8045), .B2(n8044), .A(n8048), .ZN(n9488) );
  INV_X1 U9800 ( .A(n8046), .ZN(n9326) );
  INV_X1 U9801 ( .A(n9328), .ZN(n8047) );
  INV_X1 U9802 ( .A(n8048), .ZN(n9387) );
  NAND2_X1 U9803 ( .A1(n10240), .A2(n8137), .ZN(n8050) );
  NAND2_X1 U9804 ( .A1(n9829), .A2(n4427), .ZN(n8049) );
  NAND2_X1 U9805 ( .A1(n8050), .A2(n8049), .ZN(n8051) );
  XNOR2_X1 U9806 ( .A(n8051), .B(n8141), .ZN(n8053) );
  NOR2_X1 U9807 ( .A1(n9605), .A2(n8165), .ZN(n8052) );
  AOI21_X1 U9808 ( .B1(n10240), .B2(n4427), .A(n8052), .ZN(n8054) );
  NAND2_X1 U9809 ( .A1(n8053), .A2(n8054), .ZN(n8058) );
  INV_X1 U9810 ( .A(n8053), .ZN(n8056) );
  INV_X1 U9811 ( .A(n8054), .ZN(n8055) );
  NAND2_X1 U9812 ( .A1(n8056), .A2(n8055), .ZN(n8057) );
  AND2_X1 U9813 ( .A1(n8058), .A2(n8057), .ZN(n9386) );
  NAND2_X1 U9814 ( .A1(n10235), .A2(n8137), .ZN(n8060) );
  NAND2_X1 U9815 ( .A1(n9828), .A2(n4427), .ZN(n8059) );
  NAND2_X1 U9816 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  XNOR2_X1 U9817 ( .A(n8061), .B(n9345), .ZN(n8069) );
  NOR2_X1 U9818 ( .A1(n8062), .A2(n8165), .ZN(n8063) );
  AOI21_X1 U9819 ( .B1(n10235), .B2(n4427), .A(n8063), .ZN(n8070) );
  XNOR2_X1 U9820 ( .A(n8069), .B(n8070), .ZN(n9464) );
  OAI22_X1 U9821 ( .A1(n8066), .A2(n8163), .B1(n8064), .B2(n5421), .ZN(n8065)
         );
  XNOR2_X1 U9822 ( .A(n8065), .B(n9345), .ZN(n9316) );
  OR2_X1 U9823 ( .A1(n8066), .A2(n5421), .ZN(n8068) );
  NAND2_X1 U9824 ( .A1(n9827), .A2(n9342), .ZN(n8067) );
  NAND2_X1 U9825 ( .A1(n8068), .A2(n8067), .ZN(n9315) );
  INV_X1 U9826 ( .A(n8069), .ZN(n8071) );
  NAND2_X1 U9827 ( .A1(n8071), .A2(n8070), .ZN(n9314) );
  INV_X1 U9828 ( .A(n9316), .ZN(n8074) );
  INV_X1 U9829 ( .A(n9315), .ZN(n8073) );
  NAND2_X1 U9830 ( .A1(n10225), .A2(n4427), .ZN(n8076) );
  NAND2_X1 U9831 ( .A1(n9342), .A2(n9826), .ZN(n8075) );
  NAND2_X1 U9832 ( .A1(n8076), .A2(n8075), .ZN(n8085) );
  INV_X1 U9833 ( .A(n8085), .ZN(n9549) );
  NAND2_X1 U9834 ( .A1(n10225), .A2(n8137), .ZN(n8078) );
  NAND2_X1 U9835 ( .A1(n9826), .A2(n4427), .ZN(n8077) );
  NAND2_X1 U9836 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  XNOR2_X1 U9837 ( .A(n8079), .B(n9345), .ZN(n9410) );
  INV_X1 U9838 ( .A(n9410), .ZN(n8084) );
  NAND2_X1 U9839 ( .A1(n10220), .A2(n8137), .ZN(n8081) );
  NAND2_X1 U9840 ( .A1(n9825), .A2(n4427), .ZN(n8080) );
  NAND2_X1 U9841 ( .A1(n8081), .A2(n8080), .ZN(n8082) );
  XNOR2_X1 U9842 ( .A(n8082), .B(n8141), .ZN(n8088) );
  INV_X1 U9843 ( .A(n8088), .ZN(n9409) );
  OAI22_X1 U9844 ( .A1(n10144), .A2(n5421), .B1(n8083), .B2(n8165), .ZN(n9408)
         );
  NAND2_X1 U9845 ( .A1(n9409), .A2(n9408), .ZN(n9407) );
  OAI21_X1 U9846 ( .B1(n9549), .B2(n8084), .A(n9407), .ZN(n8090) );
  OAI21_X1 U9847 ( .B1(n9410), .B2(n8085), .A(n9408), .ZN(n8087) );
  NOR3_X1 U9848 ( .A1(n9408), .A2(n8085), .A3(n9410), .ZN(n8086) );
  AOI21_X1 U9849 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8089) );
  OAI22_X1 U9850 ( .A1(n10116), .A2(n8163), .B1(n9506), .B2(n5421), .ZN(n8091)
         );
  XNOR2_X1 U9851 ( .A(n8091), .B(n9345), .ZN(n8095) );
  OR2_X1 U9852 ( .A1(n10116), .A2(n5421), .ZN(n8093) );
  INV_X1 U9853 ( .A(n9506), .ZN(n9824) );
  NAND2_X1 U9854 ( .A1(n9824), .A2(n9342), .ZN(n8092) );
  NAND2_X1 U9855 ( .A1(n8093), .A2(n8092), .ZN(n8096) );
  NAND2_X1 U9856 ( .A1(n8095), .A2(n8096), .ZN(n9497) );
  AOI22_X1 U9857 ( .A1(n6067), .A2(n4427), .B1(n9342), .B2(n9823), .ZN(n9503)
         );
  INV_X1 U9858 ( .A(n9503), .ZN(n8099) );
  AOI22_X1 U9859 ( .A1(n6067), .A2(n8137), .B1(n4427), .B2(n9823), .ZN(n8094)
         );
  XNOR2_X1 U9860 ( .A(n8094), .B(n9345), .ZN(n8100) );
  INV_X1 U9861 ( .A(n8100), .ZN(n8101) );
  INV_X1 U9862 ( .A(n8095), .ZN(n8098) );
  INV_X1 U9863 ( .A(n8096), .ZN(n8097) );
  NAND2_X1 U9864 ( .A1(n8098), .A2(n8097), .ZN(n9419) );
  AND2_X1 U9865 ( .A1(n8101), .A2(n9419), .ZN(n9499) );
  AND2_X1 U9866 ( .A1(n9497), .A2(n8100), .ZN(n8102) );
  AOI22_X1 U9867 ( .A1(n10206), .A2(n8137), .B1(n4427), .B2(n9822), .ZN(n8103)
         );
  XNOR2_X1 U9868 ( .A(n8103), .B(n9345), .ZN(n8104) );
  AOI22_X1 U9869 ( .A1(n10206), .A2(n4427), .B1(n9342), .B2(n9822), .ZN(n8105)
         );
  XNOR2_X1 U9870 ( .A(n8104), .B(n8105), .ZN(n9336) );
  INV_X1 U9871 ( .A(n8104), .ZN(n8107) );
  INV_X1 U9872 ( .A(n8105), .ZN(n8106) );
  AOI22_X1 U9873 ( .A1(n10197), .A2(n8137), .B1(n8108), .B2(n9821), .ZN(n8109)
         );
  XNOR2_X1 U9874 ( .A(n8109), .B(n9345), .ZN(n8110) );
  AOI22_X1 U9875 ( .A1(n10197), .A2(n4427), .B1(n9342), .B2(n9821), .ZN(n8111)
         );
  NAND2_X1 U9876 ( .A1(n8110), .A2(n8111), .ZN(n9453) );
  INV_X1 U9877 ( .A(n8110), .ZN(n8113) );
  INV_X1 U9878 ( .A(n8111), .ZN(n8112) );
  NAND2_X1 U9879 ( .A1(n8113), .A2(n8112), .ZN(n9454) );
  NAND2_X1 U9880 ( .A1(n8114), .A2(n9454), .ZN(n9379) );
  INV_X1 U9881 ( .A(n9377), .ZN(n8116) );
  INV_X1 U9882 ( .A(n8115), .ZN(n9376) );
  AOI22_X1 U9883 ( .A1(n9562), .A2(n8137), .B1(n4427), .B2(n9819), .ZN(n8117)
         );
  XOR2_X1 U9884 ( .A(n9345), .B(n8117), .Z(n9474) );
  OAI22_X1 U9885 ( .A1(n8118), .A2(n5421), .B1(n9561), .B2(n8165), .ZN(n9475)
         );
  OAI21_X1 U9886 ( .B1(n8120), .B2(n8119), .A(n8136), .ZN(n8121) );
  NAND2_X1 U9887 ( .A1(n8121), .A2(n9533), .ZN(n8125) );
  OAI22_X1 U9888 ( .A1(n8122), .A2(n9537), .B1(n9561), .B2(n9535), .ZN(n10049)
         );
  OAI22_X1 U9889 ( .A1(n10039), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8716), .ZN(n8123) );
  AOI21_X1 U9890 ( .B1(n10049), .B2(n9542), .A(n8123), .ZN(n8124) );
  OAI211_X1 U9891 ( .C1(n10042), .C2(n9545), .A(n8125), .B(n8124), .ZN(
        P1_U3216) );
  NOR2_X1 U9892 ( .A1(n8127), .A2(n9087), .ZN(n8809) );
  AOI21_X1 U9893 ( .B1(n8981), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8809), .ZN(
        n8128) );
  OAI21_X1 U9894 ( .B1(n8129), .B2(n9090), .A(n8128), .ZN(n8130) );
  AOI21_X1 U9895 ( .B1(n8131), .B2(n10520), .A(n8130), .ZN(n8132) );
  OAI21_X1 U9896 ( .B1(n8126), .B2(n8981), .A(n8132), .ZN(P2_U3204) );
  INV_X1 U9897 ( .A(n8133), .ZN(n10330) );
  OAI222_X1 U9898 ( .A1(n6680), .A2(P2_U3151), .B1(n9307), .B2(n10330), .C1(
        n8135), .C2(n8134), .ZN(P2_U3270) );
  NAND2_X1 U9899 ( .A1(n6074), .A2(n8137), .ZN(n8140) );
  NAND2_X1 U9900 ( .A1(n9818), .A2(n4427), .ZN(n8139) );
  NAND2_X1 U9901 ( .A1(n8140), .A2(n8139), .ZN(n8142) );
  XNOR2_X1 U9902 ( .A(n8142), .B(n8141), .ZN(n8144) );
  AND2_X1 U9903 ( .A1(n9818), .A2(n9342), .ZN(n8143) );
  AOI21_X1 U9904 ( .B1(n6074), .B2(n4427), .A(n8143), .ZN(n8145) );
  NAND2_X1 U9905 ( .A1(n8144), .A2(n8145), .ZN(n8149) );
  INV_X1 U9906 ( .A(n8144), .ZN(n8147) );
  INV_X1 U9907 ( .A(n8145), .ZN(n8146) );
  NAND2_X1 U9908 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  OAI22_X1 U9909 ( .A1(n9406), .A2(n5421), .B1(n9536), .B2(n8165), .ZN(n8156)
         );
  OAI22_X1 U9910 ( .A1(n9406), .A2(n8163), .B1(n9536), .B2(n5421), .ZN(n8150)
         );
  XNOR2_X1 U9911 ( .A(n8150), .B(n9345), .ZN(n8155) );
  XOR2_X1 U9912 ( .A(n8156), .B(n8155), .Z(n9398) );
  NAND2_X1 U9913 ( .A1(n10016), .A2(n8137), .ZN(n8152) );
  NAND2_X1 U9914 ( .A1(n9816), .A2(n4427), .ZN(n8151) );
  NAND2_X1 U9915 ( .A1(n8152), .A2(n8151), .ZN(n8153) );
  XNOR2_X1 U9916 ( .A(n8153), .B(n9345), .ZN(n8162) );
  AND2_X1 U9917 ( .A1(n9816), .A2(n9342), .ZN(n8154) );
  AOI21_X1 U9918 ( .B1(n10016), .B2(n4427), .A(n8154), .ZN(n8160) );
  XNOR2_X1 U9919 ( .A(n8162), .B(n8160), .ZN(n9534) );
  INV_X1 U9920 ( .A(n8155), .ZN(n8158) );
  INV_X1 U9921 ( .A(n8156), .ZN(n8157) );
  NAND2_X1 U9922 ( .A1(n8158), .A2(n8157), .ZN(n9530) );
  INV_X1 U9923 ( .A(n8160), .ZN(n8161) );
  NAND2_X1 U9924 ( .A1(n8162), .A2(n8161), .ZN(n8169) );
  OAI22_X1 U9925 ( .A1(n10175), .A2(n8163), .B1(n9538), .B2(n5421), .ZN(n8164)
         );
  XNOR2_X1 U9926 ( .A(n8164), .B(n9345), .ZN(n8167) );
  OAI22_X1 U9927 ( .A1(n10175), .A2(n5421), .B1(n9538), .B2(n8165), .ZN(n8166)
         );
  NOR2_X1 U9928 ( .A1(n8167), .A2(n8166), .ZN(n9357) );
  AOI21_X1 U9929 ( .B1(n8167), .B2(n8166), .A(n9357), .ZN(n8168) );
  AOI21_X1 U9930 ( .B1(n9532), .B2(n8169), .A(n8168), .ZN(n8173) );
  INV_X1 U9931 ( .A(n8168), .ZN(n8171) );
  INV_X1 U9932 ( .A(n8169), .ZN(n8170) );
  NOR2_X1 U9933 ( .A1(n8171), .A2(n8170), .ZN(n8172) );
  AOI22_X1 U9934 ( .A1(n9815), .A2(n9522), .B1(n4420), .B2(n9816), .ZN(n9999)
         );
  INV_X1 U9935 ( .A(n10002), .ZN(n8174) );
  OAI22_X1 U9936 ( .A1(n8174), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8723), .ZN(n8175) );
  AOI21_X1 U9937 ( .B1(n5009), .B2(n9542), .A(n8175), .ZN(n8176) );
  OAI222_X1 U9938 ( .A1(n10332), .A2(n8178), .B1(n10335), .B2(n8177), .C1(
        P1_U3086), .C2(n7066), .ZN(P1_U3333) );
  XOR2_X1 U9939 ( .A(n8180), .B(n8179), .Z(n8185) );
  AOI22_X1 U9940 ( .A1(n8310), .A2(n8976), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8182) );
  NAND2_X1 U9941 ( .A1(n8329), .A2(n8979), .ZN(n8181) );
  OAI211_X1 U9942 ( .C1(n6722), .C2(n8313), .A(n8182), .B(n8181), .ZN(n8183)
         );
  AOI21_X1 U9943 ( .B1(n9260), .B2(n8316), .A(n8183), .ZN(n8184) );
  OAI21_X1 U9944 ( .B1(n8185), .B2(n8318), .A(n8184), .ZN(P2_U3155) );
  INV_X1 U9945 ( .A(n8187), .ZN(n8188) );
  AOI22_X1 U9946 ( .A1(n8896), .A2(n8324), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8191) );
  NAND2_X1 U9947 ( .A1(n8874), .A2(n8329), .ZN(n8190) );
  OAI211_X1 U9948 ( .C1(n8232), .C2(n8326), .A(n8191), .B(n8190), .ZN(n8192)
         );
  AOI21_X1 U9949 ( .B1(n9216), .B2(n8316), .A(n8192), .ZN(n8193) );
  OAI21_X1 U9950 ( .B1(n8194), .B2(n8318), .A(n8193), .ZN(P2_U3156) );
  XNOR2_X1 U9951 ( .A(n8286), .B(n9066), .ZN(n8288) );
  XOR2_X1 U9952 ( .A(n8287), .B(n8288), .Z(n8200) );
  NAND2_X1 U9953 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8348) );
  OAI21_X1 U9954 ( .B1(n8326), .B2(n9009), .A(n8348), .ZN(n8195) );
  AOI21_X1 U9955 ( .B1(n8324), .B2(n9047), .A(n8195), .ZN(n8196) );
  OAI21_X1 U9956 ( .B1(n9036), .B2(n8294), .A(n8196), .ZN(n8197) );
  AOI21_X1 U9957 ( .B1(n8198), .B2(n8316), .A(n8197), .ZN(n8199) );
  OAI21_X1 U9958 ( .B1(n8200), .B2(n8318), .A(n8199), .ZN(P2_U3157) );
  XOR2_X1 U9959 ( .A(n8201), .B(n8202), .Z(n8208) );
  NAND2_X1 U9960 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8793) );
  NAND2_X1 U9961 ( .A1(n8324), .A2(n8943), .ZN(n8203) );
  OAI211_X1 U9962 ( .C1(n8204), .C2(n8326), .A(n8793), .B(n8203), .ZN(n8205)
         );
  AOI21_X1 U9963 ( .B1(n8921), .B2(n8329), .A(n8205), .ZN(n8207) );
  NAND2_X1 U9964 ( .A1(n9238), .A2(n8316), .ZN(n8206) );
  OAI211_X1 U9965 ( .C1(n8208), .C2(n8318), .A(n8207), .B(n8206), .ZN(P2_U3159) );
  XOR2_X1 U9966 ( .A(n8210), .B(n4899), .Z(n8216) );
  AOI22_X1 U9967 ( .A1(n8918), .A2(n8324), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8212) );
  NAND2_X1 U9968 ( .A1(n8899), .A2(n8329), .ZN(n8211) );
  OAI211_X1 U9969 ( .C1(n8213), .C2(n8326), .A(n8212), .B(n8211), .ZN(n8214)
         );
  AOI21_X1 U9970 ( .B1(n9226), .B2(n8316), .A(n8214), .ZN(n8215) );
  OAI21_X1 U9971 ( .B1(n8216), .B2(n8318), .A(n8215), .ZN(P2_U3163) );
  OAI211_X1 U9972 ( .C1(n8219), .C2(n8218), .A(n8217), .B(n8320), .ZN(n8223)
         );
  NAND2_X1 U9973 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8387) );
  OAI21_X1 U9974 ( .B1(n8326), .B2(n6722), .A(n8387), .ZN(n8221) );
  NOR2_X1 U9975 ( .A1(n8294), .A2(n9012), .ZN(n8220) );
  AOI211_X1 U9976 ( .C1(n8324), .C2(n9046), .A(n8221), .B(n8220), .ZN(n8222)
         );
  OAI211_X1 U9977 ( .C1(n8224), .C2(n8332), .A(n8223), .B(n8222), .ZN(P2_U3164) );
  INV_X1 U9978 ( .A(n8225), .ZN(n8254) );
  NOR3_X1 U9979 ( .A1(n8254), .A2(n5312), .A3(n8227), .ZN(n8230) );
  INV_X1 U9980 ( .A(n8228), .ZN(n8229) );
  OAI21_X1 U9981 ( .B1(n8230), .B2(n8229), .A(n8320), .ZN(n8235) );
  AOI22_X1 U9982 ( .A1(n8843), .A2(n8329), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8231) );
  OAI21_X1 U9983 ( .B1(n8232), .B2(n8313), .A(n8231), .ZN(n8233) );
  AOI21_X1 U9984 ( .B1(n8841), .B2(n8310), .A(n8233), .ZN(n8234) );
  OAI211_X1 U9985 ( .C1(n8236), .C2(n8332), .A(n8235), .B(n8234), .ZN(P2_U3165) );
  AOI21_X1 U9986 ( .B1(n8238), .B2(n8237), .A(n4462), .ZN(n8243) );
  OAI22_X1 U9987 ( .A1(n8326), .A2(n8954), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8738), .ZN(n8240) );
  NOR2_X1 U9988 ( .A1(n8313), .A2(n8953), .ZN(n8239) );
  AOI211_X1 U9989 ( .C1(n8959), .C2(n8329), .A(n8240), .B(n8239), .ZN(n8242)
         );
  NAND2_X1 U9990 ( .A1(n9253), .A2(n8316), .ZN(n8241) );
  OAI211_X1 U9991 ( .C1(n8243), .C2(n8318), .A(n8242), .B(n8241), .ZN(P2_U3166) );
  INV_X1 U9992 ( .A(n8948), .ZN(n9247) );
  NOR3_X1 U9993 ( .A1(n4462), .A2(n4555), .A3(n8244), .ZN(n8247) );
  INV_X1 U9994 ( .A(n8245), .ZN(n8246) );
  OAI21_X1 U9995 ( .B1(n8247), .B2(n8246), .A(n8320), .ZN(n8251) );
  NAND2_X1 U9996 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U9997 ( .A1(n8324), .A2(n8964), .ZN(n8248) );
  OAI211_X1 U9998 ( .C1(n6733), .C2(n8326), .A(n8492), .B(n8248), .ZN(n8249)
         );
  AOI21_X1 U9999 ( .B1(n8947), .B2(n8329), .A(n8249), .ZN(n8250) );
  OAI211_X1 U10000 ( .C1(n9247), .C2(n8332), .A(n8251), .B(n8250), .ZN(
        P2_U3168) );
  INV_X1 U10001 ( .A(n8860), .ZN(n8256) );
  AOI22_X1 U10002 ( .A1(n8857), .A2(n8324), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8255) );
  OAI21_X1 U10003 ( .B1(n8256), .B2(n8294), .A(n8255), .ZN(n8257) );
  AOI21_X1 U10004 ( .B1(n8858), .B2(n8310), .A(n8257), .ZN(n8258) );
  XOR2_X1 U10005 ( .A(n8260), .B(n8259), .Z(n8265) );
  AOI22_X1 U10006 ( .A1(n8908), .A2(n8310), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8262) );
  NAND2_X1 U10007 ( .A1(n8329), .A2(n8911), .ZN(n8261) );
  OAI211_X1 U10008 ( .C1(n8926), .C2(n8313), .A(n8262), .B(n8261), .ZN(n8263)
         );
  AOI21_X1 U10009 ( .B1(n9232), .B2(n8316), .A(n8263), .ZN(n8264) );
  OAI21_X1 U10010 ( .B1(n8265), .B2(n8318), .A(n8264), .ZN(P2_U3173) );
  INV_X1 U10011 ( .A(n8266), .ZN(n8267) );
  AOI21_X1 U10012 ( .B1(n8269), .B2(n8268), .A(n8267), .ZN(n8274) );
  AOI22_X1 U10013 ( .A1(n8310), .A2(n8991), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8271) );
  NAND2_X1 U10014 ( .A1(n8324), .A2(n9024), .ZN(n8270) );
  OAI211_X1 U10015 ( .C1(n8294), .C2(n8994), .A(n8271), .B(n8270), .ZN(n8272)
         );
  AOI21_X1 U10016 ( .B1(n9266), .B2(n8316), .A(n8272), .ZN(n8273) );
  OAI21_X1 U10017 ( .B1(n8274), .B2(n8318), .A(n8273), .ZN(P2_U3174) );
  NAND2_X1 U10018 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  XNOR2_X1 U10019 ( .A(n8275), .B(n8278), .ZN(n8285) );
  INV_X1 U10020 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8279) );
  OAI22_X1 U10021 ( .A1(n8882), .A2(n8313), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8279), .ZN(n8281) );
  NOR2_X1 U10022 ( .A1(n8881), .A2(n8326), .ZN(n8280) );
  AOI211_X1 U10023 ( .C1(n8886), .C2(n8329), .A(n8281), .B(n8280), .ZN(n8284)
         );
  NAND2_X1 U10024 ( .A1(n8282), .A2(n8316), .ZN(n8283) );
  OAI211_X1 U10025 ( .C1(n8285), .C2(n8318), .A(n8284), .B(n8283), .ZN(
        P2_U3175) );
  OAI22_X1 U10026 ( .A1(n8288), .A2(n8287), .B1(n9066), .B2(n8286), .ZN(n8289)
         );
  XOR2_X1 U10027 ( .A(n8290), .B(n8289), .Z(n8297) );
  NAND2_X1 U10028 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8364) );
  OAI21_X1 U10029 ( .B1(n8326), .B2(n8291), .A(n8364), .ZN(n8292) );
  AOI21_X1 U10030 ( .B1(n8324), .B2(n9066), .A(n8292), .ZN(n8293) );
  OAI21_X1 U10031 ( .B1(n9027), .B2(n8294), .A(n8293), .ZN(n8295) );
  AOI21_X1 U10032 ( .B1(n9276), .B2(n8316), .A(n8295), .ZN(n8296) );
  OAI21_X1 U10033 ( .B1(n8297), .B2(n8318), .A(n8296), .ZN(P2_U3176) );
  XOR2_X1 U10034 ( .A(n8299), .B(n8298), .Z(n8304) );
  NAND2_X1 U10035 ( .A1(n8335), .A2(n8324), .ZN(n8300) );
  NAND2_X1 U10036 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8776) );
  OAI211_X1 U10037 ( .C1(n8926), .C2(n8326), .A(n8300), .B(n8776), .ZN(n8302)
         );
  NOR2_X1 U10038 ( .A1(n9245), .A2(n8332), .ZN(n8301) );
  AOI211_X1 U10039 ( .C1(n8931), .C2(n8329), .A(n8302), .B(n8301), .ZN(n8303)
         );
  OAI21_X1 U10040 ( .B1(n8304), .B2(n8318), .A(n8303), .ZN(P2_U3178) );
  INV_X1 U10041 ( .A(n8306), .ZN(n8308) );
  NAND2_X1 U10042 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  XNOR2_X1 U10043 ( .A(n8305), .B(n8309), .ZN(n8319) );
  NAND2_X1 U10044 ( .A1(n8834), .A2(n8310), .ZN(n8312) );
  AOI22_X1 U10045 ( .A1(n8837), .A2(n8329), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8311) );
  OAI211_X1 U10046 ( .C1(n8314), .C2(n8313), .A(n8312), .B(n8311), .ZN(n8315)
         );
  AOI21_X1 U10047 ( .B1(n9198), .B2(n8316), .A(n8315), .ZN(n8317) );
  OAI21_X1 U10048 ( .B1(n8319), .B2(n8318), .A(n8317), .ZN(P2_U3180) );
  INV_X1 U10049 ( .A(n9144), .ZN(n8333) );
  OAI211_X1 U10050 ( .C1(n8323), .C2(n8322), .A(n8321), .B(n8320), .ZN(n8331)
         );
  NAND2_X1 U10051 ( .A1(n8324), .A2(n8991), .ZN(n8325) );
  NAND2_X1 U10052 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8447) );
  OAI211_X1 U10053 ( .C1(n8327), .C2(n8326), .A(n8325), .B(n8447), .ZN(n8328)
         );
  AOI21_X1 U10054 ( .B1(n8968), .B2(n8329), .A(n8328), .ZN(n8330) );
  OAI211_X1 U10055 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8330), .ZN(
        P2_U3181) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8334), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10057 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8817), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8826), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10059 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8834), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10060 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8841), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10061 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8858), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10062 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8871), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10063 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8896), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10064 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8908), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10065 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8918), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10066 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8907), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10067 ( .A(n8943), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8774), .Z(
        P2_U3509) );
  MUX2_X1 U10068 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8335), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10069 ( .A(n8964), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8774), .Z(
        P2_U3507) );
  MUX2_X1 U10070 ( .A(n8976), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8774), .Z(
        P2_U3506) );
  MUX2_X1 U10071 ( .A(n8991), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8774), .Z(
        P2_U3505) );
  MUX2_X1 U10072 ( .A(n8975), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8774), .Z(
        P2_U3504) );
  MUX2_X1 U10073 ( .A(n9024), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8774), .Z(
        P2_U3503) );
  MUX2_X1 U10074 ( .A(n9046), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8774), .Z(
        P2_U3502) );
  MUX2_X1 U10075 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9066), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10076 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n9047), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10077 ( .A(n9063), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8774), .Z(
        P2_U3499) );
  MUX2_X1 U10078 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8336), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10079 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8337), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10080 ( .A(n8338), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8774), .Z(
        P2_U3496) );
  MUX2_X1 U10081 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n7367), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10082 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n6694), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10083 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8339), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U10084 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8340), .S(P2_U3893), .Z(
        P2_U3492) );
  MUX2_X1 U10085 ( .A(n6239), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8774), .Z(
        P2_U3491) );
  XNOR2_X1 U10086 ( .A(n8367), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8358) );
  XOR2_X1 U10087 ( .A(n8358), .B(n8359), .Z(n8357) );
  INV_X1 U10088 ( .A(n8342), .ZN(n8343) );
  MUX2_X1 U10089 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8770), .Z(n8361) );
  XOR2_X1 U10090 ( .A(n8361), .B(n8367), .Z(n8362) );
  XNOR2_X1 U10091 ( .A(n8363), .B(n8362), .ZN(n8355) );
  NAND2_X1 U10092 ( .A1(n10513), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n8347) );
  OAI211_X1 U10093 ( .C1(n8795), .C2(n8360), .A(n8348), .B(n8347), .ZN(n8354)
         );
  XNOR2_X1 U10094 ( .A(n8367), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8349) );
  OR3_X1 U10095 ( .A1(n8351), .A2(n8350), .A3(n8349), .ZN(n8352) );
  AOI21_X1 U10096 ( .B1(n8369), .B2(n8352), .A(n10503), .ZN(n8353) );
  AOI211_X1 U10097 ( .C1(n8797), .C2(n8355), .A(n8354), .B(n8353), .ZN(n8356)
         );
  OAI21_X1 U10098 ( .B1(n8357), .B2(n8781), .A(n8356), .ZN(P2_U3192) );
  XNOR2_X1 U10099 ( .A(n8380), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n8378) );
  MUX2_X1 U10100 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8770), .Z(n8381) );
  XNOR2_X1 U10101 ( .A(n8381), .B(n8383), .ZN(n8384) );
  XNOR2_X1 U10102 ( .A(n8385), .B(n8384), .ZN(n8376) );
  NAND2_X1 U10103 ( .A1(n10513), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8365) );
  OAI211_X1 U10104 ( .C1(n8795), .C2(n8370), .A(n8365), .B(n8364), .ZN(n8375)
         );
  AOI21_X1 U10105 ( .B1(n9026), .B2(n8372), .A(n8389), .ZN(n8373) );
  NOR2_X1 U10106 ( .A1(n8373), .A2(n10503), .ZN(n8374) );
  AOI211_X1 U10107 ( .C1(n8376), .C2(n8797), .A(n8375), .B(n8374), .ZN(n8377)
         );
  OAI21_X1 U10108 ( .B1(n8781), .B2(n8378), .A(n8377), .ZN(P2_U3193) );
  XNOR2_X1 U10109 ( .A(n8408), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8398) );
  INV_X1 U10110 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9158) );
  XOR2_X1 U10111 ( .A(n8398), .B(n8399), .Z(n8397) );
  INV_X1 U10112 ( .A(n8381), .ZN(n8382) );
  MUX2_X1 U10113 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8770), .Z(n8401) );
  XOR2_X1 U10114 ( .A(n8401), .B(n8408), .Z(n8402) );
  XNOR2_X1 U10115 ( .A(n8403), .B(n8402), .ZN(n8395) );
  NAND2_X1 U10116 ( .A1(n10513), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n8386) );
  OAI211_X1 U10117 ( .C1(n8795), .C2(n8400), .A(n8387), .B(n8386), .ZN(n8394)
         );
  INV_X1 U10118 ( .A(n8388), .ZN(n8391) );
  XNOR2_X1 U10119 ( .A(n8408), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8390) );
  OR3_X1 U10120 ( .A1(n8389), .A2(n8391), .A3(n8390), .ZN(n8392) );
  AOI21_X1 U10121 ( .B1(n8406), .B2(n8392), .A(n10503), .ZN(n8393) );
  AOI211_X1 U10122 ( .C1(n8797), .C2(n8395), .A(n8394), .B(n8393), .ZN(n8396)
         );
  OAI21_X1 U10123 ( .B1(n8397), .B2(n8781), .A(n8396), .ZN(P2_U3194) );
  INV_X1 U10124 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9151) );
  XNOR2_X1 U10125 ( .A(n8421), .B(n9151), .ZN(n8417) );
  MUX2_X1 U10126 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8770), .Z(n8422) );
  XNOR2_X1 U10127 ( .A(n8424), .B(n8422), .ZN(n8425) );
  XNOR2_X1 U10128 ( .A(n8426), .B(n8425), .ZN(n8415) );
  NAND2_X1 U10129 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n8405) );
  NAND2_X1 U10130 ( .A1(n10513), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8404) );
  OAI211_X1 U10131 ( .C1(n8795), .C2(n8420), .A(n8405), .B(n8404), .ZN(n8414)
         );
  NAND2_X1 U10132 ( .A1(n8411), .A2(n8410), .ZN(n8412) );
  AOI21_X1 U10133 ( .B1(n8433), .B2(n8412), .A(n10503), .ZN(n8413) );
  AOI211_X1 U10134 ( .C1(n8797), .C2(n8415), .A(n8414), .B(n8413), .ZN(n8416)
         );
  OAI21_X1 U10135 ( .B1(n8417), .B2(n8781), .A(n8416), .ZN(P2_U3195) );
  XOR2_X1 U10136 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8448), .Z(n8440) );
  INV_X1 U10137 ( .A(n8418), .ZN(n8419) );
  XOR2_X1 U10138 ( .A(n8440), .B(n8441), .Z(n8439) );
  INV_X1 U10139 ( .A(n8422), .ZN(n8423) );
  MUX2_X1 U10140 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8770), .Z(n8443) );
  XOR2_X1 U10141 ( .A(n8443), .B(n8448), .Z(n8444) );
  XNOR2_X1 U10142 ( .A(n8445), .B(n8444), .ZN(n8437) );
  NAND2_X1 U10143 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3151), .ZN(n8428) );
  NAND2_X1 U10144 ( .A1(n10513), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8427) );
  OAI211_X1 U10145 ( .C1(n8795), .C2(n8442), .A(n8428), .B(n8427), .ZN(n8436)
         );
  XNOR2_X1 U10146 ( .A(n8448), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8430) );
  NAND2_X1 U10147 ( .A1(n8429), .A2(n8430), .ZN(n8450) );
  INV_X1 U10148 ( .A(n8430), .ZN(n8432) );
  NAND3_X1 U10149 ( .A1(n8433), .A2(n8432), .A3(n8431), .ZN(n8434) );
  AOI21_X1 U10150 ( .B1(n8450), .B2(n8434), .A(n10503), .ZN(n8435) );
  AOI211_X1 U10151 ( .C1(n8797), .C2(n8437), .A(n8436), .B(n8435), .ZN(n8438)
         );
  OAI21_X1 U10152 ( .B1(n8439), .B2(n8781), .A(n8438), .ZN(P2_U3196) );
  XOR2_X1 U10153 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8460), .Z(n8459) );
  MUX2_X1 U10154 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8770), .Z(n8461) );
  XNOR2_X1 U10155 ( .A(n8463), .B(n8461), .ZN(n8464) );
  XNOR2_X1 U10156 ( .A(n8465), .B(n8464), .ZN(n8457) );
  NAND2_X1 U10157 ( .A1(n10513), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8446) );
  OAI211_X1 U10158 ( .C1(n8795), .C2(n5101), .A(n8447), .B(n8446), .ZN(n8456)
         );
  INV_X1 U10159 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8453) );
  OR2_X1 U10160 ( .A1(n8448), .A2(n8985), .ZN(n8449) );
  NAND2_X1 U10161 ( .A1(n8451), .A2(n5101), .ZN(n8469) );
  AOI21_X1 U10162 ( .B1(n8453), .B2(n8452), .A(n8472), .ZN(n8454) );
  NOR2_X1 U10163 ( .A1(n8454), .A2(n10503), .ZN(n8455) );
  AOI211_X1 U10164 ( .C1(n8797), .C2(n8457), .A(n8456), .B(n8455), .ZN(n8458)
         );
  OAI21_X1 U10165 ( .B1(n8459), .B2(n8781), .A(n8458), .ZN(P2_U3197) );
  XOR2_X1 U10166 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8479), .Z(n8480) );
  XOR2_X1 U10167 ( .A(n8480), .B(n8481), .Z(n8478) );
  INV_X1 U10168 ( .A(n8461), .ZN(n8462) );
  MUX2_X1 U10169 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8770), .Z(n8488) );
  XOR2_X1 U10170 ( .A(n8479), .B(n8488), .Z(n8489) );
  XNOR2_X1 U10171 ( .A(n8490), .B(n8489), .ZN(n8476) );
  NAND2_X1 U10172 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n8468) );
  NAND2_X1 U10173 ( .A1(n10513), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8467) );
  OAI211_X1 U10174 ( .C1(n8795), .C2(n8487), .A(n8468), .B(n8467), .ZN(n8475)
         );
  INV_X1 U10175 ( .A(n8469), .ZN(n8471) );
  XNOR2_X1 U10176 ( .A(n8479), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n8470) );
  OR3_X1 U10177 ( .A1(n8472), .A2(n8471), .A3(n8470), .ZN(n8473) );
  AOI21_X1 U10178 ( .B1(n8482), .B2(n8473), .A(n10503), .ZN(n8474) );
  AOI211_X1 U10179 ( .C1(n8797), .C2(n8476), .A(n8475), .B(n8474), .ZN(n8477)
         );
  OAI21_X1 U10180 ( .B1(n8478), .B2(n8781), .A(n8477), .ZN(P2_U3198) );
  XNOR2_X1 U10181 ( .A(n8757), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8496) );
  NAND2_X1 U10182 ( .A1(n8484), .A2(n4879), .ZN(n8761) );
  MUX2_X1 U10183 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8770), .Z(n8765) );
  XNOR2_X1 U10184 ( .A(n8765), .B(n8767), .ZN(n8768) );
  XNOR2_X1 U10185 ( .A(n8769), .B(n8768), .ZN(n8494) );
  NAND2_X1 U10186 ( .A1(n10513), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8491) );
  OAI211_X1 U10187 ( .C1(n8795), .C2(n4879), .A(n8492), .B(n8491), .ZN(n8493)
         );
  AOI21_X1 U10188 ( .B1(n8494), .B2(n8797), .A(n8493), .ZN(n8495) );
  AOI22_X1 U10189 ( .A1(n9102), .A2(keyinput108), .B1(n6146), .B2(keyinput25), 
        .ZN(n8497) );
  OAI221_X1 U10190 ( .B1(n9102), .B2(keyinput108), .C1(n6146), .C2(keyinput25), 
        .A(n8497), .ZN(n8506) );
  AOI22_X1 U10191 ( .A1(n6950), .A2(keyinput83), .B1(keyinput6), .B2(n8847), 
        .ZN(n8498) );
  OAI221_X1 U10192 ( .B1(n6950), .B2(keyinput83), .C1(n8847), .C2(keyinput6), 
        .A(n8498), .ZN(n8505) );
  INV_X1 U10193 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n8500) );
  AOI22_X1 U10194 ( .A1(n9351), .A2(keyinput1), .B1(keyinput104), .B2(n8500), 
        .ZN(n8499) );
  OAI221_X1 U10195 ( .B1(n9351), .B2(keyinput1), .C1(n8500), .C2(keyinput104), 
        .A(n8499), .ZN(n8504) );
  AOI22_X1 U10196 ( .A1(n7895), .A2(keyinput47), .B1(n8502), .B2(keyinput27), 
        .ZN(n8501) );
  OAI221_X1 U10197 ( .B1(n7895), .B2(keyinput47), .C1(n8502), .C2(keyinput27), 
        .A(n8501), .ZN(n8503) );
  OR4_X1 U10198 ( .A1(n8506), .A2(n8505), .A3(n8504), .A4(n8503), .ZN(n8522)
         );
  AOI22_X1 U10199 ( .A1(n8716), .A2(keyinput84), .B1(keyinput55), .B2(n8508), 
        .ZN(n8507) );
  OAI221_X1 U10200 ( .B1(n8716), .B2(keyinput84), .C1(n8508), .C2(keyinput55), 
        .A(n8507), .ZN(n8521) );
  AOI22_X1 U10201 ( .A1(n7159), .A2(keyinput5), .B1(keyinput121), .B2(n7259), 
        .ZN(n8509) );
  OAI221_X1 U10202 ( .B1(n7159), .B2(keyinput5), .C1(n7259), .C2(keyinput121), 
        .A(n8509), .ZN(n8520) );
  INV_X1 U10203 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8511) );
  AOI22_X1 U10204 ( .A1(n9400), .A2(keyinput50), .B1(keyinput8), .B2(n8511), 
        .ZN(n8510) );
  OAI221_X1 U10205 ( .B1(n9400), .B2(keyinput50), .C1(n8511), .C2(keyinput8), 
        .A(n8510), .ZN(n8518) );
  AOI22_X1 U10206 ( .A1(n8701), .A2(keyinput109), .B1(n8513), .B2(keyinput52), 
        .ZN(n8512) );
  OAI221_X1 U10207 ( .B1(n8701), .B2(keyinput109), .C1(n8513), .C2(keyinput52), 
        .A(n8512), .ZN(n8517) );
  INV_X1 U10208 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n8514) );
  XNOR2_X1 U10209 ( .A(keyinput76), .B(n8514), .ZN(n8516) );
  INV_X1 U10210 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n10582) );
  XNOR2_X1 U10211 ( .A(keyinput13), .B(n10582), .ZN(n8515) );
  OR4_X1 U10212 ( .A1(n8518), .A2(n8517), .A3(n8516), .A4(n8515), .ZN(n8519)
         );
  NOR4_X1 U10213 ( .A1(n8522), .A2(n8521), .A3(n8520), .A4(n8519), .ZN(n8535)
         );
  INV_X1 U10214 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10397) );
  XOR2_X1 U10215 ( .A(keyinput15), .B(n10397), .Z(n8534) );
  INV_X1 U10216 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10402) );
  XOR2_X1 U10217 ( .A(keyinput12), .B(n10402), .Z(n8533) );
  AOI22_X1 U10218 ( .A1(n6958), .A2(keyinput56), .B1(keyinput90), .B2(n8958), 
        .ZN(n8523) );
  OAI221_X1 U10219 ( .B1(n6958), .B2(keyinput56), .C1(n8958), .C2(keyinput90), 
        .A(n8523), .ZN(n8531) );
  INV_X1 U10220 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U10221 ( .A1(n10295), .A2(keyinput24), .B1(n10399), .B2(keyinput7), 
        .ZN(n8524) );
  OAI221_X1 U10222 ( .B1(n10295), .B2(keyinput24), .C1(n10399), .C2(keyinput7), 
        .A(n8524), .ZN(n8530) );
  AOI22_X1 U10223 ( .A1(n9098), .A2(keyinput79), .B1(n5664), .B2(keyinput48), 
        .ZN(n8525) );
  OAI221_X1 U10224 ( .B1(n9098), .B2(keyinput79), .C1(n5664), .C2(keyinput48), 
        .A(n8525), .ZN(n8529) );
  INV_X1 U10225 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8527) );
  AOI22_X1 U10226 ( .A1(n10320), .A2(keyinput66), .B1(n8527), .B2(keyinput116), 
        .ZN(n8526) );
  OAI221_X1 U10227 ( .B1(n10320), .B2(keyinput66), .C1(n8527), .C2(keyinput116), .A(n8526), .ZN(n8528) );
  NOR4_X1 U10228 ( .A1(n8531), .A2(n8530), .A3(n8529), .A4(n8528), .ZN(n8532)
         );
  NAND4_X1 U10229 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .ZN(n8649)
         );
  INV_X1 U10230 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U10231 ( .A1(n10403), .A2(keyinput89), .B1(keyinput122), .B2(n9458), 
        .ZN(n8536) );
  OAI221_X1 U10232 ( .B1(n10403), .B2(keyinput89), .C1(n9458), .C2(keyinput122), .A(n8536), .ZN(n8545) );
  INV_X1 U10233 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U10234 ( .A1(n10396), .A2(keyinput42), .B1(keyinput51), .B2(n9252), 
        .ZN(n8537) );
  OAI221_X1 U10235 ( .B1(n10396), .B2(keyinput42), .C1(n9252), .C2(keyinput51), 
        .A(n8537), .ZN(n8544) );
  AOI22_X1 U10236 ( .A1(n8539), .A2(keyinput2), .B1(keyinput33), .B2(n10496), 
        .ZN(n8538) );
  OAI221_X1 U10237 ( .B1(n8539), .B2(keyinput2), .C1(n10496), .C2(keyinput33), 
        .A(n8538), .ZN(n8543) );
  AOI22_X1 U10238 ( .A1(n8541), .A2(keyinput37), .B1(keyinput106), .B2(n8827), 
        .ZN(n8540) );
  OAI221_X1 U10239 ( .B1(n8541), .B2(keyinput37), .C1(n8827), .C2(keyinput106), 
        .A(n8540), .ZN(n8542) );
  NOR4_X1 U10240 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n8571)
         );
  INV_X1 U10241 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10338) );
  AOI22_X1 U10242 ( .A1(n8836), .A2(keyinput57), .B1(keyinput77), .B2(n10338), 
        .ZN(n8546) );
  OAI221_X1 U10243 ( .B1(n8836), .B2(keyinput57), .C1(n10338), .C2(keyinput77), 
        .A(n8546), .ZN(n8553) );
  AOI22_X1 U10244 ( .A1(n8549), .A2(keyinput71), .B1(keyinput80), .B2(n8548), 
        .ZN(n8547) );
  OAI221_X1 U10245 ( .B1(n8549), .B2(keyinput71), .C1(n8548), .C2(keyinput80), 
        .A(n8547), .ZN(n8552) );
  AOI22_X1 U10246 ( .A1(n9106), .A2(keyinput10), .B1(n8724), .B2(keyinput28), 
        .ZN(n8550) );
  OAI221_X1 U10247 ( .B1(n9106), .B2(keyinput10), .C1(n8724), .C2(keyinput28), 
        .A(n8550), .ZN(n8551) );
  NOR3_X1 U10248 ( .A1(n8553), .A2(n8552), .A3(n8551), .ZN(n8570) );
  AOI22_X1 U10249 ( .A1(n8818), .A2(keyinput70), .B1(keyinput17), .B2(n6246), 
        .ZN(n8554) );
  OAI221_X1 U10250 ( .B1(n8818), .B2(keyinput70), .C1(n6246), .C2(keyinput17), 
        .A(n8554), .ZN(n8560) );
  AOI22_X1 U10251 ( .A1(n8556), .A2(keyinput34), .B1(keyinput110), .B2(n9265), 
        .ZN(n8555) );
  OAI221_X1 U10252 ( .B1(n8556), .B2(keyinput34), .C1(n9265), .C2(keyinput110), 
        .A(n8555), .ZN(n8559) );
  AOI22_X1 U10253 ( .A1(n10211), .A2(keyinput102), .B1(keyinput101), .B2(n9124), .ZN(n8557) );
  OAI221_X1 U10254 ( .B1(n10211), .B2(keyinput102), .C1(n9124), .C2(
        keyinput101), .A(n8557), .ZN(n8558) );
  NOR3_X1 U10255 ( .A1(n8560), .A2(n8559), .A3(n8558), .ZN(n8569) );
  INV_X1 U10256 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9243) );
  AOI22_X1 U10257 ( .A1(n8713), .A2(keyinput99), .B1(keyinput124), .B2(n9243), 
        .ZN(n8561) );
  OAI221_X1 U10258 ( .B1(n8713), .B2(keyinput99), .C1(n9243), .C2(keyinput124), 
        .A(n8561), .ZN(n8567) );
  AOI22_X1 U10259 ( .A1(n8563), .A2(keyinput30), .B1(keyinput65), .B2(n9026), 
        .ZN(n8562) );
  OAI221_X1 U10260 ( .B1(n8563), .B2(keyinput30), .C1(n9026), .C2(keyinput65), 
        .A(n8562), .ZN(n8566) );
  XNOR2_X1 U10261 ( .A(n8564), .B(keyinput120), .ZN(n8565) );
  NOR3_X1 U10262 ( .A1(n8567), .A2(n8566), .A3(n8565), .ZN(n8568) );
  NAND4_X1 U10263 ( .A1(n8571), .A2(n8570), .A3(n8569), .A4(n8568), .ZN(n8648)
         );
  XNOR2_X1 U10264 ( .A(n8572), .B(keyinput26), .ZN(n8577) );
  XOR2_X1 U10265 ( .A(P2_REG0_REG_7__SCAN_IN), .B(keyinput61), .Z(n8576) );
  XNOR2_X1 U10266 ( .A(n8573), .B(keyinput36), .ZN(n8575) );
  XNOR2_X1 U10267 ( .A(n9275), .B(keyinput105), .ZN(n8574) );
  NOR4_X1 U10268 ( .A1(n8577), .A2(n8576), .A3(n8575), .A4(n8574), .ZN(n8597)
         );
  XNOR2_X1 U10269 ( .A(n8712), .B(keyinput115), .ZN(n8583) );
  XOR2_X1 U10270 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput112), .Z(n8582) );
  XNOR2_X1 U10271 ( .A(n8578), .B(keyinput118), .ZN(n8581) );
  XNOR2_X1 U10272 ( .A(n8579), .B(keyinput94), .ZN(n8580) );
  NOR4_X1 U10273 ( .A1(n8583), .A2(n8582), .A3(n8581), .A4(n8580), .ZN(n8596)
         );
  XOR2_X1 U10274 ( .A(P2_REG0_REG_9__SCAN_IN), .B(keyinput127), .Z(n8587) );
  XOR2_X1 U10275 ( .A(P2_REG1_REG_2__SCAN_IN), .B(keyinput46), .Z(n8586) );
  XNOR2_X1 U10276 ( .A(n9271), .B(keyinput93), .ZN(n8585) );
  XNOR2_X1 U10277 ( .A(n9221), .B(keyinput21), .ZN(n8584) );
  NOR4_X1 U10278 ( .A1(n8587), .A2(n8586), .A3(n8585), .A4(n8584), .ZN(n8595)
         );
  XOR2_X1 U10279 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput31), .Z(n8593) );
  XNOR2_X1 U10280 ( .A(n8588), .B(keyinput96), .ZN(n8592) );
  INV_X1 U10281 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10583) );
  XNOR2_X1 U10282 ( .A(keyinput91), .B(n10583), .ZN(n8591) );
  INV_X1 U10283 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8589) );
  XNOR2_X1 U10284 ( .A(keyinput72), .B(n8589), .ZN(n8590) );
  NOR4_X1 U10285 ( .A1(n8593), .A2(n8592), .A3(n8591), .A4(n8590), .ZN(n8594)
         );
  NAND4_X1 U10286 ( .A1(n8597), .A2(n8596), .A3(n8595), .A4(n8594), .ZN(n8603)
         );
  INV_X1 U10287 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n8720) );
  AOI22_X1 U10288 ( .A1(n8720), .A2(keyinput16), .B1(n8723), .B2(keyinput0), 
        .ZN(n8598) );
  OAI221_X1 U10289 ( .B1(n8720), .B2(keyinput16), .C1(n8723), .C2(keyinput0), 
        .A(n8598), .ZN(n8602) );
  INV_X1 U10290 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U10291 ( .A1(n10552), .A2(keyinput86), .B1(n9170), .B2(keyinput49), 
        .ZN(n8599) );
  OAI221_X1 U10292 ( .B1(n10552), .B2(keyinput86), .C1(n9170), .C2(keyinput49), 
        .A(n8599), .ZN(n8601) );
  XNOR2_X1 U10293 ( .A(n8698), .B(keyinput3), .ZN(n8600) );
  NOR4_X1 U10294 ( .A1(n8603), .A2(n8602), .A3(n8601), .A4(n8600), .ZN(n8646)
         );
  AOI22_X1 U10295 ( .A1(n8605), .A2(keyinput11), .B1(n8722), .B2(keyinput63), 
        .ZN(n8604) );
  OAI221_X1 U10296 ( .B1(n8605), .B2(keyinput11), .C1(n8722), .C2(keyinput63), 
        .A(n8604), .ZN(n8610) );
  XNOR2_X1 U10297 ( .A(keyinput14), .B(n5485), .ZN(n8609) );
  XNOR2_X1 U10298 ( .A(SI_23_), .B(keyinput69), .ZN(n8607) );
  NAND2_X1 U10299 ( .A1(n5969), .A2(keyinput103), .ZN(n8606) );
  OAI211_X1 U10300 ( .C1(keyinput103), .C2(n5969), .A(n8607), .B(n8606), .ZN(
        n8608) );
  NOR3_X1 U10301 ( .A1(n8610), .A2(n8609), .A3(n8608), .ZN(n8645) );
  XNOR2_X1 U10302 ( .A(SI_7_), .B(keyinput38), .ZN(n8614) );
  XNOR2_X1 U10303 ( .A(SI_9_), .B(keyinput113), .ZN(n8613) );
  XNOR2_X1 U10304 ( .A(SI_1_), .B(keyinput75), .ZN(n8612) );
  XNOR2_X1 U10305 ( .A(SI_3_), .B(keyinput81), .ZN(n8611) );
  NAND4_X1 U10306 ( .A1(n8614), .A2(n8613), .A3(n8612), .A4(n8611), .ZN(n8620)
         );
  XNOR2_X1 U10307 ( .A(SI_0_), .B(keyinput123), .ZN(n8618) );
  XNOR2_X1 U10308 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput117), .ZN(n8617) );
  XNOR2_X1 U10309 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput45), .ZN(n8616) );
  XNOR2_X1 U10310 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput53), .ZN(n8615) );
  NAND4_X1 U10311 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n8619)
         );
  NOR2_X1 U10312 ( .A1(n8620), .A2(n8619), .ZN(n8644) );
  XNOR2_X1 U10313 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput125), .ZN(n8624) );
  XNOR2_X1 U10314 ( .A(P1_IR_REG_22__SCAN_IN), .B(keyinput58), .ZN(n8623) );
  XNOR2_X1 U10315 ( .A(P1_REG1_REG_17__SCAN_IN), .B(keyinput107), .ZN(n8622)
         );
  XNOR2_X1 U10316 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput60), .ZN(n8621) );
  NAND4_X1 U10317 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n8630)
         );
  XNOR2_X1 U10318 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput88), .ZN(n8628) );
  XNOR2_X1 U10319 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput22), .ZN(n8627) );
  XNOR2_X1 U10320 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput82), .ZN(n8626) );
  XNOR2_X1 U10321 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(keyinput111), .ZN(n8625)
         );
  NAND4_X1 U10322 ( .A1(n8628), .A2(n8627), .A3(n8626), .A4(n8625), .ZN(n8629)
         );
  NOR2_X1 U10323 ( .A1(n8630), .A2(n8629), .ZN(n8642) );
  XNOR2_X1 U10324 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput32), .ZN(n8634) );
  XNOR2_X1 U10325 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput40), .ZN(n8633) );
  XNOR2_X1 U10326 ( .A(P1_REG3_REG_2__SCAN_IN), .B(keyinput4), .ZN(n8632) );
  XNOR2_X1 U10327 ( .A(P1_REG3_REG_7__SCAN_IN), .B(keyinput41), .ZN(n8631) );
  NAND4_X1 U10328 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), .ZN(n8640)
         );
  XNOR2_X1 U10329 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput67), .ZN(n8638) );
  XNOR2_X1 U10330 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput64), .ZN(n8637) );
  XNOR2_X1 U10331 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput9), .ZN(n8636) );
  XNOR2_X1 U10332 ( .A(P2_IR_REG_10__SCAN_IN), .B(keyinput97), .ZN(n8635) );
  NAND4_X1 U10333 ( .A1(n8638), .A2(n8637), .A3(n8636), .A4(n8635), .ZN(n8639)
         );
  NOR2_X1 U10334 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  AND2_X1 U10335 ( .A1(n8642), .A2(n8641), .ZN(n8643) );
  NAND4_X1 U10336 ( .A1(n8646), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n8647)
         );
  NOR3_X1 U10337 ( .A1(n8649), .A2(n8648), .A3(n8647), .ZN(n8683) );
  AOI22_X1 U10338 ( .A1(n10241), .A2(keyinput18), .B1(keyinput98), .B2(n8651), 
        .ZN(n8650) );
  OAI221_X1 U10339 ( .B1(n10241), .B2(keyinput18), .C1(n8651), .C2(keyinput98), 
        .A(n8650), .ZN(n8659) );
  INV_X1 U10340 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10401) );
  INV_X1 U10341 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U10342 ( .A1(n10401), .A2(keyinput114), .B1(keyinput78), .B2(n10418), .ZN(n8652) );
  OAI221_X1 U10343 ( .B1(n10401), .B2(keyinput114), .C1(n10418), .C2(
        keyinput78), .A(n8652), .ZN(n8658) );
  INV_X1 U10344 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8732) );
  AOI22_X1 U10345 ( .A1(n8732), .A2(keyinput59), .B1(n8654), .B2(keyinput54), 
        .ZN(n8653) );
  OAI221_X1 U10346 ( .B1(n8732), .B2(keyinput59), .C1(n8654), .C2(keyinput54), 
        .A(n8653), .ZN(n8657) );
  INV_X1 U10347 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U10348 ( .A1(n9113), .A2(keyinput100), .B1(n10398), .B2(keyinput29), 
        .ZN(n8655) );
  OAI221_X1 U10349 ( .B1(n9113), .B2(keyinput100), .C1(n10398), .C2(keyinput29), .A(n8655), .ZN(n8656) );
  NOR4_X1 U10350 ( .A1(n8659), .A2(n8658), .A3(n8657), .A4(n8656), .ZN(n8682)
         );
  AOI22_X1 U10351 ( .A1(n8661), .A2(keyinput119), .B1(n10275), .B2(keyinput126), .ZN(n8660) );
  OAI221_X1 U10352 ( .B1(n8661), .B2(keyinput119), .C1(n10275), .C2(
        keyinput126), .A(n8660), .ZN(n8670) );
  AOI22_X1 U10353 ( .A1(n8738), .A2(keyinput68), .B1(keyinput73), .B2(n8663), 
        .ZN(n8662) );
  OAI221_X1 U10354 ( .B1(n8738), .B2(keyinput68), .C1(n8663), .C2(keyinput73), 
        .A(n8662), .ZN(n8669) );
  INV_X1 U10355 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U10356 ( .A1(n9116), .A2(keyinput92), .B1(n10400), .B2(keyinput19), 
        .ZN(n8664) );
  OAI221_X1 U10357 ( .B1(n9116), .B2(keyinput92), .C1(n10400), .C2(keyinput19), 
        .A(n8664), .ZN(n8668) );
  AOI22_X1 U10358 ( .A1(n8666), .A2(keyinput43), .B1(n5668), .B2(keyinput20), 
        .ZN(n8665) );
  OAI221_X1 U10359 ( .B1(n8666), .B2(keyinput43), .C1(n5668), .C2(keyinput20), 
        .A(n8665), .ZN(n8667) );
  NOR4_X1 U10360 ( .A1(n8670), .A2(n8669), .A3(n8668), .A4(n8667), .ZN(n8681)
         );
  INV_X1 U10361 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8672) );
  AOI22_X1 U10362 ( .A1(n10189), .A2(keyinput95), .B1(keyinput44), .B2(n8672), 
        .ZN(n8671) );
  OAI221_X1 U10363 ( .B1(n10189), .B2(keyinput95), .C1(n8672), .C2(keyinput44), 
        .A(n8671), .ZN(n8679) );
  INV_X1 U10364 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10404) );
  AOI22_X1 U10365 ( .A1(n10404), .A2(keyinput35), .B1(keyinput39), .B2(n5990), 
        .ZN(n8673) );
  OAI221_X1 U10366 ( .B1(n10404), .B2(keyinput35), .C1(n5990), .C2(keyinput39), 
        .A(n8673), .ZN(n8678) );
  AOI22_X1 U10367 ( .A1(n9203), .A2(keyinput62), .B1(n7926), .B2(keyinput85), 
        .ZN(n8674) );
  OAI221_X1 U10368 ( .B1(n9203), .B2(keyinput62), .C1(n7926), .C2(keyinput85), 
        .A(n8674), .ZN(n8677) );
  AOI22_X1 U10369 ( .A1(n8717), .A2(keyinput23), .B1(n5888), .B2(keyinput87), 
        .ZN(n8675) );
  OAI221_X1 U10370 ( .B1(n8717), .B2(keyinput23), .C1(n5888), .C2(keyinput87), 
        .A(n8675), .ZN(n8676) );
  NOR4_X1 U10371 ( .A1(n8679), .A2(n8678), .A3(n8677), .A4(n8676), .ZN(n8680)
         );
  NAND4_X1 U10372 ( .A1(n8683), .A2(n8682), .A3(n8681), .A4(n8680), .ZN(n8752)
         );
  NOR4_X1 U10373 ( .A1(P2_REG1_REG_31__SCAN_IN), .A2(SI_31_), .A3(n9102), .A4(
        n6146), .ZN(n8684) );
  NAND3_X1 U10374 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(P2_REG0_REG_12__SCAN_IN), .A3(n8684), .ZN(n8697) );
  INV_X1 U10375 ( .A(SI_0_), .ZN(n8685) );
  NAND4_X1 U10376 ( .A1(n10320), .A2(n8686), .A3(n8685), .A4(
        P2_REG2_REG_30__SCAN_IN), .ZN(n8687) );
  NOR3_X1 U10377 ( .A1(n8687), .A2(P2_WR_REG_SCAN_IN), .A3(n8836), .ZN(n8695)
         );
  NAND4_X1 U10378 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(P2_REG0_REG_0__SCAN_IN), 
        .A3(P1_REG2_REG_30__SCAN_IN), .A4(n10552), .ZN(n8693) );
  NAND4_X1 U10379 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_DATAO_REG_2__SCAN_IN), 
        .A3(P1_REG2_REG_7__SCAN_IN), .A4(P2_REG1_REG_2__SCAN_IN), .ZN(n8692)
         );
  NAND4_X1 U10380 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P2_REG2_REG_3__SCAN_IN), 
        .A3(n8818), .A4(n6246), .ZN(n8688) );
  NOR2_X1 U10381 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(n8688), .ZN(n8690) );
  NAND4_X1 U10382 ( .A1(n8690), .A2(P2_REG0_REG_7__SCAN_IN), .A3(n8689), .A4(
        P1_ADDR_REG_10__SCAN_IN), .ZN(n8691) );
  NOR3_X1 U10383 ( .A1(n8693), .A2(n8692), .A3(n8691), .ZN(n8694) );
  NAND4_X1 U10384 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n8695), .A3(n8694), .A4(
        n9287), .ZN(n8696) );
  NOR4_X1 U10385 ( .A1(SI_7_), .A2(P1_REG0_REG_11__SCAN_IN), .A3(n8697), .A4(
        n8696), .ZN(n8748) );
  NOR4_X1 U10386 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_REG3_REG_5__SCAN_IN), 
        .A3(P2_D_REG_17__SCAN_IN), .A4(n9221), .ZN(n8747) );
  INV_X1 U10387 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8710) );
  NAND4_X1 U10388 ( .A1(SI_3_), .A2(SI_23_), .A3(P2_ADDR_REG_14__SCAN_IN), 
        .A4(n8698), .ZN(n8700) );
  NOR2_X1 U10389 ( .A1(n8700), .A2(n8699), .ZN(n8708) );
  NOR4_X1 U10390 ( .A1(SI_1_), .A2(P2_REG2_REG_27__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .A4(P1_ADDR_REG_13__SCAN_IN), .ZN(n8703) );
  NOR4_X1 U10391 ( .A1(SI_19_), .A2(P1_IR_REG_30__SCAN_IN), .A3(n8701), .A4(
        n9243), .ZN(n8702) );
  AND2_X1 U10392 ( .A1(n8703), .A2(n8702), .ZN(n8707) );
  NOR4_X1 U10393 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(P1_REG2_REG_25__SCAN_IN), 
        .A3(P1_REG1_REG_17__SCAN_IN), .A4(n9203), .ZN(n8706) );
  INV_X1 U10394 ( .A(n8704), .ZN(n8705) );
  NAND4_X1 U10395 ( .A1(n8708), .A2(n8707), .A3(n8706), .A4(n8705), .ZN(n8709)
         );
  NOR4_X1 U10396 ( .A1(n9400), .A2(n8710), .A3(SI_6_), .A4(n8709), .ZN(n8711)
         );
  NAND3_X1 U10397 ( .A1(n8711), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P1_ADDR_REG_2__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U10398 ( .A1(n8713), .A2(n8712), .ZN(n8714) );
  NOR4_X1 U10399 ( .A1(n8715), .A2(P2_REG0_REG_13__SCAN_IN), .A3(n9124), .A4(
        n8714), .ZN(n8721) );
  NOR4_X1 U10400 ( .A1(n8717), .A2(n8716), .A3(n10211), .A4(
        P1_REG2_REG_15__SCAN_IN), .ZN(n8719) );
  NOR4_X1 U10401 ( .A1(n5325), .A2(P2_IR_REG_22__SCAN_IN), .A3(
        P2_IR_REG_2__SCAN_IN), .A4(P2_REG3_REG_28__SCAN_IN), .ZN(n8718) );
  NAND4_X1 U10402 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n8736)
         );
  NOR2_X1 U10403 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8730) );
  NAND4_X1 U10404 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(P1_REG2_REG_26__SCAN_IN), .A3(P2_IR_REG_25__SCAN_IN), .A4(n8722), .ZN(n8728) );
  NAND4_X1 U10405 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), 
        .A3(P2_IR_REG_16__SCAN_IN), .A4(P2_IR_REG_24__SCAN_IN), .ZN(n8727) );
  NAND4_X1 U10406 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_REG1_REG_29__SCAN_IN), 
        .A3(P1_REG3_REG_7__SCAN_IN), .A4(P1_REG2_REG_23__SCAN_IN), .ZN(n8726)
         );
  NAND4_X1 U10407 ( .A1(n8724), .A2(n9351), .A3(n8723), .A4(n9106), .ZN(n8725)
         );
  NOR4_X1 U10408 ( .A1(n8728), .A2(n8727), .A3(n8726), .A4(n8725), .ZN(n8729)
         );
  NAND4_X1 U10409 ( .A1(n8731), .A2(n8730), .A3(n8729), .A4(n9252), .ZN(n8735)
         );
  NOR4_X1 U10410 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(P1_REG1_REG_23__SCAN_IN), .A4(n8732), .ZN(n8733) );
  NAND3_X1 U10411 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P2_REG1_REG_24__SCAN_IN), 
        .A3(n8733), .ZN(n8734) );
  NOR3_X1 U10412 ( .A1(n8736), .A2(n8735), .A3(n8734), .ZN(n8746) );
  NAND4_X1 U10413 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P1_REG1_REG_5__SCAN_IN), 
        .A3(P2_REG2_REG_11__SCAN_IN), .A4(n8958), .ZN(n8737) );
  NOR3_X1 U10414 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(P2_REG2_REG_25__SCAN_IN), 
        .A3(n8737), .ZN(n8744) );
  NAND4_X1 U10415 ( .A1(P2_REG0_REG_11__SCAN_IN), .A2(P1_DATAO_REG_31__SCAN_IN), .A3(n10295), .A4(n8738), .ZN(n8742) );
  NAND4_X1 U10416 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .A3(
        P1_REG3_REG_20__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n8741) );
  NAND4_X1 U10417 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P2_REG1_REG_29__SCAN_IN), 
        .A3(n10418), .A4(n10241), .ZN(n8740) );
  NAND4_X1 U10418 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10275), .A3(n5668), .A4(
        n9116), .ZN(n8739) );
  NOR4_X1 U10419 ( .A1(n8742), .A2(n8741), .A3(n8740), .A4(n8739), .ZN(n8743)
         );
  AND4_X1 U10420 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_REG1_REG_1__SCAN_IN), 
        .A3(n8744), .A4(n8743), .ZN(n8745) );
  NAND4_X1 U10421 ( .A1(n8748), .A2(n8747), .A3(n8746), .A4(n8745), .ZN(n8749)
         );
  NAND2_X1 U10422 ( .A1(n8749), .A2(keyinput74), .ZN(n8750) );
  MUX2_X1 U10423 ( .A(keyinput74), .B(n8750), .S(P2_REG2_REG_1__SCAN_IN), .Z(
        n8751) );
  OR2_X1 U10424 ( .A1(n8752), .A2(n8751), .ZN(n8753) );
  XNOR2_X1 U10425 ( .A(n8786), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8800) );
  INV_X1 U10426 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8756) );
  INV_X1 U10427 ( .A(n8754), .ZN(n8755) );
  NAND2_X1 U10428 ( .A1(n8799), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8782) );
  NAND2_X1 U10429 ( .A1(n8786), .A2(n8758), .ZN(n8759) );
  NAND2_X1 U10430 ( .A1(n8782), .A2(n8759), .ZN(n8760) );
  AND3_X1 U10431 ( .A1(n8762), .A2(n8761), .A3(n8760), .ZN(n8764) );
  INV_X1 U10432 ( .A(n8765), .ZN(n8766) );
  MUX2_X1 U10433 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8770), .Z(n8771) );
  NAND2_X1 U10434 ( .A1(n8772), .A2(n8771), .ZN(n8785) );
  NAND2_X1 U10435 ( .A1(n8773), .A2(n8785), .ZN(n8775) );
  OAI21_X1 U10436 ( .B1(n8775), .B2(n8774), .A(n8795), .ZN(n8779) );
  INV_X1 U10437 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8777) );
  XNOR2_X1 U10438 ( .A(n8794), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8789) );
  XNOR2_X1 U10439 ( .A(n8784), .B(n8789), .ZN(n8805) );
  OAI21_X1 U10440 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8791) );
  XNOR2_X1 U10441 ( .A(n8794), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8802) );
  MUX2_X1 U10442 ( .A(n8802), .B(n8789), .S(n8788), .Z(n8790) );
  XNOR2_X1 U10443 ( .A(n8791), .B(n8790), .ZN(n8798) );
  NAND2_X1 U10444 ( .A1(n10513), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8792) );
  OAI211_X1 U10445 ( .C1(n8795), .C2(n8794), .A(n8793), .B(n8792), .ZN(n8796)
         );
  AOI21_X1 U10446 ( .B1(n8798), .B2(n8797), .A(n8796), .ZN(n8804) );
  OAI211_X1 U10447 ( .C1(n8805), .C2(n10503), .A(n8804), .B(n8803), .ZN(
        P2_U3201) );
  NAND2_X1 U10448 ( .A1(n9177), .A2(n9029), .ZN(n8810) );
  INV_X1 U10449 ( .A(n8806), .ZN(n8807) );
  NOR2_X1 U10450 ( .A1(n8808), .A2(n8807), .ZN(n9178) );
  AOI21_X1 U10451 ( .B1(n9178), .B2(n9091), .A(n8809), .ZN(n8813) );
  OAI211_X1 U10452 ( .C1(n9091), .C2(n8811), .A(n8810), .B(n8813), .ZN(
        P2_U3202) );
  NAND2_X1 U10453 ( .A1(n8981), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8812) );
  OAI211_X1 U10454 ( .C1(n9183), .C2(n9090), .A(n8813), .B(n8812), .ZN(
        P2_U3203) );
  XNOR2_X1 U10455 ( .A(n8814), .B(n8815), .ZN(n9189) );
  MUX2_X1 U10456 ( .A(n8818), .B(n9184), .S(n9091), .Z(n8821) );
  AOI22_X1 U10457 ( .A1(n9186), .A2(n9029), .B1(n10518), .B2(n8819), .ZN(n8820) );
  XNOR2_X1 U10458 ( .A(n8822), .B(n8823), .ZN(n9195) );
  MUX2_X1 U10459 ( .A(n8827), .B(n9190), .S(n9091), .Z(n8830) );
  AOI22_X1 U10460 ( .A1(n9192), .A2(n9029), .B1(n10518), .B2(n8828), .ZN(n8829) );
  OAI211_X1 U10461 ( .C1(n9195), .C2(n9086), .A(n8830), .B(n8829), .ZN(
        P2_U3206) );
  XNOR2_X1 U10462 ( .A(n8831), .B(n8832), .ZN(n9201) );
  XNOR2_X1 U10463 ( .A(n8833), .B(n6507), .ZN(n8835) );
  AOI222_X1 U10464 ( .A1(n9061), .A2(n8835), .B1(n8858), .B2(n9064), .C1(n8834), .C2(n9065), .ZN(n9196) );
  MUX2_X1 U10465 ( .A(n8836), .B(n4425), .S(n9091), .Z(n8839) );
  AOI22_X1 U10466 ( .A1(n9198), .A2(n9029), .B1(n10518), .B2(n8837), .ZN(n8838) );
  OAI211_X1 U10467 ( .C1(n9201), .C2(n9086), .A(n8839), .B(n8838), .ZN(
        P2_U3207) );
  XOR2_X1 U10468 ( .A(n8846), .B(n8840), .Z(n8842) );
  AOI222_X1 U10469 ( .A1(n9061), .A2(n8842), .B1(n8871), .B2(n9064), .C1(n8841), .C2(n9065), .ZN(n9202) );
  AOI22_X1 U10470 ( .A1(n9204), .A2(n8980), .B1(n10518), .B2(n8843), .ZN(n8844) );
  AOI21_X1 U10471 ( .B1(n9202), .B2(n8844), .A(n8981), .ZN(n8849) );
  XNOR2_X1 U10472 ( .A(n8845), .B(n8846), .ZN(n9207) );
  OAI22_X1 U10473 ( .A1(n9207), .A2(n9086), .B1(n8847), .B2(n9091), .ZN(n8848)
         );
  OR2_X1 U10474 ( .A1(n8849), .A2(n8848), .ZN(P2_U3208) );
  NAND2_X1 U10475 ( .A1(n8851), .A2(n8850), .ZN(n8884) );
  NAND2_X1 U10476 ( .A1(n8884), .A2(n8883), .ZN(n9122) );
  NAND2_X1 U10477 ( .A1(n9122), .A2(n8852), .ZN(n8864) );
  OAI21_X1 U10478 ( .B1(n8864), .B2(n8854), .A(n8853), .ZN(n8855) );
  XOR2_X1 U10479 ( .A(n8856), .B(n8855), .Z(n9213) );
  XNOR2_X1 U10480 ( .A(n4475), .B(n8856), .ZN(n8859) );
  AOI22_X1 U10481 ( .A1(n9210), .A2(n8980), .B1(n10518), .B2(n8860), .ZN(n8861) );
  AOI21_X1 U10482 ( .B1(n8981), .B2(P2_REG2_REG_24__SCAN_IN), .A(n8862), .ZN(
        n8863) );
  OAI21_X1 U10483 ( .B1(n9086), .B2(n9213), .A(n8863), .ZN(P2_U3209) );
  XOR2_X1 U10484 ( .A(n8869), .B(n8864), .Z(n9219) );
  INV_X1 U10485 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8873) );
  AOI21_X1 U10486 ( .B1(n8866), .B2(n8865), .A(n8883), .ZN(n8878) );
  INV_X1 U10487 ( .A(n8878), .ZN(n8868) );
  NAND2_X1 U10488 ( .A1(n8868), .A2(n8867), .ZN(n8870) );
  XNOR2_X1 U10489 ( .A(n8870), .B(n8869), .ZN(n8872) );
  AOI222_X1 U10490 ( .A1(n9061), .A2(n8872), .B1(n8871), .B2(n9065), .C1(n8896), .C2(n9064), .ZN(n9214) );
  MUX2_X1 U10491 ( .A(n8873), .B(n9214), .S(n9091), .Z(n8876) );
  AOI22_X1 U10492 ( .A1(n9216), .A2(n9029), .B1(n10518), .B2(n8874), .ZN(n8875) );
  OAI211_X1 U10493 ( .C1(n9219), .C2(n9086), .A(n8876), .B(n8875), .ZN(
        P2_U3210) );
  NOR2_X1 U10494 ( .A1(n5156), .A2(n8877), .ZN(n8879) );
  AND2_X1 U10495 ( .A1(n8906), .A2(n8905), .ZN(n8903) );
  OAI21_X1 U10496 ( .B1(n8903), .B2(n8893), .A(n8892), .ZN(n8895) );
  AOI21_X1 U10497 ( .B1(n8879), .B2(n8895), .A(n8878), .ZN(n8880) );
  OAI222_X1 U10498 ( .A1(n9010), .A2(n8882), .B1(n9008), .B2(n8881), .C1(n9007), .C2(n8880), .ZN(n9121) );
  NOR2_X1 U10499 ( .A1(n8884), .A2(n8883), .ZN(n9120) );
  INV_X1 U10500 ( .A(n9122), .ZN(n8885) );
  NOR3_X1 U10501 ( .A1(n9120), .A2(n8885), .A3(n9086), .ZN(n8889) );
  AOI22_X1 U10502 ( .A1(n8886), .A2(n10518), .B1(n8981), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8887) );
  OAI21_X1 U10503 ( .B1(n9223), .B2(n9090), .A(n8887), .ZN(n8888) );
  AOI211_X1 U10504 ( .C1(n9121), .C2(n9091), .A(n8889), .B(n8888), .ZN(n8890)
         );
  INV_X1 U10505 ( .A(n8890), .ZN(P2_U3211) );
  XNOR2_X1 U10506 ( .A(n8891), .B(n8892), .ZN(n9229) );
  OR3_X1 U10507 ( .A1(n8903), .A2(n8893), .A3(n8892), .ZN(n8894) );
  NAND2_X1 U10508 ( .A1(n8895), .A2(n8894), .ZN(n8897) );
  AOI222_X1 U10509 ( .A1(n9061), .A2(n8897), .B1(n8896), .B2(n9065), .C1(n8918), .C2(n9064), .ZN(n9224) );
  MUX2_X1 U10510 ( .A(n8898), .B(n9224), .S(n9091), .Z(n8901) );
  AOI22_X1 U10511 ( .A1(n9226), .A2(n9029), .B1(n10518), .B2(n8899), .ZN(n8900) );
  OAI211_X1 U10512 ( .C1(n9229), .C2(n9086), .A(n8901), .B(n8900), .ZN(
        P2_U3212) );
  XNOR2_X1 U10513 ( .A(n8902), .B(n8905), .ZN(n9235) );
  INV_X1 U10514 ( .A(n8903), .ZN(n8904) );
  OAI21_X1 U10515 ( .B1(n8906), .B2(n8905), .A(n8904), .ZN(n8909) );
  AOI222_X1 U10516 ( .A1(n9061), .A2(n8909), .B1(n8908), .B2(n9065), .C1(n8907), .C2(n9064), .ZN(n9230) );
  MUX2_X1 U10517 ( .A(n8910), .B(n9230), .S(n9091), .Z(n8913) );
  AOI22_X1 U10518 ( .A1(n9232), .A2(n9029), .B1(n10518), .B2(n8911), .ZN(n8912) );
  OAI211_X1 U10519 ( .C1(n9235), .C2(n9086), .A(n8913), .B(n8912), .ZN(
        P2_U3213) );
  XNOR2_X1 U10520 ( .A(n8914), .B(n8915), .ZN(n9241) );
  INV_X1 U10521 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U10522 ( .A(n8917), .B(n8916), .ZN(n8919) );
  AOI222_X1 U10523 ( .A1(n9061), .A2(n8919), .B1(n8918), .B2(n9065), .C1(n8943), .C2(n9064), .ZN(n9236) );
  MUX2_X1 U10524 ( .A(n8920), .B(n9236), .S(n9091), .Z(n8923) );
  AOI22_X1 U10525 ( .A1(n9238), .A2(n9029), .B1(n10518), .B2(n8921), .ZN(n8922) );
  OAI211_X1 U10526 ( .C1(n9241), .C2(n9086), .A(n8923), .B(n8922), .ZN(
        P2_U3214) );
  XOR2_X1 U10527 ( .A(n8924), .B(n8930), .Z(n8925) );
  OAI222_X1 U10528 ( .A1(n9008), .A2(n8926), .B1(n9010), .B2(n8954), .C1(n8925), .C2(n9007), .ZN(n9135) );
  INV_X1 U10529 ( .A(n9135), .ZN(n8935) );
  NAND2_X1 U10530 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  XOR2_X1 U10531 ( .A(n8930), .B(n8929), .Z(n9136) );
  AOI22_X1 U10532 ( .A1(n8981), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n10518), 
        .B2(n8931), .ZN(n8932) );
  OAI21_X1 U10533 ( .B1(n9245), .B2(n9090), .A(n8932), .ZN(n8933) );
  AOI21_X1 U10534 ( .B1(n9136), .B2(n9080), .A(n8933), .ZN(n8934) );
  OAI21_X1 U10535 ( .B1(n8935), .B2(n8981), .A(n8934), .ZN(P2_U3215) );
  XNOR2_X1 U10536 ( .A(n8936), .B(n8940), .ZN(n9248) );
  INV_X1 U10537 ( .A(n8938), .ZN(n8939) );
  NAND2_X1 U10538 ( .A1(n8956), .A2(n8939), .ZN(n8941) );
  XNOR2_X1 U10539 ( .A(n8941), .B(n8940), .ZN(n8942) );
  NAND2_X1 U10540 ( .A1(n8942), .A2(n9061), .ZN(n8945) );
  AOI22_X1 U10541 ( .A1(n8943), .A2(n9065), .B1(n9064), .B2(n8964), .ZN(n8944)
         );
  NAND2_X1 U10542 ( .A1(n8945), .A2(n8944), .ZN(n9246) );
  MUX2_X1 U10543 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n9246), .S(n9091), .Z(n8946) );
  INV_X1 U10544 ( .A(n8946), .ZN(n8950) );
  AOI22_X1 U10545 ( .A1(n8948), .A2(n9029), .B1(n10518), .B2(n8947), .ZN(n8949) );
  OAI211_X1 U10546 ( .C1(n9248), .C2(n9086), .A(n8950), .B(n8949), .ZN(
        P2_U3216) );
  XNOR2_X1 U10547 ( .A(n8951), .B(n8952), .ZN(n9256) );
  AOI21_X1 U10548 ( .B1(n8937), .B2(n8952), .A(n9007), .ZN(n8957) );
  OAI22_X1 U10549 ( .A1(n8954), .A2(n9008), .B1(n8953), .B2(n9010), .ZN(n8955)
         );
  AOI21_X1 U10550 ( .B1(n8957), .B2(n8956), .A(n8955), .ZN(n9251) );
  MUX2_X1 U10551 ( .A(n9251), .B(n8958), .S(n8981), .Z(n8961) );
  AOI22_X1 U10552 ( .A1(n9253), .A2(n9029), .B1(n10518), .B2(n8959), .ZN(n8960) );
  OAI211_X1 U10553 ( .C1(n9256), .C2(n9086), .A(n8961), .B(n8960), .ZN(
        P2_U3217) );
  XNOR2_X1 U10554 ( .A(n8962), .B(n8963), .ZN(n8965) );
  AOI222_X1 U10555 ( .A1(n9061), .A2(n8965), .B1(n8964), .B2(n9065), .C1(n8991), .C2(n9064), .ZN(n9147) );
  XNOR2_X1 U10556 ( .A(n8966), .B(n8967), .ZN(n9145) );
  NAND2_X1 U10557 ( .A1(n9144), .A2(n9029), .ZN(n8970) );
  AOI22_X1 U10558 ( .A1(n8981), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10518), 
        .B2(n8968), .ZN(n8969) );
  NAND2_X1 U10559 ( .A1(n8970), .A2(n8969), .ZN(n8971) );
  AOI21_X1 U10560 ( .B1(n9145), .B2(n9080), .A(n8971), .ZN(n8972) );
  OAI21_X1 U10561 ( .B1(n9147), .B2(n8981), .A(n8972), .ZN(P2_U3218) );
  XNOR2_X1 U10562 ( .A(n8973), .B(n8984), .ZN(n8974) );
  NAND2_X1 U10563 ( .A1(n8974), .A2(n9061), .ZN(n8978) );
  AOI22_X1 U10564 ( .A1(n9065), .A2(n8976), .B1(n9064), .B2(n8975), .ZN(n8977)
         );
  AOI22_X1 U10565 ( .A1(n9260), .A2(n8980), .B1(n10518), .B2(n8979), .ZN(n8982) );
  AOI21_X1 U10566 ( .B1(n9258), .B2(n8982), .A(n8981), .ZN(n8987) );
  XNOR2_X1 U10567 ( .A(n8983), .B(n8984), .ZN(n9263) );
  OAI22_X1 U10568 ( .A1(n9263), .A2(n9086), .B1(n8985), .B2(n9091), .ZN(n8986)
         );
  OR2_X1 U10569 ( .A1(n8987), .A2(n8986), .ZN(P2_U3219) );
  XNOR2_X1 U10570 ( .A(n8988), .B(n4539), .ZN(n9269) );
  XNOR2_X1 U10571 ( .A(n8989), .B(n4539), .ZN(n8990) );
  NAND2_X1 U10572 ( .A1(n8990), .A2(n9061), .ZN(n8993) );
  AOI22_X1 U10573 ( .A1(n9065), .A2(n8991), .B1(n9064), .B2(n9024), .ZN(n8992)
         );
  INV_X1 U10574 ( .A(n9264), .ZN(n8998) );
  INV_X1 U10575 ( .A(n9266), .ZN(n8996) );
  OAI22_X1 U10576 ( .A1(n8996), .A2(n8995), .B1(n8994), .B2(n9087), .ZN(n8997)
         );
  OAI21_X1 U10577 ( .B1(n8998), .B2(n8997), .A(n9091), .ZN(n9000) );
  NAND2_X1 U10578 ( .A1(n8981), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8999) );
  OAI211_X1 U10579 ( .C1(n9269), .C2(n9086), .A(n9000), .B(n8999), .ZN(
        P2_U3220) );
  NAND2_X1 U10580 ( .A1(n9001), .A2(n9005), .ZN(n9002) );
  NAND2_X1 U10581 ( .A1(n9003), .A2(n9002), .ZN(n9273) );
  XOR2_X1 U10582 ( .A(n9005), .B(n9004), .Z(n9006) );
  OAI222_X1 U10583 ( .A1(n9010), .A2(n9009), .B1(n9008), .B2(n6722), .C1(n9007), .C2(n9006), .ZN(n9154) );
  NAND2_X1 U10584 ( .A1(n9154), .A2(n9091), .ZN(n9015) );
  NAND2_X1 U10585 ( .A1(n8981), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n9011) );
  OAI21_X1 U10586 ( .B1(n9012), .B2(n9087), .A(n9011), .ZN(n9013) );
  AOI21_X1 U10587 ( .B1(n9155), .B2(n9029), .A(n9013), .ZN(n9014) );
  OAI211_X1 U10588 ( .C1(n9273), .C2(n9086), .A(n9015), .B(n9014), .ZN(
        P2_U3221) );
  AOI21_X1 U10589 ( .B1(n7659), .B2(n9017), .A(n9016), .ZN(n9019) );
  NOR2_X1 U10590 ( .A1(n9019), .A2(n4842), .ZN(n9021) );
  XNOR2_X1 U10591 ( .A(n9021), .B(n9020), .ZN(n9281) );
  XNOR2_X1 U10592 ( .A(n9023), .B(n9022), .ZN(n9025) );
  AOI222_X1 U10593 ( .A1(n9061), .A2(n9025), .B1(n9024), .B2(n9065), .C1(n9066), .C2(n9064), .ZN(n9274) );
  MUX2_X1 U10594 ( .A(n9026), .B(n9274), .S(n9091), .Z(n9031) );
  INV_X1 U10595 ( .A(n9027), .ZN(n9028) );
  AOI22_X1 U10596 ( .A1(n9276), .A2(n9029), .B1(n10518), .B2(n9028), .ZN(n9030) );
  OAI211_X1 U10597 ( .C1(n9281), .C2(n9086), .A(n9031), .B(n9030), .ZN(
        P2_U3222) );
  NAND2_X1 U10598 ( .A1(n9081), .A2(n9032), .ZN(n9054) );
  INV_X1 U10599 ( .A(n9033), .ZN(n9058) );
  NAND2_X1 U10600 ( .A1(n9054), .A2(n9058), .ZN(n9056) );
  NAND2_X1 U10601 ( .A1(n9056), .A2(n9034), .ZN(n9035) );
  XNOR2_X1 U10602 ( .A(n9035), .B(n9042), .ZN(n9050) );
  INV_X1 U10603 ( .A(n9050), .ZN(n9164) );
  OAI22_X1 U10604 ( .A1(n9285), .A2(n9090), .B1(n9036), .B2(n9087), .ZN(n9052)
         );
  OR2_X1 U10605 ( .A1(n9037), .A2(n9058), .ZN(n9060) );
  INV_X1 U10606 ( .A(n9038), .ZN(n9041) );
  NAND2_X1 U10607 ( .A1(n9060), .A2(n9041), .ZN(n9040) );
  NAND2_X1 U10608 ( .A1(n9040), .A2(n9039), .ZN(n9044) );
  NAND3_X1 U10609 ( .A1(n9060), .A2(n9042), .A3(n9041), .ZN(n9043) );
  NAND2_X1 U10610 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  NAND2_X1 U10611 ( .A1(n9045), .A2(n9061), .ZN(n9049) );
  AOI22_X1 U10612 ( .A1(n9047), .A2(n9064), .B1(n9065), .B2(n9046), .ZN(n9048)
         );
  OAI211_X1 U10613 ( .C1(n9050), .C2(n9069), .A(n9049), .B(n9048), .ZN(n9163)
         );
  MUX2_X1 U10614 ( .A(n9163), .B(P2_REG2_REG_10__SCAN_IN), .S(n8981), .Z(n9051) );
  AOI211_X1 U10615 ( .C1(n10520), .C2(n9164), .A(n9052), .B(n9051), .ZN(n9053)
         );
  INV_X1 U10616 ( .A(n9053), .ZN(P2_U3223) );
  OR2_X1 U10617 ( .A1(n9054), .A2(n9058), .ZN(n9055) );
  NAND2_X1 U10618 ( .A1(n9056), .A2(n9055), .ZN(n9070) );
  INV_X1 U10619 ( .A(n9070), .ZN(n9168) );
  OAI22_X1 U10620 ( .A1(n9090), .A2(n9290), .B1(n9057), .B2(n9087), .ZN(n9072)
         );
  NAND2_X1 U10621 ( .A1(n9037), .A2(n9058), .ZN(n9059) );
  NAND2_X1 U10622 ( .A1(n9060), .A2(n9059), .ZN(n9062) );
  NAND2_X1 U10623 ( .A1(n9062), .A2(n9061), .ZN(n9068) );
  AOI22_X1 U10624 ( .A1(n9066), .A2(n9065), .B1(n9064), .B2(n9063), .ZN(n9067)
         );
  OAI211_X1 U10625 ( .C1(n9070), .C2(n9069), .A(n9068), .B(n9067), .ZN(n9167)
         );
  MUX2_X1 U10626 ( .A(n9167), .B(P2_REG2_REG_9__SCAN_IN), .S(n8981), .Z(n9071)
         );
  AOI211_X1 U10627 ( .C1(n9168), .C2(n10520), .A(n9072), .B(n9071), .ZN(n9073)
         );
  INV_X1 U10628 ( .A(n9073), .ZN(P2_U3224) );
  MUX2_X1 U10629 ( .A(n9075), .B(n9074), .S(n9091), .Z(n9085) );
  INV_X1 U10630 ( .A(n9076), .ZN(n9078) );
  OAI22_X1 U10631 ( .A1(n9090), .A2(n9078), .B1(n9077), .B2(n9087), .ZN(n9079)
         );
  INV_X1 U10632 ( .A(n9079), .ZN(n9084) );
  NAND3_X1 U10633 ( .A1(n9082), .A2(n9081), .A3(n9080), .ZN(n9083) );
  NAND3_X1 U10634 ( .A1(n9085), .A2(n9084), .A3(n9083), .ZN(P2_U3225) );
  OAI22_X1 U10635 ( .A1(n9090), .A2(n9089), .B1(n9088), .B2(n9087), .ZN(n9094)
         );
  MUX2_X1 U10636 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n9092), .S(n9091), .Z(n9093)
         );
  AOI211_X1 U10637 ( .C1(n9095), .C2(n9080), .A(n9094), .B(n9093), .ZN(n9096)
         );
  INV_X1 U10638 ( .A(n9096), .ZN(P2_U3226) );
  NAND2_X1 U10639 ( .A1(n9177), .A2(n9159), .ZN(n9097) );
  NAND2_X1 U10640 ( .A1(n9178), .A2(n10557), .ZN(n9100) );
  OAI211_X1 U10641 ( .C1(n10557), .C2(n9098), .A(n9097), .B(n9100), .ZN(
        P2_U3490) );
  NAND2_X1 U10642 ( .A1(n9099), .A2(n9159), .ZN(n9101) );
  OAI211_X1 U10643 ( .C1(n10557), .C2(n9102), .A(n9101), .B(n9100), .ZN(
        P2_U3489) );
  INV_X1 U10644 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U10645 ( .A1(n9186), .A2(n9159), .ZN(n9104) );
  OAI211_X1 U10646 ( .C1(n9189), .C2(n9162), .A(n9105), .B(n9104), .ZN(
        P2_U3487) );
  INV_X1 U10647 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9107) );
  MUX2_X1 U10648 ( .A(n9107), .B(n4425), .S(n10557), .Z(n9109) );
  NAND2_X1 U10649 ( .A1(n9198), .A2(n9159), .ZN(n9108) );
  OAI211_X1 U10650 ( .C1(n9162), .C2(n9201), .A(n9109), .B(n9108), .ZN(
        P2_U3485) );
  INV_X1 U10651 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9110) );
  MUX2_X1 U10652 ( .A(n9110), .B(n9202), .S(n10557), .Z(n9112) );
  NAND2_X1 U10653 ( .A1(n9204), .A2(n9159), .ZN(n9111) );
  OAI211_X1 U10654 ( .C1(n9207), .C2(n9162), .A(n9112), .B(n9111), .ZN(
        P2_U3484) );
  MUX2_X1 U10655 ( .A(n9113), .B(n9208), .S(n10557), .Z(n9115) );
  NAND2_X1 U10656 ( .A1(n9210), .A2(n9159), .ZN(n9114) );
  OAI211_X1 U10657 ( .C1(n9162), .C2(n9213), .A(n9115), .B(n9114), .ZN(
        P2_U3483) );
  MUX2_X1 U10658 ( .A(n9116), .B(n9214), .S(n10557), .Z(n9118) );
  NAND2_X1 U10659 ( .A1(n9216), .A2(n9159), .ZN(n9117) );
  OAI211_X1 U10660 ( .C1(n9219), .C2(n9162), .A(n9118), .B(n9117), .ZN(
        P2_U3482) );
  NOR2_X1 U10661 ( .A1(n9120), .A2(n9119), .ZN(n9123) );
  AOI21_X1 U10662 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9220) );
  MUX2_X1 U10663 ( .A(n9124), .B(n9220), .S(n10557), .Z(n9125) );
  OAI21_X1 U10664 ( .B1(n9223), .B2(n9172), .A(n9125), .ZN(P2_U3481) );
  INV_X1 U10665 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9126) );
  MUX2_X1 U10666 ( .A(n9126), .B(n9224), .S(n10557), .Z(n9128) );
  NAND2_X1 U10667 ( .A1(n9226), .A2(n9159), .ZN(n9127) );
  OAI211_X1 U10668 ( .C1(n9162), .C2(n9229), .A(n9128), .B(n9127), .ZN(
        P2_U3480) );
  INV_X1 U10669 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9129) );
  MUX2_X1 U10670 ( .A(n9129), .B(n9230), .S(n10557), .Z(n9131) );
  NAND2_X1 U10671 ( .A1(n9232), .A2(n9159), .ZN(n9130) );
  OAI211_X1 U10672 ( .C1(n9162), .C2(n9235), .A(n9131), .B(n9130), .ZN(
        P2_U3479) );
  MUX2_X1 U10673 ( .A(n9132), .B(n9236), .S(n10557), .Z(n9134) );
  NAND2_X1 U10674 ( .A1(n9238), .A2(n9159), .ZN(n9133) );
  OAI211_X1 U10675 ( .C1(n9162), .C2(n9241), .A(n9134), .B(n9133), .ZN(
        P2_U3478) );
  INV_X1 U10676 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9137) );
  AOI21_X1 U10677 ( .B1(n10544), .B2(n9136), .A(n9135), .ZN(n9242) );
  MUX2_X1 U10678 ( .A(n9137), .B(n9242), .S(n10557), .Z(n9138) );
  OAI21_X1 U10679 ( .B1(n9245), .B2(n9172), .A(n9138), .ZN(P2_U3477) );
  MUX2_X1 U10680 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9246), .S(n10557), .Z(
        n9140) );
  OAI22_X1 U10681 ( .A1(n9248), .A2(n9162), .B1(n9247), .B2(n9172), .ZN(n9139)
         );
  OR2_X1 U10682 ( .A1(n9140), .A2(n9139), .ZN(P2_U3476) );
  MUX2_X1 U10683 ( .A(n9141), .B(n9251), .S(n10557), .Z(n9143) );
  NAND2_X1 U10684 ( .A1(n9253), .A2(n9159), .ZN(n9142) );
  OAI211_X1 U10685 ( .C1(n9256), .C2(n9162), .A(n9143), .B(n9142), .ZN(
        P2_U3475) );
  AOI22_X1 U10686 ( .A1(n9145), .A2(n10544), .B1(n10543), .B2(n9144), .ZN(
        n9146) );
  NAND2_X1 U10687 ( .A1(n9147), .A2(n9146), .ZN(n9257) );
  MUX2_X1 U10688 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9257), .S(n10557), .Z(
        P2_U3474) );
  MUX2_X1 U10689 ( .A(n9148), .B(n9258), .S(n10557), .Z(n9150) );
  NAND2_X1 U10690 ( .A1(n9260), .A2(n9159), .ZN(n9149) );
  OAI211_X1 U10691 ( .C1(n9263), .C2(n9162), .A(n9150), .B(n9149), .ZN(
        P2_U3473) );
  MUX2_X1 U10692 ( .A(n9151), .B(n9264), .S(n10557), .Z(n9153) );
  NAND2_X1 U10693 ( .A1(n9266), .A2(n9159), .ZN(n9152) );
  OAI211_X1 U10694 ( .C1(n9162), .C2(n9269), .A(n9153), .B(n9152), .ZN(
        P2_U3472) );
  INV_X1 U10695 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9156) );
  AOI21_X1 U10696 ( .B1(n10543), .B2(n9155), .A(n9154), .ZN(n9270) );
  MUX2_X1 U10697 ( .A(n9156), .B(n9270), .S(n10557), .Z(n9157) );
  OAI21_X1 U10698 ( .B1(n9162), .B2(n9273), .A(n9157), .ZN(P2_U3471) );
  MUX2_X1 U10699 ( .A(n9158), .B(n9274), .S(n10557), .Z(n9161) );
  NAND2_X1 U10700 ( .A1(n9276), .A2(n9159), .ZN(n9160) );
  OAI211_X1 U10701 ( .C1(n9281), .C2(n9162), .A(n9161), .B(n9160), .ZN(
        P2_U3470) );
  AOI21_X1 U10702 ( .B1(n9169), .B2(n9164), .A(n9163), .ZN(n9282) );
  MUX2_X1 U10703 ( .A(n9165), .B(n9282), .S(n10557), .Z(n9166) );
  OAI21_X1 U10704 ( .B1(n9285), .B2(n9172), .A(n9166), .ZN(P2_U3469) );
  AOI21_X1 U10705 ( .B1(n9169), .B2(n9168), .A(n9167), .ZN(n9286) );
  MUX2_X1 U10706 ( .A(n9170), .B(n9286), .S(n10557), .Z(n9171) );
  OAI21_X1 U10707 ( .B1(n9290), .B2(n9172), .A(n9171), .ZN(P2_U3468) );
  INV_X1 U10708 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9174) );
  MUX2_X1 U10709 ( .A(n9174), .B(n9173), .S(n10557), .Z(n9175) );
  INV_X1 U10710 ( .A(n9175), .ZN(P2_U3467) );
  MUX2_X1 U10711 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9176), .S(n10557), .Z(
        P2_U3459) );
  INV_X1 U10712 ( .A(n9177), .ZN(n9180) );
  NAND2_X1 U10713 ( .A1(n10550), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9179) );
  NAND2_X1 U10714 ( .A1(n9178), .A2(n10548), .ZN(n9182) );
  OAI211_X1 U10715 ( .C1(n9180), .C2(n9289), .A(n9179), .B(n9182), .ZN(
        P2_U3458) );
  NAND2_X1 U10716 ( .A1(n10550), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9181) );
  OAI211_X1 U10717 ( .C1(n9183), .C2(n9289), .A(n9182), .B(n9181), .ZN(
        P2_U3457) );
  INV_X1 U10718 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9185) );
  MUX2_X1 U10719 ( .A(n9185), .B(n9184), .S(n10548), .Z(n9188) );
  NAND2_X1 U10720 ( .A1(n9186), .A2(n9277), .ZN(n9187) );
  INV_X1 U10721 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9191) );
  MUX2_X1 U10722 ( .A(n9191), .B(n9190), .S(n10548), .Z(n9194) );
  NAND2_X1 U10723 ( .A1(n9192), .A2(n9277), .ZN(n9193) );
  OAI211_X1 U10724 ( .C1(n9195), .C2(n9280), .A(n9194), .B(n9193), .ZN(
        P2_U3454) );
  INV_X1 U10725 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9197) );
  MUX2_X1 U10726 ( .A(n9197), .B(n4425), .S(n10548), .Z(n9200) );
  NAND2_X1 U10727 ( .A1(n9198), .A2(n9277), .ZN(n9199) );
  OAI211_X1 U10728 ( .C1(n9201), .C2(n9280), .A(n9200), .B(n9199), .ZN(
        P2_U3453) );
  MUX2_X1 U10729 ( .A(n9203), .B(n9202), .S(n10548), .Z(n9206) );
  NAND2_X1 U10730 ( .A1(n9204), .A2(n9277), .ZN(n9205) );
  OAI211_X1 U10731 ( .C1(n9207), .C2(n9280), .A(n9206), .B(n9205), .ZN(
        P2_U3452) );
  INV_X1 U10732 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9209) );
  MUX2_X1 U10733 ( .A(n9209), .B(n9208), .S(n10548), .Z(n9212) );
  NAND2_X1 U10734 ( .A1(n9210), .A2(n9277), .ZN(n9211) );
  OAI211_X1 U10735 ( .C1(n9213), .C2(n9280), .A(n9212), .B(n9211), .ZN(
        P2_U3451) );
  INV_X1 U10736 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9215) );
  MUX2_X1 U10737 ( .A(n9215), .B(n9214), .S(n10548), .Z(n9218) );
  NAND2_X1 U10738 ( .A1(n9216), .A2(n9277), .ZN(n9217) );
  OAI211_X1 U10739 ( .C1(n9219), .C2(n9280), .A(n9218), .B(n9217), .ZN(
        P2_U3450) );
  MUX2_X1 U10740 ( .A(n9221), .B(n9220), .S(n10548), .Z(n9222) );
  OAI21_X1 U10741 ( .B1(n9223), .B2(n9289), .A(n9222), .ZN(P2_U3449) );
  INV_X1 U10742 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9225) );
  MUX2_X1 U10743 ( .A(n9225), .B(n9224), .S(n10548), .Z(n9228) );
  NAND2_X1 U10744 ( .A1(n9226), .A2(n9277), .ZN(n9227) );
  OAI211_X1 U10745 ( .C1(n9229), .C2(n9280), .A(n9228), .B(n9227), .ZN(
        P2_U3448) );
  INV_X1 U10746 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9231) );
  MUX2_X1 U10747 ( .A(n9231), .B(n9230), .S(n10548), .Z(n9234) );
  NAND2_X1 U10748 ( .A1(n9232), .A2(n9277), .ZN(n9233) );
  OAI211_X1 U10749 ( .C1(n9235), .C2(n9280), .A(n9234), .B(n9233), .ZN(
        P2_U3447) );
  INV_X1 U10750 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9237) );
  MUX2_X1 U10751 ( .A(n9237), .B(n9236), .S(n10548), .Z(n9240) );
  NAND2_X1 U10752 ( .A1(n9238), .A2(n9277), .ZN(n9239) );
  OAI211_X1 U10753 ( .C1(n9241), .C2(n9280), .A(n9240), .B(n9239), .ZN(
        P2_U3446) );
  MUX2_X1 U10754 ( .A(n9243), .B(n9242), .S(n10548), .Z(n9244) );
  OAI21_X1 U10755 ( .B1(n9245), .B2(n9289), .A(n9244), .ZN(P2_U3444) );
  MUX2_X1 U10756 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9246), .S(n10548), .Z(
        n9250) );
  OAI22_X1 U10757 ( .A1(n9248), .A2(n9280), .B1(n9247), .B2(n9289), .ZN(n9249)
         );
  OR2_X1 U10758 ( .A1(n9250), .A2(n9249), .ZN(P2_U3441) );
  MUX2_X1 U10759 ( .A(n9252), .B(n9251), .S(n10548), .Z(n9255) );
  NAND2_X1 U10760 ( .A1(n9253), .A2(n9277), .ZN(n9254) );
  OAI211_X1 U10761 ( .C1(n9256), .C2(n9280), .A(n9255), .B(n9254), .ZN(
        P2_U3438) );
  MUX2_X1 U10762 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9257), .S(n10548), .Z(
        P2_U3435) );
  MUX2_X1 U10763 ( .A(n9259), .B(n9258), .S(n10548), .Z(n9262) );
  NAND2_X1 U10764 ( .A1(n9260), .A2(n9277), .ZN(n9261) );
  OAI211_X1 U10765 ( .C1(n9263), .C2(n9280), .A(n9262), .B(n9261), .ZN(
        P2_U3432) );
  MUX2_X1 U10766 ( .A(n9265), .B(n9264), .S(n10548), .Z(n9268) );
  NAND2_X1 U10767 ( .A1(n9266), .A2(n9277), .ZN(n9267) );
  OAI211_X1 U10768 ( .C1(n9269), .C2(n9280), .A(n9268), .B(n9267), .ZN(
        P2_U3429) );
  MUX2_X1 U10769 ( .A(n9271), .B(n9270), .S(n10548), .Z(n9272) );
  OAI21_X1 U10770 ( .B1(n9273), .B2(n9280), .A(n9272), .ZN(P2_U3426) );
  MUX2_X1 U10771 ( .A(n9275), .B(n9274), .S(n10548), .Z(n9279) );
  NAND2_X1 U10772 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  OAI211_X1 U10773 ( .C1(n9281), .C2(n9280), .A(n9279), .B(n9278), .ZN(
        P2_U3423) );
  INV_X1 U10774 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9283) );
  MUX2_X1 U10775 ( .A(n9283), .B(n9282), .S(n10548), .Z(n9284) );
  OAI21_X1 U10776 ( .B1(n9285), .B2(n9289), .A(n9284), .ZN(P2_U3420) );
  MUX2_X1 U10777 ( .A(n9287), .B(n9286), .S(n10548), .Z(n9288) );
  OAI21_X1 U10778 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(P2_U3417) );
  INV_X1 U10779 ( .A(n9291), .ZN(n10317) );
  NOR4_X1 U10780 ( .A1(n9292), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n4693), .ZN(n9293) );
  AOI21_X1 U10781 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n9309), .A(n9293), .ZN(
        n9294) );
  OAI21_X1 U10782 ( .B1(n10317), .B2(n9307), .A(n9294), .ZN(P2_U3264) );
  INV_X1 U10783 ( .A(n9295), .ZN(n10319) );
  AOI22_X1 U10784 ( .A1(n9296), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9309), .ZN(n9297) );
  OAI21_X1 U10785 ( .B1(n10319), .B2(n9307), .A(n9297), .ZN(P2_U3265) );
  INV_X1 U10786 ( .A(n9298), .ZN(n10321) );
  AOI22_X1 U10787 ( .A1(n9299), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9309), .ZN(n9300) );
  OAI21_X1 U10788 ( .B1(n10321), .B2(n9307), .A(n9300), .ZN(P2_U3266) );
  NAND2_X1 U10789 ( .A1(n9309), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9301) );
  OAI211_X1 U10790 ( .C1(n9303), .C2(n9307), .A(n9302), .B(n9301), .ZN(
        P2_U3267) );
  INV_X1 U10791 ( .A(n9304), .ZN(n10324) );
  NAND2_X1 U10792 ( .A1(n9309), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n9305) );
  OAI211_X1 U10793 ( .C1(n10324), .C2(n9307), .A(n9306), .B(n9305), .ZN(
        P2_U3268) );
  INV_X1 U10794 ( .A(n9308), .ZN(n10334) );
  AOI22_X1 U10795 ( .A1(n9310), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9309), .ZN(n9311) );
  OAI21_X1 U10796 ( .B1(n10334), .B2(n9307), .A(n9311), .ZN(P2_U3271) );
  MUX2_X1 U10797 ( .A(n9312), .B(n4848), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10798 ( .A1(n9313), .A2(n9314), .ZN(n9318) );
  XNOR2_X1 U10799 ( .A(n9316), .B(n9315), .ZN(n9317) );
  XNOR2_X1 U10800 ( .A(n9318), .B(n9317), .ZN(n9325) );
  NOR2_X1 U10801 ( .A1(n9552), .A2(n9319), .ZN(n9323) );
  OAI21_X1 U10802 ( .B1(n9554), .B2(n9321), .A(n9320), .ZN(n9322) );
  AOI211_X1 U10803 ( .C1(n10230), .C2(n9557), .A(n9323), .B(n9322), .ZN(n9324)
         );
  OAI21_X1 U10804 ( .B1(n9325), .B2(n9559), .A(n9324), .ZN(P1_U3215) );
  NOR2_X1 U10805 ( .A1(n4463), .A2(n9326), .ZN(n9486) );
  AOI21_X1 U10806 ( .B1(n4463), .B2(n9326), .A(n9486), .ZN(n9327) );
  NAND2_X1 U10807 ( .A1(n9327), .A2(n9328), .ZN(n9489) );
  OAI21_X1 U10808 ( .B1(n9328), .B2(n9327), .A(n9489), .ZN(n9329) );
  NAND2_X1 U10809 ( .A1(n9329), .A2(n9533), .ZN(n9335) );
  NAND2_X1 U10810 ( .A1(n9832), .A2(n4420), .ZN(n9331) );
  NAND2_X1 U10811 ( .A1(n9830), .A2(n9551), .ZN(n9330) );
  NAND2_X1 U10812 ( .A1(n9331), .A2(n9330), .ZN(n10341) );
  OAI21_X1 U10813 ( .B1(n9554), .B2(n10343), .A(n9332), .ZN(n9333) );
  AOI21_X1 U10814 ( .B1(n9542), .B2(n10341), .A(n9333), .ZN(n9334) );
  OAI211_X1 U10815 ( .C1(n10469), .C2(n9545), .A(n9335), .B(n9334), .ZN(
        P1_U3217) );
  XNOR2_X1 U10816 ( .A(n9337), .B(n9336), .ZN(n9341) );
  AOI22_X1 U10817 ( .A1(n9821), .A2(n9551), .B1(n4420), .B2(n9823), .ZN(n10094) );
  NOR2_X1 U10818 ( .A1(n10094), .A2(n9552), .ZN(n9339) );
  NAND2_X1 U10819 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9992) );
  OAI21_X1 U10820 ( .B1(n9554), .B2(n10088), .A(n9992), .ZN(n9338) );
  AOI211_X1 U10821 ( .C1(n10206), .C2(n9557), .A(n9339), .B(n9338), .ZN(n9340)
         );
  OAI21_X1 U10822 ( .B1(n9341), .B2(n9559), .A(n9340), .ZN(P1_U3219) );
  NAND2_X1 U10823 ( .A1(n9347), .A2(n4427), .ZN(n9344) );
  NAND2_X1 U10824 ( .A1(n9815), .A2(n9342), .ZN(n9343) );
  NAND2_X1 U10825 ( .A1(n9344), .A2(n9343), .ZN(n9346) );
  XNOR2_X1 U10826 ( .A(n9346), .B(n9345), .ZN(n9349) );
  AOI22_X1 U10827 ( .A1(n9347), .A2(n8137), .B1(n4427), .B2(n9815), .ZN(n9348)
         );
  XNOR2_X1 U10828 ( .A(n9349), .B(n9348), .ZN(n9358) );
  NAND3_X1 U10829 ( .A1(n9350), .A2(n9533), .A3(n9358), .ZN(n9361) );
  OAI22_X1 U10830 ( .A1(n9352), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9351), .ZN(n9355) );
  NOR2_X1 U10831 ( .A1(n9353), .A2(n9545), .ZN(n9354) );
  AOI211_X1 U10832 ( .C1(n9542), .C2(n9356), .A(n9355), .B(n9354), .ZN(n9360)
         );
  NAND3_X1 U10833 ( .A1(n9358), .A2(n9357), .A3(n9533), .ZN(n9359) );
  NAND4_X1 U10834 ( .A1(n9362), .A2(n9361), .A3(n9360), .A4(n9359), .ZN(
        P1_U3220) );
  NOR2_X1 U10835 ( .A1(n9364), .A2(n9363), .ZN(n9437) );
  XNOR2_X1 U10836 ( .A(n9437), .B(n9365), .ZN(n9367) );
  NOR2_X1 U10837 ( .A1(n9367), .A2(n9366), .ZN(n9438) );
  AOI21_X1 U10838 ( .B1(n9367), .B2(n9366), .A(n9438), .ZN(n9375) );
  OAI21_X1 U10839 ( .B1(n9554), .B2(n9369), .A(n9368), .ZN(n9372) );
  NOR2_X1 U10840 ( .A1(n9545), .A2(n9370), .ZN(n9371) );
  AOI211_X1 U10841 ( .C1(n9542), .C2(n9373), .A(n9372), .B(n9371), .ZN(n9374)
         );
  OAI21_X1 U10842 ( .B1(n9375), .B2(n9559), .A(n9374), .ZN(P1_U3221) );
  XNOR2_X1 U10843 ( .A(n9377), .B(n9376), .ZN(n9378) );
  XNOR2_X1 U10844 ( .A(n9379), .B(n9378), .ZN(n9383) );
  AOI22_X1 U10845 ( .A1(n9819), .A2(n9551), .B1(n4420), .B2(n9821), .ZN(n10055) );
  INV_X1 U10846 ( .A(n9554), .ZN(n9480) );
  AOI22_X1 U10847 ( .A1(n9480), .A2(n10062), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(n10311), .ZN(n9380) );
  OAI21_X1 U10848 ( .B1(n10055), .B2(n9552), .A(n9380), .ZN(n9381) );
  AOI21_X1 U10849 ( .B1(n10194), .B2(n9557), .A(n9381), .ZN(n9382) );
  OAI21_X1 U10850 ( .B1(n9383), .B2(n9559), .A(n9382), .ZN(P1_U3223) );
  INV_X1 U10851 ( .A(n9384), .ZN(n9389) );
  NOR3_X1 U10852 ( .A1(n9385), .A2(n9387), .A3(n9386), .ZN(n9388) );
  OAI21_X1 U10853 ( .B1(n9389), .B2(n9388), .A(n9533), .ZN(n9396) );
  INV_X1 U10854 ( .A(n9390), .ZN(n9394) );
  OAI21_X1 U10855 ( .B1(n9554), .B2(n9392), .A(n9391), .ZN(n9393) );
  AOI21_X1 U10856 ( .B1(n9542), .B2(n9394), .A(n9393), .ZN(n9395) );
  OAI211_X1 U10857 ( .C1(n5390), .C2(n9545), .A(n9396), .B(n9395), .ZN(
        P1_U3224) );
  OAI21_X1 U10858 ( .B1(n9398), .B2(n9397), .A(n9531), .ZN(n9399) );
  NAND2_X1 U10859 ( .A1(n9399), .A2(n9533), .ZN(n9405) );
  OAI22_X1 U10860 ( .A1(n9401), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9400), .ZN(n9402) );
  AOI21_X1 U10861 ( .B1(n9403), .B2(n9542), .A(n9402), .ZN(n9404) );
  OAI211_X1 U10862 ( .C1(n9406), .C2(n9545), .A(n9405), .B(n9404), .ZN(
        P1_U3225) );
  OAI21_X1 U10863 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9413) );
  NAND2_X1 U10864 ( .A1(n9411), .A2(n9410), .ZN(n9547) );
  NOR2_X1 U10865 ( .A1(n9411), .A2(n9410), .ZN(n9546) );
  AOI21_X1 U10866 ( .B1(n9549), .B2(n9547), .A(n9546), .ZN(n9412) );
  XOR2_X1 U10867 ( .A(n9413), .B(n9412), .Z(n9418) );
  AOI22_X1 U10868 ( .A1(n9824), .A2(n9551), .B1(n4420), .B2(n9826), .ZN(n10137) );
  NOR2_X1 U10869 ( .A1(n10137), .A2(n9552), .ZN(n9416) );
  OAI22_X1 U10870 ( .A1(n9554), .A2(n10140), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9414), .ZN(n9415) );
  AOI211_X1 U10871 ( .C1(n10220), .C2(n9557), .A(n9416), .B(n9415), .ZN(n9417)
         );
  OAI21_X1 U10872 ( .B1(n9418), .B2(n9559), .A(n9417), .ZN(P1_U3226) );
  NAND2_X1 U10873 ( .A1(n9419), .A2(n9497), .ZN(n9420) );
  XNOR2_X1 U10874 ( .A(n9498), .B(n9420), .ZN(n9424) );
  AOI22_X1 U10875 ( .A1(n9823), .A2(n9551), .B1(n4420), .B2(n9825), .ZN(n10127) );
  NOR2_X1 U10876 ( .A1(n10127), .A2(n9552), .ZN(n9422) );
  NAND2_X1 U10877 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9950) );
  OAI21_X1 U10878 ( .B1(n9554), .B2(n10118), .A(n9950), .ZN(n9421) );
  AOI211_X1 U10879 ( .C1(n10215), .C2(n9557), .A(n9422), .B(n9421), .ZN(n9423)
         );
  OAI21_X1 U10880 ( .B1(n9424), .B2(n9559), .A(n9423), .ZN(P1_U3228) );
  INV_X1 U10881 ( .A(n6074), .ZN(n10033) );
  INV_X1 U10882 ( .A(n8136), .ZN(n9427) );
  NOR3_X1 U10883 ( .A1(n9427), .A2(n9426), .A3(n9425), .ZN(n9430) );
  INV_X1 U10884 ( .A(n9428), .ZN(n9429) );
  OAI21_X1 U10885 ( .B1(n9430), .B2(n9429), .A(n9533), .ZN(n9436) );
  OAI22_X1 U10886 ( .A1(n9536), .A2(n9537), .B1(n9431), .B2(n9535), .ZN(n10026) );
  INV_X1 U10887 ( .A(n10030), .ZN(n9433) );
  OAI22_X1 U10888 ( .A1(n9433), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9432), .ZN(n9434) );
  AOI21_X1 U10889 ( .B1(n10026), .B2(n9542), .A(n9434), .ZN(n9435) );
  OAI211_X1 U10890 ( .C1(n10033), .C2(n9545), .A(n9436), .B(n9435), .ZN(
        P1_U3229) );
  INV_X1 U10891 ( .A(n9437), .ZN(n9439) );
  AOI21_X1 U10892 ( .B1(n9440), .B2(n9439), .A(n9438), .ZN(n9443) );
  OAI211_X1 U10893 ( .C1(n9443), .C2(n9442), .A(n9533), .B(n9441), .ZN(n9452)
         );
  AND2_X1 U10894 ( .A1(n9445), .A2(n9444), .ZN(n9449) );
  OR2_X1 U10895 ( .A1(n9554), .A2(n9446), .ZN(n9447) );
  OAI211_X1 U10896 ( .C1(n9552), .C2(n9449), .A(n9448), .B(n9447), .ZN(n9450)
         );
  INV_X1 U10897 ( .A(n9450), .ZN(n9451) );
  OAI211_X1 U10898 ( .C1(n10462), .C2(n9545), .A(n9452), .B(n9451), .ZN(
        P1_U3231) );
  NAND2_X1 U10899 ( .A1(n9454), .A2(n9453), .ZN(n9456) );
  XOR2_X1 U10900 ( .A(n9456), .B(n9455), .Z(n9462) );
  AND2_X1 U10901 ( .A1(n9822), .A2(n4420), .ZN(n9457) );
  AOI21_X1 U10902 ( .B1(n9820), .B2(n9522), .A(n9457), .ZN(n10072) );
  NOR2_X1 U10903 ( .A1(n10072), .A2(n9552), .ZN(n9460) );
  OAI22_X1 U10904 ( .A1(n9554), .A2(n10077), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9458), .ZN(n9459) );
  AOI211_X1 U10905 ( .C1(n10197), .C2(n9557), .A(n9460), .B(n9459), .ZN(n9461)
         );
  OAI21_X1 U10906 ( .B1(n9462), .B2(n9559), .A(n9461), .ZN(P1_U3233) );
  OAI21_X1 U10907 ( .B1(n9464), .B2(n9463), .A(n9313), .ZN(n9465) );
  NAND2_X1 U10908 ( .A1(n9465), .A2(n9533), .ZN(n9472) );
  INV_X1 U10909 ( .A(n9466), .ZN(n9470) );
  OAI21_X1 U10910 ( .B1(n9554), .B2(n9468), .A(n9467), .ZN(n9469) );
  AOI21_X1 U10911 ( .B1(n9542), .B2(n9470), .A(n9469), .ZN(n9471) );
  OAI211_X1 U10912 ( .C1(n9473), .C2(n9545), .A(n9472), .B(n9471), .ZN(
        P1_U3234) );
  XOR2_X1 U10913 ( .A(n9475), .B(n9474), .Z(n9476) );
  XNOR2_X1 U10914 ( .A(n9477), .B(n9476), .ZN(n9485) );
  INV_X1 U10915 ( .A(n9478), .ZN(n9482) );
  AOI22_X1 U10916 ( .A1(n9480), .A2(n9479), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9481) );
  OAI21_X1 U10917 ( .B1(n9482), .B2(n9552), .A(n9481), .ZN(n9483) );
  AOI21_X1 U10918 ( .B1(n9562), .B2(n9557), .A(n9483), .ZN(n9484) );
  OAI21_X1 U10919 ( .B1(n9485), .B2(n9559), .A(n9484), .ZN(P1_U3235) );
  INV_X1 U10920 ( .A(n9486), .ZN(n9487) );
  AND3_X1 U10921 ( .A1(n9489), .A2(n9488), .A3(n9487), .ZN(n9490) );
  OAI21_X1 U10922 ( .B1(n9490), .B2(n9385), .A(n9533), .ZN(n9496) );
  OAI21_X1 U10923 ( .B1(n9554), .B2(n9492), .A(n9491), .ZN(n9493) );
  AOI21_X1 U10924 ( .B1(n9542), .B2(n9494), .A(n9493), .ZN(n9495) );
  OAI211_X1 U10925 ( .C1(n10474), .C2(n9545), .A(n9496), .B(n9495), .ZN(
        P1_U3236) );
  NAND2_X1 U10926 ( .A1(n9498), .A2(n9497), .ZN(n9500) );
  NAND2_X1 U10927 ( .A1(n9500), .A2(n9499), .ZN(n9501) );
  NAND2_X1 U10928 ( .A1(n9502), .A2(n9501), .ZN(n9504) );
  XNOR2_X1 U10929 ( .A(n9504), .B(n9503), .ZN(n9512) );
  NAND2_X1 U10930 ( .A1(n9822), .A2(n9522), .ZN(n9505) );
  OAI21_X1 U10931 ( .B1(n9506), .B2(n9535), .A(n9505), .ZN(n10102) );
  INV_X1 U10932 ( .A(n10109), .ZN(n9508) );
  OAI22_X1 U10933 ( .A1(n9554), .A2(n9508), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9507), .ZN(n9510) );
  NOR2_X1 U10934 ( .A1(n10112), .A2(n9545), .ZN(n9509) );
  AOI211_X1 U10935 ( .C1(n9542), .C2(n10102), .A(n9510), .B(n9509), .ZN(n9511)
         );
  OAI21_X1 U10936 ( .B1(n9512), .B2(n9559), .A(n9511), .ZN(P1_U3238) );
  INV_X1 U10937 ( .A(n9513), .ZN(n9515) );
  AOI21_X1 U10938 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(n9521) );
  OAI21_X1 U10939 ( .B1(n9519), .B2(n9518), .A(n9517), .ZN(n9520) );
  XOR2_X1 U10940 ( .A(n9521), .B(n9520), .Z(n9529) );
  NAND2_X1 U10941 ( .A1(n9836), .A2(n4420), .ZN(n9524) );
  NAND2_X1 U10942 ( .A1(n9834), .A2(n9522), .ZN(n9523) );
  AND2_X1 U10943 ( .A1(n9524), .A2(n9523), .ZN(n10357) );
  NAND2_X1 U10944 ( .A1(n10311), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9894) );
  OR2_X1 U10945 ( .A1(n9554), .A2(n10360), .ZN(n9525) );
  OAI211_X1 U10946 ( .C1(n9552), .C2(n10357), .A(n9894), .B(n9525), .ZN(n9526)
         );
  AOI21_X1 U10947 ( .B1(n9527), .B2(n9557), .A(n9526), .ZN(n9528) );
  OAI21_X1 U10948 ( .B1(n9529), .B2(n9559), .A(n9528), .ZN(P1_U3239) );
  OAI22_X1 U10949 ( .A1(n9538), .A2(n9537), .B1(n9536), .B2(n9535), .ZN(n10009) );
  INV_X1 U10950 ( .A(n10015), .ZN(n9540) );
  OAI22_X1 U10951 ( .A1(n9540), .A2(n9554), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9539), .ZN(n9541) );
  AOI21_X1 U10952 ( .B1(n10009), .B2(n9542), .A(n9541), .ZN(n9543) );
  OAI211_X1 U10953 ( .C1(n10180), .C2(n9545), .A(n9544), .B(n9543), .ZN(
        P1_U3240) );
  INV_X1 U10954 ( .A(n9546), .ZN(n9548) );
  NAND2_X1 U10955 ( .A1(n9548), .A2(n9547), .ZN(n9550) );
  XNOR2_X1 U10956 ( .A(n9550), .B(n9549), .ZN(n9560) );
  AOI22_X1 U10957 ( .A1(n9827), .A2(n4420), .B1(n9551), .B2(n9825), .ZN(n10151) );
  NOR2_X1 U10958 ( .A1(n9552), .A2(n10151), .ZN(n9556) );
  OAI22_X1 U10959 ( .A1(n9554), .A2(n10156), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9553), .ZN(n9555) );
  AOI211_X1 U10960 ( .C1(n10225), .C2(n9557), .A(n9556), .B(n9555), .ZN(n9558)
         );
  OAI21_X1 U10961 ( .B1(n9560), .B2(n9559), .A(n9558), .ZN(P1_U3241) );
  NAND2_X1 U10962 ( .A1(n9562), .A2(n9561), .ZN(n9563) );
  INV_X1 U10963 ( .A(n9699), .ZN(n9565) );
  INV_X1 U10964 ( .A(n9769), .ZN(n9564) );
  NOR2_X1 U10965 ( .A1(n9565), .A2(n9564), .ZN(n9622) );
  NAND2_X1 U10966 ( .A1(n6054), .A2(n9792), .ZN(n9566) );
  AND2_X1 U10967 ( .A1(n9567), .A2(n6054), .ZN(n9749) );
  NAND4_X1 U10968 ( .A1(n9568), .A2(n9571), .A3(n9577), .A4(n9791), .ZN(n9569)
         );
  AOI21_X1 U10969 ( .B1(n9570), .B2(n9749), .A(n9569), .ZN(n9579) );
  INV_X1 U10970 ( .A(n9571), .ZN(n9573) );
  NAND3_X1 U10971 ( .A1(n9573), .A2(n9572), .A3(n9792), .ZN(n9576) );
  NAND3_X1 U10972 ( .A1(n9574), .A2(n9577), .A3(n9791), .ZN(n9575) );
  NAND2_X1 U10973 ( .A1(n9591), .A2(n9583), .ZN(n9586) );
  INV_X1 U10974 ( .A(n9584), .ZN(n9585) );
  MUX2_X1 U10975 ( .A(n9586), .B(n9585), .S(n9792), .Z(n9587) );
  INV_X1 U10976 ( .A(n9587), .ZN(n9588) );
  INV_X1 U10977 ( .A(n9594), .ZN(n9592) );
  OAI211_X1 U10978 ( .C1(n9592), .C2(n9591), .A(n9792), .B(n9597), .ZN(n9593)
         );
  NAND2_X1 U10979 ( .A1(n9594), .A2(n9596), .ZN(n9600) );
  INV_X1 U10980 ( .A(n9751), .ZN(n9598) );
  AND2_X1 U10981 ( .A1(n9601), .A2(n9792), .ZN(n9602) );
  NAND2_X1 U10982 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  OAI21_X1 U10983 ( .B1(n9791), .B2(n9829), .A(n9604), .ZN(n9607) );
  INV_X1 U10984 ( .A(n9604), .ZN(n9606) );
  AOI22_X1 U10985 ( .A1(n9607), .A2(n10240), .B1(n9606), .B2(n9605), .ZN(n9608) );
  AND2_X1 U10986 ( .A1(n9621), .A2(n9613), .ZN(n9762) );
  INV_X1 U10987 ( .A(n9616), .ZN(n9610) );
  AOI21_X1 U10988 ( .B1(n9611), .B2(n9762), .A(n9610), .ZN(n9612) );
  INV_X1 U10989 ( .A(n9758), .ZN(n9614) );
  AND2_X1 U10990 ( .A1(n9617), .A2(n9616), .ZN(n9760) );
  NAND3_X1 U10991 ( .A1(n9618), .A2(n9760), .A3(n10148), .ZN(n9620) );
  AND2_X1 U10992 ( .A1(n9768), .A2(n9791), .ZN(n9623) );
  AND2_X1 U10993 ( .A1(n9769), .A2(n9623), .ZN(n9627) );
  INV_X1 U10994 ( .A(n9627), .ZN(n9630) );
  NAND2_X1 U10995 ( .A1(n9625), .A2(n9624), .ZN(n9765) );
  NOR2_X1 U10996 ( .A1(n9822), .A2(n9792), .ZN(n9626) );
  AOI22_X1 U10997 ( .A1(n9627), .A2(n9765), .B1(n9626), .B2(n10206), .ZN(n9629) );
  OAI211_X1 U10998 ( .C1(n9631), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9635)
         );
  INV_X1 U10999 ( .A(n9688), .ZN(n9638) );
  NAND3_X1 U11000 ( .A1(n9700), .A2(n9699), .A3(n9791), .ZN(n9632) );
  OAI21_X1 U11001 ( .B1(n9633), .B2(n9791), .A(n9632), .ZN(n9634) );
  INV_X1 U11002 ( .A(n9700), .ZN(n9639) );
  NAND2_X1 U11003 ( .A1(n9636), .A2(n9791), .ZN(n9637) );
  OAI211_X1 U11004 ( .C1(n9639), .C2(n9791), .A(n9638), .B(n9637), .ZN(n9640)
         );
  NAND2_X1 U11005 ( .A1(n9641), .A2(n10045), .ZN(n9703) );
  INV_X1 U11006 ( .A(n10025), .ZN(n10021) );
  OAI21_X1 U11007 ( .B1(n9702), .B2(n9791), .A(n10021), .ZN(n9643) );
  MUX2_X1 U11008 ( .A(n9705), .B(n9713), .S(n9791), .Z(n9642) );
  NOR2_X1 U11009 ( .A1(n9714), .A2(n9791), .ZN(n9644) );
  OAI211_X1 U11010 ( .C1(n9656), .C2(n9645), .A(n9644), .B(n9653), .ZN(n9650)
         );
  NOR3_X1 U11011 ( .A1(n10016), .A2(n9654), .A3(n9791), .ZN(n9646) );
  NOR2_X1 U11012 ( .A1(n9720), .A2(n9646), .ZN(n9649) );
  NAND2_X1 U11013 ( .A1(n9648), .A2(n9647), .ZN(n9659) );
  AOI21_X1 U11014 ( .B1(n9650), .B2(n9649), .A(n9659), .ZN(n9651) );
  NOR3_X1 U11015 ( .A1(n10180), .A2(n9792), .A3(n9816), .ZN(n9652) );
  INV_X1 U11016 ( .A(n9653), .ZN(n9716) );
  OR2_X1 U11017 ( .A1(n10016), .A2(n9654), .ZN(n9715) );
  AND2_X1 U11018 ( .A1(n9715), .A2(n9655), .ZN(n9707) );
  INV_X1 U11019 ( .A(n9659), .ZN(n9723) );
  AOI21_X1 U11020 ( .B1(n9723), .B2(n9720), .A(n9660), .ZN(n9661) );
  INV_X1 U11021 ( .A(n9726), .ZN(n9664) );
  INV_X1 U11022 ( .A(n9698), .ZN(n9663) );
  MUX2_X1 U11023 ( .A(n9664), .B(n9663), .S(n9791), .Z(n9665) );
  INV_X1 U11024 ( .A(n9734), .ZN(n9667) );
  NAND2_X1 U11025 ( .A1(n9666), .A2(n9667), .ZN(n9790) );
  INV_X1 U11026 ( .A(n9814), .ZN(n9692) );
  NOR2_X1 U11027 ( .A1(n9692), .A2(n9667), .ZN(n9728) );
  INV_X1 U11028 ( .A(n9798), .ZN(n9669) );
  OR2_X1 U11029 ( .A1(n9730), .A2(n9692), .ZN(n9670) );
  NAND2_X1 U11030 ( .A1(n9790), .A2(n9670), .ZN(n9782) );
  INV_X1 U11031 ( .A(n10386), .ZN(n9673) );
  INV_X1 U11032 ( .A(n9672), .ZN(n10387) );
  NAND4_X1 U11033 ( .A1(n9674), .A2(n9673), .A3(n10387), .A4(n7063), .ZN(n9676) );
  NOR4_X1 U11034 ( .A1(n9676), .A2(n9675), .A3(n10250), .A4(n7798), .ZN(n9679)
         );
  INV_X1 U11035 ( .A(n10356), .ZN(n10365) );
  NAND4_X1 U11036 ( .A1(n9679), .A2(n9678), .A3(n10365), .A4(n9677), .ZN(n9680) );
  NOR4_X1 U11037 ( .A1(n9682), .A2(n9681), .A3(n5224), .A4(n9680), .ZN(n9683)
         );
  NAND4_X1 U11038 ( .A1(n10149), .A2(n9685), .A3(n9684), .A4(n9683), .ZN(n9686) );
  NOR4_X1 U11039 ( .A1(n10101), .A2(n10123), .A3(n10135), .A4(n9686), .ZN(
        n9687) );
  NAND4_X1 U11040 ( .A1(n10047), .A2(n6072), .A3(n10093), .A4(n9687), .ZN(
        n9690) );
  NOR4_X1 U11041 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n10058), .ZN(n9691)
         );
  AND4_X1 U11042 ( .A1(n9691), .A2(n9996), .A3(n10021), .A4(n10012), .ZN(n9693) );
  NAND2_X1 U11043 ( .A1(n9730), .A2(n9692), .ZN(n9727) );
  NAND4_X1 U11044 ( .A1(n9695), .A2(n9694), .A3(n9693), .A4(n9727), .ZN(n9696)
         );
  NOR3_X1 U11045 ( .A1(n9732), .A2(n9782), .A3(n9696), .ZN(n9697) );
  OAI21_X1 U11046 ( .B1(n9697), .B2(n9800), .A(n4613), .ZN(n9740) );
  INV_X1 U11047 ( .A(n9697), .ZN(n9738) );
  NAND2_X1 U11048 ( .A1(n9698), .A2(n7888), .ZN(n9778) );
  NAND2_X1 U11049 ( .A1(n9700), .A2(n9699), .ZN(n9701) );
  OR2_X1 U11050 ( .A1(n9720), .A2(n9701), .ZN(n9709) );
  NAND2_X1 U11051 ( .A1(n9703), .A2(n9702), .ZN(n9704) );
  NAND2_X1 U11052 ( .A1(n9705), .A2(n9704), .ZN(n9706) );
  NAND2_X1 U11053 ( .A1(n9706), .A2(n9713), .ZN(n9708) );
  NAND2_X1 U11054 ( .A1(n9708), .A2(n9707), .ZN(n9719) );
  NOR2_X1 U11055 ( .A1(n9709), .A2(n9719), .ZN(n9742) );
  AND3_X1 U11056 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n9718) );
  AOI21_X1 U11057 ( .B1(n9716), .B2(n9715), .A(n9714), .ZN(n9717) );
  OAI21_X1 U11058 ( .B1(n9719), .B2(n9718), .A(n9717), .ZN(n9722) );
  INV_X1 U11059 ( .A(n9720), .ZN(n9721) );
  NAND2_X1 U11060 ( .A1(n9722), .A2(n9721), .ZN(n9724) );
  NAND2_X1 U11061 ( .A1(n9724), .A2(n9723), .ZN(n9775) );
  AOI21_X1 U11062 ( .B1(n9742), .B2(n9710), .A(n9775), .ZN(n9725) );
  NOR2_X1 U11063 ( .A1(n9778), .A2(n9725), .ZN(n9731) );
  NAND2_X1 U11064 ( .A1(n9727), .A2(n9726), .ZN(n9779) );
  INV_X1 U11065 ( .A(n9728), .ZN(n9729) );
  OAI22_X1 U11066 ( .A1(n9731), .A2(n9779), .B1(n9730), .B2(n9729), .ZN(n9733)
         );
  OAI211_X1 U11067 ( .C1(n10168), .C2(n9734), .A(n9733), .B(n9801), .ZN(n9736)
         );
  NAND3_X1 U11068 ( .A1(n9736), .A2(n9735), .A3(n9790), .ZN(n9737) );
  AOI21_X1 U11069 ( .B1(n9738), .B2(n9737), .A(n9991), .ZN(n9739) );
  AOI21_X1 U11070 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9813) );
  INV_X1 U11071 ( .A(n9742), .ZN(n9774) );
  AOI21_X1 U11072 ( .B1(n5482), .B2(n10421), .A(n7063), .ZN(n9748) );
  NAND2_X1 U11073 ( .A1(n9840), .A2(n10253), .ZN(n9744) );
  AND2_X1 U11074 ( .A1(n9745), .A2(n9744), .ZN(n9747) );
  AND4_X1 U11075 ( .A1(n9749), .A2(n9748), .A3(n9747), .A4(n9746), .ZN(n9750)
         );
  OAI21_X1 U11076 ( .B1(n9743), .B2(n9750), .A(n10339), .ZN(n9752) );
  NAND2_X1 U11077 ( .A1(n9752), .A2(n9751), .ZN(n9754) );
  NAND2_X1 U11078 ( .A1(n9754), .A2(n9753), .ZN(n9757) );
  NAND3_X1 U11079 ( .A1(n9757), .A2(n9756), .A3(n9755), .ZN(n9759) );
  NAND3_X1 U11080 ( .A1(n9759), .A2(n10148), .A3(n9758), .ZN(n9763) );
  INV_X1 U11081 ( .A(n9760), .ZN(n9761) );
  AOI21_X1 U11082 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  OAI21_X1 U11083 ( .B1(n9764), .B2(n10124), .A(n10099), .ZN(n9767) );
  INV_X1 U11084 ( .A(n9765), .ZN(n9766) );
  NAND2_X1 U11085 ( .A1(n9767), .A2(n9766), .ZN(n9770) );
  NAND3_X1 U11086 ( .A1(n9770), .A2(n9769), .A3(n9768), .ZN(n9772) );
  AND2_X1 U11087 ( .A1(n9772), .A2(n9771), .ZN(n9773) );
  NOR2_X1 U11088 ( .A1(n9774), .A2(n9773), .ZN(n9776) );
  NOR2_X1 U11089 ( .A1(n9776), .A2(n9775), .ZN(n9777) );
  NOR2_X1 U11090 ( .A1(n9778), .A2(n9777), .ZN(n9780) );
  NOR2_X1 U11091 ( .A1(n9780), .A2(n9779), .ZN(n9781) );
  OR2_X1 U11092 ( .A1(n9782), .A2(n9781), .ZN(n9783) );
  NAND2_X1 U11093 ( .A1(n9783), .A2(n9801), .ZN(n9788) );
  NAND3_X1 U11094 ( .A1(n9788), .A2(n9991), .A3(n9784), .ZN(n9786) );
  INV_X1 U11095 ( .A(n9797), .ZN(n9785) );
  OAI211_X1 U11096 ( .C1(n9788), .C2(n9787), .A(n9786), .B(n9785), .ZN(n9812)
         );
  INV_X1 U11097 ( .A(n9789), .ZN(n9795) );
  INV_X1 U11098 ( .A(n9790), .ZN(n9793) );
  NAND2_X1 U11099 ( .A1(n9793), .A2(n9792), .ZN(n9794) );
  OR2_X1 U11100 ( .A1(n9797), .A2(n9796), .ZN(n9808) );
  NOR2_X1 U11101 ( .A1(n9808), .A2(n9798), .ZN(n9799) );
  NAND4_X1 U11102 ( .A1(n10409), .A2(n9807), .A3(n9806), .A4(n4420), .ZN(n9809) );
  NAND3_X1 U11103 ( .A1(n9809), .A2(P1_B_REG_SCAN_IN), .A3(n9808), .ZN(n9810)
         );
  OAI211_X1 U11104 ( .C1(n9813), .C2(n9812), .A(n9811), .B(n9810), .ZN(
        P1_U3242) );
  MUX2_X1 U11105 ( .A(n9814), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9839), .Z(
        P1_U3584) );
  MUX2_X1 U11106 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9815), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U11107 ( .A(n9816), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9839), .Z(
        P1_U3580) );
  MUX2_X1 U11108 ( .A(n9817), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9839), .Z(
        P1_U3579) );
  MUX2_X1 U11109 ( .A(n9818), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9839), .Z(
        P1_U3578) );
  MUX2_X1 U11110 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9819), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U11111 ( .A(n9820), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9839), .Z(
        P1_U3575) );
  MUX2_X1 U11112 ( .A(n9821), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9839), .Z(
        P1_U3574) );
  MUX2_X1 U11113 ( .A(n9822), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9839), .Z(
        P1_U3573) );
  MUX2_X1 U11114 ( .A(n9823), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9839), .Z(
        P1_U3572) );
  MUX2_X1 U11115 ( .A(n9824), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9839), .Z(
        P1_U3571) );
  MUX2_X1 U11116 ( .A(n9825), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9839), .Z(
        P1_U3570) );
  MUX2_X1 U11117 ( .A(n9826), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9839), .Z(
        P1_U3569) );
  MUX2_X1 U11118 ( .A(n9827), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9839), .Z(
        P1_U3568) );
  MUX2_X1 U11119 ( .A(n9828), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9839), .Z(
        P1_U3567) );
  MUX2_X1 U11120 ( .A(n9829), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9839), .Z(
        P1_U3566) );
  MUX2_X1 U11121 ( .A(n9830), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9839), .Z(
        P1_U3565) );
  MUX2_X1 U11122 ( .A(n9831), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9839), .Z(
        P1_U3564) );
  MUX2_X1 U11123 ( .A(n9832), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9839), .Z(
        P1_U3563) );
  MUX2_X1 U11124 ( .A(n9833), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9839), .Z(
        P1_U3562) );
  MUX2_X1 U11125 ( .A(n9834), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9839), .Z(
        P1_U3561) );
  MUX2_X1 U11126 ( .A(n9835), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9839), .Z(
        P1_U3560) );
  MUX2_X1 U11127 ( .A(n9836), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9839), .Z(
        P1_U3559) );
  MUX2_X1 U11128 ( .A(n9837), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9839), .Z(
        P1_U3558) );
  MUX2_X1 U11129 ( .A(n9838), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9839), .Z(
        P1_U3557) );
  MUX2_X1 U11130 ( .A(n5482), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9839), .Z(
        P1_U3556) );
  MUX2_X1 U11131 ( .A(n5464), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9839), .Z(
        P1_U3555) );
  MUX2_X1 U11132 ( .A(n9840), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9839), .Z(
        P1_U3554) );
  OAI211_X1 U11133 ( .C1(n9843), .C2(n9842), .A(n9990), .B(n9841), .ZN(n9851)
         );
  AOI22_X1 U11134 ( .A1(n9965), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9850) );
  NAND2_X1 U11135 ( .A1(n9988), .A2(n9844), .ZN(n9849) );
  OAI211_X1 U11136 ( .C1(n9847), .C2(n9846), .A(n9984), .B(n9845), .ZN(n9848)
         );
  NAND4_X1 U11137 ( .A1(n9851), .A2(n9850), .A3(n9849), .A4(n9848), .ZN(
        P1_U3244) );
  AND2_X1 U11138 ( .A1(n10311), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9854) );
  NOR2_X1 U11139 ( .A1(n9975), .A2(n9852), .ZN(n9853) );
  AOI211_X1 U11140 ( .C1(n9965), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n9854), .B(
        n9853), .ZN(n9862) );
  OAI211_X1 U11141 ( .C1(n9857), .C2(n9856), .A(n9984), .B(n9855), .ZN(n9861)
         );
  OAI211_X1 U11142 ( .C1(n9859), .C2(n9858), .A(n9990), .B(n9873), .ZN(n9860)
         );
  NAND3_X1 U11143 ( .A1(n9862), .A2(n9861), .A3(n9860), .ZN(P1_U3246) );
  INV_X1 U11144 ( .A(n9870), .ZN(n9866) );
  INV_X1 U11145 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9864) );
  OAI21_X1 U11146 ( .B1(n9994), .B2(n9864), .A(n9863), .ZN(n9865) );
  AOI21_X1 U11147 ( .B1(n9866), .B2(n9988), .A(n9865), .ZN(n9877) );
  OAI211_X1 U11148 ( .C1(n9869), .C2(n9868), .A(n9984), .B(n9867), .ZN(n9876)
         );
  MUX2_X1 U11149 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6955), .S(n9870), .Z(n9871)
         );
  NAND3_X1 U11150 ( .A1(n9873), .A2(n9872), .A3(n9871), .ZN(n9874) );
  NAND3_X1 U11151 ( .A1(n9990), .A2(n9889), .A3(n9874), .ZN(n9875) );
  NAND4_X1 U11152 ( .A1(n9878), .A2(n9877), .A3(n9876), .A4(n9875), .ZN(
        P1_U3247) );
  INV_X1 U11153 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9880) );
  OAI21_X1 U11154 ( .B1(n9994), .B2(n9880), .A(n9879), .ZN(n9881) );
  AOI21_X1 U11155 ( .B1(n9882), .B2(n9988), .A(n9881), .ZN(n9893) );
  OAI211_X1 U11156 ( .C1(n9885), .C2(n9884), .A(n9984), .B(n9883), .ZN(n9892)
         );
  MUX2_X1 U11157 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6958), .S(n9886), .Z(n9887)
         );
  NAND3_X1 U11158 ( .A1(n9889), .A2(n9888), .A3(n9887), .ZN(n9890) );
  NAND3_X1 U11159 ( .A1(n9990), .A2(n9903), .A3(n9890), .ZN(n9891) );
  NAND3_X1 U11160 ( .A1(n9893), .A2(n9892), .A3(n9891), .ZN(P1_U3248) );
  INV_X1 U11161 ( .A(n9894), .ZN(n9896) );
  NOR2_X1 U11162 ( .A1(n9975), .A2(n9900), .ZN(n9895) );
  AOI211_X1 U11163 ( .C1(n9965), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n9896), .B(
        n9895), .ZN(n9907) );
  OAI211_X1 U11164 ( .C1(n9899), .C2(n9898), .A(n9984), .B(n9897), .ZN(n9906)
         );
  MUX2_X1 U11165 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6963), .S(n9900), .Z(n9901)
         );
  NAND3_X1 U11166 ( .A1(n9903), .A2(n9902), .A3(n9901), .ZN(n9904) );
  NAND3_X1 U11167 ( .A1(n9990), .A2(n9910), .A3(n9904), .ZN(n9905) );
  NAND3_X1 U11168 ( .A1(n9907), .A2(n9906), .A3(n9905), .ZN(P1_U3249) );
  NAND3_X1 U11169 ( .A1(n9910), .A2(n9909), .A3(n9908), .ZN(n9911) );
  NAND3_X1 U11170 ( .A1(n9990), .A2(n9912), .A3(n9911), .ZN(n9922) );
  INV_X1 U11171 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9914) );
  OAI21_X1 U11172 ( .B1(n9994), .B2(n9914), .A(n9913), .ZN(n9915) );
  AOI21_X1 U11173 ( .B1(n9988), .B2(n9916), .A(n9915), .ZN(n9921) );
  OAI211_X1 U11174 ( .C1(n9919), .C2(n9918), .A(n9984), .B(n9917), .ZN(n9920)
         );
  NAND3_X1 U11175 ( .A1(n9922), .A2(n9921), .A3(n9920), .ZN(P1_U3250) );
  XNOR2_X1 U11176 ( .A(n9942), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9926) );
  OAI22_X1 U11177 ( .A1(n9924), .A2(n10226), .B1(n9923), .B2(n9928), .ZN(n9925) );
  NOR2_X1 U11178 ( .A1(n9925), .A2(n9926), .ZN(n9944) );
  AOI21_X1 U11179 ( .B1(n9926), .B2(n9925), .A(n9944), .ZN(n9940) );
  OAI21_X1 U11180 ( .B1(n9929), .B2(n9928), .A(n9927), .ZN(n9930) );
  INV_X1 U11181 ( .A(n9930), .ZN(n9933) );
  NAND2_X1 U11182 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9942), .ZN(n9931) );
  OAI21_X1 U11183 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9942), .A(n9931), .ZN(
        n9932) );
  AOI211_X1 U11184 ( .C1(n9933), .C2(n9932), .A(n9941), .B(n9960), .ZN(n9934)
         );
  INV_X1 U11185 ( .A(n9934), .ZN(n9938) );
  AND2_X1 U11186 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9936) );
  NOR2_X1 U11187 ( .A1(n9975), .A2(n9945), .ZN(n9935) );
  AOI211_X1 U11188 ( .C1(n9965), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9936), .B(
        n9935), .ZN(n9937) );
  OAI211_X1 U11189 ( .C1(n9940), .C2(n9939), .A(n9938), .B(n9937), .ZN(
        P1_U3259) );
  INV_X1 U11190 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10119) );
  XNOR2_X1 U11191 ( .A(n9943), .B(n10119), .ZN(n9955) );
  XOR2_X1 U11192 ( .A(n9955), .B(n9956), .Z(n9954) );
  INV_X1 U11193 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n10216) );
  XNOR2_X1 U11194 ( .A(n9943), .B(n10216), .ZN(n9948) );
  AOI21_X1 U11195 ( .B1(n9945), .B2(n10221), .A(n9944), .ZN(n9946) );
  INV_X1 U11196 ( .A(n9946), .ZN(n9947) );
  NAND2_X1 U11197 ( .A1(n9948), .A2(n9947), .ZN(n9968) );
  OAI21_X1 U11198 ( .B1(n9948), .B2(n9947), .A(n9968), .ZN(n9952) );
  NAND2_X1 U11199 ( .A1(n9965), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9949) );
  OAI211_X1 U11200 ( .C1(n9975), .C2(n9966), .A(n9950), .B(n9949), .ZN(n9951)
         );
  AOI21_X1 U11201 ( .B1(n9990), .B2(n9952), .A(n9951), .ZN(n9953) );
  OAI21_X1 U11202 ( .B1(n9954), .B2(n9960), .A(n9953), .ZN(P1_U3260) );
  INV_X1 U11203 ( .A(n9979), .ZN(n9974) );
  AND2_X1 U11204 ( .A1(n10311), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11205 ( .A1(n9956), .A2(n9955), .ZN(n9958) );
  NAND2_X1 U11206 ( .A1(n9966), .A2(n10119), .ZN(n9957) );
  NAND2_X1 U11207 ( .A1(n9958), .A2(n9957), .ZN(n9962) );
  INV_X1 U11208 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9959) );
  MUX2_X1 U11209 ( .A(n9959), .B(P1_REG2_REG_18__SCAN_IN), .S(n9979), .Z(n9961) );
  NOR2_X1 U11210 ( .A1(n9962), .A2(n9961), .ZN(n9977) );
  AOI211_X1 U11211 ( .C1(n9962), .C2(n9961), .A(n9977), .B(n9960), .ZN(n9963)
         );
  AOI211_X1 U11212 ( .C1(n9965), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9964), .B(
        n9963), .ZN(n9973) );
  NAND2_X1 U11213 ( .A1(n9966), .A2(n10216), .ZN(n9967) );
  NAND2_X1 U11214 ( .A1(n9968), .A2(n9967), .ZN(n9970) );
  XNOR2_X1 U11215 ( .A(n9979), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U11216 ( .A1(n9970), .A2(n9969), .ZN(n9971) );
  NAND3_X1 U11217 ( .A1(n9990), .A2(n9981), .A3(n9971), .ZN(n9972) );
  OAI211_X1 U11218 ( .C1(n9975), .C2(n9974), .A(n9973), .B(n9972), .ZN(
        P1_U3261) );
  INV_X1 U11219 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9995) );
  AND2_X1 U11220 ( .A1(n9979), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9976) );
  OR2_X1 U11221 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  INV_X1 U11222 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10089) );
  XNOR2_X1 U11223 ( .A(n9978), .B(n10089), .ZN(n9986) );
  NAND2_X1 U11224 ( .A1(n9979), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9980) );
  NAND2_X1 U11225 ( .A1(n9981), .A2(n9980), .ZN(n9982) );
  XNOR2_X1 U11226 ( .A(n9982), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9989) );
  INV_X1 U11227 ( .A(n9989), .ZN(n9983) );
  NOR3_X1 U11228 ( .A1(n9986), .A2(n6924), .A3(n9985), .ZN(n9987) );
  OAI211_X1 U11229 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(
        P1_U3262) );
  XNOR2_X1 U11230 ( .A(n9997), .B(n10005), .ZN(n9998) );
  AOI21_X1 U11231 ( .B1(n10013), .B2(n10174), .A(n10475), .ZN(n10001) );
  NAND2_X1 U11232 ( .A1(n10173), .A2(n10392), .ZN(n10004) );
  AOI22_X1 U11233 ( .A1(n10002), .A2(n10380), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n7610), .ZN(n10003) );
  OAI211_X1 U11234 ( .C1(n10175), .C2(n10383), .A(n10004), .B(n10003), .ZN(
        n10007) );
  XOR2_X1 U11235 ( .A(n10012), .B(n10011), .Z(n10260) );
  OAI211_X1 U11236 ( .C1(n10014), .C2(n10180), .A(n10390), .B(n10013), .ZN(
        n10178) );
  AOI22_X1 U11237 ( .A1(n10015), .A2(n10380), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n7610), .ZN(n10018) );
  NAND2_X1 U11238 ( .A1(n10016), .A2(n10079), .ZN(n10017) );
  OAI211_X1 U11239 ( .C1(n10178), .C2(n10082), .A(n10018), .B(n10017), .ZN(
        n10019) );
  AOI21_X1 U11240 ( .B1(n10260), .B2(n10393), .A(n10019), .ZN(n10020) );
  OAI21_X1 U11241 ( .B1(n7610), .B2(n10179), .A(n10020), .ZN(P1_U3267) );
  XNOR2_X1 U11242 ( .A(n10022), .B(n10021), .ZN(n10265) );
  AOI211_X1 U11243 ( .C1(n10025), .C2(n10024), .A(n10152), .B(n10023), .ZN(
        n10027) );
  INV_X1 U11244 ( .A(n10028), .ZN(n10029) );
  AOI211_X1 U11245 ( .C1(n6074), .C2(n10037), .A(n10475), .B(n10029), .ZN(
        n10183) );
  NAND2_X1 U11246 ( .A1(n10183), .A2(n10392), .ZN(n10032) );
  AOI22_X1 U11247 ( .A1(n10030), .A2(n10380), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n7610), .ZN(n10031) );
  OAI211_X1 U11248 ( .C1(n10033), .C2(n10383), .A(n10032), .B(n10031), .ZN(
        n10034) );
  AOI21_X1 U11249 ( .B1(n10182), .B2(n10162), .A(n10034), .ZN(n10035) );
  OAI21_X1 U11250 ( .B1(n10265), .B2(n10164), .A(n10035), .ZN(P1_U3269) );
  XOR2_X1 U11251 ( .A(n10036), .B(n10047), .Z(n10269) );
  AOI21_X1 U11252 ( .B1(n7935), .B2(n10188), .A(n10475), .ZN(n10038) );
  AND2_X1 U11253 ( .A1(n10038), .A2(n10037), .ZN(n10187) );
  INV_X1 U11254 ( .A(n10039), .ZN(n10040) );
  AOI22_X1 U11255 ( .A1(n10040), .A2(n10380), .B1(n7610), .B2(
        P1_REG2_REG_23__SCAN_IN), .ZN(n10041) );
  OAI21_X1 U11256 ( .B1(n10042), .B2(n10383), .A(n10041), .ZN(n10043) );
  AOI21_X1 U11257 ( .B1(n10187), .B2(n10392), .A(n10043), .ZN(n10053) );
  INV_X1 U11258 ( .A(n10044), .ZN(n10046) );
  NAND2_X1 U11259 ( .A1(n10046), .A2(n10045), .ZN(n10048) );
  XNOR2_X1 U11260 ( .A(n10048), .B(n10047), .ZN(n10051) );
  INV_X1 U11261 ( .A(n10049), .ZN(n10050) );
  OAI21_X1 U11262 ( .B1(n10051), .B2(n10152), .A(n10050), .ZN(n10186) );
  NAND2_X1 U11263 ( .A1(n10186), .A2(n10162), .ZN(n10052) );
  OAI211_X1 U11264 ( .C1(n10269), .C2(n10164), .A(n10053), .B(n10052), .ZN(
        P1_U3270) );
  XOR2_X1 U11265 ( .A(n10054), .B(n10058), .Z(n10056) );
  OAI21_X1 U11266 ( .B1(n10056), .B2(n10152), .A(n10055), .ZN(n10192) );
  INV_X1 U11267 ( .A(n10192), .ZN(n10068) );
  XOR2_X1 U11268 ( .A(n10057), .B(n10058), .Z(n10273) );
  INV_X1 U11269 ( .A(n10273), .ZN(n10066) );
  OAI21_X1 U11270 ( .B1(n10075), .B2(n10059), .A(n10390), .ZN(n10061) );
  OR2_X1 U11271 ( .A1(n10061), .A2(n10060), .ZN(n10191) );
  AOI22_X1 U11272 ( .A1(n7610), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n10062), 
        .B2(n10380), .ZN(n10064) );
  NAND2_X1 U11273 ( .A1(n10194), .A2(n10079), .ZN(n10063) );
  OAI211_X1 U11274 ( .C1(n10191), .C2(n10082), .A(n10064), .B(n10063), .ZN(
        n10065) );
  AOI21_X1 U11275 ( .B1(n10066), .B2(n10393), .A(n10065), .ZN(n10067) );
  OAI21_X1 U11276 ( .B1(n7610), .B2(n10068), .A(n10067), .ZN(P1_U3272) );
  XNOR2_X1 U11277 ( .A(n10069), .B(n6072), .ZN(n10277) );
  NAND2_X1 U11278 ( .A1(n9710), .A2(n5011), .ZN(n10070) );
  NAND3_X1 U11279 ( .A1(n10071), .A2(n10377), .A3(n10070), .ZN(n10073) );
  NAND2_X1 U11280 ( .A1(n10073), .A2(n10072), .ZN(n10201) );
  NAND2_X1 U11281 ( .A1(n10086), .A2(n10197), .ZN(n10074) );
  NAND2_X1 U11282 ( .A1(n10074), .A2(n10390), .ZN(n10076) );
  OR2_X1 U11283 ( .A1(n10076), .A2(n10075), .ZN(n10199) );
  INV_X1 U11284 ( .A(n10077), .ZN(n10078) );
  AOI22_X1 U11285 ( .A1(n7610), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n10078), 
        .B2(n10380), .ZN(n10081) );
  NAND2_X1 U11286 ( .A1(n10197), .A2(n10079), .ZN(n10080) );
  OAI211_X1 U11287 ( .C1(n10199), .C2(n10082), .A(n10081), .B(n10080), .ZN(
        n10083) );
  AOI21_X1 U11288 ( .B1(n10201), .B2(n10162), .A(n10083), .ZN(n10084) );
  OAI21_X1 U11289 ( .B1(n10277), .B2(n10164), .A(n10084), .ZN(P1_U3273) );
  XNOR2_X1 U11290 ( .A(n10093), .B(n10085), .ZN(n10281) );
  AOI211_X1 U11291 ( .C1(n10206), .C2(n10106), .A(n10475), .B(n6087), .ZN(
        n10205) );
  INV_X1 U11292 ( .A(n10206), .ZN(n10087) );
  NOR2_X1 U11293 ( .A1(n10087), .A2(n10383), .ZN(n10091) );
  OAI22_X1 U11294 ( .A1(n10162), .A2(n10089), .B1(n10088), .B2(n10117), .ZN(
        n10090) );
  AOI211_X1 U11295 ( .C1(n10205), .C2(n10392), .A(n10091), .B(n10090), .ZN(
        n10097) );
  XOR2_X1 U11296 ( .A(n10093), .B(n10092), .Z(n10095) );
  OAI21_X1 U11297 ( .B1(n10095), .B2(n10152), .A(n10094), .ZN(n10204) );
  NAND2_X1 U11298 ( .A1(n10204), .A2(n10162), .ZN(n10096) );
  OAI211_X1 U11299 ( .C1(n10281), .C2(n10164), .A(n10097), .B(n10096), .ZN(
        P1_U3274) );
  XOR2_X1 U11300 ( .A(n10101), .B(n10098), .Z(n10285) );
  NAND2_X1 U11301 ( .A1(n10125), .A2(n10099), .ZN(n10100) );
  XOR2_X1 U11302 ( .A(n10101), .B(n10100), .Z(n10104) );
  INV_X1 U11303 ( .A(n10102), .ZN(n10103) );
  OAI21_X1 U11304 ( .B1(n10104), .B2(n10152), .A(n10103), .ZN(n10209) );
  INV_X1 U11305 ( .A(n10105), .ZN(n10108) );
  INV_X1 U11306 ( .A(n10106), .ZN(n10107) );
  AOI211_X1 U11307 ( .C1(n6067), .C2(n10108), .A(n10475), .B(n10107), .ZN(
        n10210) );
  NAND2_X1 U11308 ( .A1(n10210), .A2(n10392), .ZN(n10111) );
  AOI22_X1 U11309 ( .A1(n7610), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10109), 
        .B2(n10380), .ZN(n10110) );
  OAI211_X1 U11310 ( .C1(n10112), .C2(n10383), .A(n10111), .B(n10110), .ZN(
        n10113) );
  AOI21_X1 U11311 ( .B1(n10162), .B2(n10209), .A(n10113), .ZN(n10114) );
  OAI21_X1 U11312 ( .B1(n10285), .B2(n10164), .A(n10114), .ZN(P1_U3275) );
  XNOR2_X1 U11313 ( .A(n10115), .B(n10123), .ZN(n10289) );
  AOI211_X1 U11314 ( .C1(n10215), .C2(n4459), .A(n10475), .B(n10105), .ZN(
        n10214) );
  NOR2_X1 U11315 ( .A1(n10116), .A2(n10383), .ZN(n10121) );
  OAI22_X1 U11316 ( .A1(n10162), .A2(n10119), .B1(n10118), .B2(n10117), .ZN(
        n10120) );
  AOI211_X1 U11317 ( .C1(n10214), .C2(n10392), .A(n10121), .B(n10120), .ZN(
        n10130) );
  INV_X1 U11318 ( .A(n10122), .ZN(n10134) );
  OAI21_X1 U11319 ( .B1(n10134), .B2(n10124), .A(n10123), .ZN(n10126) );
  NAND3_X1 U11320 ( .A1(n10126), .A2(n10125), .A3(n10377), .ZN(n10128) );
  NAND2_X1 U11321 ( .A1(n10128), .A2(n10127), .ZN(n10213) );
  NAND2_X1 U11322 ( .A1(n10213), .A2(n10162), .ZN(n10129) );
  OAI211_X1 U11323 ( .C1(n10289), .C2(n10164), .A(n10130), .B(n10129), .ZN(
        P1_U3276) );
  OAI21_X1 U11324 ( .B1(n10132), .B2(n10135), .A(n10131), .ZN(n10293) );
  INV_X1 U11325 ( .A(n10133), .ZN(n10136) );
  AOI21_X1 U11326 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(n10138) );
  OAI21_X1 U11327 ( .B1(n10138), .B2(n10152), .A(n10137), .ZN(n10218) );
  AOI21_X1 U11328 ( .B1(n10154), .B2(n10220), .A(n10475), .ZN(n10139) );
  AND2_X1 U11329 ( .A1(n10139), .A2(n4459), .ZN(n10219) );
  NAND2_X1 U11330 ( .A1(n10219), .A2(n10392), .ZN(n10143) );
  INV_X1 U11331 ( .A(n10140), .ZN(n10141) );
  AOI22_X1 U11332 ( .A1(n7610), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n10141), 
        .B2(n10380), .ZN(n10142) );
  OAI211_X1 U11333 ( .C1(n10144), .C2(n10383), .A(n10143), .B(n10142), .ZN(
        n10145) );
  AOI21_X1 U11334 ( .B1(n10218), .B2(n10162), .A(n10145), .ZN(n10146) );
  OAI21_X1 U11335 ( .B1(n10293), .B2(n10164), .A(n10146), .ZN(P1_U3277) );
  XNOR2_X1 U11336 ( .A(n10147), .B(n10149), .ZN(n10297) );
  NAND2_X1 U11337 ( .A1(n7850), .A2(n10148), .ZN(n10150) );
  XNOR2_X1 U11338 ( .A(n10150), .B(n10149), .ZN(n10153) );
  OAI21_X1 U11339 ( .B1(n10153), .B2(n10152), .A(n10151), .ZN(n10223) );
  OR2_X1 U11340 ( .A1(n7853), .A2(n10160), .ZN(n10155) );
  AND3_X1 U11341 ( .A1(n10155), .A2(n10154), .A3(n10390), .ZN(n10224) );
  NAND2_X1 U11342 ( .A1(n10224), .A2(n10392), .ZN(n10159) );
  INV_X1 U11343 ( .A(n10156), .ZN(n10157) );
  AOI22_X1 U11344 ( .A1(n7610), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n10157), 
        .B2(n10380), .ZN(n10158) );
  OAI211_X1 U11345 ( .C1(n10160), .C2(n10383), .A(n10159), .B(n10158), .ZN(
        n10161) );
  AOI21_X1 U11346 ( .B1(n10223), .B2(n10162), .A(n10161), .ZN(n10163) );
  OAI21_X1 U11347 ( .B1(n10297), .B2(n10164), .A(n10163), .ZN(P1_U3278) );
  MUX2_X1 U11348 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10255), .S(n10494), .Z(
        P1_U3553) );
  INV_X1 U11349 ( .A(n10169), .ZN(n10170) );
  MUX2_X1 U11350 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10256), .S(n10494), .Z(
        P1_U3552) );
  INV_X1 U11351 ( .A(n10480), .ZN(n10249) );
  INV_X1 U11352 ( .A(n10173), .ZN(n10176) );
  INV_X1 U11353 ( .A(n10174), .ZN(n10175) );
  MUX2_X1 U11354 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10257), .S(n10494), .Z(
        P1_U3549) );
  INV_X1 U11355 ( .A(n10243), .ZN(n10181) );
  AOI211_X1 U11356 ( .C1(n6090), .C2(n6074), .A(n10183), .B(n10182), .ZN(
        n10262) );
  MUX2_X1 U11357 ( .A(n10184), .B(n10262), .S(n10494), .Z(n10185) );
  OAI21_X1 U11358 ( .B1(n10265), .B2(n10243), .A(n10185), .ZN(P1_U3546) );
  AOI211_X1 U11359 ( .C1(n6090), .C2(n10188), .A(n10187), .B(n10186), .ZN(
        n10266) );
  MUX2_X1 U11360 ( .A(n10189), .B(n10266), .S(n10494), .Z(n10190) );
  OAI21_X1 U11361 ( .B1(n10269), .B2(n10243), .A(n10190), .ZN(P1_U3545) );
  INV_X1 U11362 ( .A(n10191), .ZN(n10193) );
  AOI211_X1 U11363 ( .C1(n6090), .C2(n10194), .A(n10193), .B(n10192), .ZN(
        n10270) );
  MUX2_X1 U11364 ( .A(n10195), .B(n10270), .S(n10494), .Z(n10196) );
  OAI21_X1 U11365 ( .B1(n10273), .B2(n10243), .A(n10196), .ZN(P1_U3543) );
  INV_X1 U11366 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10202) );
  NAND2_X1 U11367 ( .A1(n10197), .A2(n6090), .ZN(n10198) );
  NAND2_X1 U11368 ( .A1(n10199), .A2(n10198), .ZN(n10200) );
  NOR2_X1 U11369 ( .A1(n10201), .A2(n10200), .ZN(n10274) );
  MUX2_X1 U11370 ( .A(n10202), .B(n10274), .S(n10494), .Z(n10203) );
  OAI21_X1 U11371 ( .B1(n10277), .B2(n10243), .A(n10203), .ZN(P1_U3542) );
  AOI211_X1 U11372 ( .C1(n6090), .C2(n10206), .A(n10205), .B(n10204), .ZN(
        n10278) );
  MUX2_X1 U11373 ( .A(n10207), .B(n10278), .S(n10494), .Z(n10208) );
  OAI21_X1 U11374 ( .B1(n10281), .B2(n10243), .A(n10208), .ZN(P1_U3541) );
  AOI211_X1 U11375 ( .C1(n6090), .C2(n6067), .A(n10210), .B(n10209), .ZN(
        n10282) );
  MUX2_X1 U11376 ( .A(n10211), .B(n10282), .S(n10494), .Z(n10212) );
  OAI21_X1 U11377 ( .B1(n10285), .B2(n10243), .A(n10212), .ZN(P1_U3540) );
  AOI211_X1 U11378 ( .C1(n6090), .C2(n10215), .A(n10214), .B(n10213), .ZN(
        n10286) );
  MUX2_X1 U11379 ( .A(n10216), .B(n10286), .S(n10494), .Z(n10217) );
  OAI21_X1 U11380 ( .B1(n10289), .B2(n10243), .A(n10217), .ZN(P1_U3539) );
  AOI211_X1 U11381 ( .C1(n6090), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10290) );
  MUX2_X1 U11382 ( .A(n10221), .B(n10290), .S(n10494), .Z(n10222) );
  OAI21_X1 U11383 ( .B1(n10243), .B2(n10293), .A(n10222), .ZN(P1_U3538) );
  AOI211_X1 U11384 ( .C1(n6090), .C2(n10225), .A(n10224), .B(n10223), .ZN(
        n10294) );
  MUX2_X1 U11385 ( .A(n10226), .B(n10294), .S(n10494), .Z(n10227) );
  OAI21_X1 U11386 ( .B1(n10243), .B2(n10297), .A(n10227), .ZN(P1_U3537) );
  AOI211_X1 U11387 ( .C1(n6090), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10231) );
  OAI21_X1 U11388 ( .B1(n10232), .B2(n10249), .A(n10231), .ZN(n10298) );
  MUX2_X1 U11389 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10298), .S(n10494), .Z(
        P1_U3536) );
  AOI211_X1 U11390 ( .C1(n6090), .C2(n10235), .A(n10234), .B(n10233), .ZN(
        n10299) );
  MUX2_X1 U11391 ( .A(n10236), .B(n10299), .S(n10494), .Z(n10237) );
  OAI21_X1 U11392 ( .B1(n10302), .B2(n10243), .A(n10237), .ZN(P1_U3535) );
  AOI211_X1 U11393 ( .C1(n6090), .C2(n10240), .A(n10239), .B(n10238), .ZN(
        n10303) );
  MUX2_X1 U11394 ( .A(n10241), .B(n10303), .S(n10494), .Z(n10242) );
  OAI21_X1 U11395 ( .B1(n10307), .B2(n10243), .A(n10242), .ZN(P1_U3534) );
  AOI21_X1 U11396 ( .B1(n6090), .B2(n10245), .A(n10244), .ZN(n10246) );
  OAI211_X1 U11397 ( .C1(n10249), .C2(n10248), .A(n10247), .B(n10246), .ZN(
        n10308) );
  MUX2_X1 U11398 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10308), .S(n10494), .Z(
        P1_U3530) );
  OAI21_X1 U11399 ( .B1(n10480), .B2(n10377), .A(n10250), .ZN(n10252) );
  OAI211_X1 U11400 ( .C1(n10254), .C2(n10253), .A(n10252), .B(n10251), .ZN(
        n10309) );
  MUX2_X1 U11401 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10309), .S(n10494), .Z(
        P1_U3522) );
  MUX2_X1 U11402 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10256), .S(n10482), .Z(
        P1_U3520) );
  MUX2_X1 U11403 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10257), .S(n10482), .Z(
        P1_U3517) );
  MUX2_X1 U11404 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10258), .S(n10482), .Z(
        n10259) );
  AOI21_X1 U11405 ( .B1(n10260), .B2(n6050), .A(n10259), .ZN(n10261) );
  INV_X1 U11406 ( .A(n10261), .ZN(P1_U3516) );
  INV_X1 U11407 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10263) );
  MUX2_X1 U11408 ( .A(n10263), .B(n10262), .S(n10482), .Z(n10264) );
  OAI21_X1 U11409 ( .B1(n10265), .B2(n10306), .A(n10264), .ZN(P1_U3514) );
  INV_X1 U11410 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10267) );
  MUX2_X1 U11411 ( .A(n10267), .B(n10266), .S(n10482), .Z(n10268) );
  OAI21_X1 U11412 ( .B1(n10269), .B2(n10306), .A(n10268), .ZN(P1_U3513) );
  INV_X1 U11413 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10271) );
  MUX2_X1 U11414 ( .A(n10271), .B(n10270), .S(n10482), .Z(n10272) );
  OAI21_X1 U11415 ( .B1(n10273), .B2(n10306), .A(n10272), .ZN(P1_U3511) );
  MUX2_X1 U11416 ( .A(n10275), .B(n10274), .S(n10482), .Z(n10276) );
  OAI21_X1 U11417 ( .B1(n10277), .B2(n10306), .A(n10276), .ZN(P1_U3510) );
  INV_X1 U11418 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10279) );
  MUX2_X1 U11419 ( .A(n10279), .B(n10278), .S(n10482), .Z(n10280) );
  OAI21_X1 U11420 ( .B1(n10281), .B2(n10306), .A(n10280), .ZN(P1_U3509) );
  INV_X1 U11421 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10283) );
  MUX2_X1 U11422 ( .A(n10283), .B(n10282), .S(n10482), .Z(n10284) );
  OAI21_X1 U11423 ( .B1(n10285), .B2(n10306), .A(n10284), .ZN(P1_U3507) );
  INV_X1 U11424 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10287) );
  MUX2_X1 U11425 ( .A(n10287), .B(n10286), .S(n10482), .Z(n10288) );
  OAI21_X1 U11426 ( .B1(n10289), .B2(n10306), .A(n10288), .ZN(P1_U3504) );
  INV_X1 U11427 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10291) );
  MUX2_X1 U11428 ( .A(n10291), .B(n10290), .S(n10482), .Z(n10292) );
  OAI21_X1 U11429 ( .B1(n10293), .B2(n10306), .A(n10292), .ZN(P1_U3501) );
  MUX2_X1 U11430 ( .A(n10295), .B(n10294), .S(n10482), .Z(n10296) );
  OAI21_X1 U11431 ( .B1(n10297), .B2(n10306), .A(n10296), .ZN(P1_U3498) );
  MUX2_X1 U11432 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10298), .S(n10482), .Z(
        P1_U3495) );
  MUX2_X1 U11433 ( .A(n10300), .B(n10299), .S(n10482), .Z(n10301) );
  OAI21_X1 U11434 ( .B1(n10302), .B2(n10306), .A(n10301), .ZN(P1_U3492) );
  INV_X1 U11435 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10304) );
  MUX2_X1 U11436 ( .A(n10304), .B(n10303), .S(n10482), .Z(n10305) );
  OAI21_X1 U11437 ( .B1(n10307), .B2(n10306), .A(n10305), .ZN(P1_U3489) );
  MUX2_X1 U11438 ( .A(P1_REG0_REG_8__SCAN_IN), .B(n10308), .S(n10482), .Z(
        P1_U3477) );
  MUX2_X1 U11439 ( .A(P1_REG0_REG_0__SCAN_IN), .B(n10309), .S(n10482), .Z(
        P1_U3453) );
  INV_X1 U11440 ( .A(n10310), .ZN(n10313) );
  NOR4_X1 U11441 ( .A1(n10313), .A2(P1_IR_REG_30__SCAN_IN), .A3(n10312), .A4(
        n10311), .ZN(n10314) );
  AOI21_X1 U11442 ( .B1(n10315), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10314), 
        .ZN(n10316) );
  OAI21_X1 U11443 ( .B1(n10317), .B2(n10335), .A(n10316), .ZN(P1_U3324) );
  OAI222_X1 U11444 ( .A1(n10332), .A2(n10320), .B1(n10335), .B2(n10319), .C1(
        n10318), .C2(P1_U3086), .ZN(P1_U3325) );
  OAI222_X1 U11445 ( .A1(n10332), .A2(n10323), .B1(P1_U3086), .B2(n10322), 
        .C1(n10335), .C2(n10321), .ZN(P1_U3326) );
  OAI222_X1 U11446 ( .A1(n10328), .A2(P1_U3086), .B1(n10335), .B2(n10327), 
        .C1(n10326), .C2(n10332), .ZN(P1_U3329) );
  OAI222_X1 U11447 ( .A1(n10331), .A2(n10311), .B1(n10335), .B2(n10330), .C1(
        n10329), .C2(n10332), .ZN(P1_U3330) );
  OAI222_X1 U11448 ( .A1(n10336), .A2(P1_U3086), .B1(n10335), .B2(n10334), 
        .C1(n10333), .C2(n10332), .ZN(P1_U3331) );
  MUX2_X1 U11449 ( .A(n10337), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XOR2_X1 U11450 ( .A(n10338), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  NAND2_X1 U11451 ( .A1(n9743), .A2(n10339), .ZN(n10340) );
  XNOR2_X1 U11452 ( .A(n10340), .B(n5224), .ZN(n10342) );
  AOI21_X1 U11453 ( .B1(n10342), .B2(n10377), .A(n10341), .ZN(n10468) );
  INV_X1 U11454 ( .A(n10343), .ZN(n10344) );
  AOI22_X1 U11455 ( .A1(n7610), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n10344), 
        .B2(n10380), .ZN(n10345) );
  OAI21_X1 U11456 ( .B1(n10383), .B2(n10469), .A(n10345), .ZN(n10346) );
  INV_X1 U11457 ( .A(n10346), .ZN(n10354) );
  XNOR2_X1 U11458 ( .A(n10348), .B(n10347), .ZN(n10471) );
  INV_X1 U11459 ( .A(n10349), .ZN(n10350) );
  OAI211_X1 U11460 ( .C1(n10469), .C2(n10351), .A(n10350), .B(n10390), .ZN(
        n10467) );
  INV_X1 U11461 ( .A(n10467), .ZN(n10352) );
  AOI22_X1 U11462 ( .A1(n10471), .A2(n10393), .B1(n10392), .B2(n10352), .ZN(
        n10353) );
  OAI211_X1 U11463 ( .C1(n7610), .C2(n10468), .A(n10354), .B(n10353), .ZN(
        P1_U3283) );
  XNOR2_X1 U11464 ( .A(n10355), .B(n10356), .ZN(n10359) );
  INV_X1 U11465 ( .A(n10357), .ZN(n10358) );
  AOI21_X1 U11466 ( .B1(n10359), .B2(n10377), .A(n10358), .ZN(n10446) );
  INV_X1 U11467 ( .A(n10360), .ZN(n10361) );
  AOI22_X1 U11468 ( .A1(n7610), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n10361), .B2(
        n10380), .ZN(n10362) );
  OAI21_X1 U11469 ( .B1(n10383), .B2(n10445), .A(n10362), .ZN(n10363) );
  INV_X1 U11470 ( .A(n10363), .ZN(n10373) );
  AOI21_X1 U11471 ( .B1(n7803), .B2(n7798), .A(n10364), .ZN(n10366) );
  XNOR2_X1 U11472 ( .A(n10366), .B(n10365), .ZN(n10449) );
  INV_X1 U11473 ( .A(n10367), .ZN(n10370) );
  INV_X1 U11474 ( .A(n10368), .ZN(n10369) );
  OAI211_X1 U11475 ( .C1(n10445), .C2(n10370), .A(n10369), .B(n10390), .ZN(
        n10444) );
  INV_X1 U11476 ( .A(n10444), .ZN(n10371) );
  AOI22_X1 U11477 ( .A1(n10449), .A2(n10393), .B1(n10371), .B2(n10392), .ZN(
        n10372) );
  OAI211_X1 U11478 ( .C1(n7610), .C2(n10446), .A(n10373), .B(n10372), .ZN(
        P1_U3287) );
  XNOR2_X1 U11479 ( .A(n10374), .B(n9672), .ZN(n10378) );
  INV_X1 U11480 ( .A(n10375), .ZN(n10376) );
  AOI21_X1 U11481 ( .B1(n10378), .B2(n10377), .A(n10376), .ZN(n10433) );
  INV_X1 U11482 ( .A(n10379), .ZN(n10381) );
  AOI22_X1 U11483 ( .A1(n7610), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n10381), .B2(
        n10380), .ZN(n10382) );
  OAI21_X1 U11484 ( .B1(n10383), .B2(n10432), .A(n10382), .ZN(n10384) );
  INV_X1 U11485 ( .A(n10384), .ZN(n10395) );
  AOI21_X1 U11486 ( .B1(n7637), .B2(n10386), .A(n10385), .ZN(n10388) );
  XNOR2_X1 U11487 ( .A(n10388), .B(n10387), .ZN(n10436) );
  OAI211_X1 U11488 ( .C1(n4797), .C2(n10432), .A(n10390), .B(n10389), .ZN(
        n10431) );
  INV_X1 U11489 ( .A(n10431), .ZN(n10391) );
  AOI22_X1 U11490 ( .A1(n10436), .A2(n10393), .B1(n10392), .B2(n10391), .ZN(
        n10394) );
  OAI211_X1 U11491 ( .C1(n7610), .C2(n10433), .A(n10395), .B(n10394), .ZN(
        P1_U3289) );
  AND2_X1 U11492 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10406), .ZN(P1_U3294) );
  NOR2_X1 U11493 ( .A1(n10405), .A2(n10396), .ZN(P1_U3295) );
  AND2_X1 U11494 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10406), .ZN(P1_U3296) );
  AND2_X1 U11495 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10406), .ZN(P1_U3297) );
  AND2_X1 U11496 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10406), .ZN(P1_U3298) );
  AND2_X1 U11497 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10406), .ZN(P1_U3299) );
  NOR2_X1 U11498 ( .A1(n10405), .A2(n10397), .ZN(P1_U3300) );
  NOR2_X1 U11499 ( .A1(n10405), .A2(n10398), .ZN(P1_U3301) );
  AND2_X1 U11500 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10406), .ZN(P1_U3302) );
  AND2_X1 U11501 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10406), .ZN(P1_U3303) );
  NOR2_X1 U11502 ( .A1(n10405), .A2(n10399), .ZN(P1_U3304) );
  NOR2_X1 U11503 ( .A1(n10405), .A2(n10400), .ZN(P1_U3305) );
  AND2_X1 U11504 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10406), .ZN(P1_U3306) );
  AND2_X1 U11505 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10406), .ZN(P1_U3307) );
  AND2_X1 U11506 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10406), .ZN(P1_U3308) );
  AND2_X1 U11507 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10406), .ZN(P1_U3309) );
  AND2_X1 U11508 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10406), .ZN(P1_U3310) );
  AND2_X1 U11509 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10406), .ZN(P1_U3311) );
  NOR2_X1 U11510 ( .A1(n10405), .A2(n10401), .ZN(P1_U3312) );
  AND2_X1 U11511 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10406), .ZN(P1_U3313) );
  AND2_X1 U11512 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10406), .ZN(P1_U3314) );
  AND2_X1 U11513 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10406), .ZN(P1_U3315) );
  AND2_X1 U11514 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10406), .ZN(P1_U3316) );
  NOR2_X1 U11515 ( .A1(n10405), .A2(n10402), .ZN(P1_U3317) );
  AND2_X1 U11516 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10406), .ZN(P1_U3318) );
  NOR2_X1 U11517 ( .A1(n10405), .A2(n10403), .ZN(P1_U3319) );
  AND2_X1 U11518 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10406), .ZN(P1_U3320) );
  NOR2_X1 U11519 ( .A1(n10405), .A2(n10404), .ZN(P1_U3321) );
  AND2_X1 U11520 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10406), .ZN(P1_U3322) );
  AND2_X1 U11521 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10406), .ZN(P1_U3323) );
  OAI21_X1 U11522 ( .B1(n10409), .B2(n10408), .A(n10407), .ZN(P1_U3439) );
  INV_X1 U11523 ( .A(n10410), .ZN(n10460) );
  INV_X1 U11524 ( .A(n10411), .ZN(n10417) );
  NOR2_X1 U11525 ( .A1(n10411), .A2(n10451), .ZN(n10416) );
  OAI211_X1 U11526 ( .C1(n10414), .C2(n10473), .A(n10413), .B(n10412), .ZN(
        n10415) );
  AOI211_X1 U11527 ( .C1(n10460), .C2(n10417), .A(n10416), .B(n10415), .ZN(
        n10483) );
  AOI22_X1 U11528 ( .A1(n10482), .A2(n10483), .B1(n10418), .B2(n10481), .ZN(
        P1_U3456) );
  OAI211_X1 U11529 ( .C1(n10421), .C2(n10473), .A(n10420), .B(n10419), .ZN(
        n10422) );
  AOI21_X1 U11530 ( .B1(n10423), .B2(n10480), .A(n10422), .ZN(n10484) );
  INV_X1 U11531 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10424) );
  AOI22_X1 U11532 ( .A1(n10482), .A2(n10484), .B1(n10424), .B2(n10481), .ZN(
        P1_U3459) );
  OAI21_X1 U11533 ( .B1(n10426), .B2(n10473), .A(n10425), .ZN(n10429) );
  INV_X1 U11534 ( .A(n10427), .ZN(n10428) );
  AOI211_X1 U11535 ( .C1(n10480), .C2(n10430), .A(n10429), .B(n10428), .ZN(
        n10485) );
  AOI22_X1 U11536 ( .A1(n10482), .A2(n10485), .B1(n5485), .B2(n10481), .ZN(
        P1_U3462) );
  OAI21_X1 U11537 ( .B1(n10432), .B2(n10473), .A(n10431), .ZN(n10435) );
  INV_X1 U11538 ( .A(n10433), .ZN(n10434) );
  AOI211_X1 U11539 ( .C1(n10480), .C2(n10436), .A(n10435), .B(n10434), .ZN(
        n10486) );
  INV_X1 U11540 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U11541 ( .A1(n10482), .A2(n10486), .B1(n10437), .B2(n10481), .ZN(
        P1_U3465) );
  OAI21_X1 U11542 ( .B1(n10439), .B2(n10473), .A(n10438), .ZN(n10441) );
  AOI211_X1 U11543 ( .C1(n10480), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10487) );
  INV_X1 U11544 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U11545 ( .A1(n10482), .A2(n10487), .B1(n10443), .B2(n10481), .ZN(
        P1_U3468) );
  OAI21_X1 U11546 ( .B1(n10445), .B2(n10473), .A(n10444), .ZN(n10448) );
  INV_X1 U11547 ( .A(n10446), .ZN(n10447) );
  AOI211_X1 U11548 ( .C1(n10480), .C2(n10449), .A(n10448), .B(n10447), .ZN(
        n10488) );
  INV_X1 U11549 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U11550 ( .A1(n10482), .A2(n10488), .B1(n10450), .B2(n10481), .ZN(
        P1_U3471) );
  INV_X1 U11551 ( .A(n10451), .ZN(n10452) );
  NAND2_X1 U11552 ( .A1(n10459), .A2(n10452), .ZN(n10454) );
  OAI211_X1 U11553 ( .C1(n10455), .C2(n10473), .A(n10454), .B(n10453), .ZN(
        n10458) );
  INV_X1 U11554 ( .A(n10456), .ZN(n10457) );
  AOI211_X1 U11555 ( .C1(n10460), .C2(n10459), .A(n10458), .B(n10457), .ZN(
        n10489) );
  AOI22_X1 U11556 ( .A1(n10482), .A2(n10489), .B1(n5577), .B2(n10481), .ZN(
        P1_U3474) );
  OAI21_X1 U11557 ( .B1(n10462), .B2(n10473), .A(n10461), .ZN(n10464) );
  AOI211_X1 U11558 ( .C1(n10480), .C2(n10465), .A(n10464), .B(n10463), .ZN(
        n10490) );
  INV_X1 U11559 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U11560 ( .A1(n10482), .A2(n10490), .B1(n10466), .B2(n10481), .ZN(
        P1_U3480) );
  OAI211_X1 U11561 ( .C1(n10469), .C2(n10473), .A(n10468), .B(n10467), .ZN(
        n10470) );
  AOI21_X1 U11562 ( .B1(n10480), .B2(n10471), .A(n10470), .ZN(n10491) );
  INV_X1 U11563 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U11564 ( .A1(n10482), .A2(n10491), .B1(n10472), .B2(n10481), .ZN(
        P1_U3483) );
  OAI22_X1 U11565 ( .A1(n10476), .A2(n10475), .B1(n10474), .B2(n10473), .ZN(
        n10478) );
  AOI211_X1 U11566 ( .C1(n10480), .C2(n10479), .A(n10478), .B(n10477), .ZN(
        n10493) );
  AOI22_X1 U11567 ( .A1(n10482), .A2(n10493), .B1(n5664), .B2(n10481), .ZN(
        P1_U3486) );
  AOI22_X1 U11568 ( .A1(n10494), .A2(n10483), .B1(n6950), .B2(n10492), .ZN(
        P1_U3523) );
  AOI22_X1 U11569 ( .A1(n10494), .A2(n10484), .B1(n6949), .B2(n10492), .ZN(
        P1_U3524) );
  AOI22_X1 U11570 ( .A1(n10494), .A2(n10485), .B1(n6954), .B2(n10492), .ZN(
        P1_U3525) );
  AOI22_X1 U11571 ( .A1(n10494), .A2(n10486), .B1(n6955), .B2(n10492), .ZN(
        P1_U3526) );
  AOI22_X1 U11572 ( .A1(n10494), .A2(n10487), .B1(n6958), .B2(n10492), .ZN(
        P1_U3527) );
  AOI22_X1 U11573 ( .A1(n10494), .A2(n10488), .B1(n6963), .B2(n10492), .ZN(
        P1_U3528) );
  AOI22_X1 U11574 ( .A1(n10494), .A2(n10489), .B1(n5571), .B2(n10492), .ZN(
        P1_U3529) );
  AOI22_X1 U11575 ( .A1(n10494), .A2(n10490), .B1(n7003), .B2(n10492), .ZN(
        P1_U3531) );
  AOI22_X1 U11576 ( .A1(n10494), .A2(n10491), .B1(n5646), .B2(n10492), .ZN(
        P1_U3532) );
  AOI22_X1 U11577 ( .A1(n10494), .A2(n10493), .B1(n5668), .B2(n10492), .ZN(
        P1_U3533) );
  AOI21_X1 U11578 ( .B1(n10496), .B2(n10495), .A(n4573), .ZN(n10502) );
  XNOR2_X1 U11579 ( .A(n10497), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n10498) );
  NAND2_X1 U11580 ( .A1(n10499), .A2(n10498), .ZN(n10501) );
  OAI211_X1 U11581 ( .C1(n10503), .C2(n10502), .A(n10501), .B(n10500), .ZN(
        n10504) );
  AOI21_X1 U11582 ( .B1(n10506), .B2(n10505), .A(n10504), .ZN(n10515) );
  AOI21_X1 U11583 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(n10511) );
  NOR2_X1 U11584 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  AOI21_X1 U11585 ( .B1(n10513), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n10512), .ZN(
        n10514) );
  NAND2_X1 U11586 ( .A1(n10515), .A2(n10514), .ZN(P2_U3185) );
  AOI22_X1 U11587 ( .A1(n10518), .A2(P2_REG3_REG_2__SCAN_IN), .B1(n10517), 
        .B2(n10516), .ZN(n10522) );
  AOI22_X1 U11588 ( .A1(n10520), .A2(n10519), .B1(P2_REG2_REG_2__SCAN_IN), 
        .B2(n8981), .ZN(n10521) );
  OAI221_X1 U11589 ( .B1(n8981), .B2(n10523), .C1(n8981), .C2(n10522), .A(
        n10521), .ZN(P2_U3231) );
  INV_X1 U11590 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10529) );
  INV_X1 U11591 ( .A(n10524), .ZN(n10528) );
  OAI22_X1 U11592 ( .A1(n10526), .A2(n10525), .B1(n6803), .B2(n10537), .ZN(
        n10527) );
  NOR2_X1 U11593 ( .A1(n10528), .A2(n10527), .ZN(n10551) );
  AOI22_X1 U11594 ( .A1(n10550), .A2(n10529), .B1(n10551), .B2(n10548), .ZN(
        P2_U3393) );
  INV_X1 U11595 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U11596 ( .A1(n10550), .A2(n10531), .B1(n10530), .B2(n10548), .ZN(
        P2_U3396) );
  OAI21_X1 U11597 ( .B1(n10533), .B2(n10537), .A(n10532), .ZN(n10534) );
  AOI21_X1 U11598 ( .B1(n10535), .B2(n10544), .A(n10534), .ZN(n10553) );
  AOI22_X1 U11599 ( .A1(n10550), .A2(n6261), .B1(n10553), .B2(n10548), .ZN(
        P2_U3399) );
  INV_X1 U11600 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10541) );
  OAI21_X1 U11601 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(n10539) );
  AOI21_X1 U11602 ( .B1(n10540), .B2(n10544), .A(n10539), .ZN(n10555) );
  AOI22_X1 U11603 ( .A1(n10550), .A2(n10541), .B1(n10555), .B2(n10548), .ZN(
        P2_U3402) );
  INV_X1 U11604 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U11605 ( .A1(n10545), .A2(n10544), .B1(n10543), .B2(n10542), .ZN(
        n10546) );
  AND2_X1 U11606 ( .A1(n10547), .A2(n10546), .ZN(n10556) );
  AOI22_X1 U11607 ( .A1(n10550), .A2(n10549), .B1(n10556), .B2(n10548), .ZN(
        P2_U3405) );
  AOI22_X1 U11608 ( .A1(n10557), .A2(n10551), .B1(n7174), .B2(n6883), .ZN(
        P2_U3460) );
  AOI22_X1 U11609 ( .A1(n10557), .A2(n10553), .B1(n10552), .B2(n6883), .ZN(
        P2_U3462) );
  AOI22_X1 U11610 ( .A1(n10557), .A2(n10555), .B1(n10554), .B2(n6883), .ZN(
        P2_U3463) );
  AOI22_X1 U11611 ( .A1(n10557), .A2(n10556), .B1(n7270), .B2(n6883), .ZN(
        P2_U3464) );
  OAI222_X1 U11612 ( .A1(n10562), .A2(n10561), .B1(n10562), .B2(n10560), .C1(
        n10559), .C2(n10558), .ZN(ADD_1068_U5) );
  XOR2_X1 U11613 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11614 ( .B1(n10565), .B2(n10564), .A(n10563), .ZN(n10566) );
  XNOR2_X1 U11615 ( .A(n10566), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11616 ( .B1(n10569), .B2(n10568), .A(n10567), .ZN(ADD_1068_U56) );
  OAI21_X1 U11617 ( .B1(n10572), .B2(n10571), .A(n10570), .ZN(ADD_1068_U57) );
  OAI21_X1 U11618 ( .B1(n10575), .B2(n10574), .A(n10573), .ZN(ADD_1068_U58) );
  OAI21_X1 U11619 ( .B1(n10578), .B2(n10577), .A(n10576), .ZN(ADD_1068_U59) );
  OAI21_X1 U11620 ( .B1(n10581), .B2(n10580), .A(n10579), .ZN(ADD_1068_U60) );
  AOI22_X1 U11621 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .B1(n10583), .B2(n10582), .ZN(n10586) );
  OAI21_X1 U11622 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(ADD_1068_U61) );
  OAI21_X1 U11623 ( .B1(n10589), .B2(n10588), .A(n10587), .ZN(ADD_1068_U62) );
  OAI21_X1 U11624 ( .B1(n10592), .B2(n10591), .A(n10590), .ZN(ADD_1068_U63) );
  OAI21_X1 U11625 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(ADD_1068_U50) );
  OAI21_X1 U11626 ( .B1(n10598), .B2(n10597), .A(n10596), .ZN(ADD_1068_U51) );
  OAI21_X1 U11627 ( .B1(n10601), .B2(n10600), .A(n10599), .ZN(ADD_1068_U47) );
  OAI21_X1 U11628 ( .B1(n10604), .B2(n10603), .A(n10602), .ZN(ADD_1068_U49) );
  OAI21_X1 U11629 ( .B1(n10607), .B2(n10606), .A(n10605), .ZN(ADD_1068_U48) );
  AOI21_X1 U11630 ( .B1(n10610), .B2(n10609), .A(n10608), .ZN(ADD_1068_U54) );
  AOI21_X1 U11631 ( .B1(n10613), .B2(n10612), .A(n10611), .ZN(ADD_1068_U53) );
  OAI21_X1 U11632 ( .B1(n10616), .B2(n10615), .A(n10614), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4947 ( .A(n6454), .Z(n4776) );
  OR2_X2 U4952 ( .A1(n8026), .A2(n7668), .ZN(n9591) );
  NOR2_X1 U4953 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5513) );
  AOI21_X1 U4967 ( .B1(n7132), .B2(n5637), .A(n5018), .ZN(n8066) );
  CLKBUF_X1 U4993 ( .A(n5449), .Z(n4431) );
  AND2_X1 U5309 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n7743) );
endmodule

