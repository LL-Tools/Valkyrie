

module b21_C_gen_AntiSAT_k_128_5 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2, 
        keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7, 
        keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12, 
        keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17, 
        keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22, 
        keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27, 
        keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32, 
        keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37, 
        keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42, 
        keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47, 
        keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52, 
        keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57, 
        keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62, 
        keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, 
        keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, 
        keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, 
        keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, 
        keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, 
        keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, 
        keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, 
        keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, 
        keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, 
        keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, 
        keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, 
        keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, 
        keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167;

  NAND2_X1 U4816 ( .A1(n4429), .A2(n5195), .ZN(n5217) );
  INV_X2 U4817 ( .A(n5090), .ZN(n5100) );
  INV_X1 U4818 ( .A(n5505), .ZN(n5300) );
  CLKBUF_X1 U4820 ( .A(n5811), .Z(n6456) );
  AND3_X1 U4821 ( .A1(n5843), .A2(n5842), .A3(n5841), .ZN(n7089) );
  CLKBUF_X1 U4822 ( .A(n5462), .Z(n4312) );
  NAND2_X1 U4823 ( .A1(n4575), .A2(n4977), .ZN(n7054) );
  INV_X2 U4824 ( .A(n6639), .ZN(n6198) );
  INV_X2 U4825 ( .A(n7030), .ZN(n5751) );
  INV_X2 U4826 ( .A(n6496), .ZN(n6495) );
  INV_X1 U4827 ( .A(n5935), .ZN(n4508) );
  INV_X1 U4828 ( .A(n5662), .ZN(n5677) );
  NOR2_X2 U4829 ( .A1(n5724), .A2(n5705), .ZN(n5706) );
  INV_X2 U4830 ( .A(n5814), .ZN(n6157) );
  OAI21_X1 U4831 ( .B1(n6210), .B2(n4766), .A(n4763), .ZN(n8977) );
  AND2_X1 U4832 ( .A1(n8633), .A2(n8831), .ZN(n8634) );
  NOR2_X1 U4833 ( .A1(n9190), .A2(n9390), .ZN(n9422) );
  XNOR2_X1 U4834 ( .A(n5217), .B(n5214), .ZN(n6660) );
  XNOR2_X1 U4835 ( .A(n4975), .B(n4563), .ZN(n8248) );
  NOR3_X2 U4836 ( .A1(n4913), .A2(n4571), .A3(n4632), .ZN(n4570) );
  INV_X2 U4837 ( .A(n4316), .ZN(n6730) );
  INV_X2 U4838 ( .A(n5878), .ZN(n6080) );
  NAND2_X2 U4839 ( .A1(n4517), .A2(n4828), .ZN(n5046) );
  CLKBUF_X1 U4840 ( .A(n5462), .Z(n4311) );
  BUF_X2 U4841 ( .A(n5462), .Z(n4313) );
  NAND2_X1 U4842 ( .A1(n4934), .A2(n4933), .ZN(n5462) );
  NAND4_X4 U4843 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n5771)
         );
  NAND2_X2 U4844 ( .A1(n8256), .A2(n6859), .ZN(n7098) );
  XNOR2_X2 U4845 ( .A(n8304), .B(n8305), .ZN(n8357) );
  OR2_X2 U4846 ( .A1(n4920), .A2(n4919), .ZN(n4921) );
  NAND2_X2 U4847 ( .A1(n6804), .A2(n6495), .ZN(n5090) );
  AOI211_X2 U4848 ( .C1(n5599), .C2(n5598), .A(n5597), .B(n7657), .ZN(n5606)
         );
  OAI21_X2 U4849 ( .B1(n6900), .B2(n6899), .A(n6864), .ZN(n8250) );
  NAND2_X2 U4850 ( .A1(n6858), .A2(n6857), .ZN(n6900) );
  INV_X1 U4851 ( .A(n6934), .ZN(n8342) );
  AND2_X2 U4852 ( .A1(n7597), .A2(n7587), .ZN(n7588) );
  NAND2_X1 U4853 ( .A1(n4887), .A2(n4886), .ZN(n8676) );
  NAND2_X1 U4854 ( .A1(n8687), .A2(n4652), .ZN(n4887) );
  NAND2_X1 U4855 ( .A1(n8786), .A2(n8787), .ZN(n8785) );
  OR2_X1 U4856 ( .A1(n9264), .A2(n9248), .ZN(n9227) );
  NAND2_X1 U4857 ( .A1(n8267), .A2(n4737), .ZN(n8467) );
  NAND2_X1 U4858 ( .A1(n7165), .A2(n5574), .ZN(n5071) );
  NAND2_X1 U4859 ( .A1(n8502), .A2(n7148), .ZN(n7152) );
  INV_X2 U4860 ( .A(n5033), .ZN(n10044) );
  NAND2_X2 U4861 ( .A1(n5520), .A2(n5522), .ZN(n7110) );
  INV_X1 U4862 ( .A(n7149), .ZN(n8502) );
  INV_X1 U4863 ( .A(n4996), .ZN(n10037) );
  NAND2_X2 U4864 ( .A1(n8342), .A2(n7387), .ZN(n10016) );
  AND4_X1 U4865 ( .A1(n4985), .A2(n4984), .A3(n4983), .A4(n4982), .ZN(n7063)
         );
  INV_X4 U4866 ( .A(n5000), .ZN(n5074) );
  INV_X4 U4867 ( .A(n8828), .ZN(n8583) );
  NAND2_X2 U4868 ( .A1(n9891), .A2(n9886), .ZN(n5814) );
  INV_X1 U4869 ( .A(n4923), .ZN(n4934) );
  NOR2_X1 U4870 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4633) );
  NOR2_X1 U4871 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4634) );
  INV_X2 U4872 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR3_X1 U4873 ( .A1(n9075), .A2(n6474), .A3(n6473), .ZN(n6475) );
  AOI211_X1 U4874 ( .C1(n8882), .C2(n8856), .A(n8664), .B(n8663), .ZN(n8665)
         );
  OR2_X1 U4875 ( .A1(n7955), .A2(n4526), .ZN(n4522) );
  AND2_X1 U4876 ( .A1(n5486), .A2(n5485), .ZN(n5494) );
  OAI21_X1 U4877 ( .B1(n7952), .B2(n7951), .A(n4386), .ZN(n7955) );
  NAND2_X1 U4878 ( .A1(n4713), .A2(n4717), .ZN(n8349) );
  NOR2_X1 U4879 ( .A1(n4388), .A2(n4387), .ZN(n4386) );
  NOR2_X1 U4880 ( .A1(n7950), .A2(n7948), .ZN(n4388) );
  NOR2_X1 U4881 ( .A1(n7949), .A2(n7929), .ZN(n4387) );
  AND2_X1 U4882 ( .A1(n7932), .A2(n4552), .ZN(n7943) );
  AND2_X1 U4883 ( .A1(n7931), .A2(n7930), .ZN(n7932) );
  NAND2_X1 U4884 ( .A1(n8365), .A2(n4739), .ZN(n8431) );
  NAND2_X1 U4885 ( .A1(n8768), .A2(n8767), .ZN(n8917) );
  OAI21_X1 U4886 ( .B1(n7485), .B2(n4726), .A(n4724), .ZN(n7717) );
  OAI21_X1 U4887 ( .B1(n8508), .B2(P2_REG1_REG_14__SCAN_IN), .A(n8506), .ZN(
        n8519) );
  OR2_X1 U4888 ( .A1(n9388), .A2(n9378), .ZN(n9376) );
  NAND2_X1 U4889 ( .A1(n7541), .A2(n5584), .ZN(n7561) );
  OR2_X1 U4890 ( .A1(n7739), .A2(n9100), .ZN(n7814) );
  NAND2_X1 U4891 ( .A1(n5071), .A2(n4883), .ZN(n7420) );
  OAI21_X1 U4892 ( .B1(n6424), .B2(n4790), .A(n4788), .ZN(n7314) );
  OAI21_X1 U4893 ( .B1(n7822), .B2(n4334), .A(n4389), .ZN(n7829) );
  NAND2_X1 U4894 ( .A1(n6905), .A2(n6906), .ZN(n6904) );
  OR2_X1 U4895 ( .A1(n7155), .A2(n7154), .ZN(n10053) );
  INV_X2 U4896 ( .A(n8831), .ZN(n4314) );
  NAND2_X1 U4897 ( .A1(n4792), .A2(n8089), .ZN(n7822) );
  AND2_X1 U4898 ( .A1(n5931), .A2(n5930), .ZN(n7308) );
  NAND2_X1 U4899 ( .A1(n5092), .A2(n5091), .ZN(n10064) );
  AND3_X1 U4900 ( .A1(n5891), .A2(n5890), .A3(n5889), .ZN(n7008) );
  INV_X1 U4901 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U4902 ( .A1(n4658), .A2(n5032), .ZN(n7189) );
  AND3_X1 U4903 ( .A1(n5786), .A2(n5785), .A3(n5784), .ZN(n6839) );
  AND4_X2 U4904 ( .A1(n4970), .A2(n4972), .A3(n4969), .A4(n4971), .ZN(n4316)
         );
  BUF_X2 U4905 ( .A(n5025), .Z(n5505) );
  AND2_X2 U4906 ( .A1(n6361), .A2(n6412), .ZN(n7030) );
  XNOR2_X1 U4907 ( .A(n4932), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6731) );
  XNOR2_X1 U4908 ( .A(n5513), .B(n5512), .ZN(n8257) );
  INV_X1 U4909 ( .A(n4311), .ZN(n4315) );
  CLKBUF_X2 U4910 ( .A(n5803), .Z(n6639) );
  NAND2_X1 U4911 ( .A1(n4923), .A2(n4922), .ZN(n5001) );
  NAND2_X2 U4912 ( .A1(n8136), .A2(n4923), .ZN(n5000) );
  NAND2_X1 U4914 ( .A1(n4514), .A2(n4512), .ZN(n9891) );
  XNOR2_X1 U4915 ( .A(n5715), .B(n5714), .ZN(n8338) );
  NAND2_X1 U4916 ( .A1(n8960), .A2(n4918), .ZN(n4923) );
  XNOR2_X1 U4917 ( .A(n5734), .B(n5735), .ZN(n7749) );
  XNOR2_X1 U4918 ( .A(n5727), .B(n5726), .ZN(n8122) );
  MUX2_X1 U4919 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4917), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n4918) );
  NAND2_X1 U4920 ( .A1(n5691), .A2(n4661), .ZN(n4943) );
  XNOR2_X1 U4921 ( .A(n5010), .B(n4993), .ZN(n5008) );
  AND2_X1 U4922 ( .A1(n4780), .A2(n5698), .ZN(n4504) );
  NAND2_X2 U4923 ( .A1(n6496), .A2(P1_U3084), .ZN(n9537) );
  NOR2_X1 U4924 ( .A1(n4632), .A2(n4631), .ZN(n4897) );
  NAND2_X1 U4925 ( .A1(n9759), .A2(n4948), .ZN(n4865) );
  AND2_X1 U4926 ( .A1(n5697), .A2(n5898), .ZN(n5698) );
  NAND2_X1 U4927 ( .A1(n9758), .A2(n4947), .ZN(n4866) );
  NAND4_X1 U4928 ( .A1(n4635), .A2(n4634), .A3(n4633), .A4(n5162), .ZN(n4632)
         );
  NAND2_X1 U4929 ( .A1(n4915), .A2(n4891), .ZN(n4890) );
  INV_X1 U4930 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5162) );
  INV_X4 U4931 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X2 U4932 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9758) );
  AND2_X1 U4933 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9759) );
  INV_X1 U4934 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5063) );
  INV_X1 U4935 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4698) );
  NOR2_X1 U4936 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4781) );
  INV_X1 U4937 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5749) );
  NOR2_X1 U4938 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5699) );
  NOR2_X1 U4939 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5700) );
  NOR2_X1 U4940 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5701) );
  NOR3_X1 U4941 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n4912) );
  NOR2_X1 U4942 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4635) );
  INV_X1 U4943 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4697) );
  INV_X1 U4944 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4891) );
  INV_X1 U4945 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4915) );
  AND3_X2 U4946 ( .A1(n5821), .A2(n5820), .A3(n5819), .ZN(n9969) );
  NOR2_X2 U4947 ( .A1(n7814), .A2(n9017), .ZN(n9387) );
  NAND2_X1 U4948 ( .A1(n4520), .A2(n4992), .ZN(n5009) );
  AND4_X2 U4949 ( .A1(n4940), .A2(n4939), .A3(n4938), .A4(n4937), .ZN(n8256)
         );
  NAND2_X1 U4950 ( .A1(n4316), .A2(n7054), .ZN(n5543) );
  NAND2_X1 U4951 ( .A1(n4894), .A2(n4893), .ZN(n8627) );
  AOI21_X2 U4952 ( .B1(n8250), .B2(n8249), .A(n6868), .ZN(n6905) );
  OR2_X1 U4953 ( .A1(n8659), .A2(n8652), .ZN(n4895) );
  NAND2_X1 U4954 ( .A1(n8659), .A2(n4336), .ZN(n4894) );
  NAND2_X1 U4955 ( .A1(n4943), .A2(n4942), .ZN(n6803) );
  NAND3_X2 U4956 ( .A1(n5766), .A2(n5767), .A3(n5765), .ZN(n5774) );
  INV_X2 U4957 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4945) );
  INV_X2 U4958 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4988) );
  NAND2_X2 U4959 ( .A1(n7101), .A2(n5520), .ZN(n7127) );
  INV_X8 U4960 ( .A(n8308), .ZN(n8318) );
  NAND2_X1 U4961 ( .A1(n8757), .A2(n5337), .ZN(n8740) );
  OR2_X4 U4962 ( .A1(n8338), .A2(n8131), .ZN(n5804) );
  NOR2_X2 U4963 ( .A1(n4943), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4920) );
  AOI21_X2 U4964 ( .B1(n7138), .B2(n7154), .A(n5053), .ZN(n7165) );
  AOI211_X2 U4965 ( .C1(n10088), .C2(n8888), .A(n8887), .B(n8886), .ZN(n8889)
         );
  AOI21_X2 U4966 ( .B1(n8679), .B2(n8678), .A(n8677), .ZN(n8680) );
  AOI21_X2 U4967 ( .B1(n8785), .B2(n5327), .A(n5326), .ZN(n8757) );
  NAND2_X1 U4968 ( .A1(n5178), .A2(n9623), .ZN(n5195) );
  NAND2_X1 U4969 ( .A1(n4482), .A2(n4481), .ZN(n5744) );
  AOI21_X1 U4970 ( .B1(n4484), .B2(n5899), .A(n5899), .ZN(n4481) );
  AOI21_X1 U4971 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_20__SCAN_IN), .ZN(n4484) );
  AND2_X1 U4972 ( .A1(n8257), .A2(n8828), .ZN(n6760) );
  AND2_X1 U4973 ( .A1(n5534), .A2(n5669), .ZN(n5675) );
  AND3_X1 U4974 ( .A1(n7387), .A2(n8828), .A3(n8257), .ZN(n4740) );
  NAND2_X1 U4975 ( .A1(n6492), .A2(n4750), .ZN(n5935) );
  OAI21_X1 U4976 ( .B1(n5606), .B2(n5605), .A(n4344), .ZN(n4641) );
  OR2_X1 U4977 ( .A1(n5635), .A2(n4656), .ZN(n4655) );
  NAND2_X1 U4978 ( .A1(n8727), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U4979 ( .A1(n5636), .A2(n5637), .ZN(n4657) );
  INV_X1 U4980 ( .A(n4372), .ZN(n4489) );
  INV_X1 U4981 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5177) );
  OR2_X1 U4982 ( .A1(n8881), .A2(n8888), .ZN(n4585) );
  AND2_X1 U4983 ( .A1(n5646), .A2(n5643), .ZN(n8613) );
  OR2_X1 U4984 ( .A1(n5372), .A2(n9724), .ZN(n5386) );
  OR2_X1 U4985 ( .A1(n8907), .A2(n8612), .ZN(n5360) );
  OR2_X1 U4986 ( .A1(n8925), .A2(n8929), .ZN(n4590) );
  OR2_X1 U4987 ( .A1(n5186), .A2(n6989), .ZN(n5205) );
  OR2_X1 U4988 ( .A1(n8398), .A2(n7660), .ZN(n7514) );
  NOR2_X1 U4989 ( .A1(n4462), .A2(n4458), .ZN(n4455) );
  NOR2_X1 U4990 ( .A1(n4458), .A2(n4460), .ZN(n4454) );
  NAND2_X1 U4991 ( .A1(n5244), .A2(n4930), .ZN(n5279) );
  INV_X1 U4992 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4930) );
  OR2_X1 U4993 ( .A1(n5103), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5140) );
  INV_X1 U4994 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4696) );
  XNOR2_X1 U4995 ( .A(n5794), .B(n7030), .ZN(n5798) );
  NAND2_X1 U4996 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  OR2_X1 U4997 ( .A1(n6839), .A2(n5935), .ZN(n5793) );
  OAI21_X1 U4998 ( .B1(n5773), .B2(n4748), .A(n5796), .ZN(n5799) );
  NAND2_X1 U4999 ( .A1(n7987), .A2(n4403), .ZN(n4402) );
  INV_X1 U5000 ( .A(n8060), .ZN(n4403) );
  NAND2_X1 U5001 ( .A1(n6265), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6282) );
  OR2_X1 U5002 ( .A1(n9267), .A2(n9280), .ZN(n9237) );
  NOR2_X1 U5003 ( .A1(n6405), .A2(n4624), .ZN(n4623) );
  INV_X1 U5004 ( .A(n4625), .ZN(n4624) );
  OR2_X1 U5005 ( .A1(n9328), .A2(n9306), .ZN(n7998) );
  OR2_X1 U5006 ( .A1(n9126), .A2(n9969), .ZN(n8089) );
  NAND2_X1 U5007 ( .A1(n6350), .A2(n8122), .ZN(n4750) );
  NAND2_X1 U5008 ( .A1(n4846), .A2(n4845), .ZN(n5498) );
  AOI21_X1 U5009 ( .B1(n4848), .B2(n4850), .A(n4376), .ZN(n4845) );
  NAND2_X1 U5010 ( .A1(n5470), .A2(n4848), .ZN(n4846) );
  AOI21_X1 U5011 ( .B1(n5434), .B2(n4836), .A(n4835), .ZN(n4834) );
  INV_X1 U5012 ( .A(n5436), .ZN(n4835) );
  INV_X1 U5013 ( .A(n5416), .ZN(n4836) );
  INV_X1 U5014 ( .A(n5434), .ZN(n4837) );
  NAND2_X1 U5015 ( .A1(n5400), .A2(n5399), .ZN(n5415) );
  NAND2_X1 U5016 ( .A1(n4863), .A2(n4371), .ZN(n5400) );
  AOI21_X1 U5017 ( .B1(n4546), .B2(n4544), .A(n4366), .ZN(n4543) );
  AND2_X1 U5018 ( .A1(n5330), .A2(n5317), .ZN(n5328) );
  AND2_X1 U5019 ( .A1(n5698), .A2(n4356), .ZN(n4502) );
  INV_X1 U5020 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4503) );
  OAI21_X1 U5021 ( .B1(n5175), .B2(n5174), .A(n5176), .ZN(n5194) );
  NAND2_X1 U5022 ( .A1(n5121), .A2(n9670), .ZN(n5138) );
  INV_X1 U5023 ( .A(SI_11_), .ZN(n5139) );
  AND2_X1 U5024 ( .A1(n5120), .A2(n5099), .ZN(n5118) );
  OAI21_X1 U5025 ( .B1(n6496), .B2(n4565), .A(n4564), .ZN(n5024) );
  NAND2_X1 U5026 ( .A1(n6496), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5027 ( .A1(n8290), .A2(n8376), .ZN(n8379) );
  INV_X1 U5028 ( .A(n8305), .ZN(n4390) );
  NOR2_X1 U5029 ( .A1(n6759), .A2(n6751), .ZN(n6761) );
  NAND2_X1 U5030 ( .A1(n6934), .A2(n8583), .ZN(n6944) );
  NAND2_X1 U5031 ( .A1(n7209), .A2(n7210), .ZN(n8506) );
  NAND2_X1 U5032 ( .A1(n8618), .A2(n8681), .ZN(n8619) );
  INV_X1 U5033 ( .A(n8619), .ZN(n4682) );
  XNOR2_X1 U5034 ( .A(n8881), .B(n8681), .ZN(n8652) );
  AND2_X1 U5035 ( .A1(n5433), .A2(n5641), .ZN(n4886) );
  INV_X1 U5036 ( .A(n8679), .ZN(n5433) );
  OR2_X1 U5037 ( .A1(n8893), .A2(n8714), .ZN(n5641) );
  OR2_X1 U5038 ( .A1(n8897), .A2(n8729), .ZN(n4471) );
  NOR2_X1 U5039 ( .A1(n8613), .A2(n4473), .ZN(n4470) );
  AOI21_X1 U5040 ( .B1(n8917), .B2(n4331), .A(n4684), .ZN(n4683) );
  NAND2_X1 U5041 ( .A1(n4687), .A2(n4685), .ZN(n4684) );
  AND2_X1 U5042 ( .A1(n8721), .A2(n4693), .ZN(n4687) );
  OR2_X1 U5043 ( .A1(n8750), .A2(n8907), .ZN(n8734) );
  AND2_X1 U5044 ( .A1(n4317), .A2(n5539), .ZN(n4877) );
  NAND2_X1 U5045 ( .A1(n8605), .A2(n8604), .ZN(n4464) );
  INV_X1 U5046 ( .A(n6804), .ZN(n5299) );
  AOI21_X1 U5047 ( .B1(n4699), .B2(n7117), .A(n4904), .ZN(n7155) );
  AND2_X1 U5048 ( .A1(n7116), .A2(n7153), .ZN(n4699) );
  AND2_X1 U5049 ( .A1(n4741), .A2(n6752), .ZN(n10088) );
  MUX2_X1 U5050 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4941), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n4942) );
  OAI21_X1 U5051 ( .B1(n5689), .B2(n4890), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4941) );
  AND2_X1 U5052 ( .A1(n5756), .A2(n5755), .ZN(n6614) );
  OR2_X1 U5053 ( .A1(n6177), .A2(n9043), .ZN(n6196) );
  AND2_X1 U5054 ( .A1(n8122), .A2(n8070), .ZN(n8121) );
  INV_X1 U5055 ( .A(n5805), .ZN(n6462) );
  AOI21_X1 U5056 ( .B1(n9907), .B2(n4449), .A(n9926), .ZN(n4447) );
  INV_X1 U5057 ( .A(n6535), .ZN(n4449) );
  NOR2_X1 U5058 ( .A1(n5713), .A2(n4513), .ZN(n4512) );
  OR2_X1 U5059 ( .A1(n4862), .A2(n4515), .ZN(n4514) );
  NOR2_X1 U5060 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4513) );
  NAND2_X1 U5061 ( .A1(n4662), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U5062 ( .A1(n9302), .A2(n4623), .ZN(n4620) );
  INV_X1 U5063 ( .A(n7900), .ZN(n4804) );
  OR2_X1 U5064 ( .A1(n9458), .A2(n9322), .ZN(n4625) );
  INV_X1 U5065 ( .A(n6395), .ZN(n4842) );
  AND2_X1 U5066 ( .A1(n6440), .A2(n6439), .ZN(n9400) );
  XNOR2_X1 U5067 ( .A(n5771), .B(n8079), .ZN(n6707) );
  AND2_X1 U5068 ( .A1(n5814), .A2(n6496), .ZN(n5812) );
  NOR2_X1 U5069 ( .A1(n4323), .A2(n4860), .ZN(n4859) );
  NAND2_X1 U5070 ( .A1(n5729), .A2(n4861), .ZN(n4860) );
  INV_X1 U5071 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4861) );
  XNOR2_X1 U5072 ( .A(n5733), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U5073 ( .A1(n4533), .A2(n4534), .ZN(n5278) );
  NAND2_X1 U5074 ( .A1(n5217), .A2(n4537), .ZN(n4533) );
  AOI21_X1 U5075 ( .B1(n4426), .B2(n5065), .A(n4347), .ZN(n4425) );
  MUX2_X1 U5076 ( .A(n5668), .B(n5677), .S(n5667), .Z(n5676) );
  XNOR2_X1 U5077 ( .A(n4875), .B(n8583), .ZN(n5516) );
  OAI21_X1 U5078 ( .B1(n5494), .B2(n4871), .A(n4868), .ZN(n4875) );
  NOR2_X1 U5079 ( .A1(n8073), .A2(n8122), .ZN(n8074) );
  INV_X1 U5080 ( .A(n8070), .ZN(n9184) );
  MUX2_X1 U5081 ( .A(n5554), .B(n5553), .S(n5671), .Z(n5562) );
  OR2_X1 U5082 ( .A1(n5551), .A2(n5544), .ZN(n5554) );
  INV_X1 U5083 ( .A(n4646), .ZN(n4645) );
  AOI22_X1 U5084 ( .A1(n5578), .A2(n5671), .B1(n4649), .B2(n10064), .ZN(n4646)
         );
  AND2_X1 U5085 ( .A1(n5587), .A2(n5581), .ZN(n4647) );
  NAND2_X1 U5086 ( .A1(n4638), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5087 ( .A1(n4640), .A2(n5612), .ZN(n4639) );
  NAND2_X1 U5088 ( .A1(n5275), .A2(n5677), .ZN(n4637) );
  NAND2_X1 U5089 ( .A1(n4557), .A2(n4554), .ZN(n7909) );
  OAI21_X1 U5090 ( .B1(n7904), .B2(n9307), .A(n4337), .ZN(n4557) );
  NOR2_X1 U5091 ( .A1(n5639), .A2(n5640), .ZN(n4654) );
  NOR2_X1 U5092 ( .A1(n4545), .A2(n4542), .ZN(n4541) );
  INV_X1 U5093 ( .A(n5313), .ZN(n4542) );
  INV_X1 U5094 ( .A(n4546), .ZN(n4545) );
  INV_X1 U5095 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n4747) );
  INV_X1 U5096 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4745) );
  AND2_X1 U5097 ( .A1(n4858), .A2(n5257), .ZN(n4857) );
  NAND2_X1 U5098 ( .A1(n5236), .A2(n5238), .ZN(n4858) );
  INV_X1 U5099 ( .A(n4857), .ZN(n4856) );
  INV_X1 U5100 ( .A(n5214), .ZN(n4539) );
  NAND2_X1 U5101 ( .A1(n5159), .A2(n9726), .ZN(n5176) );
  AOI21_X1 U5102 ( .B1(n5093), .B2(n5095), .A(n4416), .ZN(n4415) );
  INV_X1 U5103 ( .A(n5118), .ZN(n4416) );
  INV_X1 U5104 ( .A(SI_9_), .ZN(n5096) );
  AOI21_X1 U5105 ( .B1(n7588), .B2(n4725), .A(n4325), .ZN(n4724) );
  INV_X1 U5106 ( .A(n7588), .ZN(n4726) );
  AND2_X1 U5107 ( .A1(n8869), .A2(n5484), .ZN(n5664) );
  OR2_X1 U5108 ( .A1(n8888), .A2(n8404), .ZN(n5653) );
  OR2_X1 U5109 ( .A1(n5304), .A2(n5303), .ZN(n5320) );
  OR2_X1 U5110 ( .A1(n8919), .A2(n8610), .ZN(n5629) );
  OR2_X1 U5111 ( .A1(n8603), .A2(n8841), .ZN(n5608) );
  NAND2_X1 U5112 ( .A1(n5167), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5186) );
  OR2_X1 U5113 ( .A1(n5146), .A2(n5145), .ZN(n5168) );
  AOI21_X1 U5114 ( .B1(n10012), .B2(n6750), .A(n10014), .ZN(n7183) );
  NAND2_X1 U5115 ( .A1(n5683), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5686) );
  NAND2_X1 U5116 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  INV_X1 U5117 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5681) );
  OR2_X1 U5118 ( .A1(n5079), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5103) );
  INV_X1 U5119 ( .A(n6209), .ZN(n4765) );
  AOI21_X1 U5120 ( .B1(n4769), .B2(n4770), .A(n4359), .ZN(n4767) );
  INV_X1 U5121 ( .A(n6174), .ZN(n4761) );
  XNOR2_X1 U5122 ( .A(n5824), .B(n7030), .ZN(n5828) );
  INV_X1 U5123 ( .A(n5799), .ZN(n5797) );
  NOR2_X1 U5124 ( .A1(n4494), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U5125 ( .A1(n4485), .A2(n6090), .ZN(n4490) );
  NAND2_X1 U5126 ( .A1(n4493), .A2(n4497), .ZN(n4485) );
  INV_X1 U5127 ( .A(n4498), .ZN(n4493) );
  NAND2_X1 U5128 ( .A1(n6068), .A2(n7793), .ZN(n4498) );
  AND2_X1 U5129 ( .A1(n7932), .A2(n4553), .ZN(n7947) );
  NOR2_X1 U5130 ( .A1(n7945), .A2(n7944), .ZN(n4553) );
  OR2_X1 U5131 ( .A1(n5805), .A2(n6533), .ZN(n5791) );
  NAND2_X1 U5132 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  NAND2_X1 U5133 ( .A1(n4604), .A2(n4606), .ZN(n4601) );
  NOR2_X1 U5134 ( .A1(n9225), .A2(n4603), .ZN(n4602) );
  INV_X1 U5135 ( .A(n4604), .ZN(n4603) );
  NAND2_X1 U5136 ( .A1(n9225), .A2(n7987), .ZN(n4404) );
  NOR2_X1 U5137 ( .A1(n7985), .A2(n4608), .ZN(n4607) );
  INV_X1 U5138 ( .A(n6408), .ZN(n4608) );
  OR2_X1 U5139 ( .A1(n6479), .A2(n9243), .ZN(n8060) );
  OAI22_X1 U5140 ( .A1(n6402), .A2(n4824), .B1(n9342), .B2(n9365), .ZN(n4823)
         );
  NAND2_X1 U5141 ( .A1(n4352), .A2(n6401), .ZN(n4824) );
  AND2_X1 U5142 ( .A1(n4825), .A2(n4615), .ZN(n4614) );
  NAND2_X1 U5143 ( .A1(n4616), .A2(n6400), .ZN(n4615) );
  NOR2_X1 U5144 ( .A1(n6402), .A2(n4826), .ZN(n4825) );
  INV_X1 U5145 ( .A(n9375), .ZN(n4616) );
  NAND2_X1 U5146 ( .A1(n4614), .A2(n4617), .ZN(n4612) );
  INV_X1 U5147 ( .A(n6400), .ZN(n4617) );
  AND2_X1 U5148 ( .A1(n7878), .A2(n9368), .ZN(n7960) );
  NOR2_X1 U5149 ( .A1(n7978), .A2(n4802), .ZN(n4801) );
  INV_X1 U5150 ( .A(n7856), .ZN(n4802) );
  OR2_X1 U5151 ( .A1(n7646), .A2(n9844), .ZN(n4679) );
  INV_X1 U5152 ( .A(n7968), .ZN(n4791) );
  NAND2_X1 U5153 ( .A1(n8082), .A2(n8084), .ZN(n4838) );
  AOI21_X1 U5154 ( .B1(n4784), .B2(n4787), .A(n7852), .ZN(n4783) );
  INV_X1 U5155 ( .A(n7857), .ZN(n4787) );
  NAND2_X1 U5156 ( .A1(n5454), .A2(n5453), .ZN(n5470) );
  AOI21_X1 U5157 ( .B1(n4834), .B2(n4837), .A(n4833), .ZN(n4832) );
  AND2_X1 U5158 ( .A1(n5453), .A2(n5440), .ZN(n5451) );
  AND2_X1 U5159 ( .A1(n5436), .A2(n5421), .ZN(n5434) );
  OR2_X1 U5160 ( .A1(n5415), .A2(n5414), .ZN(n5417) );
  NAND2_X1 U5161 ( .A1(n4528), .A2(n4527), .ZN(n4843) );
  AOI21_X1 U5162 ( .B1(n4529), .B2(n4532), .A(n5291), .ZN(n4527) );
  OAI21_X1 U5163 ( .B1(n5217), .B2(n4539), .A(n5216), .ZN(n5237) );
  AND2_X1 U5164 ( .A1(n5195), .A2(n5180), .ZN(n5193) );
  NAND2_X1 U5165 ( .A1(n5158), .A2(n5157), .ZN(n5175) );
  AND2_X1 U5166 ( .A1(n5138), .A2(n5123), .ZN(n5136) );
  INV_X1 U5167 ( .A(n4819), .ZN(n4780) );
  NAND2_X1 U5168 ( .A1(n5087), .A2(n9638), .ZN(n5095) );
  NAND2_X1 U5169 ( .A1(n5086), .A2(n5085), .ZN(n5094) );
  INV_X1 U5170 ( .A(SI_5_), .ZN(n9636) );
  INV_X1 U5171 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5696) );
  NAND2_X1 U5172 ( .A1(n4820), .A2(n5696), .ZN(n4819) );
  INV_X1 U5173 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4820) );
  INV_X1 U5174 ( .A(SI_8_), .ZN(n9638) );
  NAND2_X1 U5175 ( .A1(n8300), .A2(n8299), .ZN(n8304) );
  OR2_X1 U5176 ( .A1(n5000), .A2(n4936), .ZN(n4937) );
  NOR2_X1 U5177 ( .A1(n7284), .A2(n7283), .ZN(n4902) );
  NOR2_X1 U5178 ( .A1(n4902), .A2(n4733), .ZN(n4730) );
  XNOR2_X1 U5179 ( .A(n8308), .B(n7054), .ZN(n6733) );
  OAI21_X1 U5180 ( .B1(n8421), .B2(n8729), .A(n8356), .ZN(n8301) );
  AND2_X1 U5181 ( .A1(n8288), .A2(n8283), .ZN(n4739) );
  INV_X1 U5182 ( .A(n8434), .ZN(n8288) );
  INV_X1 U5183 ( .A(n6736), .ZN(n4391) );
  AND2_X1 U5184 ( .A1(n7184), .A2(n7183), .ZN(n6756) );
  OR2_X1 U5185 ( .A1(n8865), .A2(n5533), .ZN(n5669) );
  AND2_X1 U5186 ( .A1(n8625), .A2(n8491), .ZN(n5667) );
  AND2_X1 U5187 ( .A1(n5393), .A2(n5392), .ZN(n8423) );
  AND2_X1 U5188 ( .A1(n5359), .A2(n5358), .ZN(n8612) );
  AND4_X1 U5189 ( .A1(n5005), .A2(n5004), .A3(n5003), .A4(n5002), .ZN(n7118)
         );
  NOR2_X1 U5190 ( .A1(n8239), .A2(n4562), .ZN(n8238) );
  NAND2_X1 U5191 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n4562) );
  NOR2_X1 U5192 ( .A1(n8229), .A2(n8228), .ZN(n8227) );
  INV_X1 U5193 ( .A(n8865), .ZN(n8596) );
  NOR2_X1 U5194 ( .A1(n8690), .A2(n4583), .ZN(n8621) );
  NAND2_X1 U5195 ( .A1(n8620), .A2(n4584), .ZN(n4583) );
  NOR2_X1 U5196 ( .A1(n8869), .A2(n4585), .ZN(n4584) );
  OR2_X1 U5197 ( .A1(n8645), .A2(n4312), .ZN(n5467) );
  OR2_X1 U5198 ( .A1(n8652), .A2(n4682), .ZN(n4681) );
  NAND2_X1 U5199 ( .A1(n5658), .A2(n5661), .ZN(n8641) );
  NAND2_X1 U5200 ( .A1(n8666), .A2(n8616), .ZN(n8653) );
  NAND2_X1 U5201 ( .A1(n8671), .A2(n8404), .ZN(n8616) );
  OR2_X1 U5202 ( .A1(n8690), .A2(n8888), .ZN(n8669) );
  NAND2_X1 U5203 ( .A1(n5653), .A2(n5651), .ZN(n8679) );
  NAND2_X1 U5204 ( .A1(n8667), .A2(n8679), .ZN(n8666) );
  INV_X1 U5205 ( .A(n4468), .ZN(n4467) );
  OAI21_X1 U5206 ( .B1(n4470), .B2(n4469), .A(n8686), .ZN(n4468) );
  INV_X1 U5207 ( .A(n4471), .ZN(n4469) );
  AND2_X1 U5208 ( .A1(n5413), .A2(n5412), .ZN(n8714) );
  NAND2_X1 U5209 ( .A1(n8739), .A2(n8612), .ZN(n4693) );
  INV_X1 U5210 ( .A(n4690), .ZN(n4689) );
  NOR2_X1 U5211 ( .A1(n8917), .A2(n4318), .ZN(n4692) );
  NOR2_X1 U5212 ( .A1(n4588), .A2(n8919), .ZN(n4587) );
  NAND2_X1 U5213 ( .A1(n4589), .A2(n8755), .ZN(n4588) );
  OAI22_X1 U5214 ( .A1(n8795), .A2(n8608), .B1(n8801), .B2(n8819), .ZN(n8779)
         );
  OR2_X1 U5215 ( .A1(n8822), .A2(n8934), .ZN(n8823) );
  NOR2_X1 U5216 ( .A1(n8823), .A2(n8929), .ZN(n8796) );
  NAND2_X1 U5217 ( .A1(n8842), .A2(n4333), .ZN(n4456) );
  AND2_X1 U5218 ( .A1(n4464), .A2(n4333), .ZN(n8843) );
  AND4_X1 U5219 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n8820)
         );
  AOI21_X1 U5220 ( .B1(n5213), .B2(n7657), .A(n4881), .ZN(n4880) );
  INV_X1 U5221 ( .A(n5602), .ZN(n4881) );
  INV_X1 U5222 ( .A(n4703), .ZN(n4702) );
  OAI21_X1 U5223 ( .B1(n4705), .B2(n7657), .A(n7776), .ZN(n4703) );
  NAND2_X1 U5224 ( .A1(n7656), .A2(n5213), .ZN(n7685) );
  NAND2_X1 U5225 ( .A1(n7683), .A2(n4706), .ZN(n4705) );
  INV_X1 U5226 ( .A(n4899), .ZN(n4706) );
  NOR2_X1 U5227 ( .A1(n7652), .A2(n7653), .ZN(n7682) );
  OR2_X1 U5228 ( .A1(n7528), .A2(n8398), .ZN(n7665) );
  NAND2_X1 U5229 ( .A1(n10053), .A2(n4707), .ZN(n7415) );
  NOR2_X1 U5230 ( .A1(n7166), .A2(n4708), .ZN(n4707) );
  INV_X1 U5231 ( .A(n7162), .ZN(n4708) );
  NAND2_X1 U5232 ( .A1(n4577), .A2(n4576), .ZN(n7142) );
  NOR2_X1 U5233 ( .A1(n5033), .A2(n7189), .ZN(n4576) );
  INV_X1 U5234 ( .A(n7120), .ZN(n4577) );
  AND2_X1 U5235 ( .A1(n7110), .A2(n7113), .ZN(n7111) );
  OR2_X1 U5236 ( .A1(n6797), .A2(n6762), .ZN(n8838) );
  NAND2_X1 U5237 ( .A1(n5406), .A2(n5405), .ZN(n8893) );
  NAND2_X1 U5238 ( .A1(n5384), .A2(n5383), .ZN(n8897) );
  AND2_X1 U5239 ( .A1(n5106), .A2(n5105), .ZN(n10072) );
  NAND2_X1 U5240 ( .A1(n4741), .A2(n8257), .ZN(n10096) );
  OAI21_X1 U5241 ( .B1(n6749), .B2(n6748), .A(n6750), .ZN(n7194) );
  OAI21_X1 U5242 ( .B1(n7746), .B2(n6738), .A(n7801), .ZN(n10007) );
  XOR2_X1 U5243 ( .A(n7702), .B(P2_B_REG_SCAN_IN), .Z(n6738) );
  AND2_X1 U5244 ( .A1(n6878), .A2(n10013), .ZN(n10008) );
  NOR2_X1 U5245 ( .A1(n4888), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4661) );
  NAND2_X1 U5246 ( .A1(n4889), .A2(n4916), .ZN(n4888) );
  INV_X1 U5247 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4916) );
  NAND2_X1 U5248 ( .A1(n4572), .A2(n4914), .ZN(n4571) );
  INV_X1 U5249 ( .A(n5279), .ZN(n4736) );
  AOI21_X1 U5250 ( .B1(P2_IR_REG_31__SCAN_IN), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_19__SCAN_IN), .ZN(n4735) );
  AND2_X2 U5251 ( .A1(n5028), .A2(n4907), .ZN(n5062) );
  INV_X1 U5252 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4907) );
  NAND2_X1 U5253 ( .A1(n4755), .A2(n5897), .ZN(n4753) );
  INV_X1 U5254 ( .A(n4756), .ZN(n4755) );
  AOI21_X1 U5255 ( .B1(n4776), .B2(n9000), .A(n6474), .ZN(n4775) );
  OR2_X1 U5256 ( .A1(n6282), .A2(n6281), .ZN(n6313) );
  INV_X1 U5257 ( .A(n4495), .ZN(n4496) );
  AND2_X1 U5258 ( .A1(n9050), .A2(n6226), .ZN(n4770) );
  OR2_X1 U5259 ( .A1(n9050), .A2(n6226), .ZN(n4769) );
  NAND2_X1 U5260 ( .A1(n9088), .A2(n9091), .ZN(n4742) );
  NAND2_X1 U5261 ( .A1(n5742), .A2(n5741), .ZN(n6611) );
  AOI21_X1 U5262 ( .B1(n5740), .B2(n6920), .A(n5739), .ZN(n5741) );
  INV_X1 U5263 ( .A(n8986), .ZN(n4762) );
  NAND2_X1 U5264 ( .A1(n9058), .A2(n9059), .ZN(n9057) );
  NOR2_X1 U5265 ( .A1(n6366), .A2(n6521), .ZN(n6362) );
  OR2_X1 U5266 ( .A1(n5805), .A2(n5717), .ZN(n5723) );
  INV_X1 U5267 ( .A(n4451), .ZN(n7375) );
  OR2_X1 U5268 ( .A1(n7499), .A2(n7498), .ZN(n4440) );
  AOI21_X1 U5269 ( .B1(n4607), .B2(n4605), .A(n4326), .ZN(n4604) );
  INV_X1 U5270 ( .A(n4607), .ZN(n4606) );
  NOR2_X1 U5271 ( .A1(n4364), .A2(n4619), .ZN(n4618) );
  AOI21_X1 U5272 ( .B1(n4358), .B2(n4623), .A(n4622), .ZN(n4621) );
  INV_X1 U5273 ( .A(n7905), .ZN(n4622) );
  NAND2_X1 U5274 ( .A1(n4803), .A2(n4338), .ZN(n9275) );
  AOI21_X1 U5275 ( .B1(n4420), .B2(n6432), .A(n4419), .ZN(n4418) );
  INV_X1 U5276 ( .A(n9304), .ZN(n4419) );
  NAND2_X1 U5277 ( .A1(n6404), .A2(n6403), .ZN(n9302) );
  AND2_X1 U5278 ( .A1(n8002), .A2(n7900), .ZN(n9304) );
  INV_X1 U5279 ( .A(n6162), .ZN(n6160) );
  INV_X1 U5280 ( .A(n8000), .ZN(n4796) );
  AOI21_X1 U5281 ( .B1(n8000), .B2(n4795), .A(n4794), .ZN(n4793) );
  INV_X1 U5282 ( .A(n8013), .ZN(n4794) );
  INV_X1 U5283 ( .A(n4613), .ZN(n9355) );
  AOI21_X1 U5284 ( .B1(n9374), .B2(n9375), .A(n4617), .ZN(n4613) );
  NOR2_X1 U5285 ( .A1(n8012), .A2(n4798), .ZN(n4797) );
  AND4_X1 U5286 ( .A1(n6103), .A2(n6102), .A3(n6101), .A4(n6100), .ZN(n9402)
         );
  NAND2_X1 U5287 ( .A1(n7811), .A2(n7981), .ZN(n6430) );
  INV_X1 U5288 ( .A(n7960), .ZN(n9398) );
  NAND2_X1 U5289 ( .A1(n4432), .A2(n4430), .ZN(n7811) );
  AOI21_X1 U5290 ( .B1(n6429), .B2(n4800), .A(n4799), .ZN(n4432) );
  NAND2_X1 U5291 ( .A1(n4431), .A2(n6429), .ZN(n4430) );
  INV_X1 U5292 ( .A(n8043), .ZN(n4799) );
  INV_X1 U5293 ( .A(n4840), .ZN(n4596) );
  AOI21_X1 U5294 ( .B1(n4841), .B2(n4322), .A(n4339), .ZN(n4840) );
  OR2_X1 U5295 ( .A1(n6077), .A2(n6076), .ZN(n6098) );
  AND2_X1 U5296 ( .A1(n4433), .A2(n7869), .ZN(n6429) );
  NAND2_X1 U5297 ( .A1(n6428), .A2(n4801), .ZN(n7723) );
  NAND2_X1 U5298 ( .A1(n6010), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6033) );
  OAI21_X1 U5299 ( .B1(n7440), .B2(n6389), .A(n6388), .ZN(n7615) );
  NOR2_X1 U5300 ( .A1(n7447), .A2(n9844), .ZN(n7616) );
  NAND2_X1 U5301 ( .A1(n6427), .A2(n8033), .ZN(n7441) );
  OR2_X1 U5302 ( .A1(n9122), .A2(n7352), .ZN(n8017) );
  AND2_X1 U5303 ( .A1(n7969), .A2(n6383), .ZN(n4851) );
  NAND2_X1 U5304 ( .A1(n6424), .A2(n4332), .ZN(n7245) );
  NAND2_X1 U5305 ( .A1(n6999), .A2(n6382), .ZN(n7029) );
  NAND2_X1 U5306 ( .A1(n7029), .A2(n7968), .ZN(n7028) );
  OAI21_X1 U5307 ( .B1(n7822), .B2(n6420), .A(n8024), .ZN(n7218) );
  NAND2_X1 U5308 ( .A1(n6887), .A2(n4844), .ZN(n7225) );
  AND2_X1 U5309 ( .A1(n7217), .A2(n6380), .ZN(n4844) );
  NAND2_X1 U5310 ( .A1(n6888), .A2(n6890), .ZN(n6887) );
  INV_X1 U5311 ( .A(n4838), .ZN(n7964) );
  NAND2_X1 U5312 ( .A1(n6706), .A2(n6707), .ZN(n6709) );
  NAND2_X1 U5313 ( .A1(n7967), .A2(n6711), .ZN(n6710) );
  OR2_X1 U5314 ( .A1(n6493), .A2(n9861), .ZN(n9405) );
  OR2_X1 U5315 ( .A1(n6917), .A2(n6438), .ZN(n9390) );
  NOR2_X1 U5316 ( .A1(n7749), .A2(n7705), .ZN(n4480) );
  XNOR2_X1 U5317 ( .A(n5503), .B(n5502), .ZN(n8959) );
  NAND2_X1 U5318 ( .A1(n5500), .A2(n5499), .ZN(n5503) );
  XNOR2_X1 U5319 ( .A(n5498), .B(n5491), .ZN(n8134) );
  AND2_X1 U5320 ( .A1(n5706), .A2(n4807), .ZN(n4628) );
  XNOR2_X1 U5321 ( .A(n5746), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U5322 ( .A1(n5745), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U5323 ( .A1(n4548), .A2(n5330), .ZN(n5342) );
  NAND2_X1 U5324 ( .A1(n5329), .A2(n5328), .ZN(n4548) );
  XNOR2_X1 U5325 ( .A(n5237), .B(n5236), .ZN(n6688) );
  NAND2_X1 U5326 ( .A1(n4852), .A2(n5138), .ZN(n5154) );
  XNOR2_X1 U5327 ( .A(n5137), .B(n5136), .ZN(n6560) );
  NAND2_X1 U5328 ( .A1(n4406), .A2(n4410), .ZN(n5137) );
  OR2_X1 U5329 ( .A1(n5094), .A2(n4413), .ZN(n4406) );
  AOI21_X1 U5330 ( .B1(n4829), .B2(n5022), .A(n4342), .ZN(n4828) );
  NAND2_X1 U5331 ( .A1(n4518), .A2(n5009), .ZN(n4517) );
  NAND2_X1 U5332 ( .A1(n5442), .A2(n5441), .ZN(n8881) );
  NAND2_X1 U5333 ( .A1(n5371), .A2(n5370), .ZN(n8902) );
  NAND2_X1 U5334 ( .A1(n4712), .A2(n4711), .ZN(n8331) );
  AOI21_X1 U5335 ( .B1(n4714), .B2(n4716), .A(n4341), .ZN(n4711) );
  INV_X1 U5336 ( .A(n8755), .ZN(n8912) );
  AND2_X1 U5337 ( .A1(n5379), .A2(n5378), .ZN(n8713) );
  INV_X2 U5338 ( .A(n8295), .ZN(n8319) );
  AND4_X1 U5339 ( .A1(n5274), .A2(n5273), .A3(n5272), .A4(n5271), .ZN(n8839)
         );
  INV_X1 U5340 ( .A(n8459), .ZN(n8490) );
  NAND2_X1 U5341 ( .A1(n6761), .A2(n6754), .ZN(n8477) );
  AOI21_X1 U5342 ( .B1(n5679), .B2(n8257), .A(n4330), .ZN(n4817) );
  OR2_X1 U5343 ( .A1(n5537), .A2(n6731), .ZN(n4814) );
  INV_X1 U5344 ( .A(n8423), .ZN(n8729) );
  INV_X1 U5345 ( .A(n7167), .ZN(n8501) );
  OR2_X1 U5346 ( .A1(n5000), .A2(n4958), .ZN(n4961) );
  AND2_X1 U5347 ( .A1(n5202), .A2(n5222), .ZN(n8508) );
  XNOR2_X1 U5348 ( .A(n4474), .B(n8628), .ZN(n8874) );
  AOI21_X1 U5349 ( .B1(n8653), .B2(n4319), .A(n4475), .ZN(n4474) );
  INV_X1 U5350 ( .A(n4680), .ZN(n4475) );
  AOI21_X1 U5351 ( .B1(n4319), .B2(n4682), .A(n4343), .ZN(n4680) );
  OR2_X1 U5352 ( .A1(n5298), .A2(n4919), .ZN(n5510) );
  NAND2_X1 U5353 ( .A1(n6159), .A2(n6158), .ZN(n9473) );
  OR2_X1 U5354 ( .A1(n5814), .A2(n5764), .ZN(n5765) );
  NAND2_X1 U5355 ( .A1(n6264), .A2(n6263), .ZN(n9267) );
  NAND2_X1 U5356 ( .A1(n6096), .A2(n6095), .ZN(n9017) );
  AND4_X1 U5357 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n9404)
         );
  NAND2_X1 U5358 ( .A1(n6119), .A2(n6118), .ZN(n9483) );
  NAND2_X1 U5359 ( .A1(n6212), .A2(n6211), .ZN(n9458) );
  AND2_X1 U5360 ( .A1(n6273), .A2(n6272), .ZN(n9280) );
  NOR2_X1 U5361 ( .A1(n8130), .A2(n8119), .ZN(n4523) );
  NAND4_X1 U5362 ( .A1(n5837), .A2(n5836), .A3(n5835), .A4(n5834), .ZN(n9125)
         );
  OR2_X1 U5363 ( .A1(n5804), .A2(n7073), .ZN(n5760) );
  AND2_X1 U5364 ( .A1(n4450), .A2(n4335), .ZN(n9132) );
  NAND2_X1 U5365 ( .A1(n4444), .A2(n4443), .ZN(n4442) );
  OR2_X1 U5366 ( .A1(n9182), .A2(n4380), .ZN(n4444) );
  AOI21_X1 U5367 ( .B1(n9183), .B2(n9959), .A(n9951), .ZN(n4443) );
  OAI21_X1 U5368 ( .B1(n4321), .B2(n4405), .A(n4395), .ZN(n4394) );
  NAND2_X1 U5369 ( .A1(n6349), .A2(n8066), .ZN(n6917) );
  NOR2_X1 U5370 ( .A1(n9208), .A2(n4434), .ZN(n6490) );
  NAND2_X1 U5371 ( .A1(n4435), .A2(n6471), .ZN(n4434) );
  INV_X1 U5372 ( .A(n9201), .ZN(n6471) );
  NAND2_X1 U5373 ( .A1(n9200), .A2(n9986), .ZN(n4435) );
  NAND2_X1 U5374 ( .A1(n4812), .A2(n4630), .ZN(n4811) );
  NAND2_X1 U5375 ( .A1(n9211), .A2(n9986), .ZN(n4812) );
  NOR2_X1 U5376 ( .A1(n9217), .A2(n9212), .ZN(n4630) );
  NAND2_X1 U5377 ( .A1(n9988), .A2(n6450), .ZN(n4629) );
  NAND2_X1 U5378 ( .A1(n6335), .A2(n6334), .ZN(n6507) );
  AND2_X1 U5379 ( .A1(n4807), .A2(n5711), .ZN(n4627) );
  NAND2_X1 U5380 ( .A1(n4483), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U5381 ( .A(n5750), .B(n5749), .ZN(n8070) );
  OAI22_X1 U5382 ( .A1(n5562), .A2(n5561), .B1(n5560), .B2(n5662), .ZN(n5569)
         );
  OAI21_X1 U5383 ( .B1(n5565), .B2(n5564), .A(n5563), .ZN(n5566) );
  INV_X1 U5384 ( .A(n4648), .ZN(n4644) );
  NAND2_X1 U5385 ( .A1(n5579), .A2(n5671), .ZN(n4643) );
  INV_X1 U5386 ( .A(n5613), .ZN(n4638) );
  NAND2_X1 U5387 ( .A1(n4559), .A2(n4558), .ZN(n7904) );
  INV_X1 U5388 ( .A(n7821), .ZN(n4558) );
  OAI21_X1 U5389 ( .B1(n7904), .B2(n4671), .A(n4555), .ZN(n4554) );
  NOR2_X1 U5390 ( .A1(n4556), .A2(n7929), .ZN(n4555) );
  INV_X1 U5391 ( .A(n8107), .ZN(n4556) );
  AOI211_X1 U5392 ( .C1(n5630), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5633)
         );
  OAI21_X1 U5393 ( .B1(n7923), .B2(n7915), .A(n7914), .ZN(n7925) );
  AOI21_X1 U5394 ( .B1(n5645), .B2(n5643), .A(n5642), .ZN(n5644) );
  NAND2_X1 U5395 ( .A1(n4908), .A2(n5063), .ZN(n4631) );
  INV_X1 U5396 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4908) );
  INV_X1 U5397 ( .A(n6401), .ZN(n4826) );
  NOR2_X1 U5398 ( .A1(n9458), .A2(n9328), .ZN(n4672) );
  AND2_X1 U5399 ( .A1(n7853), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5400 ( .A1(n7857), .A2(n4786), .ZN(n4785) );
  INV_X1 U5401 ( .A(n4849), .ZN(n4848) );
  OAI21_X1 U5402 ( .B1(n5469), .B2(n4850), .A(n5487), .ZN(n4849) );
  INV_X1 U5403 ( .A(n5474), .ZN(n4850) );
  INV_X1 U5404 ( .A(n5451), .ZN(n4833) );
  INV_X1 U5405 ( .A(n5328), .ZN(n4544) );
  NOR2_X1 U5406 ( .A1(n5341), .A2(n4547), .ZN(n4546) );
  INV_X1 U5407 ( .A(n5330), .ZN(n4547) );
  INV_X1 U5408 ( .A(n5238), .ZN(n4855) );
  INV_X1 U5409 ( .A(n5259), .ZN(n4854) );
  INV_X1 U5410 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n4505) );
  INV_X1 U5411 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5697) );
  BUF_X1 U5412 ( .A(n8295), .Z(n8309) );
  INV_X1 U5413 ( .A(n6756), .ZN(n6759) );
  OR2_X1 U5414 ( .A1(n8897), .A2(n8423), .ZN(n5646) );
  NAND2_X1 U5415 ( .A1(n4331), .A2(n4318), .ZN(n4685) );
  INV_X1 U5416 ( .A(n4590), .ZN(n4589) );
  NOR2_X1 U5417 ( .A1(n8603), .A2(n4581), .ZN(n4579) );
  INV_X1 U5418 ( .A(n7665), .ZN(n4580) );
  INV_X1 U5419 ( .A(n4705), .ZN(n4704) );
  NAND2_X1 U5420 ( .A1(n9801), .A2(n4578), .ZN(n4581) );
  NAND2_X1 U5421 ( .A1(n5587), .A2(n5585), .ZN(n7523) );
  AND2_X1 U5422 ( .A1(n7125), .A2(n7109), .ZN(n5556) );
  INV_X1 U5423 ( .A(n10007), .ZN(n6750) );
  INV_X1 U5424 ( .A(n4890), .ZN(n4889) );
  INV_X1 U5425 ( .A(n4631), .ZN(n4572) );
  OAI21_X2 U5426 ( .B1(n5514), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5682) );
  NOR2_X1 U5427 ( .A1(n5140), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5163) );
  OAI21_X1 U5428 ( .B1(n5876), .B2(n5897), .A(n6847), .ZN(n4756) );
  NAND2_X1 U5429 ( .A1(n4756), .A2(n4754), .ZN(n4752) );
  NAND2_X1 U5430 ( .A1(n5876), .A2(n5897), .ZN(n4754) );
  NAND2_X1 U5431 ( .A1(n5920), .A2(n6954), .ZN(n5937) );
  INV_X1 U5432 ( .A(n6492), .ZN(n5738) );
  INV_X1 U5433 ( .A(n6413), .ZN(n4393) );
  OR2_X1 U5434 ( .A1(n6968), .A2(n4452), .ZN(n4451) );
  AND2_X1 U5435 ( .A1(n6969), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4452) );
  NOR2_X1 U5436 ( .A1(n5731), .A2(n4323), .ZN(n4862) );
  NAND2_X1 U5437 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n4515) );
  AND2_X1 U5438 ( .A1(n4807), .A2(n5729), .ZN(n4806) );
  INV_X1 U5439 ( .A(n5709), .ZN(n4805) );
  INV_X1 U5440 ( .A(n4621), .ZN(n4619) );
  INV_X1 U5441 ( .A(n4797), .ZN(n4795) );
  AND2_X1 U5442 ( .A1(n7883), .A2(n8008), .ZN(n7959) );
  INV_X1 U5443 ( .A(n6428), .ZN(n4431) );
  INV_X1 U5444 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5445 ( .A1(n4678), .A2(n7762), .ZN(n4677) );
  INV_X1 U5446 ( .A(n4679), .ZN(n4678) );
  NAND2_X1 U5447 ( .A1(n5989), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6012) );
  INV_X1 U5448 ( .A(n5991), .ZN(n5989) );
  NAND2_X1 U5449 ( .A1(n4748), .A2(n4839), .ZN(n8082) );
  NAND2_X1 U5450 ( .A1(n6710), .A2(n6418), .ZN(n8086) );
  NOR2_X1 U5451 ( .A1(n9227), .A2(n4665), .ZN(n6468) );
  OR2_X1 U5452 ( .A1(n9227), .A2(n6479), .ZN(n9229) );
  AND2_X1 U5453 ( .A1(n9336), .A2(n4668), .ZN(n9281) );
  NOR2_X1 U5454 ( .A1(n9282), .A2(n4670), .ZN(n4668) );
  NAND2_X1 U5455 ( .A1(n9336), .A2(n4672), .ZN(n9308) );
  NAND2_X1 U5456 ( .A1(n9336), .A2(n9518), .ZN(n9325) );
  NAND2_X1 U5457 ( .A1(n4675), .A2(n4674), .ZN(n7739) );
  NOR2_X1 U5458 ( .A1(n4677), .A2(n7797), .ZN(n4674) );
  INV_X1 U5459 ( .A(n7447), .ZN(n4675) );
  NAND2_X1 U5460 ( .A1(n7225), .A2(n4626), .ZN(n6999) );
  AND2_X1 U5461 ( .A1(n7824), .A2(n6381), .ZN(n4626) );
  AOI21_X1 U5462 ( .B1(n4531), .B2(n4530), .A(n4365), .ZN(n4529) );
  INV_X1 U5463 ( .A(n4537), .ZN(n4530) );
  NOR2_X1 U5464 ( .A1(n4856), .A2(n4538), .ZN(n4537) );
  INV_X1 U5465 ( .A(n5216), .ZN(n4538) );
  INV_X1 U5466 ( .A(n4535), .ZN(n4534) );
  OAI21_X1 U5467 ( .B1(n4856), .B2(n4536), .A(n4853), .ZN(n4535) );
  NAND2_X1 U5468 ( .A1(n4539), .A2(n5216), .ZN(n4536) );
  AOI21_X1 U5469 ( .B1(n4857), .B2(n4855), .A(n4854), .ZN(n4853) );
  AND2_X1 U5470 ( .A1(n5259), .A2(n5241), .ZN(n5257) );
  INV_X1 U5471 ( .A(SI_14_), .ZN(n5196) );
  NAND2_X1 U5472 ( .A1(n5194), .A2(n5193), .ZN(n4429) );
  NAND2_X1 U5473 ( .A1(n4409), .A2(n4407), .ZN(n4852) );
  AOI21_X1 U5474 ( .B1(n4410), .B2(n4413), .A(n4408), .ZN(n4407) );
  INV_X1 U5475 ( .A(n5136), .ZN(n4408) );
  INV_X1 U5476 ( .A(n4415), .ZN(n4413) );
  AOI21_X1 U5477 ( .B1(n4415), .B2(n4412), .A(n4411), .ZN(n4410) );
  INV_X1 U5478 ( .A(n5120), .ZN(n4411) );
  INV_X1 U5479 ( .A(n5095), .ZN(n4412) );
  NOR2_X1 U5480 ( .A1(n4427), .A2(n4424), .ZN(n4423) );
  INV_X1 U5481 ( .A(n5065), .ZN(n4427) );
  INV_X1 U5482 ( .A(n5045), .ZN(n4424) );
  INV_X1 U5483 ( .A(n5048), .ZN(n4426) );
  NOR2_X1 U5484 ( .A1(n4519), .A2(n4827), .ZN(n4518) );
  INV_X1 U5485 ( .A(n5008), .ZN(n4827) );
  INV_X1 U5486 ( .A(n5011), .ZN(n4829) );
  NAND2_X1 U5487 ( .A1(n4438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5816) );
  INV_X1 U5488 ( .A(n5783), .ZN(n4438) );
  INV_X1 U5489 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4947) );
  INV_X1 U5490 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4948) );
  INV_X1 U5491 ( .A(SI_20_), .ZN(n9633) );
  INV_X1 U5492 ( .A(SI_16_), .ZN(n9738) );
  NAND2_X1 U5493 ( .A1(n8479), .A2(n4719), .ZN(n4713) );
  AND2_X1 U5494 ( .A1(n4718), .A2(n8346), .ZN(n4717) );
  NAND2_X1 U5495 ( .A1(n4719), .A2(n8478), .ZN(n4718) );
  AOI21_X1 U5496 ( .B1(n4717), .B2(n4720), .A(n4715), .ZN(n4714) );
  INV_X1 U5497 ( .A(n8325), .ZN(n4715) );
  INV_X1 U5498 ( .A(n4717), .ZN(n4716) );
  OR2_X1 U5499 ( .A1(n5072), .A2(n9719), .ZN(n5109) );
  INV_X1 U5500 ( .A(n5386), .ZN(n5385) );
  INV_X1 U5501 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9735) );
  INV_X1 U5502 ( .A(n5350), .ZN(n5352) );
  NOR2_X1 U5503 ( .A1(n8413), .A2(n4738), .ZN(n4737) );
  INV_X1 U5504 ( .A(n8266), .ZN(n4738) );
  OR2_X1 U5505 ( .A1(n5283), .A2(n9650), .ZN(n5304) );
  OR2_X1 U5506 ( .A1(n5205), .A2(n9582), .ZN(n5229) );
  AOI21_X1 U5507 ( .B1(n4724), .B2(n4726), .A(n4723), .ZN(n4722) );
  INV_X1 U5508 ( .A(n7716), .ZN(n4723) );
  NAND2_X1 U5509 ( .A1(n4876), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U5510 ( .A1(n4874), .A2(n4873), .ZN(n4872) );
  INV_X1 U5511 ( .A(n5673), .ZN(n4876) );
  NOR2_X1 U5512 ( .A1(n8596), .A2(n4329), .ZN(n4874) );
  INV_X1 U5513 ( .A(n4869), .ZN(n4868) );
  OAI21_X1 U5514 ( .B1(n4871), .B2(n4873), .A(n5670), .ZN(n4869) );
  NOR2_X1 U5515 ( .A1(n5678), .A2(n4864), .ZN(n5535) );
  AND4_X1 U5516 ( .A1(n5061), .A2(n5060), .A3(n5059), .A4(n5058), .ZN(n7413)
         );
  AND4_X1 U5517 ( .A1(n5043), .A2(n5042), .A3(n5041), .A4(n5040), .ZN(n7167)
         );
  AOI21_X1 U5518 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6809), .A(n8238), .ZN(
        n9778) );
  NOR2_X1 U5519 ( .A1(n8216), .A2(n4549), .ZN(n8207) );
  NOR2_X1 U5520 ( .A1(n8226), .A2(n6814), .ZN(n4549) );
  NOR2_X1 U5521 ( .A1(n8183), .A2(n4361), .ZN(n8174) );
  NOR2_X1 U5522 ( .A1(n8174), .A2(n8173), .ZN(n8172) );
  NOR2_X1 U5523 ( .A1(n8152), .A2(n8151), .ZN(n8150) );
  NOR2_X1 U5524 ( .A1(n8150), .A2(n4561), .ZN(n6826) );
  AND2_X1 U5525 ( .A1(n6825), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4561) );
  NOR2_X1 U5526 ( .A1(n6826), .A2(n6827), .ZN(n6982) );
  NOR2_X1 U5527 ( .A1(n6982), .A2(n4560), .ZN(n8141) );
  AND2_X1 U5528 ( .A1(n6983), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4560) );
  NAND2_X1 U5529 ( .A1(n8140), .A2(n4551), .ZN(n6986) );
  OR2_X1 U5530 ( .A1(n6985), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4551) );
  NAND2_X1 U5531 ( .A1(n6986), .A2(n6987), .ZN(n7207) );
  NAND2_X1 U5532 ( .A1(n7207), .A2(n4550), .ZN(n7209) );
  OR2_X1 U5533 ( .A1(n7208), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4550) );
  INV_X1 U5534 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5197) );
  INV_X1 U5535 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U5536 ( .A1(n8546), .A2(n8547), .ZN(n8548) );
  NOR2_X1 U5537 ( .A1(n8548), .A2(n8549), .ZN(n8558) );
  AOI21_X1 U5538 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8559), .A(n8558), .ZN(
        n8562) );
  NAND2_X1 U5539 ( .A1(n4348), .A2(n5658), .ZN(n4893) );
  NAND2_X1 U5540 ( .A1(n8652), .A2(n5656), .ZN(n4896) );
  NOR3_X1 U5541 ( .A1(n8690), .A2(n8876), .A3(n4585), .ZN(n8643) );
  NOR2_X1 U5542 ( .A1(n8690), .A2(n4585), .ZN(n8655) );
  NAND2_X1 U5543 ( .A1(n8684), .A2(n8615), .ZN(n8667) );
  OR2_X1 U5544 ( .A1(n8893), .A2(n8614), .ZN(n8615) );
  AND2_X1 U5545 ( .A1(n8723), .A2(n8706), .ZN(n8701) );
  NOR2_X1 U5546 ( .A1(n8734), .A2(n8902), .ZN(n8723) );
  OAI21_X1 U5547 ( .B1(n4903), .B2(n4318), .A(n4691), .ZN(n4690) );
  AOI21_X1 U5548 ( .B1(n4478), .B2(n4477), .A(n4476), .ZN(n8768) );
  NAND2_X1 U5549 ( .A1(n8925), .A2(n8807), .ZN(n4477) );
  NOR2_X1 U5550 ( .A1(n8925), .A2(n8807), .ZN(n4476) );
  INV_X1 U5551 ( .A(n8779), .ZN(n4478) );
  NOR3_X1 U5552 ( .A1(n8823), .A2(n4590), .A3(n8919), .ZN(n8772) );
  NOR2_X1 U5553 ( .A1(n8823), .A2(n4590), .ZN(n8780) );
  AND2_X1 U5554 ( .A1(n5623), .A2(n8763), .ZN(n8787) );
  OR2_X1 U5555 ( .A1(n5249), .A2(n9735), .ZN(n5269) );
  NAND2_X1 U5556 ( .A1(n5268), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5283) );
  INV_X1 U5557 ( .A(n5269), .ZN(n5268) );
  AND4_X1 U5558 ( .A1(n5234), .A2(n5233), .A3(n5232), .A4(n5231), .ZN(n8841)
         );
  NAND2_X1 U5559 ( .A1(n4580), .A2(n4579), .ZN(n8855) );
  NOR2_X1 U5560 ( .A1(n7665), .A2(n4581), .ZN(n7782) );
  NOR2_X1 U5561 ( .A1(n7665), .A2(n7681), .ZN(n7692) );
  AND4_X1 U5562 ( .A1(n5211), .A2(n5210), .A3(n5209), .A4(n5208), .ZN(n7781)
         );
  NAND2_X1 U5563 ( .A1(n4882), .A2(n7653), .ZN(n7656) );
  AND2_X1 U5564 ( .A1(n7609), .A2(n7525), .ZN(n7527) );
  NAND2_X1 U5565 ( .A1(n4479), .A2(n7522), .ZN(n7607) );
  NAND2_X1 U5566 ( .A1(n7523), .A2(n7557), .ZN(n4479) );
  AND4_X1 U5567 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n8451)
         );
  AND2_X1 U5568 ( .A1(n7566), .A2(n10079), .ZN(n7603) );
  INV_X1 U5569 ( .A(n7523), .ZN(n7560) );
  AND4_X1 U5570 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n8390)
         );
  OR2_X1 U5571 ( .A1(n7425), .A2(n10064), .ZN(n7548) );
  NOR2_X1 U5572 ( .A1(n7548), .A2(n7554), .ZN(n7566) );
  NOR2_X1 U5573 ( .A1(n4885), .A2(n4884), .ZN(n4883) );
  INV_X1 U5574 ( .A(n5573), .ZN(n4884) );
  OR2_X1 U5575 ( .A1(n7417), .A2(n7416), .ZN(n7538) );
  OR2_X1 U5576 ( .A1(n5056), .A2(n5055), .ZN(n5072) );
  NAND2_X1 U5577 ( .A1(n7171), .A2(n10059), .ZN(n7425) );
  NOR2_X1 U5578 ( .A1(n7142), .A2(n10049), .ZN(n7171) );
  NAND2_X1 U5579 ( .A1(n7128), .A2(n7125), .ZN(n7113) );
  NOR2_X1 U5580 ( .A1(n7069), .A2(n10022), .ZN(n7094) );
  OR2_X1 U5581 ( .A1(n5090), .A2(n6514), .ZN(n4956) );
  NAND2_X1 U5582 ( .A1(n5423), .A2(n5422), .ZN(n8888) );
  NAND2_X1 U5583 ( .A1(n5348), .A2(n5347), .ZN(n8907) );
  NAND2_X1 U5584 ( .A1(n5282), .A2(n5281), .ZN(n8929) );
  NAND2_X1 U5585 ( .A1(n4457), .A2(n4459), .ZN(n8814) );
  NAND2_X1 U5586 ( .A1(n4456), .A2(n8607), .ZN(n4459) );
  NAND2_X1 U5587 ( .A1(n8605), .A2(n4461), .ZN(n4457) );
  XNOR2_X1 U5588 ( .A(n5688), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U5589 ( .A1(n5687), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U5590 ( .A1(n5686), .A2(n5685), .ZN(n5687) );
  XNOR2_X1 U5591 ( .A(n5686), .B(P2_IR_REG_23__SCAN_IN), .ZN(n6875) );
  INV_X1 U5592 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5101) );
  AND2_X1 U5593 ( .A1(n5030), .A2(n5029), .ZN(n6816) );
  NOR2_X1 U5594 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n4867) );
  AND2_X1 U5595 ( .A1(n4975), .A2(n4697), .ZN(n4944) );
  INV_X1 U5596 ( .A(n4769), .ZN(n4766) );
  AND2_X1 U5597 ( .A1(n4767), .A2(n4764), .ZN(n4763) );
  NAND2_X1 U5598 ( .A1(n4769), .A2(n4765), .ZN(n4764) );
  CLKBUF_X1 U5599 ( .A(n5825), .Z(n6326) );
  NAND2_X1 U5600 ( .A1(n5774), .A2(n5740), .ZN(n5768) );
  AND2_X1 U5601 ( .A1(n4760), .A2(n9040), .ZN(n4758) );
  NAND2_X1 U5602 ( .A1(n9039), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5603 ( .A1(n5868), .A2(n4507), .ZN(n5869) );
  NAND2_X1 U5604 ( .A1(n4509), .A2(n4508), .ZN(n4507) );
  OR2_X1 U5605 ( .A1(n6245), .A2(n9034), .ZN(n6267) );
  XNOR2_X1 U5606 ( .A(n5846), .B(n7030), .ZN(n5849) );
  INV_X1 U5607 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5948) );
  INV_X1 U5608 ( .A(n6214), .ZN(n6213) );
  INV_X1 U5609 ( .A(n5798), .ZN(n5800) );
  AOI21_X1 U5610 ( .B1(n9033), .B2(n4778), .A(n4516), .ZN(n9075) );
  NAND2_X1 U5611 ( .A1(n4497), .A2(n4501), .ZN(n4491) );
  NOR2_X1 U5612 ( .A1(n4490), .A2(n4488), .ZN(n4487) );
  NAND2_X1 U5613 ( .A1(n4500), .A2(n4498), .ZN(n4492) );
  AOI211_X1 U5614 ( .C1(n8068), .C2(n8067), .A(n8066), .B(n8119), .ZN(n8069)
         );
  AND4_X1 U5615 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n7442)
         );
  OR2_X1 U5616 ( .A1(n5804), .A2(n5787), .ZN(n5790) );
  NAND2_X1 U5617 ( .A1(n5878), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5788) );
  OR2_X1 U5618 ( .A1(n5805), .A2(n6534), .ZN(n5761) );
  NAND2_X1 U5619 ( .A1(n4437), .A2(n4436), .ZN(n9894) );
  OR2_X1 U5620 ( .A1(n6548), .A2(n6533), .ZN(n4437) );
  NAND2_X1 U5621 ( .A1(n6548), .A2(n6533), .ZN(n4436) );
  NAND2_X1 U5622 ( .A1(n9895), .A2(n9894), .ZN(n9893) );
  NOR2_X1 U5623 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  INV_X1 U5624 ( .A(n5944), .ZN(n5984) );
  NOR2_X1 U5625 ( .A1(n6696), .A2(n4453), .ZN(n6700) );
  AND2_X1 U5626 ( .A1(n6697), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4453) );
  NOR2_X1 U5627 ( .A1(n6700), .A2(n6699), .ZN(n6968) );
  XNOR2_X1 U5628 ( .A(n4451), .B(n7380), .ZN(n6970) );
  AND2_X1 U5629 ( .A1(n4440), .A2(n4439), .ZN(n9158) );
  NAND2_X1 U5630 ( .A1(n9160), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4439) );
  NOR2_X1 U5631 ( .A1(n9158), .A2(n9157), .ZN(n9170) );
  NAND2_X1 U5632 ( .A1(n4664), .A2(n9497), .ZN(n4663) );
  INV_X1 U5633 ( .A(n4665), .ZN(n4664) );
  NOR3_X1 U5634 ( .A1(n9227), .A2(n6470), .A3(n4665), .ZN(n9195) );
  NAND2_X1 U5635 ( .A1(n4321), .A2(n4396), .ZN(n4395) );
  NAND2_X1 U5636 ( .A1(n4404), .A2(n7989), .ZN(n4396) );
  NAND2_X1 U5637 ( .A1(n4400), .A2(n4405), .ZN(n4399) );
  INV_X1 U5638 ( .A(n4404), .ZN(n4400) );
  NAND2_X1 U5639 ( .A1(n4599), .A2(n4597), .ZN(n6410) );
  INV_X1 U5640 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5641 ( .B1(n4601), .B2(n9225), .A(n6409), .ZN(n4598) );
  NOR2_X1 U5642 ( .A1(n6410), .A2(n7987), .ZN(n6454) );
  AND2_X1 U5643 ( .A1(n6360), .A2(n6359), .ZN(n7944) );
  NAND2_X1 U5644 ( .A1(n4401), .A2(n4402), .ZN(n6460) );
  AND2_X1 U5645 ( .A1(n6321), .A2(n6320), .ZN(n9222) );
  AND2_X1 U5646 ( .A1(n6313), .A2(n6283), .ZN(n9249) );
  AND2_X1 U5647 ( .A1(n6304), .A2(n6303), .ZN(n9243) );
  AND2_X1 U5648 ( .A1(n4822), .A2(n4612), .ZN(n4611) );
  INV_X1 U5649 ( .A(n4823), .ZN(n4822) );
  NAND2_X1 U5650 ( .A1(n9343), .A2(n7889), .ZN(n9319) );
  AND2_X1 U5651 ( .A1(n9356), .A2(n9342), .ZN(n9336) );
  INV_X1 U5652 ( .A(n6141), .ZN(n6139) );
  NOR2_X1 U5653 ( .A1(n9376), .A2(n9473), .ZN(n9356) );
  INV_X1 U5654 ( .A(n7959), .ZN(n9362) );
  INV_X1 U5655 ( .A(n6098), .ZN(n6097) );
  OR2_X1 U5656 ( .A1(n6121), .A2(n9024), .ZN(n6141) );
  AOI21_X1 U5657 ( .B1(n4594), .B2(n4596), .A(n4363), .ZN(n4592) );
  INV_X1 U5658 ( .A(n6057), .ZN(n6055) );
  INV_X1 U5659 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6032) );
  OR2_X1 U5660 ( .A1(n6033), .A2(n6032), .ZN(n6057) );
  NOR2_X1 U5661 ( .A1(n7447), .A2(n4679), .ZN(n7753) );
  OR2_X1 U5662 ( .A1(n7394), .A2(n7398), .ZN(n7447) );
  OR2_X1 U5663 ( .A1(n5949), .A2(n5948), .ZN(n5968) );
  INV_X1 U5664 ( .A(n4789), .ZN(n4788) );
  OAI21_X1 U5665 ( .B1(n4332), .B2(n4790), .A(n7841), .ZN(n4789) );
  INV_X1 U5666 ( .A(n6426), .ZN(n4790) );
  AND2_X1 U5667 ( .A1(n7842), .A2(n7845), .ZN(n7972) );
  NAND2_X1 U5668 ( .A1(n7245), .A2(n6426), .ZN(n7243) );
  AND2_X1 U5669 ( .A1(n7238), .A2(n7308), .ZN(n7317) );
  NOR2_X1 U5670 ( .A1(n7036), .A2(n7037), .ZN(n7238) );
  OR2_X1 U5671 ( .A1(n7226), .A2(n9413), .ZN(n7036) );
  NOR2_X1 U5672 ( .A1(n7335), .A2(n6889), .ZN(n7227) );
  NAND2_X1 U5673 ( .A1(n7227), .A2(n9976), .ZN(n7226) );
  NAND2_X1 U5674 ( .A1(n8089), .A2(n8023), .ZN(n7961) );
  INV_X1 U5675 ( .A(n6707), .ZN(n7967) );
  NAND2_X1 U5676 ( .A1(n7935), .A2(n7934), .ZN(n9189) );
  NAND2_X1 U5677 ( .A1(n7938), .A2(n7937), .ZN(n9188) );
  NAND2_X1 U5678 ( .A1(n6280), .A2(n6279), .ZN(n9248) );
  INV_X1 U5679 ( .A(n4509), .ZN(n9976) );
  INV_X1 U5680 ( .A(n9982), .ZN(n9843) );
  AND2_X1 U5681 ( .A1(n6448), .A2(n6447), .ZN(n6486) );
  XNOR2_X1 U5682 ( .A(n5488), .B(n5487), .ZN(n8132) );
  NAND2_X1 U5683 ( .A1(n4847), .A2(n5474), .ZN(n5488) );
  XNOR2_X1 U5684 ( .A(n5470), .B(n5469), .ZN(n8966) );
  XNOR2_X1 U5685 ( .A(n5452), .B(n5451), .ZN(n7807) );
  XNOR2_X1 U5686 ( .A(n5435), .B(n5434), .ZN(n7802) );
  NAND2_X1 U5687 ( .A1(n5417), .A2(n5416), .ZN(n5435) );
  NAND2_X1 U5688 ( .A1(n5731), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5734) );
  INV_X1 U5689 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5735) );
  INV_X1 U5690 ( .A(n5724), .ZN(n5725) );
  NAND2_X1 U5691 ( .A1(n4843), .A2(n5294), .ZN(n5310) );
  OR2_X1 U5692 ( .A1(n6112), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n6113) );
  OR2_X1 U5693 ( .A1(n6028), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U5694 ( .A1(n4414), .A2(n5095), .ZN(n5119) );
  OR2_X1 U5695 ( .A1(n5094), .A2(n5093), .ZN(n4414) );
  XNOR2_X1 U5696 ( .A(n5816), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6548) );
  XNOR2_X1 U5697 ( .A(n5763), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6546) );
  INV_X1 U5698 ( .A(n7252), .ZN(n10059) );
  AND2_X1 U5699 ( .A1(n5460), .A2(n5444), .ZN(n8656) );
  AND4_X1 U5700 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n7590)
         );
  OR2_X1 U5701 ( .A1(n4313), .A2(n9625), .ZN(n4939) );
  NAND2_X1 U5702 ( .A1(n8364), .A2(n8279), .ZN(n8365) );
  AND2_X1 U5703 ( .A1(n7285), .A2(n7024), .ZN(n4729) );
  NAND2_X1 U5704 ( .A1(n4382), .A2(n4381), .ZN(n6734) );
  INV_X1 U5705 ( .A(n6732), .ZN(n4381) );
  INV_X1 U5706 ( .A(n6733), .ZN(n4382) );
  NAND2_X1 U5707 ( .A1(n5166), .A2(n5165), .ZN(n8398) );
  NAND3_X1 U5708 ( .A1(n4383), .A2(n8307), .A3(n4362), .ZN(n8403) );
  NAND2_X1 U5709 ( .A1(n8267), .A2(n8266), .ZN(n8414) );
  NAND2_X1 U5710 ( .A1(n8365), .A2(n8283), .ZN(n8433) );
  AND4_X1 U5711 ( .A1(n5173), .A2(n5172), .A3(n5171), .A4(n5170), .ZN(n7660)
         );
  AND2_X1 U5712 ( .A1(n8335), .A2(n8806), .ZN(n8460) );
  AND2_X1 U5713 ( .A1(n8335), .A2(n8804), .ZN(n8461) );
  AOI21_X1 U5714 ( .B1(n6904), .B2(n4732), .A(n4731), .ZN(n7286) );
  INV_X1 U5715 ( .A(n8477), .ZN(n8441) );
  NAND2_X1 U5716 ( .A1(n6757), .A2(n8852), .ZN(n8459) );
  NOR2_X1 U5717 ( .A1(n4379), .A2(n5536), .ZN(n4818) );
  INV_X1 U5718 ( .A(P2_U3966), .ZN(n8492) );
  INV_X1 U5719 ( .A(n8612), .ZN(n8758) );
  INV_X1 U5720 ( .A(n7413), .ZN(n8500) );
  INV_X1 U5721 ( .A(n7118), .ZN(n8503) );
  AOI21_X1 U5722 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6813), .A(n8227), .ZN(
        n8218) );
  NOR2_X1 U5723 ( .A1(n8218), .A2(n8217), .ZN(n8216) );
  AOI21_X1 U5724 ( .B1(n6818), .B2(P2_REG1_REG_6__SCAN_IN), .A(n8194), .ZN(
        n8185) );
  NOR2_X1 U5725 ( .A1(n8185), .A2(n8184), .ZN(n8183) );
  AOI21_X1 U5726 ( .B1(n6821), .B2(P2_REG1_REG_8__SCAN_IN), .A(n8172), .ZN(
        n8163) );
  NOR2_X1 U5727 ( .A1(n8521), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U5728 ( .A1(n8524), .A2(n8523), .ZN(n8546) );
  AND2_X1 U5729 ( .A1(n6802), .A2(n6801), .ZN(n9997) );
  NAND2_X1 U5730 ( .A1(n5507), .A2(n5506), .ZN(n8862) );
  NAND2_X1 U5731 ( .A1(n5493), .A2(n5492), .ZN(n8865) );
  OAI21_X1 U5732 ( .B1(n8653), .B2(n4682), .A(n4319), .ZN(n8640) );
  NAND2_X1 U5733 ( .A1(n8651), .A2(n8619), .ZN(n8642) );
  NAND2_X1 U5734 ( .A1(n4895), .A2(n5656), .ZN(n8637) );
  NAND2_X1 U5735 ( .A1(n4887), .A2(n5641), .ZN(n8678) );
  NAND2_X1 U5736 ( .A1(n4466), .A2(n4471), .ZN(n8685) );
  NAND2_X1 U5737 ( .A1(n8720), .A2(n4470), .ZN(n4466) );
  NAND2_X1 U5738 ( .A1(n8720), .A2(n4472), .ZN(n8700) );
  AND2_X1 U5739 ( .A1(n4688), .A2(n4693), .ZN(n8722) );
  NAND2_X1 U5740 ( .A1(n4686), .A2(n4331), .ZN(n4688) );
  INV_X1 U5741 ( .A(n4692), .ZN(n4686) );
  AND2_X1 U5742 ( .A1(n5332), .A2(n5331), .ZN(n8755) );
  AND2_X1 U5743 ( .A1(n4878), .A2(n5539), .ZN(n8803) );
  NAND2_X1 U5744 ( .A1(n5256), .A2(n5611), .ZN(n8816) );
  NAND2_X1 U5745 ( .A1(n5265), .A2(n5264), .ZN(n8934) );
  INV_X1 U5746 ( .A(n4456), .ZN(n4463) );
  NOR2_X1 U5747 ( .A1(n7682), .A2(n4899), .ZN(n7684) );
  OR2_X1 U5748 ( .A1(n7682), .A2(n4705), .ZN(n7777) );
  NAND2_X1 U5749 ( .A1(n4465), .A2(n5125), .ZN(n7578) );
  NAND2_X1 U5750 ( .A1(n6560), .A2(n5100), .ZN(n4465) );
  INV_X1 U5751 ( .A(n10072), .ZN(n7554) );
  NAND2_X1 U5752 ( .A1(n10053), .A2(n7162), .ZN(n7164) );
  AND2_X1 U5753 ( .A1(n7116), .A2(n7117), .ZN(n4700) );
  INV_X1 U5754 ( .A(n4660), .ZN(n4658) );
  OAI21_X1 U5755 ( .B1(n5505), .B2(n6506), .A(n5031), .ZN(n4660) );
  NAND2_X1 U5756 ( .A1(n8831), .A2(n6946), .ZN(n8800) );
  NAND2_X1 U5757 ( .A1(n10008), .A2(n7180), .ZN(n8852) );
  CLKBUF_X1 U5758 ( .A(n6859), .Z(n7069) );
  NAND2_X1 U5759 ( .A1(n6804), .A2(n8975), .ZN(n4574) );
  INV_X1 U5760 ( .A(n8800), .ZN(n8854) );
  AND2_X1 U5761 ( .A1(n6947), .A2(n8319), .ZN(n8856) );
  AND2_X2 U5762 ( .A1(n7185), .A2(n7184), .ZN(n10120) );
  NAND2_X1 U5763 ( .A1(n8873), .A2(n4385), .ZN(n8945) );
  OR2_X1 U5764 ( .A1(n8874), .A2(n10085), .ZN(n4385) );
  NOR2_X1 U5765 ( .A1(n6875), .A2(P2_U3152), .ZN(n10013) );
  NAND2_X1 U5766 ( .A1(n4943), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4917) );
  XNOR2_X1 U5767 ( .A(n5690), .B(P2_IR_REG_26__SCAN_IN), .ZN(n7801) );
  INV_X1 U5768 ( .A(n6739), .ZN(n7702) );
  INV_X1 U5769 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7635) );
  INV_X1 U5770 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8344) );
  INV_X1 U5771 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7388) );
  INV_X1 U5772 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8259) );
  NAND2_X1 U5773 ( .A1(n5511), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  OAI21_X1 U5774 ( .B1(n4736), .B2(n4919), .A(n4735), .ZN(n5511) );
  INV_X1 U5775 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7179) );
  INV_X1 U5776 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6691) );
  INV_X1 U5777 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6642) );
  INV_X1 U5778 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6610) );
  INV_X1 U5779 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6531) );
  INV_X1 U5780 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6525) );
  INV_X1 U5781 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6517) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U5783 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4563) );
  NOR2_X1 U5784 ( .A1(n6492), .A2(n6491), .ZN(n9890) );
  CLKBUF_X1 U5785 ( .A(n6953), .Z(n6957) );
  AOI21_X1 U5786 ( .B1(n4775), .B2(n4516), .A(n4774), .ZN(n4773) );
  INV_X1 U5787 ( .A(n6473), .ZN(n4774) );
  NAND2_X1 U5788 ( .A1(n4495), .A2(n4499), .ZN(n7791) );
  NAND2_X1 U5789 ( .A1(n4496), .A2(n6068), .ZN(n7790) );
  INV_X1 U5790 ( .A(n6068), .ZN(n4499) );
  NAND2_X1 U5791 ( .A1(n6156), .A2(n9067), .ZN(n8985) );
  XNOR2_X1 U5792 ( .A(n5936), .B(n7030), .ZN(n7264) );
  CLKBUF_X1 U5793 ( .A(n6627), .Z(n6628) );
  CLKBUF_X1 U5794 ( .A(n8991), .Z(n8992) );
  CLKBUF_X1 U5795 ( .A(n7636), .Z(n7637) );
  NAND2_X1 U5796 ( .A1(n4749), .A2(n6005), .ZN(n7639) );
  INV_X1 U5797 ( .A(n4779), .ZN(n9001) );
  INV_X1 U5798 ( .A(n6668), .ZN(n4743) );
  CLKBUF_X1 U5799 ( .A(n6722), .Z(n6769) );
  CLKBUF_X1 U5800 ( .A(n7363), .Z(n7364) );
  NAND2_X1 U5801 ( .A1(n4759), .A2(n6174), .ZN(n9042) );
  NAND2_X1 U5802 ( .A1(n6176), .A2(n6175), .ZN(n9467) );
  AND4_X1 U5803 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n7757)
         );
  OR2_X1 U5804 ( .A1(n4768), .A2(n6226), .ZN(n9049) );
  NAND2_X1 U5805 ( .A1(n6138), .A2(n6137), .ZN(n9378) );
  NAND2_X1 U5806 ( .A1(n6363), .A2(n9861), .ZN(n9094) );
  AND2_X1 U5807 ( .A1(n6362), .A2(n6351), .ZN(n9080) );
  INV_X1 U5808 ( .A(n9222), .ZN(n9107) );
  INV_X1 U5809 ( .A(n9243), .ZN(n9108) );
  OR3_X1 U5810 ( .A1(n6184), .A2(n6183), .A3(n6182), .ZN(n9321) );
  OR2_X1 U5811 ( .A1(n5804), .A2(n6918), .ZN(n5721) );
  NOR2_X1 U5812 ( .A1(n9906), .A2(n6535), .ZN(n9927) );
  NOR2_X1 U5813 ( .A1(n7495), .A2(n7496), .ZN(n7499) );
  INV_X1 U5814 ( .A(n4440), .ZN(n9155) );
  AND2_X1 U5815 ( .A1(n9179), .A2(n6555), .ZN(n9959) );
  OAI21_X1 U5816 ( .B1(n9964), .B2(n9187), .A(n9186), .ZN(n4446) );
  NOR2_X1 U5817 ( .A1(n6454), .A2(n6411), .ZN(n9211) );
  AND2_X1 U5818 ( .A1(n6410), .A2(n7987), .ZN(n6411) );
  NAND2_X1 U5819 ( .A1(n4600), .A2(n4604), .ZN(n9226) );
  OR2_X1 U5820 ( .A1(n9255), .A2(n4606), .ZN(n4600) );
  NAND2_X1 U5821 ( .A1(n4609), .A2(n6408), .ZN(n9236) );
  NAND2_X1 U5822 ( .A1(n9255), .A2(n9257), .ZN(n4609) );
  NAND2_X1 U5823 ( .A1(n4620), .A2(n4621), .ZN(n9274) );
  NAND2_X1 U5824 ( .A1(n4803), .A2(n8003), .ZN(n9278) );
  NAND2_X1 U5825 ( .A1(n6433), .A2(n7900), .ZN(n9291) );
  OAI21_X1 U5826 ( .B1(n9302), .B2(n4358), .A(n4625), .ZN(n9289) );
  OAI21_X1 U5827 ( .B1(n9343), .B2(n6432), .A(n4420), .ZN(n9303) );
  NAND2_X1 U5828 ( .A1(n4821), .A2(n6401), .ZN(n9335) );
  OR2_X1 U5829 ( .A1(n9355), .A2(n4352), .ZN(n4821) );
  NAND2_X1 U5830 ( .A1(n6430), .A2(n4797), .ZN(n9369) );
  NAND2_X1 U5831 ( .A1(n6430), .A2(n8011), .ZN(n9399) );
  INV_X1 U5832 ( .A(n4593), .ZN(n7813) );
  AOI21_X1 U5833 ( .B1(n7727), .B2(n4841), .A(n4596), .ZN(n4593) );
  NAND2_X1 U5834 ( .A1(n7723), .A2(n6429), .ZN(n7734) );
  NAND2_X1 U5835 ( .A1(n6075), .A2(n6074), .ZN(n9100) );
  OAI21_X1 U5836 ( .B1(n7727), .B2(n4322), .A(n6395), .ZN(n7737) );
  NAND2_X1 U5837 ( .A1(n6428), .A2(n7856), .ZN(n7724) );
  NAND2_X1 U5838 ( .A1(n6031), .A2(n6030), .ZN(n9830) );
  NAND2_X1 U5839 ( .A1(n7441), .A2(n7857), .ZN(n7622) );
  NAND2_X1 U5840 ( .A1(n5987), .A2(n5986), .ZN(n9844) );
  NAND2_X1 U5841 ( .A1(n7028), .A2(n6383), .ZN(n7237) );
  NAND2_X1 U5842 ( .A1(n6424), .A2(n6423), .ZN(n7033) );
  INV_X1 U5843 ( .A(n7008), .ZN(n9413) );
  INV_X1 U5844 ( .A(n9392), .ZN(n9831) );
  INV_X1 U5845 ( .A(n9199), .ZN(n9818) );
  NAND2_X1 U5846 ( .A1(n6887), .A2(n6380), .ZN(n7223) );
  INV_X1 U5847 ( .A(n9408), .ZN(n9414) );
  NAND2_X1 U5848 ( .A1(n6709), .A2(n6377), .ZN(n6676) );
  NAND2_X1 U5849 ( .A1(n9409), .A2(n6916), .ZN(n9392) );
  OR2_X1 U5850 ( .A1(n9390), .A2(n6354), .ZN(n9820) );
  MUX2_X1 U5851 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9539), .S(n5814), .Z(n6920) );
  INV_X1 U5852 ( .A(n9189), .ZN(n9494) );
  INV_X1 U5853 ( .A(n9188), .ZN(n9497) );
  INV_X1 U5854 ( .A(n9248), .ZN(n9504) );
  INV_X1 U5855 ( .A(n9267), .ZN(n9508) );
  AND3_X1 U5856 ( .A1(n5904), .A2(n5903), .A3(n5902), .ZN(n7352) );
  INV_X1 U5857 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5714) );
  OR2_X1 U5858 ( .A1(n5713), .A2(n5899), .ZN(n5712) );
  OR2_X1 U5859 ( .A1(n5728), .A2(n5899), .ZN(n5730) );
  AND2_X1 U5860 ( .A1(n4628), .A2(n5707), .ZN(n5728) );
  XNOR2_X1 U5861 ( .A(n5381), .B(n5380), .ZN(n7632) );
  INV_X1 U5862 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7493) );
  INV_X1 U5863 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7402) );
  INV_X1 U5864 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7373) );
  INV_X1 U5865 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7177) );
  INV_X1 U5866 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6837) );
  INV_X1 U5867 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6608) );
  INV_X1 U5868 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6529) );
  INV_X1 U5869 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6527) );
  INV_X1 U5870 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6519) );
  NAND2_X1 U5871 ( .A1(n4428), .A2(n5048), .ZN(n5066) );
  NAND2_X1 U5872 ( .A1(n5046), .A2(n5045), .ZN(n4428) );
  AND2_X1 U5873 ( .A1(n5865), .A2(n5864), .ZN(n9918) );
  NAND2_X1 U5874 ( .A1(n4830), .A2(n5011), .ZN(n5023) );
  NAND2_X1 U5875 ( .A1(n5009), .A2(n5008), .ZN(n4830) );
  NAND2_X1 U5876 ( .A1(n6904), .A2(n6874), .ZN(n7019) );
  AOI21_X1 U5877 ( .B1(n4324), .B2(n5684), .A(n4375), .ZN(n4651) );
  INV_X1 U5878 ( .A(n8588), .ZN(n4566) );
  NAND2_X1 U5879 ( .A1(n8584), .A2(n8828), .ZN(n4569) );
  NAND2_X1 U5880 ( .A1(n4568), .A2(n8583), .ZN(n4567) );
  INV_X1 U5881 ( .A(n4525), .ZN(n4524) );
  OAI21_X1 U5882 ( .B1(n8074), .B2(n8130), .A(n8129), .ZN(n4525) );
  OAI211_X1 U5883 ( .C1(n9185), .C2(n9184), .A(n4445), .B(n4441), .ZN(P1_U3260) );
  INV_X1 U5884 ( .A(n4446), .ZN(n4445) );
  NAND2_X1 U5885 ( .A1(n4442), .A2(n9184), .ZN(n4441) );
  OAI22_X1 U5886 ( .A1(n9206), .A2(n9491), .B1(n9994), .B2(n6487), .ZN(n6488)
         );
  NAND2_X1 U5887 ( .A1(n4810), .A2(n4808), .ZN(P1_U3551) );
  INV_X1 U5888 ( .A(n4809), .ZN(n4808) );
  NAND2_X1 U5889 ( .A1(n4811), .A2(n9994), .ZN(n4810) );
  OAI22_X1 U5890 ( .A1(n4667), .A2(n9491), .B1(n9994), .B2(n9429), .ZN(n4809)
         );
  OAI21_X1 U5891 ( .B1(n6490), .B2(n9988), .A(n4898), .ZN(P1_U3520) );
  OAI21_X1 U5892 ( .B1(n4811), .B2(n9988), .A(n4629), .ZN(n6453) );
  INV_X1 U5893 ( .A(n5811), .ZN(n6072) );
  AND2_X1 U5894 ( .A1(n5622), .A2(n5614), .ZN(n4317) );
  AND2_X1 U5895 ( .A1(n8755), .A2(n8611), .ZN(n4318) );
  AND2_X1 U5896 ( .A1(n4681), .A2(n8641), .ZN(n4319) );
  OR2_X1 U5897 ( .A1(n8876), .A2(n8632), .ZN(n5658) );
  OR3_X1 U5898 ( .A1(n9227), .A2(n6470), .A3(n4663), .ZN(n4320) );
  OAI21_X1 U5899 ( .B1(n6804), .B2(n10005), .A(n4574), .ZN(n7158) );
  AND2_X1 U5900 ( .A1(n4402), .A2(n8062), .ZN(n4321) );
  AND2_X1 U5901 ( .A1(n7797), .A2(n9115), .ZN(n4322) );
  OR2_X1 U5902 ( .A1(n5709), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4323) );
  AND2_X1 U5903 ( .A1(n8062), .A2(n8059), .ZN(n7987) );
  INV_X1 U5904 ( .A(n5753), .ZN(n6349) );
  INV_X1 U5905 ( .A(n8815), .ZN(n4458) );
  INV_X1 U5906 ( .A(n4532), .ZN(n4531) );
  NAND2_X1 U5907 ( .A1(n4534), .A2(n5276), .ZN(n4532) );
  NOR2_X1 U5908 ( .A1(n4777), .A2(n4340), .ZN(n4776) );
  INV_X1 U5909 ( .A(n4776), .ZN(n4516) );
  INV_X1 U5910 ( .A(n9282), .ZN(n9512) );
  NAND2_X1 U5911 ( .A1(n6244), .A2(n6243), .ZN(n9282) );
  INV_X1 U5912 ( .A(n7865), .ZN(n4433) );
  NAND2_X1 U5913 ( .A1(n5783), .A2(n4781), .ZN(n5839) );
  AND2_X1 U5914 ( .A1(n5516), .A2(n5515), .ZN(n4324) );
  AND2_X1 U5915 ( .A1(n7715), .A2(n7714), .ZN(n4325) );
  AND2_X1 U5916 ( .A1(n9248), .A2(n9261), .ZN(n4326) );
  NAND2_X1 U5917 ( .A1(n8596), .A2(n4374), .ZN(n4873) );
  AND2_X1 U5918 ( .A1(n4579), .A2(n4582), .ZN(n4327) );
  AND2_X1 U5919 ( .A1(n4454), .A2(n4456), .ZN(n4328) );
  INV_X1 U5920 ( .A(n4595), .ZN(n4594) );
  OAI21_X1 U5921 ( .B1(n4596), .B2(n4841), .A(n7810), .ZN(n4595) );
  INV_X1 U5922 ( .A(n6455), .ZN(n4667) );
  NAND2_X1 U5923 ( .A1(n4506), .A2(n4504), .ZN(n5928) );
  INV_X1 U5924 ( .A(n7416), .ZN(n4885) );
  NAND2_X1 U5925 ( .A1(n6054), .A2(n6053), .ZN(n7797) );
  INV_X1 U5926 ( .A(n7797), .ZN(n4676) );
  OR2_X1 U5927 ( .A1(n8592), .A2(n7387), .ZN(n4329) );
  NOR2_X1 U5928 ( .A1(n6944), .A2(n5536), .ZN(n4330) );
  INV_X2 U5929 ( .A(n5662), .ZN(n5671) );
  AND2_X1 U5930 ( .A1(n4689), .A2(n8743), .ZN(n4331) );
  NOR2_X1 U5931 ( .A1(n5839), .A2(n4819), .ZN(n5863) );
  NAND2_X1 U5932 ( .A1(n5062), .A2(n5063), .ZN(n5079) );
  INV_X1 U5933 ( .A(n7989), .ZN(n4405) );
  NOR2_X1 U5934 ( .A1(n4842), .A2(n6396), .ZN(n4841) );
  NAND2_X1 U5935 ( .A1(n5457), .A2(n5456), .ZN(n8876) );
  AND2_X1 U5936 ( .A1(n6423), .A2(n4791), .ZN(n4332) );
  INV_X1 U5937 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5509) );
  OR2_X1 U5938 ( .A1(n8603), .A2(n8602), .ZN(n4333) );
  NAND2_X1 U5939 ( .A1(n5314), .A2(n5313), .ZN(n5329) );
  AOI21_X1 U5940 ( .B1(n8132), .B2(n5100), .A(n5475), .ZN(n8625) );
  OAI21_X1 U5941 ( .B1(n5417), .B2(n4837), .A(n4834), .ZN(n5452) );
  NOR2_X1 U5942 ( .A1(n5664), .A2(n5667), .ZN(n8626) );
  NAND2_X1 U5943 ( .A1(n6195), .A2(n6194), .ZN(n9328) );
  NAND2_X1 U5944 ( .A1(n4768), .A2(n6226), .ZN(n9048) );
  OR2_X1 U5945 ( .A1(n8934), .A2(n8839), .ZN(n5539) );
  AND2_X1 U5946 ( .A1(n8026), .A2(n7948), .ZN(n4334) );
  OR2_X1 U5947 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9918), .ZN(n4335) );
  INV_X1 U5948 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U5949 ( .A1(n4867), .A2(n4944), .ZN(n5006) );
  NAND2_X1 U5950 ( .A1(n4506), .A2(n5696), .ZN(n5861) );
  INV_X1 U5951 ( .A(n4720), .ZN(n4719) );
  OAI21_X1 U5952 ( .B1(n8478), .B2(n8316), .A(n8317), .ZN(n4720) );
  NAND2_X1 U5953 ( .A1(n5225), .A2(n5224), .ZN(n8603) );
  NAND2_X1 U5954 ( .A1(n8006), .A2(n9256), .ZN(n9277) );
  INV_X1 U5955 ( .A(n9277), .ZN(n4559) );
  INV_X1 U5956 ( .A(n6470), .ZN(n9206) );
  NAND2_X1 U5957 ( .A1(n6458), .A2(n6457), .ZN(n6470) );
  AND2_X1 U5958 ( .A1(n5658), .A2(n5656), .ZN(n4336) );
  AND3_X1 U5959 ( .A1(n9237), .A2(n8006), .A3(n7929), .ZN(n4337) );
  NAND2_X1 U5960 ( .A1(n9336), .A2(n4669), .ZN(n4673) );
  AND2_X1 U5961 ( .A1(n4559), .A2(n8003), .ZN(n4338) );
  INV_X1 U5962 ( .A(n6839), .ZN(n4839) );
  INV_X1 U5963 ( .A(n4473), .ZN(n4472) );
  AND2_X1 U5964 ( .A1(n9100), .A2(n9114), .ZN(n4339) );
  AND2_X1 U5965 ( .A1(n5574), .A2(n5573), .ZN(n7166) );
  AND2_X1 U5966 ( .A1(n4778), .A2(n6262), .ZN(n4340) );
  OR2_X1 U5967 ( .A1(n6455), .A2(n9222), .ZN(n8062) );
  NOR2_X1 U5968 ( .A1(n8329), .A2(n8328), .ZN(n4341) );
  AND2_X1 U5969 ( .A1(n5600), .A2(n7687), .ZN(n7653) );
  AND2_X1 U5970 ( .A1(n8060), .A2(n8058), .ZN(n9225) );
  AND2_X1 U5971 ( .A1(n5024), .A2(SI_4_), .ZN(n4342) );
  INV_X1 U5972 ( .A(n4462), .ZN(n4461) );
  NAND2_X1 U5973 ( .A1(n8607), .A2(n8604), .ZN(n4462) );
  AND2_X1 U5974 ( .A1(n8620), .A2(n8632), .ZN(n4343) );
  AND2_X1 U5975 ( .A1(n7778), .A2(n5604), .ZN(n4344) );
  AND2_X1 U5976 ( .A1(n4492), .A2(n4497), .ZN(n4345) );
  AND2_X1 U5977 ( .A1(n4772), .A2(n4773), .ZN(n4346) );
  INV_X1 U5978 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U5979 ( .A1(n4734), .A2(n6874), .ZN(n4733) );
  INV_X1 U5980 ( .A(n4670), .ZN(n4669) );
  NAND2_X1 U5981 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  INV_X1 U5982 ( .A(n8607), .ZN(n4460) );
  INV_X1 U5983 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4914) );
  AND2_X1 U5984 ( .A1(n5068), .A2(SI_6_), .ZN(n4347) );
  INV_X1 U5985 ( .A(n8876), .ZN(n8620) );
  INV_X1 U5986 ( .A(n4497), .ZN(n4494) );
  OR2_X1 U5987 ( .A1(n6068), .A2(n7793), .ZN(n4497) );
  INV_X1 U5988 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U5989 ( .A1(n5468), .A2(n4896), .ZN(n4348) );
  NOR2_X1 U5990 ( .A1(n4692), .A2(n4690), .ZN(n4349) );
  AND2_X1 U5991 ( .A1(n5155), .A2(n5138), .ZN(n4350) );
  NAND2_X1 U5992 ( .A1(n5641), .A2(n5647), .ZN(n8686) );
  INV_X1 U5993 ( .A(n8686), .ZN(n4652) );
  AND3_X1 U5994 ( .A1(n5021), .A2(n5020), .A3(n5019), .ZN(n4351) );
  NAND2_X1 U5995 ( .A1(n6009), .A2(n6008), .ZN(n7646) );
  AND2_X1 U5996 ( .A1(n9473), .A2(n9347), .ZN(n4352) );
  NOR2_X1 U5997 ( .A1(n7958), .A2(n4804), .ZN(n4353) );
  OR2_X1 U5998 ( .A1(n7797), .A2(n9093), .ZN(n7869) );
  AND2_X1 U5999 ( .A1(n4458), .A2(n5611), .ZN(n4354) );
  NAND2_X1 U6000 ( .A1(n8862), .A2(n5508), .ZN(n5670) );
  INV_X1 U6001 ( .A(n5670), .ZN(n4870) );
  INV_X1 U6002 ( .A(n4421), .ZN(n4420) );
  OAI21_X1 U6003 ( .B1(n6432), .B2(n7889), .A(n7896), .ZN(n4421) );
  AND2_X1 U6004 ( .A1(n6026), .A2(n6005), .ZN(n4355) );
  AND2_X1 U6005 ( .A1(n4505), .A2(n4503), .ZN(n4356) );
  AND2_X1 U6006 ( .A1(n4321), .A2(n7989), .ZN(n4357) );
  INV_X1 U6007 ( .A(n7024), .ZN(n4731) );
  INV_X1 U6008 ( .A(n7673), .ZN(n4501) );
  XNOR2_X1 U6009 ( .A(n5744), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U6010 ( .A1(n6298), .A2(n6297), .ZN(n6479) );
  INV_X1 U6011 ( .A(n6479), .ZN(n4666) );
  INV_X1 U6012 ( .A(n8919), .ZN(n8770) );
  NAND2_X1 U6013 ( .A1(n5319), .A2(n5318), .ZN(n8919) );
  NAND2_X1 U6014 ( .A1(n6228), .A2(n6227), .ZN(n9453) );
  INV_X1 U6015 ( .A(n9453), .ZN(n4671) );
  AND2_X1 U6016 ( .A1(n9458), .A2(n9322), .ZN(n4358) );
  INV_X1 U6017 ( .A(n9257), .ZN(n4605) );
  INV_X1 U6018 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n4565) );
  XOR2_X1 U6019 ( .A(n6240), .B(n5751), .Z(n4359) );
  INV_X1 U6020 ( .A(n8011), .ZN(n4798) );
  INV_X1 U6021 ( .A(n8033), .ZN(n4786) );
  OR2_X1 U6022 ( .A1(n9206), .A2(n9529), .ZN(n4360) );
  OAI21_X1 U6023 ( .B1(n7675), .B2(n4491), .A(n4487), .ZN(n9088) );
  NAND2_X1 U6024 ( .A1(n8277), .A2(n8465), .ZN(n8364) );
  NAND2_X1 U6025 ( .A1(n4742), .A2(n9089), .ZN(n9008) );
  INV_X1 U6026 ( .A(n9000), .ZN(n4778) );
  NAND2_X1 U6027 ( .A1(n5302), .A2(n5301), .ZN(n8925) );
  NAND2_X1 U6028 ( .A1(n6311), .A2(n6310), .ZN(n6455) );
  NOR2_X1 U6029 ( .A1(n8193), .A2(n6819), .ZN(n4361) );
  INV_X1 U6030 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n4746) );
  OR2_X1 U6031 ( .A1(n8302), .A2(n8425), .ZN(n4362) );
  AND2_X1 U6032 ( .A1(n9017), .A2(n9113), .ZN(n4363) );
  AND2_X1 U6033 ( .A1(n9282), .A2(n9260), .ZN(n4364) );
  INV_X1 U6034 ( .A(n8119), .ZN(n7956) );
  AND2_X1 U6035 ( .A1(n9494), .A2(n9192), .ZN(n8119) );
  AND2_X1 U6036 ( .A1(n5277), .A2(SI_17_), .ZN(n4365) );
  AND2_X1 U6037 ( .A1(n5340), .A2(SI_21_), .ZN(n4366) );
  AND2_X1 U6038 ( .A1(n4464), .A2(n4463), .ZN(n4367) );
  AND2_X1 U6039 ( .A1(n5312), .A2(n5294), .ZN(n4368) );
  AND2_X1 U6040 ( .A1(n5698), .A2(n4505), .ZN(n4369) );
  NAND2_X1 U6041 ( .A1(n5184), .A2(n5183), .ZN(n7681) );
  INV_X1 U6042 ( .A(n7681), .ZN(n4578) );
  NAND2_X1 U6043 ( .A1(n7485), .A2(n7484), .ZN(n7589) );
  NOR2_X1 U6044 ( .A1(n7447), .A2(n4677), .ZN(n4370) );
  NAND2_X1 U6045 ( .A1(n5248), .A2(n5247), .ZN(n8938) );
  INV_X1 U6046 ( .A(n8938), .ZN(n4582) );
  NAND2_X1 U6047 ( .A1(n5877), .A2(n5876), .ZN(n6846) );
  AND2_X1 U6048 ( .A1(n6052), .A2(n6069), .ZN(n7380) );
  NAND2_X1 U6049 ( .A1(n5071), .A2(n5573), .ZN(n7419) );
  AND2_X1 U6050 ( .A1(n5396), .A2(n5382), .ZN(n4371) );
  AND2_X1 U6051 ( .A1(n6046), .A2(n6045), .ZN(n4372) );
  INV_X1 U6052 ( .A(n7484), .ZN(n4725) );
  NAND2_X1 U6053 ( .A1(n5706), .A2(n5707), .ZN(n6346) );
  AND2_X1 U6054 ( .A1(n7589), .A2(n7588), .ZN(n4373) );
  AND2_X1 U6055 ( .A1(n4329), .A2(n8629), .ZN(n4374) );
  NOR2_X1 U6056 ( .A1(n5695), .A2(n5694), .ZN(n4375) );
  AND2_X1 U6057 ( .A1(n5490), .A2(n9635), .ZN(n4376) );
  AND2_X1 U6058 ( .A1(n7225), .A2(n6381), .ZN(n4377) );
  NOR2_X1 U6059 ( .A1(n6361), .A2(n6412), .ZN(n4378) );
  AND2_X1 U6060 ( .A1(n6349), .A2(n9184), .ZN(n7948) );
  NOR2_X1 U6061 ( .A1(n5517), .A2(n4741), .ZN(n4379) );
  INV_X1 U6062 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4807) );
  INV_X1 U6063 ( .A(n9127), .ZN(n4748) );
  OR2_X1 U6064 ( .A1(n9181), .A2(n9180), .ZN(n4380) );
  INV_X1 U6065 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6989) );
  INV_X1 U6066 ( .A(n8257), .ZN(n5536) );
  OAI22_X1 U6067 ( .A1(n8318), .A2(n7158), .B1(n7046), .B2(n8319), .ZN(n6736)
         );
  AOI21_X2 U6068 ( .B1(n7356), .B2(n7357), .A(n7290), .ZN(n7457) );
  AOI21_X2 U6069 ( .B1(n8480), .B2(n8347), .A(n8477), .ZN(n8351) );
  NAND2_X1 U6070 ( .A1(n5062), .A2(n4897), .ZN(n5242) );
  NAND2_X1 U6071 ( .A1(n4392), .A2(n4391), .ZN(n6858) );
  NAND2_X1 U6072 ( .A1(n8357), .A2(n8303), .ZN(n4383) );
  NAND2_X2 U6073 ( .A1(n8392), .A2(n7483), .ZN(n7485) );
  INV_X1 U6074 ( .A(n6737), .ZN(n4392) );
  AND2_X4 U6075 ( .A1(n4384), .A2(n6933), .ZN(n8308) );
  NAND3_X1 U6076 ( .A1(n10016), .A2(n6944), .A3(n7387), .ZN(n4384) );
  OR2_X1 U6077 ( .A1(n7717), .A2(n7716), .ZN(n7766) );
  NAND2_X1 U6078 ( .A1(n8728), .A2(n8727), .ZN(n8707) );
  OAI21_X2 U6079 ( .B1(n7779), .B2(n5235), .A(n5607), .ZN(n8836) );
  NAND2_X1 U6080 ( .A1(n5117), .A2(n5116), .ZN(n7541) );
  OR2_X1 U6081 ( .A1(n5001), .A2(n9996), .ZN(n4963) );
  OAI21_X2 U6082 ( .B1(n7516), .B2(n5596), .A(n7514), .ZN(n7658) );
  NAND3_X1 U6083 ( .A1(n7899), .A2(n8002), .A3(n7998), .ZN(n7901) );
  MUX2_X1 U6084 ( .A(n7903), .B(n7902), .S(n7948), .Z(n7907) );
  MUX2_X1 U6085 ( .A(n7836), .B(n7835), .S(n7929), .Z(n7844) );
  NAND2_X1 U6086 ( .A1(n8025), .A2(n6419), .ZN(n4792) );
  NAND2_X1 U6087 ( .A1(n7822), .A2(n7823), .ZN(n4389) );
  NOR2_X1 U6088 ( .A1(n8304), .A2(n4390), .ZN(n8418) );
  NAND2_X1 U6089 ( .A1(n4697), .A2(n4906), .ZN(n4694) );
  NAND2_X2 U6090 ( .A1(n8403), .A2(n8402), .ZN(n8479) );
  AOI21_X2 U6091 ( .B1(n8479), .B2(n8316), .A(n8478), .ZN(n8345) );
  NAND2_X1 U6092 ( .A1(n10032), .A2(n8505), .ZN(n5541) );
  NAND2_X2 U6093 ( .A1(n8676), .A2(n5651), .ZN(n8659) );
  AOI21_X2 U6094 ( .B1(n5035), .B2(n5556), .A(n4905), .ZN(n7138) );
  NAND2_X1 U6095 ( .A1(n4878), .A2(n4877), .ZN(n8802) );
  NAND2_X1 U6096 ( .A1(n4879), .A2(n4880), .ZN(n7779) );
  NAND2_X1 U6097 ( .A1(n6627), .A2(n5778), .ZN(n5777) );
  NAND2_X1 U6098 ( .A1(n6612), .A2(n5757), .ZN(n6627) );
  OR2_X2 U6099 ( .A1(n9033), .A2(n6262), .ZN(n4779) );
  NOR2_X2 U6100 ( .A1(n5935), .A2(n4393), .ZN(n5772) );
  NAND2_X1 U6101 ( .A1(n7435), .A2(n7434), .ZN(n4749) );
  NAND2_X1 U6102 ( .A1(n6210), .A2(n6209), .ZN(n4771) );
  INV_X1 U6103 ( .A(n4511), .ZN(n6242) );
  INV_X1 U6104 ( .A(n4486), .ZN(n4500) );
  NAND2_X1 U6105 ( .A1(n4345), .A2(n6091), .ZN(n9089) );
  OR2_X1 U6106 ( .A1(n9220), .A2(n4404), .ZN(n4401) );
  OR2_X1 U6107 ( .A1(n9220), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U6108 ( .A1(n9220), .A2(n4357), .ZN(n4397) );
  OR2_X1 U6109 ( .A1(n9220), .A2(n7915), .ZN(n6437) );
  NAND3_X1 U6110 ( .A1(n4398), .A2(n4397), .A3(n4394), .ZN(n6467) );
  NAND2_X1 U6111 ( .A1(n5094), .A2(n4410), .ZN(n4409) );
  INV_X1 U6112 ( .A(n9343), .ZN(n4417) );
  OAI21_X1 U6113 ( .B1(n4417), .B2(n4421), .A(n4418), .ZN(n6433) );
  NAND2_X1 U6114 ( .A1(n5046), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U6115 ( .A1(n4422), .A2(n4425), .ZN(n5082) );
  NAND2_X1 U6116 ( .A1(n9908), .A2(n4449), .ZN(n4448) );
  NAND2_X1 U6117 ( .A1(n4448), .A2(n4447), .ZN(n4450) );
  INV_X1 U6118 ( .A(n4450), .ZN(n9925) );
  AOI21_X1 U6119 ( .B1(n8605), .B2(n4455), .A(n4328), .ZN(n8813) );
  OAI21_X1 U6120 ( .B1(n8720), .B2(n4469), .A(n4467), .ZN(n8684) );
  NOR2_X1 U6121 ( .A1(n8726), .A2(n8713), .ZN(n4473) );
  INV_X1 U6122 ( .A(n6611), .ZN(n5752) );
  NAND2_X1 U6123 ( .A1(n6614), .A2(n6611), .ZN(n6612) );
  INV_X4 U6124 ( .A(n5825), .ZN(n5997) );
  NAND2_X2 U6125 ( .A1(n7071), .A2(n6492), .ZN(n5825) );
  INV_X2 U6126 ( .A(n4750), .ZN(n7071) );
  NAND2_X2 U6127 ( .A1(n6330), .A2(n4480), .ZN(n6492) );
  NAND2_X1 U6128 ( .A1(n5747), .A2(n4484), .ZN(n4482) );
  NAND2_X1 U6129 ( .A1(n5747), .A2(n5749), .ZN(n4483) );
  OAI21_X1 U6130 ( .B1(n7675), .B2(n7673), .A(n4489), .ZN(n4486) );
  CLKBUF_X1 U6131 ( .A(n4500), .Z(n4495) );
  NAND3_X1 U6132 ( .A1(n4506), .A2(n4369), .A3(n4780), .ZN(n5942) );
  AND3_X1 U6133 ( .A1(n4506), .A2(n4502), .A3(n4780), .ZN(n5944) );
  INV_X2 U6134 ( .A(n5839), .ZN(n4506) );
  NAND2_X1 U6135 ( .A1(n7936), .A2(n5860), .ZN(n4510) );
  NAND3_X1 U6136 ( .A1(n5867), .A2(n5866), .A3(n4510), .ZN(n4509) );
  OAI21_X2 U6137 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n4511) );
  AOI21_X2 U6138 ( .B1(n9030), .B2(n9031), .A(n9029), .ZN(n9033) );
  INV_X1 U6139 ( .A(n5022), .ZN(n4519) );
  NAND2_X1 U6140 ( .A1(n4990), .A2(n4989), .ZN(n4520) );
  NAND2_X1 U6141 ( .A1(n4524), .A2(n4521), .ZN(P1_U3240) );
  NAND3_X1 U6142 ( .A1(n7957), .A2(n4523), .A3(n4522), .ZN(n4521) );
  AND2_X1 U6143 ( .A1(n7953), .A2(n9184), .ZN(n4526) );
  NAND2_X1 U6144 ( .A1(n5217), .A2(n4529), .ZN(n4528) );
  OAI21_X1 U6145 ( .B1(n5217), .B2(n4532), .A(n4529), .ZN(n5292) );
  NAND2_X1 U6146 ( .A1(n5314), .A2(n4541), .ZN(n4540) );
  NAND2_X1 U6147 ( .A1(n4540), .A2(n4543), .ZN(n5363) );
  NOR2_X1 U6148 ( .A1(n7946), .A2(n9206), .ZN(n4552) );
  MUX2_X1 U6149 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6808), .S(n8248), .Z(n8239)
         );
  NAND2_X4 U6150 ( .A1(n4866), .A2(n4865), .ZN(n6496) );
  NAND3_X1 U6151 ( .A1(n4569), .A2(n4567), .A3(n4566), .ZN(P2_U3264) );
  NAND3_X1 U6152 ( .A1(n8581), .A2(n8582), .A3(n9998), .ZN(n4568) );
  INV_X1 U6153 ( .A(n4913), .ZN(n4573) );
  NAND2_X1 U6154 ( .A1(n4570), .A2(n5062), .ZN(n5689) );
  AND3_X2 U6155 ( .A1(n5062), .A2(n4573), .A3(n4897), .ZN(n5691) );
  NAND3_X1 U6156 ( .A1(n4575), .A2(n4977), .A3(n10015), .ZN(n10022) );
  NAND2_X4 U6157 ( .A1(n6803), .A2(n8971), .ZN(n6804) );
  INV_X1 U6158 ( .A(n4710), .ZN(n4575) );
  NAND2_X1 U6159 ( .A1(n4327), .A2(n4580), .ZN(n8822) );
  INV_X1 U6160 ( .A(n8823), .ZN(n4586) );
  NAND2_X1 U6161 ( .A1(n4586), .A2(n4587), .ZN(n8750) );
  INV_X1 U6162 ( .A(n7727), .ZN(n4591) );
  OAI21_X1 U6163 ( .B1(n4591), .B2(n4595), .A(n4592), .ZN(n9386) );
  NAND2_X1 U6164 ( .A1(n4602), .A2(n9255), .ZN(n4599) );
  NAND2_X1 U6165 ( .A1(n9374), .A2(n4614), .ZN(n4610) );
  NAND2_X1 U6166 ( .A1(n4610), .A2(n4611), .ZN(n9317) );
  NAND2_X1 U6167 ( .A1(n4620), .A2(n4618), .ZN(n6407) );
  AND3_X1 U6168 ( .A1(n4628), .A2(n5707), .A3(n4859), .ZN(n5713) );
  NAND2_X1 U6169 ( .A1(n9531), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5715) );
  NAND4_X1 U6170 ( .A1(n5707), .A2(n4859), .A3(n4627), .A4(n5706), .ZN(n9531)
         );
  NAND3_X1 U6171 ( .A1(n4838), .A2(n6377), .A3(n6709), .ZN(n6675) );
  AOI21_X1 U6172 ( .B1(n4639), .B2(n4458), .A(n4636), .ZN(n5625) );
  NAND3_X1 U6173 ( .A1(n4641), .A2(n5609), .A3(n8837), .ZN(n4640) );
  NAND2_X1 U6174 ( .A1(n5586), .A2(n4647), .ZN(n5583) );
  NAND3_X1 U6175 ( .A1(n4644), .A2(n4643), .A3(n4642), .ZN(n5586) );
  AOI21_X1 U6176 ( .B1(n5577), .B2(n4649), .A(n4645), .ZN(n4642) );
  OAI21_X1 U6177 ( .B1(n5580), .B2(n7537), .A(n5584), .ZN(n4648) );
  AND2_X1 U6178 ( .A1(n7168), .A2(n5662), .ZN(n4649) );
  NAND2_X1 U6179 ( .A1(n4650), .A2(n4651), .ZN(P2_U3244) );
  NAND3_X1 U6180 ( .A1(n4813), .A2(n4816), .A3(n5684), .ZN(n4650) );
  AND2_X1 U6181 ( .A1(n4653), .A2(n4652), .ZN(n5645) );
  OAI21_X1 U6182 ( .B1(n5634), .B2(n4655), .A(n4654), .ZN(n4653) );
  INV_X1 U6183 ( .A(n7189), .ZN(n7148) );
  NAND2_X1 U6184 ( .A1(n7149), .A2(n7189), .ZN(n7109) );
  AND2_X2 U6185 ( .A1(n4659), .A2(n4351), .ZN(n7149) );
  OR2_X1 U6186 ( .A1(n5480), .A2(n7134), .ZN(n4659) );
  OR2_X1 U6187 ( .A1(n5572), .A2(n5571), .ZN(n5576) );
  OR2_X1 U6188 ( .A1(n5363), .A2(n5362), .ZN(n5365) );
  NAND2_X1 U6189 ( .A1(n5365), .A2(n5364), .ZN(n5381) );
  AOI21_X2 U6190 ( .B1(n5676), .B2(n5675), .A(n5674), .ZN(n5680) );
  NAND2_X1 U6191 ( .A1(n5576), .A2(n5575), .ZN(n5580) );
  MUX2_X1 U6192 ( .A(n5591), .B(n5590), .S(n5671), .Z(n5599) );
  INV_X1 U6193 ( .A(n8256), .ZN(n8505) );
  OAI22_X1 U6194 ( .A1(n5025), .A2(n4976), .B1(n6804), .B2(n8248), .ZN(n4710)
         );
  MUX2_X1 U6195 ( .A(n5556), .B(n5555), .S(n5677), .Z(n5565) );
  NAND4_X1 U6196 ( .A1(n5707), .A2(n5706), .A3(n4806), .A4(n4805), .ZN(n4662)
         );
  INV_X1 U6197 ( .A(n4673), .ZN(n9295) );
  NAND2_X1 U6198 ( .A1(n8653), .A2(n8652), .ZN(n8651) );
  INV_X1 U6199 ( .A(n4683), .ZN(n8720) );
  NAND2_X1 U6200 ( .A1(n8917), .A2(n4903), .ZN(n8749) );
  NAND2_X1 U6201 ( .A1(n8912), .A2(n8765), .ZN(n4691) );
  NOR2_X2 U6202 ( .A1(n4695), .A2(n4694), .ZN(n5028) );
  NAND4_X1 U6203 ( .A1(n4698), .A2(n4945), .A3(n4988), .A4(n4696), .ZN(n4695)
         );
  NAND4_X1 U6204 ( .A1(n4867), .A2(n4697), .A3(n4698), .A4(n4906), .ZN(n5026)
         );
  NAND2_X1 U6205 ( .A1(n4700), .A2(n7151), .ZN(n7119) );
  NAND2_X1 U6206 ( .A1(n7652), .A2(n4704), .ZN(n4701) );
  NAND2_X1 U6207 ( .A1(n4701), .A2(n4702), .ZN(n8605) );
  NAND2_X1 U6208 ( .A1(n7415), .A2(n7414), .ZN(n7417) );
  XNOR2_X2 U6209 ( .A(n4709), .B(n4915), .ZN(n8971) );
  OAI21_X2 U6210 ( .B1(n5689), .B2(P2_IR_REG_26__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4709) );
  OAI21_X1 U6211 ( .B1(n8479), .B2(n4716), .A(n4714), .ZN(n8332) );
  NAND2_X1 U6212 ( .A1(n8479), .A2(n4714), .ZN(n4712) );
  NAND2_X1 U6213 ( .A1(n7485), .A2(n4724), .ZN(n4721) );
  NAND2_X1 U6214 ( .A1(n4721), .A2(n4722), .ZN(n7764) );
  NAND2_X1 U6215 ( .A1(n6904), .A2(n4730), .ZN(n4727) );
  NAND2_X1 U6216 ( .A1(n4727), .A2(n4728), .ZN(n7356) );
  OR2_X1 U6217 ( .A1(n4902), .A2(n4729), .ZN(n4728) );
  INV_X1 U6218 ( .A(n7018), .ZN(n4734) );
  NOR2_X2 U6219 ( .A1(n5279), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5298) );
  OR2_X2 U6220 ( .A1(n7768), .A2(n7769), .ZN(n8267) );
  NAND2_X1 U6221 ( .A1(n8431), .A2(n8289), .ZN(n8290) );
  NOR2_X2 U6222 ( .A1(n5242), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5244) );
  NAND2_X2 U6223 ( .A1(n8342), .A2(n4740), .ZN(n8295) );
  INV_X1 U6224 ( .A(n10016), .ZN(n4741) );
  NAND3_X1 U6225 ( .A1(n4742), .A2(n6108), .A3(n9089), .ZN(n9009) );
  INV_X1 U6226 ( .A(n4744), .ZN(n6666) );
  NAND2_X1 U6227 ( .A1(n6723), .A2(n6724), .ZN(n6722) );
  OAI21_X1 U6228 ( .B1(n4744), .B2(n4743), .A(n6667), .ZN(n6723) );
  NAND2_X1 U6229 ( .A1(n9057), .A2(n5802), .ZN(n4744) );
  AND3_X2 U6230 ( .A1(n4747), .A2(n4746), .A3(n4745), .ZN(n5702) );
  NAND2_X1 U6231 ( .A1(n4749), .A2(n4355), .ZN(n7636) );
  NAND2_X1 U6232 ( .A1(n4751), .A2(n4753), .ZN(n6953) );
  NAND2_X1 U6233 ( .A1(n5877), .A2(n4752), .ZN(n4751) );
  NAND4_X1 U6234 ( .A1(n6156), .A2(n9067), .A3(n9039), .A4(n4762), .ZN(n4757)
         );
  NAND2_X1 U6235 ( .A1(n4757), .A2(n4758), .ZN(n8991) );
  NAND3_X1 U6236 ( .A1(n6156), .A2(n9067), .A3(n4762), .ZN(n4759) );
  CLKBUF_X1 U6237 ( .A(n4771), .Z(n4768) );
  NAND2_X1 U6238 ( .A1(n9033), .A2(n4775), .ZN(n4772) );
  AND2_X2 U6239 ( .A1(n4778), .A2(n4779), .ZN(n9078) );
  OR2_X1 U6240 ( .A1(n9076), .A2(n9077), .ZN(n4777) );
  NOR2_X2 U6241 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5783) );
  NAND2_X1 U6242 ( .A1(n6427), .A2(n4784), .ZN(n4782) );
  NAND2_X1 U6243 ( .A1(n4782), .A2(n4783), .ZN(n7755) );
  OAI21_X1 U6244 ( .B1(n6430), .B2(n4796), .A(n4793), .ZN(n9363) );
  NAND2_X1 U6245 ( .A1(n6433), .A2(n4353), .ZN(n4803) );
  NAND3_X1 U6246 ( .A1(n5706), .A2(n4806), .A3(n5707), .ZN(n5731) );
  INV_X2 U6247 ( .A(n5774), .ZN(n8079) );
  NAND3_X1 U6248 ( .A1(n4815), .A2(n4814), .A3(n4817), .ZN(n4813) );
  NAND2_X1 U6249 ( .A1(n5680), .A2(n8257), .ZN(n4815) );
  OAI21_X1 U6250 ( .B1(n5680), .B2(n5679), .A(n4818), .ZN(n4816) );
  NAND2_X1 U6251 ( .A1(n5417), .A2(n4834), .ZN(n4831) );
  NAND2_X1 U6252 ( .A1(n4831), .A2(n4832), .ZN(n5454) );
  NAND2_X1 U6253 ( .A1(n4843), .A2(n4368), .ZN(n5314) );
  NAND2_X1 U6254 ( .A1(n5470), .A2(n5469), .ZN(n4847) );
  NAND2_X1 U6255 ( .A1(n7028), .A2(n4851), .ZN(n7235) );
  NAND2_X1 U6256 ( .A1(n4852), .A2(n4350), .ZN(n5158) );
  OAI21_X1 U6257 ( .B1(n5237), .B2(n5236), .A(n5238), .ZN(n5258) );
  NAND2_X1 U6258 ( .A1(n5381), .A2(n5380), .ZN(n4863) );
  NAND2_X1 U6259 ( .A1(n4863), .A2(n5382), .ZN(n5395) );
  NAND4_X1 U6260 ( .A1(n5670), .A2(n5532), .A3(n5675), .A4(n8626), .ZN(n4864)
         );
  NAND3_X1 U6261 ( .A1(n4866), .A2(n4865), .A3(n4949), .ZN(n4966) );
  NAND2_X1 U6262 ( .A1(n5256), .A2(n4354), .ZN(n4878) );
  INV_X1 U6263 ( .A(n7658), .ZN(n4882) );
  NAND2_X1 U6264 ( .A1(n7658), .A2(n5213), .ZN(n4879) );
  NAND2_X1 U6265 ( .A1(n7420), .A2(n7542), .ZN(n5117) );
  NAND3_X1 U6266 ( .A1(n4894), .A2(n4893), .A3(n4892), .ZN(n5486) );
  INV_X1 U6267 ( .A(n5664), .ZN(n4892) );
  INV_X1 U6268 ( .A(n10096), .ZN(n10089) );
  NAND2_X1 U6269 ( .A1(n5298), .A2(n4931), .ZN(n5514) );
  AND2_X1 U6270 ( .A1(n8872), .A2(n8871), .ZN(n8873) );
  AOI211_X2 U6271 ( .C1(n8870), .C2(n8856), .A(n8635), .B(n8634), .ZN(n8636)
         );
  NAND2_X1 U6272 ( .A1(n7955), .A2(n7954), .ZN(n7957) );
  NAND2_X1 U6273 ( .A1(n6479), .A2(n6480), .ZN(n6481) );
  NAND2_X1 U6274 ( .A1(n5719), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5759) );
  OR2_X1 U6275 ( .A1(n5001), .A2(n6785), .ZN(n5002) );
  XNOR2_X1 U6276 ( .A(n4952), .B(n4951), .ZN(n4974) );
  NAND2_X1 U6277 ( .A1(n4950), .A2(n4966), .ZN(n4952) );
  INV_X4 U6278 ( .A(n6495), .ZN(n5418) );
  AOI21_X2 U6279 ( .B1(n8740), .B2(n5361), .A(n5632), .ZN(n8728) );
  AND2_X4 U6280 ( .A1(n8136), .A2(n4934), .ZN(n4998) );
  AND2_X1 U6281 ( .A1(n4360), .A2(n6472), .ZN(n4898) );
  INV_X1 U6282 ( .A(n5539), .ZN(n5275) );
  AND2_X1 U6283 ( .A1(n7681), .A2(n8494), .ZN(n4899) );
  AND2_X2 U6284 ( .A1(n6486), .A2(n6915), .ZN(n9989) );
  INV_X2 U6285 ( .A(n9992), .ZN(n9994) );
  INV_X1 U6286 ( .A(n6330), .ZN(n6331) );
  NAND2_X1 U6287 ( .A1(n8338), .A2(n8131), .ZN(n5803) );
  OR2_X1 U6288 ( .A1(n6475), .A2(n6352), .ZN(n4900) );
  INV_X1 U6289 ( .A(n8881), .ZN(n8618) );
  XNOR2_X1 U6290 ( .A(n8628), .B(n8627), .ZN(n4901) );
  NAND2_X1 U6291 ( .A1(n6944), .A2(n6943), .ZN(n8848) );
  INV_X1 U6292 ( .A(n8848), .ZN(n8817) );
  NAND2_X2 U6293 ( .A1(n7057), .A2(n8852), .ZN(n8831) );
  OR2_X1 U6294 ( .A1(n7198), .A2(n7197), .ZN(n10102) );
  INV_X2 U6295 ( .A(n10102), .ZN(n10104) );
  AND2_X1 U6296 ( .A1(n6753), .A2(n6762), .ZN(n8804) );
  OR2_X1 U6297 ( .A1(n8770), .A2(n8610), .ZN(n4903) );
  AND2_X1 U6298 ( .A1(n5450), .A2(n5449), .ZN(n8681) );
  AND2_X1 U6299 ( .A1(n7152), .A2(n8502), .ZN(n4904) );
  NOR2_X1 U6300 ( .A1(n5034), .A2(n5555), .ZN(n4905) );
  INV_X1 U6301 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5055) );
  INV_X1 U6302 ( .A(n7633), .ZN(n5684) );
  INV_X1 U6303 ( .A(n8404), .ZN(n8661) );
  AND2_X1 U6304 ( .A1(n5432), .A2(n5431), .ZN(n8404) );
  INV_X1 U6305 ( .A(n8632), .ZN(n8660) );
  AND2_X1 U6306 ( .A1(n5467), .A2(n5466), .ZN(n8632) );
  INV_X1 U6307 ( .A(n5812), .ZN(n6047) );
  INV_X1 U6308 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5708) );
  INV_X1 U6309 ( .A(n5935), .ZN(n5740) );
  INV_X1 U6310 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9582) );
  INV_X1 U6311 ( .A(n8756), .ZN(n5337) );
  INV_X1 U6312 ( .A(n7060), .ZN(n4980) );
  INV_X1 U6313 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5710) );
  OR4_X1 U6314 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6341) );
  INV_X1 U6315 ( .A(n5168), .ZN(n5167) );
  INV_X1 U6316 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5145) );
  INV_X1 U6317 ( .A(n5229), .ZN(n5227) );
  INV_X1 U6318 ( .A(n5109), .ZN(n5107) );
  INV_X1 U6319 ( .A(n7653), .ZN(n7657) );
  NAND2_X1 U6320 ( .A1(n6804), .A2(n5418), .ZN(n5025) );
  INV_X1 U6321 ( .A(n5629), .ZN(n5326) );
  NAND2_X1 U6322 ( .A1(n4980), .A2(n4979), .ZN(n7099) );
  INV_X1 U6323 ( .A(n7640), .ZN(n6026) );
  INV_X1 U6324 ( .A(n6230), .ZN(n6229) );
  OR2_X1 U6325 ( .A1(n6196), .A2(n8994), .ZN(n6214) );
  NOR2_X1 U6326 ( .A1(n6048), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n6093) );
  INV_X1 U6327 ( .A(SI_10_), .ZN(n9670) );
  INV_X1 U6328 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U6329 ( .A1(n5385), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U6330 ( .A1(n5352), .A2(n5351), .ZN(n5372) );
  NAND2_X1 U6331 ( .A1(n5227), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6332 ( .A1(n5107), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5128) );
  OAI222_X1 U6333 ( .A1(n4901), .A2(n8817), .B1(n8632), .B2(n8840), .C1(n5533), 
        .C2(n8631), .ZN(n8633) );
  NOR2_X1 U6334 ( .A1(n10096), .A2(n8828), .ZN(n7180) );
  OR2_X1 U6335 ( .A1(n5181), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n5182) );
  INV_X1 U6336 ( .A(n5938), .ZN(n5939) );
  NAND2_X1 U6337 ( .A1(n6229), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U6338 ( .A1(n6213), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U6339 ( .A1(n6160), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U6340 ( .A1(n6139), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U6341 ( .A1(n6097), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U6342 ( .A1(n6055), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6077) );
  OR2_X1 U6343 ( .A1(n5968), .A2(n6592), .ZN(n5991) );
  NAND2_X1 U6344 ( .A1(n5921), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6345 ( .A1(n5732), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  OR2_X1 U6346 ( .A1(n5498), .A2(n5497), .ZN(n5499) );
  INV_X1 U6347 ( .A(SI_17_), .ZN(n5260) );
  OR2_X1 U6348 ( .A1(n6093), .A2(n5899), .ZN(n6051) );
  AND2_X1 U6349 ( .A1(n7801), .A2(n7746), .ZN(n5693) );
  NAND2_X1 U6350 ( .A1(n5127), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6351 ( .A1(n5443), .A2(n9734), .ZN(n5460) );
  OR2_X1 U6352 ( .A1(n5320), .A2(n9694), .ZN(n5350) );
  OR2_X1 U6353 ( .A1(n5407), .A2(n9712), .ZN(n5426) );
  OR2_X1 U6354 ( .A1(n8477), .A2(n8319), .ZN(n8475) );
  OR2_X1 U6355 ( .A1(n8672), .A2(n4313), .ZN(n5432) );
  INV_X1 U6356 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9719) );
  INV_X1 U6357 ( .A(n8925), .ZN(n8784) );
  AND2_X1 U6358 ( .A1(n5570), .A2(n5568), .ZN(n7154) );
  INV_X1 U6359 ( .A(n8804), .ZN(n8840) );
  AOI21_X1 U6360 ( .B1(n6750), .B2(n10009), .A(n10010), .ZN(n7196) );
  AND2_X1 U6361 ( .A1(n6296), .A2(n6295), .ZN(n6474) );
  NAND2_X1 U6362 ( .A1(n9021), .A2(n9022), .ZN(n9020) );
  INV_X1 U6363 ( .A(n9082), .ZN(n9096) );
  INV_X1 U6364 ( .A(n5804), .ZN(n6299) );
  INV_X1 U6365 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6592) );
  INV_X1 U6366 ( .A(n9110), .ZN(n9307) );
  INV_X1 U6367 ( .A(n6432), .ZN(n9318) );
  INV_X1 U6368 ( .A(n9321), .ZN(n9365) );
  OR2_X1 U6369 ( .A1(n6493), .A2(n8121), .ZN(n6913) );
  NOR2_X1 U6370 ( .A1(n9965), .A2(n6345), .ZN(n6484) );
  NAND2_X1 U6371 ( .A1(n9988), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6472) );
  INV_X1 U6372 ( .A(n9346), .ZN(n9403) );
  OR2_X1 U6373 ( .A1(n6917), .A2(n8121), .ZN(n9982) );
  AND2_X1 U6374 ( .A1(n5382), .A2(n5369), .ZN(n5380) );
  XNOR2_X1 U6375 ( .A(n5156), .B(n5139), .ZN(n5155) );
  NOR2_X1 U6376 ( .A1(n10167), .A2(n10166), .ZN(n9549) );
  NAND2_X1 U6377 ( .A1(n4935), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4938) );
  AND2_X1 U6378 ( .A1(n6761), .A2(n6760), .ZN(n8335) );
  INV_X1 U6379 ( .A(n8483), .ZN(n8472) );
  AND3_X1 U6380 ( .A1(n4929), .A2(n4928), .A3(n4927), .ZN(n5508) );
  AND3_X1 U6381 ( .A1(n5324), .A2(n5323), .A3(n5322), .ZN(n8610) );
  INV_X1 U6382 ( .A(n9995), .ZN(n10000) );
  AND2_X1 U6383 ( .A1(n6806), .A2(n6805), .ZN(n9995) );
  INV_X1 U6384 ( .A(n8613), .ZN(n8708) );
  INV_X1 U6385 ( .A(n8838), .ZN(n8806) );
  AND2_X1 U6386 ( .A1(n7655), .A2(n7654), .ZN(n9809) );
  AND2_X1 U6387 ( .A1(n7196), .A2(n7194), .ZN(n7184) );
  AND2_X1 U6388 ( .A1(n8845), .A2(n9806), .ZN(n10085) );
  OR2_X1 U6389 ( .A1(n4367), .A2(n8844), .ZN(n8942) );
  AND2_X1 U6390 ( .A1(n7538), .A2(n7418), .ZN(n10069) );
  INV_X1 U6391 ( .A(n10085), .ZN(n10101) );
  OR2_X1 U6392 ( .A1(n7183), .A2(n7182), .ZN(n7198) );
  XNOR2_X1 U6393 ( .A(n5692), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7746) );
  AND2_X1 U6394 ( .A1(n5104), .A2(n5140), .ZN(n6823) );
  INV_X1 U6395 ( .A(n9087), .ZN(n6480) );
  INV_X1 U6396 ( .A(n9094), .ZN(n9062) );
  INV_X1 U6397 ( .A(n9070), .ZN(n9099) );
  AND3_X1 U6398 ( .A1(n6201), .A2(n6200), .A3(n6199), .ZN(n9306) );
  NAND4_X1 U6399 ( .A1(n5791), .A2(n5790), .A3(n5789), .A4(n5788), .ZN(n5795)
         );
  INV_X1 U6400 ( .A(n9964), .ZN(n9866) );
  INV_X1 U6401 ( .A(n9951), .ZN(n9943) );
  AND2_X1 U6402 ( .A1(n9179), .A2(n6542), .ZN(n9951) );
  INV_X1 U6403 ( .A(n9390), .ZN(n9228) );
  AND2_X1 U6404 ( .A1(n7895), .A2(n7889), .ZN(n9345) );
  AND2_X1 U6405 ( .A1(n9409), .A2(n8070), .ZN(n9397) );
  AND2_X1 U6406 ( .A1(n7953), .A2(n9861), .ZN(n9346) );
  INV_X1 U6407 ( .A(n9400), .ZN(n9351) );
  OR2_X1 U6408 ( .A1(n9973), .A2(n9824), .ZN(n9986) );
  AND2_X1 U6409 ( .A1(n7948), .A2(n8122), .ZN(n9973) );
  INV_X1 U6410 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5729) );
  AND2_X1 U6411 ( .A1(n6117), .A2(n6135), .ZN(n9175) );
  NOR2_X1 U6412 ( .A1(n9550), .A2(n9549), .ZN(n10162) );
  INV_X1 U6413 ( .A(n8587), .ZN(n10002) );
  INV_X1 U6414 ( .A(n8461), .ZN(n8485) );
  NAND2_X1 U6415 ( .A1(n6881), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8483) );
  INV_X1 U6416 ( .A(n8714), .ZN(n8614) );
  NAND2_X1 U6417 ( .A1(n6803), .A2(n6802), .ZN(n9998) );
  INV_X1 U6418 ( .A(n9997), .ZN(n8578) );
  NAND2_X1 U6419 ( .A1(n8831), .A2(n6932), .ZN(n8859) );
  AND2_X1 U6420 ( .A1(n8859), .A2(n6935), .ZN(n8812) );
  INV_X1 U6421 ( .A(n10120), .ZN(n10118) );
  AND3_X1 U6422 ( .A1(n10093), .A2(n10092), .A3(n10091), .ZN(n10117) );
  NAND2_X1 U6423 ( .A1(n10008), .A2(n10007), .ZN(n10011) );
  INV_X1 U6424 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7701) );
  INV_X1 U6425 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6836) );
  INV_X1 U6426 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6561) );
  INV_X1 U6427 ( .A(n7631), .ZN(n8970) );
  AND2_X1 U6428 ( .A1(n6355), .A2(n9820), .ZN(n9087) );
  INV_X1 U6429 ( .A(n9080), .ZN(n9103) );
  NAND2_X1 U6430 ( .A1(n6288), .A2(n6287), .ZN(n9261) );
  INV_X1 U6431 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9916) );
  INV_X1 U6432 ( .A(n9960), .ZN(n9935) );
  OR2_X1 U6433 ( .A1(P1_U3083), .A2(n9890), .ZN(n9964) );
  NAND2_X1 U6434 ( .A1(n9409), .A2(n7031), .ZN(n9408) );
  AND2_X2 U6435 ( .A1(n7038), .A2(n9820), .ZN(n9826) );
  NAND2_X1 U6436 ( .A1(n9994), .A2(n9843), .ZN(n9491) );
  NAND2_X1 U6437 ( .A1(n6486), .A2(n6485), .ZN(n9992) );
  INV_X1 U6438 ( .A(n9830), .ZN(n7762) );
  NAND2_X1 U6439 ( .A1(n9989), .A2(n9843), .ZN(n9529) );
  INV_X1 U6440 ( .A(n9989), .ZN(n9988) );
  NAND2_X1 U6441 ( .A1(n9966), .A2(n9965), .ZN(n9967) );
  AND2_X1 U6442 ( .A1(n6492), .A2(n6348), .ZN(n9966) );
  INV_X1 U6443 ( .A(n6350), .ZN(n8066) );
  INV_X1 U6444 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6689) );
  INV_X1 U6445 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6563) );
  AND2_X2 U6446 ( .A1(n6796), .A2(n10013), .ZN(P2_U3966) );
  INV_X2 U6447 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4906) );
  NOR2_X1 U6448 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n4911) );
  NOR2_X1 U6449 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4910) );
  NOR2_X1 U6450 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4909) );
  NAND4_X1 U6451 ( .A1(n4912), .A2(n4911), .A3(n4910), .A4(n4909), .ZN(n4913)
         );
  INV_X1 U6452 ( .A(n4920), .ZN(n8960) );
  INV_X1 U6453 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4919) );
  XNOR2_X2 U6454 ( .A(n4921), .B(P2_IR_REG_30__SCAN_IN), .ZN(n4933) );
  INV_X1 U6455 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n8597) );
  INV_X2 U6456 ( .A(n4933), .ZN(n8136) );
  NAND2_X1 U6457 ( .A1(n4998), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n4925) );
  NAND2_X1 U6458 ( .A1(n5074), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n4924) );
  OAI211_X1 U6459 ( .C1(n5480), .C2(n8597), .A(n4925), .B(n4924), .ZN(n8629)
         );
  INV_X1 U6460 ( .A(n8629), .ZN(n5533) );
  NAND2_X1 U6461 ( .A1(n4998), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n4929) );
  INV_X1 U6462 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8589) );
  OR2_X1 U6463 ( .A1(n5480), .A2(n8589), .ZN(n4928) );
  INV_X1 U6464 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n4926) );
  OR2_X1 U6465 ( .A1(n5000), .A2(n4926), .ZN(n4927) );
  INV_X1 U6466 ( .A(n5508), .ZN(n8592) );
  NOR2_X1 U6467 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n4931) );
  NAND2_X1 U6468 ( .A1(n5514), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4932) );
  INV_X2 U6469 ( .A(n6731), .ZN(n7387) );
  NAND2_X1 U6470 ( .A1(n4998), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4940) );
  INV_X1 U6471 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9625) );
  INV_X1 U6472 ( .A(n5001), .ZN(n4935) );
  INV_X1 U6473 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4936) );
  OR2_X1 U6474 ( .A1(n4944), .A2(n4919), .ZN(n4946) );
  XNOR2_X1 U6475 ( .A(n4946), .B(n4945), .ZN(n6810) );
  INV_X1 U6476 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6502) );
  OR2_X1 U6477 ( .A1(n5025), .A2(n6502), .ZN(n4957) );
  NAND3_X1 U6478 ( .A1(n6496), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4950) );
  AND2_X1 U6479 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4949) );
  INV_X1 U6480 ( .A(SI_1_), .ZN(n4951) );
  MUX2_X1 U6481 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n6496), .Z(n4973) );
  NAND2_X1 U6482 ( .A1(n4974), .A2(n4973), .ZN(n4954) );
  NAND2_X1 U6483 ( .A1(n4952), .A2(SI_1_), .ZN(n4953) );
  NAND2_X1 U6484 ( .A1(n4954), .A2(n4953), .ZN(n4990) );
  MUX2_X1 U6485 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n6496), .Z(n4991) );
  INV_X1 U6486 ( .A(SI_2_), .ZN(n4955) );
  XNOR2_X1 U6487 ( .A(n4991), .B(n4955), .ZN(n4989) );
  XNOR2_X1 U6488 ( .A(n4990), .B(n4989), .ZN(n6514) );
  OAI211_X1 U6489 ( .C1(n6804), .C2(n6810), .A(n4957), .B(n4956), .ZN(n6859)
         );
  INV_X1 U6490 ( .A(n6859), .ZN(n10032) );
  NAND2_X2 U6491 ( .A1(n5541), .A2(n7098), .ZN(n7060) );
  INV_X1 U6492 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U6493 ( .A1(n4998), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4962) );
  INV_X1 U6494 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n4958) );
  INV_X1 U6495 ( .A(n4313), .ZN(n4959) );
  NAND2_X1 U6496 ( .A1(n4315), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n4960) );
  NAND4_X2 U6497 ( .A1(n4963), .A2(n4962), .A3(n4961), .A4(n4960), .ZN(n6763)
         );
  INV_X1 U6498 ( .A(n6763), .ZN(n4967) );
  INV_X1 U6499 ( .A(SI_0_), .ZN(n9659) );
  INV_X1 U6500 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4964) );
  OAI21_X1 U6501 ( .B1(n5418), .B2(n9659), .A(n4964), .ZN(n4965) );
  AND2_X1 U6502 ( .A1(n4966), .A2(n4965), .ZN(n8975) );
  NAND2_X2 U6503 ( .A1(n4967), .A2(n7158), .ZN(n5519) );
  INV_X1 U6504 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n4968) );
  OR2_X1 U6505 ( .A1(n5000), .A2(n4968), .ZN(n4972) );
  NAND2_X1 U6506 ( .A1(n4315), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n4971) );
  NAND2_X1 U6507 ( .A1(n4935), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4970) );
  NAND2_X1 U6508 ( .A1(n4998), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4969) );
  XNOR2_X1 U6509 ( .A(n4974), .B(n4973), .ZN(n6512) );
  OR2_X1 U6510 ( .A1(n5090), .A2(n6512), .ZN(n4977) );
  INV_X1 U6511 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n4976) );
  INV_X1 U6512 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6513 ( .A1(n5519), .A2(n5543), .ZN(n4978) );
  INV_X1 U6514 ( .A(n7054), .ZN(n10024) );
  NAND2_X1 U6515 ( .A1(n6730), .A2(n10024), .ZN(n5542) );
  NAND2_X1 U6516 ( .A1(n4978), .A2(n5542), .ZN(n7061) );
  INV_X1 U6517 ( .A(n7061), .ZN(n4979) );
  NAND2_X1 U6518 ( .A1(n7099), .A2(n7098), .ZN(n4997) );
  NAND2_X1 U6519 ( .A1(n4998), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4985) );
  OR2_X1 U6520 ( .A1(n4313), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4984) );
  INV_X1 U6521 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6786) );
  OR2_X1 U6522 ( .A1(n5001), .A2(n6786), .ZN(n4983) );
  INV_X1 U6523 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n4981) );
  OR2_X1 U6524 ( .A1(n5000), .A2(n4981), .ZN(n4982) );
  OR3_X1 U6525 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4986) );
  NAND2_X1 U6526 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4986), .ZN(n4987) );
  XNOR2_X1 U6527 ( .A(n4988), .B(n4987), .ZN(n8237) );
  INV_X1 U6528 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6500) );
  OR2_X1 U6529 ( .A1(n5025), .A2(n6500), .ZN(n4995) );
  NAND2_X1 U6530 ( .A1(n4991), .A2(SI_2_), .ZN(n4992) );
  MUX2_X1 U6531 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n6496), .Z(n5010) );
  INV_X1 U6532 ( .A(SI_3_), .ZN(n4993) );
  XNOR2_X1 U6533 ( .A(n5009), .B(n5008), .ZN(n6516) );
  OR2_X1 U6534 ( .A1(n5090), .A2(n6516), .ZN(n4994) );
  OAI211_X1 U6535 ( .C1(n6804), .C2(n8237), .A(n4995), .B(n4994), .ZN(n4996)
         );
  NAND2_X1 U6536 ( .A1(n7063), .A2(n4996), .ZN(n5520) );
  INV_X1 U6537 ( .A(n7063), .ZN(n8504) );
  NAND2_X1 U6538 ( .A1(n8504), .A2(n10037), .ZN(n5522) );
  INV_X1 U6539 ( .A(n7110), .ZN(n5557) );
  NAND2_X1 U6540 ( .A1(n4997), .A2(n5557), .ZN(n7101) );
  INV_X1 U6541 ( .A(n7127), .ZN(n5035) );
  NAND2_X1 U6542 ( .A1(n4998), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5005) );
  INV_X1 U6543 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n4999) );
  OR2_X1 U6544 ( .A1(n5000), .A2(n4999), .ZN(n5004) );
  NAND2_X1 U6545 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5017) );
  OAI21_X1 U6546 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5017), .ZN(n6910) );
  OR2_X1 U6547 ( .A1(n4312), .A2(n6910), .ZN(n5003) );
  INV_X1 U6548 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6785) );
  NAND2_X1 U6549 ( .A1(n5006), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5007) );
  XNOR2_X1 U6550 ( .A(n5007), .B(n4906), .ZN(n8226) );
  OR2_X1 U6551 ( .A1(n5025), .A2(n4565), .ZN(n5014) );
  NAND2_X1 U6552 ( .A1(n5010), .A2(SI_3_), .ZN(n5011) );
  INV_X1 U6553 ( .A(SI_4_), .ZN(n5012) );
  XNOR2_X1 U6554 ( .A(n5024), .B(n5012), .ZN(n5022) );
  XNOR2_X1 U6555 ( .A(n5023), .B(n5022), .ZN(n6501) );
  OR2_X1 U6556 ( .A1(n5090), .A2(n6501), .ZN(n5013) );
  OAI211_X1 U6557 ( .C1(n6804), .C2(n8226), .A(n5014), .B(n5013), .ZN(n5033)
         );
  NAND2_X1 U6558 ( .A1(n7118), .A2(n5033), .ZN(n7125) );
  INV_X1 U6559 ( .A(n5017), .ZN(n5015) );
  NAND2_X1 U6560 ( .A1(n5015), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5038) );
  INV_X1 U6561 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5016) );
  NAND2_X1 U6562 ( .A1(n5017), .A2(n5016), .ZN(n5018) );
  NAND2_X1 U6563 ( .A1(n5038), .A2(n5018), .ZN(n7123) );
  OR2_X1 U6564 ( .A1(n4312), .A2(n7123), .ZN(n5021) );
  INV_X1 U6565 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7134) );
  NAND2_X1 U6566 ( .A1(n4998), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6567 ( .A1(n5074), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5019) );
  MUX2_X1 U6568 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6496), .Z(n5047) );
  XNOR2_X1 U6569 ( .A(n5047), .B(n9636), .ZN(n5045) );
  XNOR2_X1 U6570 ( .A(n5046), .B(n5045), .ZN(n6505) );
  OR2_X1 U6571 ( .A1(n5090), .A2(n6505), .ZN(n5032) );
  INV_X1 U6572 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U6573 ( .A1(n5026), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5027) );
  MUX2_X1 U6574 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5027), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5030) );
  INV_X1 U6575 ( .A(n5028), .ZN(n5029) );
  INV_X1 U6576 ( .A(n6816), .ZN(n8215) );
  OR2_X1 U6577 ( .A1(n6804), .A2(n8215), .ZN(n5031) );
  INV_X1 U6578 ( .A(n7109), .ZN(n5034) );
  NAND2_X1 U6579 ( .A1(n8503), .A2(n10044), .ZN(n7128) );
  AND2_X2 U6580 ( .A1(n7128), .A2(n7152), .ZN(n5555) );
  NAND2_X1 U6581 ( .A1(n4998), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5043) );
  INV_X1 U6582 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5036) );
  OR2_X1 U6583 ( .A1(n5000), .A2(n5036), .ZN(n5042) );
  INV_X1 U6584 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6783) );
  OR2_X1 U6585 ( .A1(n5480), .A2(n6783), .ZN(n5041) );
  INV_X1 U6586 ( .A(n5038), .ZN(n5037) );
  NAND2_X1 U6587 ( .A1(n5037), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5056) );
  INV_X1 U6588 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9740) );
  NAND2_X1 U6589 ( .A1(n5038), .A2(n9740), .ZN(n5039) );
  NAND2_X1 U6590 ( .A1(n5056), .A2(n5039), .ZN(n7145) );
  OR2_X1 U6591 ( .A1(n4313), .A2(n7145), .ZN(n5040) );
  OR2_X1 U6592 ( .A1(n5028), .A2(n4919), .ZN(n5044) );
  XNOR2_X1 U6593 ( .A(n5044), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6818) );
  INV_X1 U6594 ( .A(n6818), .ZN(n8204) );
  NAND2_X1 U6595 ( .A1(n5047), .A2(SI_5_), .ZN(n5048) );
  INV_X1 U6596 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n5049) );
  MUX2_X1 U6597 ( .A(n6504), .B(n5049), .S(n6496), .Z(n5067) );
  XNOR2_X1 U6598 ( .A(n5067), .B(SI_6_), .ZN(n5065) );
  XNOR2_X1 U6599 ( .A(n5066), .B(n5065), .ZN(n6503) );
  OR2_X1 U6600 ( .A1(n5090), .A2(n6503), .ZN(n5051) );
  OR2_X1 U6601 ( .A1(n5505), .A2(n6504), .ZN(n5050) );
  OAI211_X1 U6602 ( .C1(n6804), .C2(n8204), .A(n5051), .B(n5050), .ZN(n10049)
         );
  NAND2_X1 U6603 ( .A1(n7167), .A2(n10049), .ZN(n5570) );
  INV_X1 U6604 ( .A(n10049), .ZN(n5052) );
  NAND2_X1 U6605 ( .A1(n8501), .A2(n5052), .ZN(n5568) );
  INV_X1 U6606 ( .A(n5570), .ZN(n5053) );
  NAND2_X1 U6607 ( .A1(n4998), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5061) );
  INV_X1 U6608 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5054) );
  OR2_X1 U6609 ( .A1(n5000), .A2(n5054), .ZN(n5060) );
  NAND2_X1 U6610 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  NAND2_X1 U6611 ( .A1(n5072), .A2(n5057), .ZN(n7260) );
  OR2_X1 U6612 ( .A1(n4312), .A2(n7260), .ZN(n5059) );
  INV_X1 U6613 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7170) );
  OR2_X1 U6614 ( .A1(n5480), .A2(n7170), .ZN(n5058) );
  OR2_X1 U6615 ( .A1(n5062), .A2(n4919), .ZN(n5064) );
  XNOR2_X1 U6616 ( .A(n5064), .B(n5063), .ZN(n8193) );
  INV_X1 U6617 ( .A(n5067), .ZN(n5068) );
  MUX2_X1 U6618 ( .A(n6517), .B(n6519), .S(n5418), .Z(n5083) );
  XNOR2_X1 U6619 ( .A(n5083), .B(SI_7_), .ZN(n5081) );
  XNOR2_X1 U6620 ( .A(n5082), .B(n5081), .ZN(n6518) );
  OR2_X1 U6621 ( .A1(n5090), .A2(n6518), .ZN(n5070) );
  OR2_X1 U6622 ( .A1(n5505), .A2(n6517), .ZN(n5069) );
  OAI211_X1 U6623 ( .C1(n6804), .C2(n8193), .A(n5070), .B(n5069), .ZN(n7252)
         );
  NAND2_X1 U6624 ( .A1(n7413), .A2(n7252), .ZN(n5574) );
  NAND2_X1 U6625 ( .A1(n8500), .A2(n10059), .ZN(n5573) );
  NAND2_X1 U6626 ( .A1(n5072), .A2(n9719), .ZN(n5073) );
  NAND2_X1 U6627 ( .A1(n5109), .A2(n5073), .ZN(n7427) );
  OR2_X1 U6628 ( .A1(n4312), .A2(n7427), .ZN(n5078) );
  NAND2_X1 U6629 ( .A1(n4998), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6630 ( .A1(n5074), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5076) );
  INV_X1 U6631 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6782) );
  OR2_X1 U6632 ( .A1(n5480), .A2(n6782), .ZN(n5075) );
  NAND4_X1 U6633 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n8499)
         );
  NAND2_X1 U6634 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6635 ( .A(n5080), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U6636 ( .A1(n5300), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5299), .B2(
        n6821), .ZN(n5092) );
  NAND2_X1 U6637 ( .A1(n5082), .A2(n5081), .ZN(n5086) );
  INV_X1 U6638 ( .A(n5083), .ZN(n5084) );
  NAND2_X1 U6639 ( .A1(n5084), .A2(SI_7_), .ZN(n5085) );
  MUX2_X1 U6640 ( .A(n6525), .B(n6527), .S(n5418), .Z(n5087) );
  INV_X1 U6641 ( .A(n5087), .ZN(n5088) );
  NAND2_X1 U6642 ( .A1(n5088), .A2(SI_8_), .ZN(n5089) );
  NAND2_X1 U6643 ( .A1(n5095), .A2(n5089), .ZN(n5093) );
  XNOR2_X1 U6644 ( .A(n5094), .B(n5093), .ZN(n6524) );
  NAND2_X1 U6645 ( .A1(n6524), .A2(n5100), .ZN(n5091) );
  NAND2_X1 U6646 ( .A1(n8499), .A2(n10064), .ZN(n7537) );
  OAI21_X1 U6647 ( .B1(n8499), .B2(n10064), .A(n7537), .ZN(n7416) );
  INV_X1 U6648 ( .A(n8499), .ZN(n7168) );
  NAND2_X1 U6649 ( .A1(n7168), .A2(n10064), .ZN(n7542) );
  MUX2_X1 U6650 ( .A(n6531), .B(n6529), .S(n6496), .Z(n5097) );
  NAND2_X1 U6651 ( .A1(n5097), .A2(n5096), .ZN(n5120) );
  INV_X1 U6652 ( .A(n5097), .ZN(n5098) );
  NAND2_X1 U6653 ( .A1(n5098), .A2(SI_9_), .ZN(n5099) );
  XNOR2_X1 U6654 ( .A(n5119), .B(n5118), .ZN(n6528) );
  NAND2_X1 U6655 ( .A1(n6528), .A2(n5100), .ZN(n5106) );
  NAND2_X1 U6656 ( .A1(n5103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  MUX2_X1 U6657 ( .A(n5102), .B(P2_IR_REG_31__SCAN_IN), .S(n5101), .Z(n5104)
         );
  AOI22_X1 U6658 ( .A1(n5300), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5299), .B2(
        n6823), .ZN(n5105) );
  INV_X1 U6659 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5108) );
  NAND2_X1 U6660 ( .A1(n5109), .A2(n5108), .ZN(n5110) );
  NAND2_X1 U6661 ( .A1(n5128), .A2(n5110), .ZN(n7550) );
  OR2_X1 U6662 ( .A1(n4313), .A2(n7550), .ZN(n5115) );
  NAND2_X1 U6663 ( .A1(n4998), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6664 ( .A1(n5074), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5113) );
  INV_X1 U6665 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5111) );
  OR2_X1 U6666 ( .A1(n5480), .A2(n5111), .ZN(n5112) );
  NAND4_X1 U6667 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n8498)
         );
  NAND2_X1 U6668 ( .A1(n10072), .A2(n8498), .ZN(n5581) );
  INV_X1 U6669 ( .A(n8498), .ZN(n7562) );
  NAND2_X1 U6670 ( .A1(n7554), .A2(n7562), .ZN(n5584) );
  NAND2_X1 U6671 ( .A1(n5581), .A2(n5584), .ZN(n7543) );
  INV_X1 U6672 ( .A(n7543), .ZN(n5116) );
  MUX2_X1 U6673 ( .A(n6561), .B(n6563), .S(n5418), .Z(n5121) );
  INV_X1 U6674 ( .A(n5121), .ZN(n5122) );
  NAND2_X1 U6675 ( .A1(n5122), .A2(SI_10_), .ZN(n5123) );
  NAND2_X1 U6676 ( .A1(n5140), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5124) );
  XNOR2_X1 U6677 ( .A(n5124), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U6678 ( .A1(n5300), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5299), .B2(
        n6825), .ZN(n5125) );
  NAND2_X1 U6679 ( .A1(n4998), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5134) );
  INV_X1 U6680 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5126) );
  OR2_X1 U6681 ( .A1(n5000), .A2(n5126), .ZN(n5133) );
  INV_X1 U6682 ( .A(n5128), .ZN(n5127) );
  INV_X1 U6683 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9725) );
  NAND2_X1 U6684 ( .A1(n5128), .A2(n9725), .ZN(n5129) );
  NAND2_X1 U6685 ( .A1(n5146), .A2(n5129), .ZN(n7581) );
  OR2_X1 U6686 ( .A1(n4313), .A2(n7581), .ZN(n5132) );
  INV_X1 U6687 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5130) );
  OR2_X1 U6688 ( .A1(n5480), .A2(n5130), .ZN(n5131) );
  OR2_X1 U6689 ( .A1(n7578), .A2(n8451), .ZN(n5587) );
  NAND2_X1 U6690 ( .A1(n7561), .A2(n5587), .ZN(n5135) );
  NAND2_X1 U6691 ( .A1(n7578), .A2(n8451), .ZN(n5585) );
  NAND2_X1 U6692 ( .A1(n5135), .A2(n5585), .ZN(n7599) );
  MUX2_X1 U6693 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5418), .Z(n5156) );
  XNOR2_X1 U6694 ( .A(n5154), .B(n5155), .ZN(n6580) );
  NAND2_X1 U6695 ( .A1(n6580), .A2(n5100), .ZN(n5143) );
  OR2_X1 U6696 ( .A1(n5163), .A2(n4919), .ZN(n5141) );
  XNOR2_X1 U6697 ( .A(n5141), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U6698 ( .A1(n5300), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5299), .B2(
        n6983), .ZN(n5142) );
  NAND2_X1 U6699 ( .A1(n5143), .A2(n5142), .ZN(n10087) );
  NAND2_X1 U6700 ( .A1(n4998), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5152) );
  INV_X1 U6701 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6702 ( .A1(n5000), .A2(n5144), .ZN(n5151) );
  NAND2_X1 U6703 ( .A1(n5146), .A2(n5145), .ZN(n5147) );
  NAND2_X1 U6704 ( .A1(n5168), .A2(n5147), .ZN(n8456) );
  OR2_X1 U6705 ( .A1(n4312), .A2(n8456), .ZN(n5150) );
  INV_X1 U6706 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5148) );
  OR2_X1 U6707 ( .A1(n5480), .A2(n5148), .ZN(n5149) );
  OR2_X1 U6708 ( .A1(n10087), .A2(n8390), .ZN(n5588) );
  NAND2_X1 U6709 ( .A1(n10087), .A2(n8390), .ZN(n5582) );
  NAND2_X1 U6710 ( .A1(n5588), .A2(n5582), .ZN(n7610) );
  INV_X1 U6711 ( .A(n7610), .ZN(n7600) );
  NAND2_X1 U6712 ( .A1(n7599), .A2(n7600), .ZN(n5153) );
  NAND2_X2 U6713 ( .A1(n5153), .A2(n5582), .ZN(n7516) );
  NAND2_X1 U6714 ( .A1(n5156), .A2(SI_11_), .ZN(n5157) );
  MUX2_X1 U6715 ( .A(n6610), .B(n6608), .S(n5418), .Z(n5159) );
  INV_X1 U6716 ( .A(n5159), .ZN(n5160) );
  NAND2_X1 U6717 ( .A1(n5160), .A2(SI_12_), .ZN(n5161) );
  NAND2_X1 U6718 ( .A1(n5176), .A2(n5161), .ZN(n5174) );
  XNOR2_X1 U6719 ( .A(n5175), .B(n5174), .ZN(n6607) );
  NAND2_X1 U6720 ( .A1(n6607), .A2(n5100), .ZN(n5166) );
  NAND2_X1 U6721 ( .A1(n5163), .A2(n5162), .ZN(n5181) );
  NAND2_X1 U6722 ( .A1(n5181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6723 ( .A(n5164), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6985) );
  AOI22_X1 U6724 ( .A1(n5300), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5299), .B2(
        n6985), .ZN(n5165) );
  NAND2_X1 U6725 ( .A1(n5074), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5173) );
  INV_X1 U6726 ( .A(n4998), .ZN(n5267) );
  INV_X1 U6727 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6984) );
  OR2_X1 U6728 ( .A1(n5267), .A2(n6984), .ZN(n5172) );
  INV_X1 U6729 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8143) );
  NAND2_X1 U6730 ( .A1(n5168), .A2(n8143), .ZN(n5169) );
  NAND2_X1 U6731 ( .A1(n5186), .A2(n5169), .ZN(n8395) );
  OR2_X1 U6732 ( .A1(n4312), .A2(n8395), .ZN(n5171) );
  INV_X1 U6733 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7530) );
  OR2_X1 U6734 ( .A1(n5480), .A2(n7530), .ZN(n5170) );
  NAND2_X1 U6735 ( .A1(n8398), .A2(n7660), .ZN(n7513) );
  INV_X1 U6736 ( .A(n7513), .ZN(n5596) );
  MUX2_X1 U6737 ( .A(n6642), .B(n5177), .S(n5418), .Z(n5178) );
  INV_X1 U6738 ( .A(n5178), .ZN(n5179) );
  NAND2_X1 U6739 ( .A1(n5179), .A2(SI_13_), .ZN(n5180) );
  XNOR2_X1 U6740 ( .A(n5194), .B(n5193), .ZN(n6620) );
  NAND2_X1 U6741 ( .A1(n6620), .A2(n5100), .ZN(n5184) );
  NAND2_X1 U6742 ( .A1(n5182), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6743 ( .A(n5198), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7208) );
  AOI22_X1 U6744 ( .A1(n5300), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5299), .B2(
        n7208), .ZN(n5183) );
  NAND2_X1 U6745 ( .A1(n5074), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5192) );
  INV_X1 U6746 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5185) );
  OR2_X1 U6747 ( .A1(n5267), .A2(n5185), .ZN(n5191) );
  NAND2_X1 U6748 ( .A1(n5186), .A2(n6989), .ZN(n5187) );
  NAND2_X1 U6749 ( .A1(n5205), .A2(n5187), .ZN(n7667) );
  OR2_X1 U6750 ( .A1(n4313), .A2(n7667), .ZN(n5190) );
  INV_X1 U6751 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n5188) );
  OR2_X1 U6752 ( .A1(n5480), .A2(n5188), .ZN(n5189) );
  OR2_X1 U6753 ( .A1(n7681), .A2(n7590), .ZN(n5600) );
  NAND2_X1 U6754 ( .A1(n7681), .A2(n7590), .ZN(n7687) );
  MUX2_X1 U6755 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n5418), .Z(n5215) );
  XNOR2_X1 U6756 ( .A(n5215), .B(n5196), .ZN(n5214) );
  NAND2_X1 U6757 ( .A1(n6660), .A2(n5100), .ZN(n5204) );
  NAND2_X1 U6758 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  NAND2_X1 U6759 ( .A1(n5199), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5201) );
  OR2_X1 U6760 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6761 ( .A1(n5201), .A2(n5200), .ZN(n5222) );
  AOI22_X1 U6762 ( .A1(n5300), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5299), .B2(
        n8508), .ZN(n5203) );
  NAND2_X1 U6763 ( .A1(n5204), .A2(n5203), .ZN(n7775) );
  NAND2_X1 U6764 ( .A1(n5074), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6765 ( .A1(n5205), .A2(n9582), .ZN(n5206) );
  NAND2_X1 U6766 ( .A1(n5229), .A2(n5206), .ZN(n7693) );
  OR2_X1 U6767 ( .A1(n4312), .A2(n7693), .ZN(n5210) );
  INV_X1 U6768 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7694) );
  OR2_X1 U6769 ( .A1(n5480), .A2(n7694), .ZN(n5209) );
  INV_X1 U6770 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5207) );
  OR2_X1 U6771 ( .A1(n5267), .A2(n5207), .ZN(n5208) );
  OR2_X1 U6772 ( .A1(n7775), .A2(n7781), .ZN(n5602) );
  NAND2_X1 U6773 ( .A1(n7775), .A2(n7781), .ZN(n5603) );
  NAND2_X1 U6774 ( .A1(n5602), .A2(n5603), .ZN(n7683) );
  INV_X1 U6775 ( .A(n7687), .ZN(n5212) );
  NOR2_X1 U6776 ( .A1(n7683), .A2(n5212), .ZN(n5213) );
  NAND2_X1 U6777 ( .A1(n5215), .A2(SI_14_), .ZN(n5216) );
  MUX2_X1 U6778 ( .A(n6691), .B(n6689), .S(n5418), .Z(n5219) );
  INV_X1 U6779 ( .A(SI_15_), .ZN(n5218) );
  NAND2_X1 U6780 ( .A1(n5219), .A2(n5218), .ZN(n5238) );
  INV_X1 U6781 ( .A(n5219), .ZN(n5220) );
  NAND2_X1 U6782 ( .A1(n5220), .A2(SI_15_), .ZN(n5221) );
  NAND2_X1 U6783 ( .A1(n5238), .A2(n5221), .ZN(n5236) );
  NAND2_X1 U6784 ( .A1(n6688), .A2(n5100), .ZN(n5225) );
  NAND2_X1 U6785 ( .A1(n5222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5223) );
  XNOR2_X1 U6786 ( .A(n5223), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8526) );
  AOI22_X1 U6787 ( .A1(n5299), .A2(n8526), .B1(n5300), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6788 ( .A1(n4998), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5234) );
  INV_X1 U6789 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5226) );
  OR2_X1 U6790 ( .A1(n5000), .A2(n5226), .ZN(n5233) );
  INV_X1 U6791 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7784) );
  OR2_X1 U6792 ( .A1(n5480), .A2(n7784), .ZN(n5232) );
  INV_X1 U6793 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6794 ( .A1(n5229), .A2(n5228), .ZN(n5230) );
  NAND2_X1 U6795 ( .A1(n5249), .A2(n5230), .ZN(n7783) );
  OR2_X1 U6796 ( .A1(n4312), .A2(n7783), .ZN(n5231) );
  INV_X1 U6797 ( .A(n5608), .ZN(n5235) );
  NAND2_X1 U6798 ( .A1(n8603), .A2(n8841), .ZN(n5607) );
  MUX2_X1 U6799 ( .A(n6836), .B(n6837), .S(n5418), .Z(n5239) );
  NAND2_X1 U6800 ( .A1(n5239), .A2(n9738), .ZN(n5259) );
  INV_X1 U6801 ( .A(n5239), .ZN(n5240) );
  NAND2_X1 U6802 ( .A1(n5240), .A2(SI_16_), .ZN(n5241) );
  XNOR2_X1 U6803 ( .A(n5258), .B(n5257), .ZN(n6835) );
  NAND2_X1 U6804 ( .A1(n6835), .A2(n5100), .ZN(n5248) );
  NAND2_X1 U6805 ( .A1(n5242), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5243) );
  MUX2_X1 U6806 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5243), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5246) );
  INV_X1 U6807 ( .A(n5244), .ZN(n5245) );
  NAND2_X1 U6808 ( .A1(n5246), .A2(n5245), .ZN(n8545) );
  INV_X1 U6809 ( .A(n8545), .ZN(n8538) );
  AOI22_X1 U6810 ( .A1(n5300), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5299), .B2(
        n8538), .ZN(n5247) );
  NAND2_X1 U6811 ( .A1(n5074), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5255) );
  INV_X1 U6812 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8544) );
  OR2_X1 U6813 ( .A1(n5267), .A2(n8544), .ZN(n5254) );
  NAND2_X1 U6814 ( .A1(n5249), .A2(n9735), .ZN(n5250) );
  NAND2_X1 U6815 ( .A1(n5269), .A2(n5250), .ZN(n8851) );
  OR2_X1 U6816 ( .A1(n4312), .A2(n8851), .ZN(n5253) );
  INV_X1 U6817 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n5251) );
  OR2_X1 U6818 ( .A1(n5480), .A2(n5251), .ZN(n5252) );
  OR2_X1 U6819 ( .A1(n8938), .A2(n8820), .ZN(n5610) );
  NAND2_X1 U6820 ( .A1(n8836), .A2(n5610), .ZN(n5256) );
  NAND2_X1 U6821 ( .A1(n8938), .A2(n8820), .ZN(n5611) );
  MUX2_X1 U6822 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n5418), .Z(n5277) );
  XNOR2_X1 U6823 ( .A(n5277), .B(n5260), .ZN(n5276) );
  XNOR2_X1 U6824 ( .A(n5278), .B(n5276), .ZN(n6778) );
  NAND2_X1 U6825 ( .A1(n6778), .A2(n5100), .ZN(n5265) );
  NOR2_X1 U6826 ( .A1(n5244), .A2(n4919), .ZN(n5261) );
  MUX2_X1 U6827 ( .A(n4919), .B(n5261), .S(P2_IR_REG_17__SCAN_IN), .Z(n5262)
         );
  INV_X1 U6828 ( .A(n5262), .ZN(n5263) );
  AND2_X1 U6829 ( .A1(n5279), .A2(n5263), .ZN(n8559) );
  AOI22_X1 U6830 ( .A1(n5300), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5299), .B2(
        n8559), .ZN(n5264) );
  NAND2_X1 U6831 ( .A1(n5074), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5274) );
  INV_X1 U6832 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5266) );
  OR2_X1 U6833 ( .A1(n5267), .A2(n5266), .ZN(n5273) );
  INV_X1 U6834 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9691) );
  NAND2_X1 U6835 ( .A1(n5269), .A2(n9691), .ZN(n5270) );
  NAND2_X1 U6836 ( .A1(n5283), .A2(n5270), .ZN(n8829) );
  OR2_X1 U6837 ( .A1(n4313), .A2(n8829), .ZN(n5272) );
  INV_X1 U6838 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8830) );
  OR2_X1 U6839 ( .A1(n5480), .A2(n8830), .ZN(n5271) );
  NAND2_X1 U6840 ( .A1(n8934), .A2(n8839), .ZN(n5540) );
  NAND2_X1 U6841 ( .A1(n5539), .A2(n5540), .ZN(n8815) );
  MUX2_X1 U6842 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n5418), .Z(n5293) );
  XNOR2_X1 U6843 ( .A(n5293), .B(SI_18_), .ZN(n5291) );
  XNOR2_X1 U6844 ( .A(n5292), .B(n5291), .ZN(n6995) );
  NAND2_X1 U6845 ( .A1(n6995), .A2(n5100), .ZN(n5282) );
  NAND2_X1 U6846 ( .A1(n5279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5280) );
  XNOR2_X1 U6847 ( .A(n5280), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8573) );
  AOI22_X1 U6848 ( .A1(n5300), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5299), .B2(
        n8573), .ZN(n5281) );
  NAND2_X1 U6849 ( .A1(n4998), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5290) );
  INV_X1 U6850 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U6851 ( .A1(n5283), .A2(n9650), .ZN(n5284) );
  AND2_X1 U6852 ( .A1(n5304), .A2(n5284), .ZN(n8798) );
  NAND2_X1 U6853 ( .A1(n4959), .A2(n8798), .ZN(n5289) );
  INV_X1 U6854 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5285) );
  OR2_X1 U6855 ( .A1(n5000), .A2(n5285), .ZN(n5288) );
  INV_X1 U6856 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5286) );
  OR2_X1 U6857 ( .A1(n5480), .A2(n5286), .ZN(n5287) );
  NAND4_X1 U6858 ( .A1(n5290), .A2(n5289), .A3(n5288), .A4(n5287), .ZN(n8788)
         );
  INV_X1 U6859 ( .A(n8788), .ZN(n8819) );
  OR2_X1 U6860 ( .A1(n8929), .A2(n8819), .ZN(n5622) );
  NAND2_X1 U6861 ( .A1(n8929), .A2(n8819), .ZN(n5614) );
  NAND2_X1 U6862 ( .A1(n8802), .A2(n5614), .ZN(n8786) );
  NAND2_X1 U6863 ( .A1(n5293), .A2(SI_18_), .ZN(n5294) );
  MUX2_X1 U6864 ( .A(n7179), .B(n7177), .S(n5418), .Z(n5295) );
  NAND2_X1 U6865 ( .A1(n5295), .A2(n9742), .ZN(n5313) );
  INV_X1 U6866 ( .A(n5295), .ZN(n5296) );
  NAND2_X1 U6867 ( .A1(n5296), .A2(SI_19_), .ZN(n5297) );
  NAND2_X1 U6868 ( .A1(n5313), .A2(n5297), .ZN(n5311) );
  XNOR2_X1 U6869 ( .A(n5310), .B(n5311), .ZN(n7176) );
  NAND2_X1 U6870 ( .A1(n7176), .A2(n5100), .ZN(n5302) );
  XNOR2_X2 U6871 ( .A(n5510), .B(n5509), .ZN(n8828) );
  AOI22_X1 U6872 ( .A1(n5300), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8583), .B2(
        n5299), .ZN(n5301) );
  INV_X1 U6873 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6874 ( .A1(n5304), .A2(n5303), .ZN(n5305) );
  NAND2_X1 U6875 ( .A1(n5320), .A2(n5305), .ZN(n8369) );
  INV_X1 U6876 ( .A(n8369), .ZN(n8782) );
  NAND2_X1 U6877 ( .A1(n8782), .A2(n4959), .ZN(n5309) );
  NAND2_X1 U6878 ( .A1(n4998), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6879 ( .A1(n5074), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5307) );
  INV_X1 U6880 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8577) );
  OR2_X1 U6881 ( .A1(n5480), .A2(n8577), .ZN(n5306) );
  NAND4_X1 U6882 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n8807)
         );
  INV_X1 U6883 ( .A(n8807), .ZN(n8609) );
  OR2_X1 U6884 ( .A1(n8925), .A2(n8609), .ZN(n5623) );
  NAND2_X1 U6885 ( .A1(n8925), .A2(n8609), .ZN(n8763) );
  INV_X1 U6886 ( .A(n5311), .ZN(n5312) );
  MUX2_X1 U6887 ( .A(n8259), .B(n7373), .S(n5418), .Z(n5315) );
  NAND2_X1 U6888 ( .A1(n5315), .A2(n9633), .ZN(n5330) );
  INV_X1 U6889 ( .A(n5315), .ZN(n5316) );
  NAND2_X1 U6890 ( .A1(n5316), .A2(SI_20_), .ZN(n5317) );
  XNOR2_X1 U6891 ( .A(n5329), .B(n5328), .ZN(n7372) );
  NAND2_X1 U6892 ( .A1(n7372), .A2(n5100), .ZN(n5319) );
  OR2_X1 U6893 ( .A1(n5505), .A2(n8259), .ZN(n5318) );
  INV_X1 U6894 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U6895 ( .A1(n5320), .A2(n9694), .ZN(n5321) );
  AND2_X1 U6896 ( .A1(n5350), .A2(n5321), .ZN(n8773) );
  NAND2_X1 U6897 ( .A1(n8773), .A2(n4959), .ZN(n5324) );
  AOI22_X1 U6898 ( .A1(n4998), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n5074), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6899 ( .A1(n4935), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6900 ( .A1(n8919), .A2(n8610), .ZN(n5626) );
  NAND2_X1 U6901 ( .A1(n5629), .A2(n5626), .ZN(n8767) );
  INV_X1 U6902 ( .A(n8763), .ZN(n5325) );
  NOR2_X1 U6903 ( .A1(n8767), .A2(n5325), .ZN(n5327) );
  MUX2_X1 U6904 ( .A(n7388), .B(n7402), .S(n5418), .Z(n5339) );
  XNOR2_X1 U6905 ( .A(n5339), .B(SI_21_), .ZN(n5338) );
  XNOR2_X1 U6906 ( .A(n5342), .B(n5338), .ZN(n7386) );
  NAND2_X1 U6907 ( .A1(n7386), .A2(n5100), .ZN(n5332) );
  OR2_X1 U6908 ( .A1(n5505), .A2(n7388), .ZN(n5331) );
  XNOR2_X1 U6909 ( .A(n5350), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8753) );
  INV_X1 U6910 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5335) );
  NAND2_X1 U6911 ( .A1(n4998), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5334) );
  NAND2_X1 U6912 ( .A1(n5074), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5333) );
  OAI211_X1 U6913 ( .C1(n5335), .C2(n5480), .A(n5334), .B(n5333), .ZN(n5336)
         );
  AOI21_X1 U6914 ( .B1(n8753), .B2(n4959), .A(n5336), .ZN(n8611) );
  OR2_X1 U6915 ( .A1(n8912), .A2(n8611), .ZN(n5617) );
  NAND2_X1 U6916 ( .A1(n8912), .A2(n8611), .ZN(n8741) );
  NAND2_X1 U6917 ( .A1(n5617), .A2(n8741), .ZN(n8756) );
  INV_X1 U6918 ( .A(n5338), .ZN(n5341) );
  INV_X1 U6919 ( .A(n5339), .ZN(n5340) );
  MUX2_X1 U6920 ( .A(n8344), .B(n7493), .S(n5418), .Z(n5344) );
  INV_X1 U6921 ( .A(SI_22_), .ZN(n5343) );
  NAND2_X1 U6922 ( .A1(n5344), .A2(n5343), .ZN(n5364) );
  INV_X1 U6923 ( .A(n5344), .ZN(n5345) );
  NAND2_X1 U6924 ( .A1(n5345), .A2(SI_22_), .ZN(n5346) );
  NAND2_X1 U6925 ( .A1(n5364), .A2(n5346), .ZN(n5362) );
  XNOR2_X1 U6926 ( .A(n5363), .B(n5362), .ZN(n7492) );
  NAND2_X1 U6927 ( .A1(n7492), .A2(n5100), .ZN(n5348) );
  OR2_X1 U6928 ( .A1(n5505), .A2(n8344), .ZN(n5347) );
  INV_X1 U6929 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9708) );
  INV_X1 U6930 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5349) );
  OAI21_X1 U6931 ( .B1(n5350), .B2(n9708), .A(n5349), .ZN(n5353) );
  AND2_X1 U6932 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5351) );
  NAND2_X1 U6933 ( .A1(n5353), .A2(n5372), .ZN(n8736) );
  OR2_X1 U6934 ( .A1(n8736), .A2(n4313), .ZN(n5359) );
  INV_X1 U6935 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U6936 ( .A1(n4998), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6937 ( .A1(n5074), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5354) );
  OAI211_X1 U6938 ( .C1(n5356), .C2(n5480), .A(n5355), .B(n5354), .ZN(n5357)
         );
  INV_X1 U6939 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6940 ( .A1(n8907), .A2(n8612), .ZN(n5618) );
  NAND2_X1 U6941 ( .A1(n5360), .A2(n5618), .ZN(n8743) );
  INV_X1 U6942 ( .A(n8741), .ZN(n5628) );
  NOR2_X1 U6943 ( .A1(n8743), .A2(n5628), .ZN(n5361) );
  INV_X1 U6944 ( .A(n5360), .ZN(n5632) );
  INV_X1 U6945 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5366) );
  MUX2_X1 U6946 ( .A(n7635), .B(n5366), .S(n5418), .Z(n5367) );
  INV_X1 U6947 ( .A(SI_23_), .ZN(n9698) );
  NAND2_X1 U6948 ( .A1(n5367), .A2(n9698), .ZN(n5382) );
  INV_X1 U6949 ( .A(n5367), .ZN(n5368) );
  NAND2_X1 U6950 ( .A1(n5368), .A2(SI_23_), .ZN(n5369) );
  NAND2_X1 U6951 ( .A1(n7632), .A2(n5100), .ZN(n5371) );
  OR2_X1 U6952 ( .A1(n5505), .A2(n7635), .ZN(n5370) );
  INV_X1 U6953 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9724) );
  NAND2_X1 U6954 ( .A1(n5372), .A2(n9724), .ZN(n5373) );
  AND2_X1 U6955 ( .A1(n5386), .A2(n5373), .ZN(n8724) );
  NAND2_X1 U6956 ( .A1(n8724), .A2(n4959), .ZN(n5379) );
  INV_X1 U6957 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6958 ( .A1(n4998), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6959 ( .A1(n5074), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5374) );
  OAI211_X1 U6960 ( .C1(n5376), .C2(n5480), .A(n5375), .B(n5374), .ZN(n5377)
         );
  INV_X1 U6961 ( .A(n5377), .ZN(n5378) );
  XNOR2_X1 U6962 ( .A(n8902), .B(n8713), .ZN(n8721) );
  INV_X1 U6963 ( .A(n8721), .ZN(n8727) );
  INV_X1 U6964 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7703) );
  MUX2_X1 U6965 ( .A(n7701), .B(n7703), .S(n5418), .Z(n5397) );
  XNOR2_X1 U6966 ( .A(n5397), .B(SI_24_), .ZN(n5396) );
  XNOR2_X1 U6967 ( .A(n5395), .B(n5396), .ZN(n7700) );
  NAND2_X1 U6968 ( .A1(n7700), .A2(n5100), .ZN(n5384) );
  OR2_X1 U6969 ( .A1(n5505), .A2(n7701), .ZN(n5383) );
  INV_X1 U6970 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9705) );
  NAND2_X1 U6971 ( .A1(n5386), .A2(n9705), .ZN(n5387) );
  NAND2_X1 U6972 ( .A1(n5407), .A2(n5387), .ZN(n8703) );
  OR2_X1 U6973 ( .A1(n8703), .A2(n4312), .ZN(n5393) );
  INV_X1 U6974 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6975 ( .A1(n4998), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5389) );
  NAND2_X1 U6976 ( .A1(n5074), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5388) );
  OAI211_X1 U6977 ( .C1(n5390), .C2(n5480), .A(n5389), .B(n5388), .ZN(n5391)
         );
  INV_X1 U6978 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6979 ( .A1(n8897), .A2(n8423), .ZN(n5643) );
  AND2_X1 U6980 ( .A1(n8902), .A2(n8713), .ZN(n8709) );
  NOR2_X1 U6981 ( .A1(n8708), .A2(n8709), .ZN(n5394) );
  NAND2_X1 U6982 ( .A1(n8707), .A2(n5394), .ZN(n8711) );
  NAND2_X1 U6983 ( .A1(n8711), .A2(n5646), .ZN(n8687) );
  INV_X1 U6984 ( .A(n5397), .ZN(n5398) );
  NAND2_X1 U6985 ( .A1(n5398), .A2(SI_24_), .ZN(n5399) );
  INV_X1 U6986 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7748) );
  INV_X1 U6987 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U6988 ( .A(n7748), .B(n7751), .S(n5418), .Z(n5402) );
  INV_X1 U6989 ( .A(SI_25_), .ZN(n5401) );
  NAND2_X1 U6990 ( .A1(n5402), .A2(n5401), .ZN(n5416) );
  INV_X1 U6991 ( .A(n5402), .ZN(n5403) );
  NAND2_X1 U6992 ( .A1(n5403), .A2(SI_25_), .ZN(n5404) );
  NAND2_X1 U6993 ( .A1(n5416), .A2(n5404), .ZN(n5414) );
  XNOR2_X1 U6994 ( .A(n5415), .B(n5414), .ZN(n7745) );
  NAND2_X1 U6995 ( .A1(n7745), .A2(n5100), .ZN(n5406) );
  OR2_X1 U6996 ( .A1(n5505), .A2(n7748), .ZN(n5405) );
  INV_X1 U6997 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U6998 ( .A1(n5407), .A2(n9712), .ZN(n5408) );
  AND2_X1 U6999 ( .A1(n5426), .A2(n5408), .ZN(n8693) );
  NAND2_X1 U7000 ( .A1(n8693), .A2(n4959), .ZN(n5413) );
  INV_X1 U7001 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U7002 ( .A1(n4998), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5410) );
  NAND2_X1 U7003 ( .A1(n5074), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5409) );
  OAI211_X1 U7004 ( .C1(n8695), .C2(n5480), .A(n5410), .B(n5409), .ZN(n5411)
         );
  INV_X1 U7005 ( .A(n5411), .ZN(n5412) );
  NAND2_X1 U7006 ( .A1(n8893), .A2(n8714), .ZN(n5647) );
  INV_X1 U7007 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7803) );
  INV_X1 U7008 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7805) );
  MUX2_X1 U7009 ( .A(n7803), .B(n7805), .S(n5418), .Z(n5419) );
  INV_X1 U7010 ( .A(SI_26_), .ZN(n9743) );
  NAND2_X1 U7011 ( .A1(n5419), .A2(n9743), .ZN(n5436) );
  INV_X1 U7012 ( .A(n5419), .ZN(n5420) );
  NAND2_X1 U7013 ( .A1(n5420), .A2(SI_26_), .ZN(n5421) );
  NAND2_X1 U7014 ( .A1(n7802), .A2(n5100), .ZN(n5423) );
  OR2_X1 U7015 ( .A1(n5505), .A2(n7803), .ZN(n5422) );
  INV_X1 U7016 ( .A(n5426), .ZN(n5424) );
  NAND2_X1 U7017 ( .A1(n5424), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5443) );
  INV_X1 U7018 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U7019 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  NAND2_X1 U7020 ( .A1(n5443), .A2(n5427), .ZN(n8672) );
  INV_X1 U7021 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U7022 ( .A1(n4998), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5429) );
  NAND2_X1 U7023 ( .A1(n5074), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5428) );
  OAI211_X1 U7024 ( .C1(n8673), .C2(n5480), .A(n5429), .B(n5428), .ZN(n5430)
         );
  INV_X1 U7025 ( .A(n5430), .ZN(n5431) );
  NAND2_X1 U7026 ( .A1(n8888), .A2(n8404), .ZN(n5651) );
  INV_X1 U7027 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8974) );
  INV_X1 U7028 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5437) );
  MUX2_X1 U7029 ( .A(n8974), .B(n5437), .S(n5418), .Z(n5438) );
  INV_X1 U7030 ( .A(SI_27_), .ZN(n9737) );
  NAND2_X1 U7031 ( .A1(n5438), .A2(n9737), .ZN(n5453) );
  INV_X1 U7032 ( .A(n5438), .ZN(n5439) );
  NAND2_X1 U7033 ( .A1(n5439), .A2(SI_27_), .ZN(n5440) );
  NAND2_X1 U7034 ( .A1(n7807), .A2(n5100), .ZN(n5442) );
  OR2_X1 U7035 ( .A1(n5505), .A2(n8974), .ZN(n5441) );
  INV_X1 U7036 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9734) );
  NAND2_X1 U7037 ( .A1(n5443), .A2(n9734), .ZN(n5444) );
  NAND2_X1 U7038 ( .A1(n8656), .A2(n4959), .ZN(n5450) );
  INV_X1 U7039 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U7040 ( .A1(n4998), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5446) );
  NAND2_X1 U7041 ( .A1(n5074), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5445) );
  OAI211_X1 U7042 ( .C1(n5447), .C2(n5480), .A(n5446), .B(n5445), .ZN(n5448)
         );
  INV_X1 U7043 ( .A(n5448), .ZN(n5449) );
  OR2_X1 U7044 ( .A1(n8881), .A2(n8681), .ZN(n5656) );
  MUX2_X1 U7045 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6496), .Z(n5471) );
  INV_X1 U7046 ( .A(SI_28_), .ZN(n5472) );
  XNOR2_X1 U7047 ( .A(n5471), .B(n5472), .ZN(n5469) );
  NAND2_X1 U7048 ( .A1(n8966), .A2(n5100), .ZN(n5457) );
  INV_X1 U7049 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5455) );
  OR2_X1 U7050 ( .A1(n5505), .A2(n5455), .ZN(n5456) );
  INV_X1 U7051 ( .A(n5460), .ZN(n5458) );
  NAND2_X1 U7052 ( .A1(n5458), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5476) );
  INV_X1 U7053 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7054 ( .A1(n5460), .A2(n5459), .ZN(n5461) );
  NAND2_X1 U7055 ( .A1(n5476), .A2(n5461), .ZN(n8645) );
  INV_X1 U7056 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8646) );
  NAND2_X1 U7057 ( .A1(n4998), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U7058 ( .A1(n5074), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U7059 ( .C1(n8646), .C2(n5480), .A(n5464), .B(n5463), .ZN(n5465)
         );
  INV_X1 U7060 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U7061 ( .A1(n8876), .A2(n8632), .ZN(n5661) );
  INV_X1 U7062 ( .A(n8641), .ZN(n5468) );
  INV_X1 U7063 ( .A(n5471), .ZN(n5473) );
  NAND2_X1 U7064 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  MUX2_X1 U7065 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6496), .Z(n5489) );
  INV_X1 U7066 ( .A(SI_29_), .ZN(n9635) );
  XNOR2_X1 U7067 ( .A(n5489), .B(n9635), .ZN(n5487) );
  INV_X1 U7068 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8964) );
  NOR2_X1 U7069 ( .A1(n5505), .A2(n8964), .ZN(n5475) );
  INV_X1 U7070 ( .A(n8625), .ZN(n8869) );
  INV_X1 U7071 ( .A(n5476), .ZN(n8623) );
  NAND2_X1 U7072 ( .A1(n8623), .A2(n4959), .ZN(n5483) );
  INV_X1 U7073 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U7074 ( .A1(n5074), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7075 ( .A1(n4998), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5477) );
  OAI211_X1 U7076 ( .C1(n5480), .C2(n5479), .A(n5478), .B(n5477), .ZN(n5481)
         );
  INV_X1 U7077 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U7078 ( .A1(n5483), .A2(n5482), .ZN(n8491) );
  INV_X1 U7079 ( .A(n8491), .ZN(n5484) );
  INV_X1 U7080 ( .A(n5667), .ZN(n5485) );
  INV_X1 U7081 ( .A(n5489), .ZN(n5490) );
  MUX2_X1 U7082 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6496), .Z(n5495) );
  INV_X1 U7083 ( .A(SI_30_), .ZN(n5497) );
  XNOR2_X1 U7084 ( .A(n5495), .B(n5497), .ZN(n5491) );
  NAND2_X1 U7085 ( .A1(n8134), .A2(n5100), .ZN(n5493) );
  INV_X1 U7086 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8135) );
  OR2_X1 U7087 ( .A1(n5505), .A2(n8135), .ZN(n5492) );
  NAND2_X1 U7088 ( .A1(n5498), .A2(n5497), .ZN(n5496) );
  NAND2_X1 U7089 ( .A1(n5496), .A2(n5495), .ZN(n5500) );
  MUX2_X1 U7090 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6496), .Z(n5501) );
  XNOR2_X1 U7091 ( .A(n5501), .B(SI_31_), .ZN(n5502) );
  NAND2_X1 U7092 ( .A1(n8959), .A2(n5100), .ZN(n5507) );
  INV_X1 U7093 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5504) );
  OR2_X1 U7094 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  OR2_X1 U7095 ( .A1(n8862), .A2(n5508), .ZN(n5518) );
  NAND2_X1 U7096 ( .A1(n8865), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U7097 ( .A1(n5518), .A2(n5534), .ZN(n5673) );
  INV_X1 U7098 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5512) );
  XNOR2_X2 U7099 ( .A(n5682), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6934) );
  NAND2_X1 U7100 ( .A1(n6731), .A2(n5536), .ZN(n6943) );
  NAND2_X1 U7101 ( .A1(n8295), .A2(n6943), .ZN(n5515) );
  INV_X1 U7102 ( .A(n6944), .ZN(n5517) );
  INV_X1 U7103 ( .A(n5518), .ZN(n5678) );
  NAND2_X1 U7104 ( .A1(n5610), .A2(n5611), .ZN(n8842) );
  NAND2_X1 U7105 ( .A1(n5608), .A2(n5607), .ZN(n8604) );
  INV_X1 U7106 ( .A(n7158), .ZN(n10015) );
  NAND2_X1 U7107 ( .A1(n6763), .A2(n10015), .ZN(n5545) );
  AND2_X1 U7108 ( .A1(n5519), .A2(n5545), .ZN(n10017) );
  NAND2_X1 U7109 ( .A1(n7125), .A2(n5520), .ZN(n5559) );
  INV_X1 U7110 ( .A(n5559), .ZN(n5521) );
  NAND4_X1 U7111 ( .A1(n10017), .A2(n5521), .A3(n5536), .A4(n7109), .ZN(n5523)
         );
  NAND2_X1 U7112 ( .A1(n5555), .A2(n5522), .ZN(n5563) );
  NAND2_X1 U7113 ( .A1(n5542), .A2(n5543), .ZN(n6936) );
  NOR4_X1 U7114 ( .A1(n5523), .A2(n5563), .A3(n7060), .A4(n6936), .ZN(n5524)
         );
  NAND4_X1 U7115 ( .A1(n5524), .A2(n7166), .A3(n7154), .A4(n7416), .ZN(n5525)
         );
  INV_X1 U7116 ( .A(n5582), .ZN(n5592) );
  NOR4_X1 U7117 ( .A1(n5525), .A2(n5592), .A3(n7523), .A4(n7543), .ZN(n5526)
         );
  AND2_X1 U7118 ( .A1(n7514), .A2(n5588), .ZN(n5594) );
  NAND4_X1 U7119 ( .A1(n5526), .A2(n7653), .A3(n5594), .A4(n7513), .ZN(n5527)
         );
  NOR4_X1 U7120 ( .A1(n8842), .A2(n8604), .A3(n7683), .A4(n5527), .ZN(n5528)
         );
  NAND4_X1 U7121 ( .A1(n8787), .A2(n4458), .A3(n4317), .A4(n5528), .ZN(n5529)
         );
  NOR4_X1 U7122 ( .A1(n8743), .A2(n8756), .A3(n8767), .A4(n5529), .ZN(n5530)
         );
  NAND4_X1 U7123 ( .A1(n4652), .A2(n8613), .A3(n5530), .A4(n8727), .ZN(n5531)
         );
  NOR4_X1 U7124 ( .A1(n8641), .A2(n8652), .A3(n8679), .A4(n5531), .ZN(n5532)
         );
  XNOR2_X1 U7125 ( .A(n5535), .B(n8583), .ZN(n5537) );
  NAND2_X1 U7126 ( .A1(n6731), .A2(n8583), .ZN(n5538) );
  OR2_X1 U7127 ( .A1(n6934), .A2(n5538), .ZN(n5552) );
  INV_X1 U7128 ( .A(n5552), .ZN(n5662) );
  OAI21_X1 U7129 ( .B1(n8758), .B2(n5677), .A(n8907), .ZN(n5637) );
  INV_X1 U7130 ( .A(n8907), .ZN(n8739) );
  OAI21_X1 U7131 ( .B1(n8612), .B2(n5662), .A(n8739), .ZN(n5636) );
  AOI22_X1 U7132 ( .A1(n4317), .A2(n5540), .B1(n5622), .B2(n5677), .ZN(n5613)
         );
  NAND2_X1 U7133 ( .A1(n5542), .A2(n5541), .ZN(n5547) );
  OAI21_X1 U7134 ( .B1(n5547), .B2(n5543), .A(n7098), .ZN(n5551) );
  INV_X1 U7135 ( .A(n5545), .ZN(n6925) );
  NOR2_X1 U7136 ( .A1(n5547), .A2(n6925), .ZN(n5544) );
  NAND2_X1 U7137 ( .A1(n5545), .A2(n6731), .ZN(n5546) );
  NAND2_X1 U7138 ( .A1(n5519), .A2(n5546), .ZN(n5549) );
  INV_X1 U7139 ( .A(n5547), .ZN(n5548) );
  AND2_X1 U7140 ( .A1(n5549), .A2(n5548), .ZN(n5550) );
  NOR2_X1 U7141 ( .A1(n5551), .A2(n5550), .ZN(n5553) );
  NAND2_X1 U7142 ( .A1(n5565), .A2(n5557), .ZN(n5561) );
  NAND2_X1 U7143 ( .A1(n5570), .A2(n7109), .ZN(n5558) );
  AOI21_X1 U7144 ( .B1(n5565), .B2(n5559), .A(n5558), .ZN(n5560) );
  INV_X1 U7145 ( .A(n7152), .ZN(n5564) );
  AOI21_X1 U7146 ( .B1(n5566), .B2(n5568), .A(n5671), .ZN(n5567) );
  AOI21_X1 U7147 ( .B1(n5569), .B2(n5568), .A(n5567), .ZN(n5572) );
  OAI21_X1 U7148 ( .B1(n5570), .B2(n5677), .A(n7166), .ZN(n5571) );
  MUX2_X1 U7149 ( .A(n5574), .B(n5573), .S(n5662), .Z(n5575) );
  INV_X1 U7150 ( .A(n5580), .ZN(n5577) );
  AOI21_X1 U7151 ( .B1(n5580), .B2(n7168), .A(n10064), .ZN(n5579) );
  INV_X1 U7152 ( .A(n5581), .ZN(n5578) );
  NAND3_X1 U7153 ( .A1(n5583), .A2(n5582), .A3(n5585), .ZN(n5591) );
  NAND3_X1 U7154 ( .A1(n5586), .A2(n5585), .A3(n5584), .ZN(n5589) );
  NAND3_X1 U7155 ( .A1(n5589), .A2(n5588), .A3(n5587), .ZN(n5590) );
  NOR2_X1 U7156 ( .A1(n5596), .A2(n5592), .ZN(n5593) );
  MUX2_X1 U7157 ( .A(n5594), .B(n5593), .S(n5671), .Z(n5598) );
  INV_X1 U7158 ( .A(n7514), .ZN(n5595) );
  MUX2_X1 U7159 ( .A(n5596), .B(n5595), .S(n5671), .Z(n5597) );
  INV_X1 U7160 ( .A(n7683), .ZN(n7686) );
  MUX2_X1 U7161 ( .A(n5600), .B(n7687), .S(n5671), .Z(n5601) );
  NAND2_X1 U7162 ( .A1(n7686), .A2(n5601), .ZN(n5605) );
  INV_X1 U7163 ( .A(n8604), .ZN(n7778) );
  MUX2_X1 U7164 ( .A(n5603), .B(n5602), .S(n5671), .Z(n5604) );
  INV_X1 U7165 ( .A(n8842), .ZN(n8837) );
  MUX2_X1 U7166 ( .A(n5608), .B(n5607), .S(n5671), .Z(n5609) );
  MUX2_X1 U7167 ( .A(n5611), .B(n5610), .S(n5671), .Z(n5612) );
  INV_X1 U7168 ( .A(n5614), .ZN(n5615) );
  OAI21_X1 U7169 ( .B1(n5625), .B2(n5615), .A(n5623), .ZN(n5616) );
  NAND4_X1 U7170 ( .A1(n5616), .A2(n5626), .A3(n8763), .A4(n5677), .ZN(n5621)
         );
  INV_X1 U7171 ( .A(n5617), .ZN(n5631) );
  OAI21_X1 U7172 ( .B1(n5631), .B2(n5326), .A(n5677), .ZN(n5620) );
  INV_X1 U7173 ( .A(n5618), .ZN(n5619) );
  AOI211_X1 U7174 ( .C1(n5621), .C2(n5620), .A(n5619), .B(n5628), .ZN(n5635)
         );
  NAND2_X1 U7175 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  OAI21_X1 U7176 ( .B1(n5625), .B2(n5624), .A(n8763), .ZN(n5630) );
  INV_X1 U7177 ( .A(n5626), .ZN(n5627) );
  NOR4_X1 U7178 ( .A1(n5633), .A2(n5632), .A3(n5631), .A4(n5677), .ZN(n5634)
         );
  INV_X1 U7179 ( .A(n5643), .ZN(n5640) );
  OAI21_X1 U7180 ( .B1(n8713), .B2(n8902), .A(n5646), .ZN(n5638) );
  MUX2_X1 U7181 ( .A(n5638), .B(n8709), .S(n5677), .Z(n5639) );
  INV_X1 U7182 ( .A(n5641), .ZN(n5642) );
  OAI21_X1 U7183 ( .B1(n5644), .B2(n5677), .A(n5653), .ZN(n5652) );
  INV_X1 U7184 ( .A(n5645), .ZN(n5649) );
  INV_X1 U7185 ( .A(n5646), .ZN(n5648) );
  OAI211_X1 U7186 ( .C1(n5649), .C2(n5648), .A(n5651), .B(n5647), .ZN(n5650)
         );
  AOI22_X1 U7187 ( .A1(n5652), .A2(n5651), .B1(n5671), .B2(n5650), .ZN(n5660)
         );
  INV_X1 U7188 ( .A(n8652), .ZN(n8658) );
  OAI21_X1 U7189 ( .B1(n5662), .B2(n5653), .A(n8658), .ZN(n5659) );
  INV_X1 U7190 ( .A(n5661), .ZN(n5654) );
  AOI21_X1 U7191 ( .B1(n8681), .B2(n8881), .A(n5654), .ZN(n5655) );
  MUX2_X1 U7192 ( .A(n5656), .B(n5655), .S(n5671), .Z(n5657) );
  OAI211_X1 U7193 ( .C1(n5660), .C2(n5659), .A(n5658), .B(n5657), .ZN(n5666)
         );
  OAI21_X1 U7194 ( .B1(n5662), .B2(n8876), .A(n5661), .ZN(n5663) );
  OAI22_X1 U7195 ( .A1(n5664), .A2(n5663), .B1(n5662), .B2(n8660), .ZN(n5665)
         );
  AOI22_X1 U7196 ( .A1(n5666), .A2(n5665), .B1(n5664), .B2(n5552), .ZN(n5668)
         );
  NAND2_X1 U7197 ( .A1(n5670), .A2(n5669), .ZN(n5672) );
  MUX2_X1 U7198 ( .A(n5673), .B(n5672), .S(n5671), .Z(n5674) );
  MUX2_X1 U7199 ( .A(n4870), .B(n5678), .S(n5677), .Z(n5679) );
  NAND2_X1 U7200 ( .A1(n6875), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7633) );
  INV_X1 U7201 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5685) );
  NAND2_X1 U7202 ( .A1(n5689), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5690) );
  OR2_X1 U7203 ( .A1(n5691), .A2(n4919), .ZN(n5692) );
  NAND2_X1 U7204 ( .A1(n6739), .A2(n5693), .ZN(n6878) );
  NAND2_X1 U7205 ( .A1(n6934), .A2(n6731), .ZN(n6797) );
  OR2_X1 U7206 ( .A1(n6797), .A2(n6760), .ZN(n6876) );
  NAND2_X1 U7207 ( .A1(n10008), .A2(n6876), .ZN(n7181) );
  INV_X1 U7208 ( .A(n6797), .ZN(n6753) );
  INV_X1 U7209 ( .A(n6803), .ZN(n6762) );
  NOR3_X1 U7210 ( .A1(n7181), .A2(n8971), .A3(n8840), .ZN(n5695) );
  OAI21_X1 U7211 ( .B1(n7633), .B2(n6934), .A(P2_B_REG_SCAN_IN), .ZN(n5694) );
  INV_X1 U7212 ( .A(n5928), .ZN(n5707) );
  NAND4_X2 U7213 ( .A1(n5702), .A2(n5701), .A3(n5700), .A4(n5699), .ZN(n5724)
         );
  NOR2_X1 U7214 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5704) );
  NOR2_X1 U7215 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5703) );
  NAND4_X1 U7216 ( .A1(n5704), .A2(n5703), .A3(n5726), .A4(n5749), .ZN(n5705)
         );
  NAND2_X1 U7217 ( .A1(n5735), .A2(n5708), .ZN(n5709) );
  XNOR2_X2 U7218 ( .A(n5712), .B(n5711), .ZN(n8131) );
  INV_X1 U7219 ( .A(n8338), .ZN(n5716) );
  NAND2_X2 U7220 ( .A1(n8131), .A2(n5716), .ZN(n5805) );
  INV_X1 U7221 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5717) );
  INV_X1 U7222 ( .A(n8131), .ZN(n5718) );
  AND2_X2 U7223 ( .A1(n5718), .A2(n8338), .ZN(n5878) );
  NAND2_X1 U7224 ( .A1(n5878), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5722) );
  INV_X1 U7225 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6918) );
  INV_X1 U7226 ( .A(n5803), .ZN(n5719) );
  NAND2_X1 U7227 ( .A1(n5719), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5720) );
  NAND4_X2 U7228 ( .A1(n5723), .A2(n5722), .A3(n5721), .A4(n5720), .ZN(n6376)
         );
  AND2_X2 U7229 ( .A1(n5944), .A2(n5725), .ZN(n5747) );
  XNOR2_X2 U7230 ( .A(n5730), .B(n5729), .ZN(n7705) );
  NAND2_X1 U7231 ( .A1(n5734), .A2(n5735), .ZN(n5732) );
  NAND2_X1 U7232 ( .A1(n6376), .A2(n5997), .ZN(n5742) );
  NAND2_X1 U7233 ( .A1(n5418), .A2(SI_0_), .ZN(n5736) );
  XNOR2_X1 U7234 ( .A(n5736), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9539) );
  XNOR2_X2 U7235 ( .A(n5737), .B(n5710), .ZN(n9886) );
  AND2_X1 U7236 ( .A1(n5738), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5739) );
  INV_X1 U7237 ( .A(n7071), .ZN(n6361) );
  INV_X1 U7238 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7239 ( .A1(n5744), .A2(n5743), .ZN(n5745) );
  INV_X1 U7240 ( .A(n5747), .ZN(n5748) );
  NAND2_X1 U7241 ( .A1(n5748), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7242 ( .A1(n5753), .A2(n8070), .ZN(n6412) );
  NAND2_X1 U7243 ( .A1(n5752), .A2(n5751), .ZN(n5757) );
  NAND2_X1 U7244 ( .A1(n6349), .A2(n8121), .ZN(n6413) );
  NAND2_X1 U7245 ( .A1(n6376), .A2(n5772), .ZN(n5756) );
  INV_X1 U7246 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9862) );
  NOR2_X1 U7247 ( .A1(n6492), .A2(n9862), .ZN(n5754) );
  AOI21_X1 U7248 ( .B1(n6920), .B2(n5997), .A(n5754), .ZN(n5755) );
  INV_X1 U7249 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6534) );
  INV_X1 U7250 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U7251 ( .A1(n5878), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U7252 ( .A1(n5771), .A2(n5997), .ZN(n5769) );
  AND2_X2 U7253 ( .A1(n5814), .A2(n6495), .ZN(n5811) );
  NAND2_X1 U7254 ( .A1(n5811), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5767) );
  INV_X1 U7255 ( .A(n6512), .ZN(n5762) );
  NAND2_X1 U7256 ( .A1(n5812), .A2(n5762), .ZN(n5766) );
  NAND2_X1 U7257 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5763) );
  INV_X1 U7258 ( .A(n6546), .ZN(n5764) );
  NAND2_X1 U7259 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  XNOR2_X1 U7260 ( .A(n5770), .B(n7030), .ZN(n5778) );
  NAND2_X1 U7261 ( .A1(n5771), .A2(n5772), .ZN(n5776) );
  OR2_X1 U7262 ( .A1(n8079), .A2(n5825), .ZN(n5775) );
  NAND2_X1 U7263 ( .A1(n5776), .A2(n5775), .ZN(n6629) );
  NAND2_X1 U7264 ( .A1(n5777), .A2(n6629), .ZN(n5781) );
  INV_X1 U7265 ( .A(n6627), .ZN(n5779) );
  INV_X1 U7266 ( .A(n5778), .ZN(n6631) );
  NAND2_X1 U7267 ( .A1(n5779), .A2(n6631), .ZN(n5780) );
  AND2_X2 U7268 ( .A1(n5781), .A2(n5780), .ZN(n9058) );
  NAND2_X1 U7269 ( .A1(n5811), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5786) );
  INV_X1 U7270 ( .A(n6514), .ZN(n5782) );
  NAND2_X1 U7271 ( .A1(n5812), .A2(n5782), .ZN(n5785) );
  INV_X1 U7272 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U7273 ( .A1(n6157), .A2(n6548), .ZN(n5784) );
  INV_X1 U7274 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6533) );
  INV_X1 U7275 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7276 ( .A1(n5719), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5789) );
  INV_X2 U7277 ( .A(n5825), .ZN(n6307) );
  NAND2_X1 U7278 ( .A1(n5795), .A2(n6307), .ZN(n5792) );
  CLKBUF_X2 U7279 ( .A(n5795), .Z(n9127) );
  OR2_X1 U7280 ( .A1(n6839), .A2(n5825), .ZN(n5796) );
  NAND2_X1 U7281 ( .A1(n5798), .A2(n5797), .ZN(n5802) );
  NAND2_X1 U7282 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  AND2_X1 U7283 ( .A1(n5802), .A2(n5801), .ZN(n9059) );
  NAND2_X1 U7284 ( .A1(n6198), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7285 ( .A1(n5804), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5809) );
  INV_X1 U7286 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6532) );
  OR2_X1 U7287 ( .A1(n5805), .A2(n6532), .ZN(n5808) );
  INV_X1 U7288 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5806) );
  OR2_X1 U7289 ( .A1(n6080), .A2(n5806), .ZN(n5807) );
  NAND4_X2 U7290 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n9126)
         );
  NAND2_X1 U7291 ( .A1(n9126), .A2(n6307), .ZN(n5823) );
  NAND2_X1 U7292 ( .A1(n5811), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5821) );
  INV_X1 U7293 ( .A(n6516), .ZN(n5813) );
  NAND2_X1 U7294 ( .A1(n5812), .A2(n5813), .ZN(n5820) );
  INV_X1 U7295 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U7296 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  NAND2_X1 U7297 ( .A1(n5817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5818) );
  XNOR2_X1 U7298 ( .A(n5818), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U7299 ( .A1(n6157), .A2(n6549), .ZN(n5819) );
  OR2_X1 U7300 ( .A1(n9969), .A2(n5935), .ZN(n5822) );
  NAND2_X1 U7301 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  INV_X2 U7302 ( .A(n5773), .ZN(n6306) );
  NAND2_X1 U7303 ( .A1(n9126), .A2(n6306), .ZN(n5827) );
  OR2_X1 U7304 ( .A1(n9969), .A2(n6326), .ZN(n5826) );
  AND2_X1 U7305 ( .A1(n5827), .A2(n5826), .ZN(n5829) );
  NAND2_X1 U7306 ( .A1(n5828), .A2(n5829), .ZN(n6668) );
  INV_X1 U7307 ( .A(n5828), .ZN(n5831) );
  INV_X1 U7308 ( .A(n5829), .ZN(n5830) );
  NAND2_X1 U7309 ( .A1(n5831), .A2(n5830), .ZN(n6667) );
  NAND2_X1 U7310 ( .A1(n6198), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5837) );
  INV_X1 U7311 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5832) );
  OR2_X1 U7312 ( .A1(n5805), .A2(n5832), .ZN(n5836) );
  XNOR2_X1 U7313 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6725) );
  OR2_X1 U7314 ( .A1(n5804), .A2(n6725), .ZN(n5835) );
  INV_X1 U7315 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5833) );
  OR2_X1 U7316 ( .A1(n6080), .A2(n5833), .ZN(n5834) );
  NAND2_X1 U7317 ( .A1(n9125), .A2(n5997), .ZN(n5845) );
  NAND2_X1 U7318 ( .A1(n5811), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5843) );
  INV_X1 U7319 ( .A(n6501), .ZN(n5838) );
  NAND2_X1 U7320 ( .A1(n7936), .A2(n5838), .ZN(n5842) );
  NAND2_X1 U7321 ( .A1(n5839), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5840) );
  XNOR2_X1 U7322 ( .A(n5840), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7323 ( .A1(n6157), .A2(n6550), .ZN(n5841) );
  OR2_X1 U7324 ( .A1(n7089), .A2(n5935), .ZN(n5844) );
  NAND2_X1 U7325 ( .A1(n5845), .A2(n5844), .ZN(n5846) );
  NAND2_X1 U7326 ( .A1(n9125), .A2(n6306), .ZN(n5848) );
  OR2_X1 U7327 ( .A1(n7089), .A2(n6326), .ZN(n5847) );
  NAND2_X1 U7328 ( .A1(n5848), .A2(n5847), .ZN(n5850) );
  XNOR2_X1 U7329 ( .A(n5849), .B(n5850), .ZN(n6724) );
  INV_X1 U7330 ( .A(n5849), .ZN(n5851) );
  NAND2_X1 U7331 ( .A1(n5851), .A2(n5850), .ZN(n6768) );
  NAND2_X1 U7332 ( .A1(n6198), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5859) );
  INV_X1 U7333 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6536) );
  OR2_X1 U7334 ( .A1(n5805), .A2(n6536), .ZN(n5858) );
  NAND3_X1 U7335 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5880) );
  INV_X1 U7336 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5853) );
  NAND2_X1 U7337 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5852) );
  NAND2_X1 U7338 ( .A1(n5853), .A2(n5852), .ZN(n5854) );
  NAND2_X1 U7339 ( .A1(n5880), .A2(n5854), .ZN(n7228) );
  OR2_X1 U7340 ( .A1(n5804), .A2(n7228), .ZN(n5857) );
  INV_X1 U7341 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7342 ( .A1(n6080), .A2(n5855), .ZN(n5856) );
  NAND4_X1 U7343 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n9124)
         );
  NAND2_X1 U7344 ( .A1(n9124), .A2(n5997), .ZN(n5868) );
  INV_X1 U7345 ( .A(n6505), .ZN(n5860) );
  NAND2_X1 U7346 ( .A1(n5811), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U7347 ( .A1(n5861), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5862) );
  MUX2_X1 U7348 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5862), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5865) );
  INV_X1 U7349 ( .A(n5863), .ZN(n5864) );
  NAND2_X1 U7350 ( .A1(n6157), .A2(n9918), .ZN(n5866) );
  XNOR2_X1 U7351 ( .A(n5869), .B(n5751), .ZN(n6771) );
  NAND2_X1 U7352 ( .A1(n9124), .A2(n6306), .ZN(n5871) );
  OR2_X1 U7353 ( .A1(n9976), .A2(n6326), .ZN(n5870) );
  NAND2_X1 U7354 ( .A1(n5871), .A2(n5870), .ZN(n5874) );
  NAND2_X1 U7355 ( .A1(n6771), .A2(n5874), .ZN(n5872) );
  AND2_X1 U7356 ( .A1(n6768), .A2(n5872), .ZN(n5873) );
  NAND2_X1 U7357 ( .A1(n6722), .A2(n5873), .ZN(n5877) );
  INV_X1 U7358 ( .A(n6771), .ZN(n5875) );
  INV_X1 U7359 ( .A(n5874), .ZN(n6770) );
  NAND2_X1 U7360 ( .A1(n5875), .A2(n6770), .ZN(n5876) );
  NAND2_X1 U7361 ( .A1(n5878), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5886) );
  INV_X1 U7362 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6537) );
  OR2_X1 U7363 ( .A1(n5805), .A2(n6537), .ZN(n5885) );
  INV_X1 U7364 ( .A(n5880), .ZN(n5879) );
  NAND2_X1 U7365 ( .A1(n5879), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5907) );
  INV_X1 U7366 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6850) );
  NAND2_X1 U7367 ( .A1(n5880), .A2(n6850), .ZN(n5881) );
  NAND2_X1 U7368 ( .A1(n5907), .A2(n5881), .ZN(n9411) );
  OR2_X1 U7369 ( .A1(n5804), .A2(n9411), .ZN(n5884) );
  INV_X1 U7370 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5882) );
  OR2_X1 U7371 ( .A1(n6639), .A2(n5882), .ZN(n5883) );
  NAND4_X1 U7372 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n9123)
         );
  NAND2_X1 U7373 ( .A1(n9123), .A2(n6306), .ZN(n5893) );
  INV_X1 U7374 ( .A(n6503), .ZN(n5887) );
  NAND2_X1 U7375 ( .A1(n7936), .A2(n5887), .ZN(n5891) );
  NAND2_X1 U7376 ( .A1(n6456), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5890) );
  OR2_X1 U7377 ( .A1(n5863), .A2(n5899), .ZN(n5888) );
  XNOR2_X1 U7378 ( .A(n5888), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9129) );
  NAND2_X1 U7379 ( .A1(n6157), .A2(n9129), .ZN(n5889) );
  OR2_X1 U7380 ( .A1(n7008), .A2(n6326), .ZN(n5892) );
  AND2_X1 U7381 ( .A1(n5893), .A2(n5892), .ZN(n6848) );
  NAND2_X1 U7382 ( .A1(n9123), .A2(n5997), .ZN(n5895) );
  OR2_X1 U7383 ( .A1(n7008), .A2(n5935), .ZN(n5894) );
  NAND2_X1 U7384 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  XNOR2_X1 U7385 ( .A(n5896), .B(n5751), .ZN(n6847) );
  INV_X1 U7386 ( .A(n6848), .ZN(n5897) );
  NAND2_X1 U7387 ( .A1(n6456), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5904) );
  OR2_X1 U7388 ( .A1(n6047), .A2(n6518), .ZN(n5903) );
  AND2_X1 U7389 ( .A1(n5863), .A2(n5898), .ZN(n5900) );
  OR2_X1 U7390 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  XNOR2_X1 U7391 ( .A(n5901), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U7392 ( .A1(n6157), .A2(n6572), .ZN(n5902) );
  INV_X1 U7393 ( .A(n7352), .ZN(n7037) );
  NAND2_X1 U7394 ( .A1(n7037), .A2(n4508), .ZN(n5915) );
  NAND2_X1 U7395 ( .A1(n6198), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5913) );
  INV_X1 U7396 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7040) );
  OR2_X1 U7397 ( .A1(n5805), .A2(n7040), .ZN(n5912) );
  INV_X1 U7398 ( .A(n5907), .ZN(n5905) );
  NAND2_X1 U7399 ( .A1(n5905), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5922) );
  INV_X1 U7400 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7401 ( .A1(n5907), .A2(n5906), .ZN(n5908) );
  NAND2_X1 U7402 ( .A1(n5922), .A2(n5908), .ZN(n7039) );
  OR2_X1 U7403 ( .A1(n5804), .A2(n7039), .ZN(n5911) );
  INV_X1 U7404 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5909) );
  OR2_X1 U7405 ( .A1(n6080), .A2(n5909), .ZN(n5910) );
  NAND4_X1 U7406 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n9122)
         );
  NAND2_X1 U7407 ( .A1(n9122), .A2(n5997), .ZN(n5914) );
  NAND2_X1 U7408 ( .A1(n5915), .A2(n5914), .ZN(n5916) );
  XNOR2_X1 U7409 ( .A(n5916), .B(n5751), .ZN(n5919) );
  NAND2_X1 U7410 ( .A1(n9122), .A2(n5772), .ZN(n5917) );
  OAI21_X1 U7411 ( .B1(n7352), .B2(n6326), .A(n5917), .ZN(n5918) );
  OR2_X1 U7412 ( .A1(n5919), .A2(n5918), .ZN(n6955) );
  NAND2_X1 U7413 ( .A1(n6953), .A2(n6955), .ZN(n5920) );
  NAND2_X1 U7414 ( .A1(n5919), .A2(n5918), .ZN(n6954) );
  NAND2_X1 U7415 ( .A1(n6198), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5927) );
  INV_X1 U7416 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7240) );
  OR2_X1 U7417 ( .A1(n5805), .A2(n7240), .ZN(n5926) );
  INV_X1 U7418 ( .A(n5922), .ZN(n5921) );
  INV_X1 U7419 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U7420 ( .A1(n5922), .A2(n6568), .ZN(n5923) );
  NAND2_X1 U7421 ( .A1(n5949), .A2(n5923), .ZN(n7267) );
  OR2_X1 U7422 ( .A1(n5804), .A2(n7267), .ZN(n5925) );
  INV_X1 U7423 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6573) );
  OR2_X1 U7424 ( .A1(n6080), .A2(n6573), .ZN(n5924) );
  NAND4_X1 U7425 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n9121)
         );
  NAND2_X1 U7426 ( .A1(n9121), .A2(n6306), .ZN(n5933) );
  NAND2_X1 U7427 ( .A1(n6524), .A2(n7936), .ZN(n5931) );
  NAND2_X1 U7428 ( .A1(n5928), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5929) );
  XNOR2_X1 U7429 ( .A(n5929), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6593) );
  AOI22_X1 U7430 ( .A1(n6456), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6157), .B2(
        n6593), .ZN(n5930) );
  OR2_X1 U7431 ( .A1(n7308), .A2(n6326), .ZN(n5932) );
  NAND2_X1 U7432 ( .A1(n5933), .A2(n5932), .ZN(n5938) );
  NAND2_X1 U7433 ( .A1(n5937), .A2(n5938), .ZN(n7261) );
  NAND2_X1 U7434 ( .A1(n9121), .A2(n5997), .ZN(n5934) );
  OAI21_X1 U7435 ( .B1(n7308), .B2(n5935), .A(n5934), .ZN(n5936) );
  NAND2_X1 U7436 ( .A1(n7261), .A2(n7264), .ZN(n5941) );
  INV_X1 U7437 ( .A(n5937), .ZN(n5940) );
  NAND2_X1 U7438 ( .A1(n5940), .A2(n5939), .ZN(n7263) );
  NAND2_X1 U7439 ( .A1(n5941), .A2(n7263), .ZN(n7363) );
  NAND2_X1 U7440 ( .A1(n6528), .A2(n7936), .ZN(n5947) );
  NAND2_X1 U7441 ( .A1(n5942), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5943) );
  MUX2_X1 U7442 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5943), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5945) );
  AND2_X1 U7443 ( .A1(n5945), .A2(n5984), .ZN(n6597) );
  AOI22_X1 U7444 ( .A1(n5811), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6157), .B2(
        n6597), .ZN(n5946) );
  NAND2_X1 U7445 ( .A1(n5947), .A2(n5946), .ZN(n7320) );
  NAND2_X1 U7446 ( .A1(n7320), .A2(n4508), .ZN(n5958) );
  NAND2_X1 U7447 ( .A1(n6462), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5956) );
  NAND2_X1 U7448 ( .A1(n5949), .A2(n5948), .ZN(n5950) );
  NAND2_X1 U7449 ( .A1(n5968), .A2(n5950), .ZN(n7368) );
  OR2_X1 U7450 ( .A1(n5804), .A2(n7368), .ZN(n5955) );
  INV_X1 U7451 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5951) );
  OR2_X1 U7452 ( .A1(n6080), .A2(n5951), .ZN(n5954) );
  INV_X1 U7453 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5952) );
  OR2_X1 U7454 ( .A1(n6639), .A2(n5952), .ZN(n5953) );
  NAND4_X1 U7455 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n9120)
         );
  NAND2_X1 U7456 ( .A1(n9120), .A2(n5997), .ZN(n5957) );
  NAND2_X1 U7457 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7458 ( .A(n5959), .B(n5751), .ZN(n5960) );
  AOI22_X1 U7459 ( .A1(n7320), .A2(n6307), .B1(n6306), .B2(n9120), .ZN(n5961)
         );
  XNOR2_X1 U7460 ( .A(n5960), .B(n5961), .ZN(n7365) );
  NAND2_X1 U7461 ( .A1(n7363), .A2(n7365), .ZN(n5964) );
  INV_X1 U7462 ( .A(n5960), .ZN(n5962) );
  NAND2_X1 U7463 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U7464 ( .A1(n5964), .A2(n5963), .ZN(n7406) );
  NAND2_X1 U7465 ( .A1(n6560), .A2(n7936), .ZN(n5967) );
  NAND2_X1 U7466 ( .A1(n5984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7467 ( .A(n5965), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6651) );
  AOI22_X1 U7468 ( .A1(n5811), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6157), .B2(
        n6651), .ZN(n5966) );
  NAND2_X1 U7469 ( .A1(n5967), .A2(n5966), .ZN(n7398) );
  NAND2_X1 U7470 ( .A1(n7398), .A2(n4508), .ZN(n5976) );
  NAND2_X1 U7471 ( .A1(n6198), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5974) );
  INV_X1 U7472 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7393) );
  OR2_X1 U7473 ( .A1(n5805), .A2(n7393), .ZN(n5973) );
  NAND2_X1 U7474 ( .A1(n5968), .A2(n6592), .ZN(n5969) );
  NAND2_X1 U7475 ( .A1(n5991), .A2(n5969), .ZN(n7408) );
  OR2_X1 U7476 ( .A1(n5804), .A2(n7408), .ZN(n5972) );
  INV_X1 U7477 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7478 ( .A1(n6080), .A2(n5970), .ZN(n5971) );
  OR2_X1 U7479 ( .A1(n7442), .A2(n6326), .ZN(n5975) );
  NAND2_X1 U7480 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  XNOR2_X1 U7481 ( .A(n5977), .B(n7030), .ZN(n7404) );
  NAND2_X1 U7482 ( .A1(n7398), .A2(n6307), .ZN(n5979) );
  OR2_X1 U7483 ( .A1(n7442), .A2(n5773), .ZN(n5978) );
  AND2_X1 U7484 ( .A1(n5979), .A2(n5978), .ZN(n5980) );
  AND2_X1 U7485 ( .A1(n7404), .A2(n5980), .ZN(n5983) );
  INV_X1 U7486 ( .A(n7404), .ZN(n5981) );
  INV_X1 U7487 ( .A(n5980), .ZN(n7403) );
  NAND2_X1 U7488 ( .A1(n5981), .A2(n7403), .ZN(n5982) );
  OAI21_X2 U7489 ( .B1(n7406), .B2(n5983), .A(n5982), .ZN(n7435) );
  NAND2_X1 U7490 ( .A1(n6580), .A2(n7936), .ZN(n5987) );
  NOR2_X1 U7491 ( .A1(n5984), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6006) );
  OR2_X1 U7492 ( .A1(n6006), .A2(n5899), .ZN(n5985) );
  XNOR2_X1 U7493 ( .A(n5985), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U7494 ( .A1(n5811), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6157), .B2(
        n6652), .ZN(n5986) );
  NAND2_X1 U7495 ( .A1(n9844), .A2(n4508), .ZN(n5999) );
  NAND2_X1 U7496 ( .A1(n6198), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5996) );
  INV_X1 U7497 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7451) );
  OR2_X1 U7498 ( .A1(n5805), .A2(n7451), .ZN(n5995) );
  INV_X1 U7499 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7500 ( .A1(n6080), .A2(n5988), .ZN(n5994) );
  INV_X1 U7501 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5990) );
  NAND2_X1 U7502 ( .A1(n5991), .A2(n5990), .ZN(n5992) );
  NAND2_X1 U7503 ( .A1(n6012), .A2(n5992), .ZN(n7450) );
  OR2_X1 U7504 ( .A1(n5804), .A2(n7450), .ZN(n5993) );
  NAND4_X1 U7505 ( .A1(n5996), .A2(n5995), .A3(n5994), .A4(n5993), .ZN(n9118)
         );
  NAND2_X1 U7506 ( .A1(n9118), .A2(n5997), .ZN(n5998) );
  NAND2_X1 U7507 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  XNOR2_X1 U7508 ( .A(n6000), .B(n5751), .ZN(n6004) );
  AND2_X1 U7509 ( .A1(n9118), .A2(n6306), .ZN(n6001) );
  AOI21_X1 U7510 ( .B1(n9844), .B2(n6307), .A(n6001), .ZN(n6002) );
  XNOR2_X1 U7511 ( .A(n6004), .B(n6002), .ZN(n7434) );
  INV_X1 U7512 ( .A(n6002), .ZN(n6003) );
  NAND2_X1 U7513 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  NAND2_X1 U7514 ( .A1(n6607), .A2(n7936), .ZN(n6009) );
  NAND2_X1 U7515 ( .A1(n6006), .A2(n4746), .ZN(n6028) );
  NAND2_X1 U7516 ( .A1(n6028), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7517 ( .A(n6007), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6697) );
  AOI22_X1 U7518 ( .A1(n5811), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6157), .B2(
        n6697), .ZN(n6008) );
  NAND2_X1 U7519 ( .A1(n7646), .A2(n4508), .ZN(n6020) );
  NAND2_X1 U7520 ( .A1(n6462), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6018) );
  INV_X1 U7521 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6644) );
  OR2_X1 U7522 ( .A1(n6080), .A2(n6644), .ZN(n6017) );
  INV_X1 U7523 ( .A(n6012), .ZN(n6010) );
  INV_X1 U7524 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7525 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7526 ( .A1(n6033), .A2(n6013), .ZN(n7643) );
  OR2_X1 U7527 ( .A1(n5804), .A2(n7643), .ZN(n6016) );
  INV_X1 U7528 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n6014) );
  OR2_X1 U7529 ( .A1(n6639), .A2(n6014), .ZN(n6015) );
  OR2_X1 U7530 ( .A1(n7757), .A2(n6326), .ZN(n6019) );
  NAND2_X1 U7531 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  XNOR2_X1 U7532 ( .A(n6021), .B(n7030), .ZN(n6024) );
  NOR2_X1 U7533 ( .A1(n7757), .A2(n5773), .ZN(n6022) );
  AOI21_X1 U7534 ( .B1(n7646), .B2(n5997), .A(n6022), .ZN(n6023) );
  NAND2_X1 U7535 ( .A1(n6024), .A2(n6023), .ZN(n6027) );
  OR2_X1 U7536 ( .A1(n6024), .A2(n6023), .ZN(n6025) );
  NAND2_X1 U7537 ( .A1(n6027), .A2(n6025), .ZN(n7640) );
  NAND2_X1 U7538 ( .A1(n7636), .A2(n6027), .ZN(n7675) );
  NAND2_X1 U7539 ( .A1(n6620), .A2(n7936), .ZN(n6031) );
  NAND2_X1 U7540 ( .A1(n6048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7541 ( .A(n6029), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6969) );
  AOI22_X1 U7542 ( .A1(n5811), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6157), .B2(
        n6969), .ZN(n6030) );
  NAND2_X1 U7543 ( .A1(n9830), .A2(n4508), .ZN(n6040) );
  NAND2_X1 U7544 ( .A1(n6198), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6038) );
  INV_X1 U7545 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9822) );
  OR2_X1 U7546 ( .A1(n5805), .A2(n9822), .ZN(n6037) );
  NAND2_X1 U7547 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7548 ( .A1(n6057), .A2(n6034), .ZN(n9821) );
  OR2_X1 U7549 ( .A1(n5804), .A2(n9821), .ZN(n6036) );
  INV_X1 U7550 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6692) );
  OR2_X1 U7551 ( .A1(n6080), .A2(n6692), .ZN(n6035) );
  NAND4_X1 U7552 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n9116)
         );
  NAND2_X1 U7553 ( .A1(n9116), .A2(n6307), .ZN(n6039) );
  NAND2_X1 U7554 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  XNOR2_X1 U7555 ( .A(n6041), .B(n7030), .ZN(n6043) );
  AND2_X1 U7556 ( .A1(n9116), .A2(n6306), .ZN(n6042) );
  AOI21_X1 U7557 ( .B1(n9830), .B2(n6307), .A(n6042), .ZN(n6044) );
  AND2_X1 U7558 ( .A1(n6043), .A2(n6044), .ZN(n7673) );
  INV_X1 U7559 ( .A(n6043), .ZN(n6046) );
  INV_X1 U7560 ( .A(n6044), .ZN(n6045) );
  INV_X4 U7561 ( .A(n6047), .ZN(n7936) );
  NAND2_X1 U7562 ( .A1(n6660), .A2(n7936), .ZN(n6054) );
  INV_X1 U7563 ( .A(n6051), .ZN(n6049) );
  NAND2_X1 U7564 ( .A1(n6049), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6052) );
  INV_X1 U7565 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7566 ( .A1(n6051), .A2(n6050), .ZN(n6069) );
  AOI22_X1 U7567 ( .A1(n6456), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7380), .B2(
        n6157), .ZN(n6053) );
  NAND2_X1 U7568 ( .A1(n7797), .A2(n4508), .ZN(n6064) );
  NAND2_X1 U7569 ( .A1(n6198), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6062) );
  INV_X1 U7570 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7728) );
  OR2_X1 U7571 ( .A1(n5805), .A2(n7728), .ZN(n6061) );
  INV_X1 U7572 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7573 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  NAND2_X1 U7574 ( .A1(n6077), .A2(n6058), .ZN(n7794) );
  OR2_X1 U7575 ( .A1(n5804), .A2(n7794), .ZN(n6060) );
  INV_X1 U7576 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6964) );
  OR2_X1 U7577 ( .A1(n6080), .A2(n6964), .ZN(n6059) );
  NAND4_X1 U7578 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n9115)
         );
  NAND2_X1 U7579 ( .A1(n9115), .A2(n6307), .ZN(n6063) );
  NAND2_X1 U7580 ( .A1(n6064), .A2(n6063), .ZN(n6065) );
  XNOR2_X1 U7581 ( .A(n6065), .B(n5751), .ZN(n6068) );
  NAND2_X1 U7582 ( .A1(n7797), .A2(n6307), .ZN(n6067) );
  NAND2_X1 U7583 ( .A1(n9115), .A2(n6306), .ZN(n6066) );
  NAND2_X1 U7584 ( .A1(n6067), .A2(n6066), .ZN(n7793) );
  NAND2_X1 U7585 ( .A1(n6688), .A2(n7936), .ZN(n6075) );
  NAND2_X1 U7586 ( .A1(n6069), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6071) );
  INV_X1 U7587 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6070) );
  XNOR2_X1 U7588 ( .A(n6071), .B(n6070), .ZN(n7501) );
  OAI22_X1 U7589 ( .A1(n7501), .A2(n5814), .B1(n6072), .B2(n6689), .ZN(n6073)
         );
  INV_X1 U7590 ( .A(n6073), .ZN(n6074) );
  NAND2_X1 U7591 ( .A1(n9100), .A2(n4508), .ZN(n6086) );
  NAND2_X1 U7592 ( .A1(n6198), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6084) );
  INV_X1 U7593 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7738) );
  OR2_X1 U7594 ( .A1(n5805), .A2(n7738), .ZN(n6083) );
  INV_X1 U7595 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7596 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  NAND2_X1 U7597 ( .A1(n6098), .A2(n6078), .ZN(n9095) );
  OR2_X1 U7598 ( .A1(n5804), .A2(n9095), .ZN(n6082) );
  INV_X1 U7599 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7600 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  NAND4_X1 U7601 ( .A1(n6084), .A2(n6083), .A3(n6082), .A4(n6081), .ZN(n9114)
         );
  NAND2_X1 U7602 ( .A1(n9114), .A2(n6307), .ZN(n6085) );
  NAND2_X1 U7603 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  XNOR2_X1 U7604 ( .A(n6087), .B(n7030), .ZN(n6090) );
  NAND2_X1 U7605 ( .A1(n9100), .A2(n5997), .ZN(n6089) );
  NAND2_X1 U7606 ( .A1(n9114), .A2(n6306), .ZN(n6088) );
  NAND2_X1 U7607 ( .A1(n6089), .A2(n6088), .ZN(n9091) );
  INV_X1 U7608 ( .A(n6090), .ZN(n6091) );
  NAND2_X1 U7609 ( .A1(n6835), .A2(n7936), .ZN(n6096) );
  NOR2_X1 U7610 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n6092) );
  NAND2_X1 U7611 ( .A1(n6093), .A2(n6092), .ZN(n6112) );
  NAND2_X1 U7612 ( .A1(n6112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6094) );
  XNOR2_X1 U7613 ( .A(n6094), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9160) );
  AOI22_X1 U7614 ( .A1(n6456), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9160), .B2(
        n6157), .ZN(n6095) );
  NAND2_X1 U7615 ( .A1(n9017), .A2(n4508), .ZN(n6105) );
  NAND2_X1 U7616 ( .A1(n6198), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6103) );
  INV_X1 U7617 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7815) );
  OR2_X1 U7618 ( .A1(n5805), .A2(n7815), .ZN(n6102) );
  INV_X1 U7619 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9012) );
  NAND2_X1 U7620 ( .A1(n6098), .A2(n9012), .ZN(n6099) );
  NAND2_X1 U7621 ( .A1(n6121), .A2(n6099), .ZN(n9014) );
  OR2_X1 U7622 ( .A1(n5804), .A2(n9014), .ZN(n6101) );
  INV_X1 U7623 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7504) );
  OR2_X1 U7624 ( .A1(n6080), .A2(n7504), .ZN(n6100) );
  OR2_X1 U7625 ( .A1(n9402), .A2(n6326), .ZN(n6104) );
  NAND2_X1 U7626 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  XNOR2_X1 U7627 ( .A(n6106), .B(n7030), .ZN(n6110) );
  NOR2_X1 U7628 ( .A1(n9402), .A2(n5773), .ZN(n6107) );
  AOI21_X1 U7629 ( .B1(n9017), .B2(n6307), .A(n6107), .ZN(n6109) );
  XNOR2_X1 U7630 ( .A(n6110), .B(n6109), .ZN(n9011) );
  INV_X1 U7631 ( .A(n9011), .ZN(n6108) );
  NAND2_X1 U7632 ( .A1(n6110), .A2(n6109), .ZN(n6111) );
  NAND2_X1 U7633 ( .A1(n9009), .A2(n6111), .ZN(n9021) );
  NAND2_X1 U7634 ( .A1(n6778), .A2(n7936), .ZN(n6119) );
  NAND2_X1 U7635 ( .A1(n6113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6116) );
  INV_X1 U7636 ( .A(n6116), .ZN(n6114) );
  NAND2_X1 U7637 ( .A1(n6114), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n6117) );
  INV_X1 U7638 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6115) );
  NAND2_X1 U7639 ( .A1(n6116), .A2(n6115), .ZN(n6135) );
  AOI22_X1 U7640 ( .A1(n9175), .A2(n6157), .B1(n6456), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7641 ( .A1(n9483), .A2(n4508), .ZN(n6128) );
  NAND2_X1 U7642 ( .A1(n6198), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6126) );
  INV_X1 U7643 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9156) );
  OR2_X1 U7644 ( .A1(n5805), .A2(n9156), .ZN(n6125) );
  INV_X1 U7645 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6120) );
  OR2_X1 U7646 ( .A1(n6080), .A2(n6120), .ZN(n6124) );
  INV_X1 U7647 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9024) );
  NAND2_X1 U7648 ( .A1(n6121), .A2(n9024), .ZN(n6122) );
  NAND2_X1 U7649 ( .A1(n6141), .A2(n6122), .ZN(n9394) );
  OR2_X1 U7650 ( .A1(n5804), .A2(n9394), .ZN(n6123) );
  NAND4_X1 U7651 ( .A1(n6126), .A2(n6125), .A3(n6124), .A4(n6123), .ZN(n9112)
         );
  NAND2_X1 U7652 ( .A1(n9112), .A2(n6307), .ZN(n6127) );
  NAND2_X1 U7653 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  XNOR2_X1 U7654 ( .A(n6129), .B(n5751), .ZN(n6131) );
  AND2_X1 U7655 ( .A1(n9112), .A2(n6306), .ZN(n6130) );
  AOI21_X1 U7656 ( .B1(n9483), .B2(n6307), .A(n6130), .ZN(n6132) );
  XNOR2_X1 U7657 ( .A(n6131), .B(n6132), .ZN(n9022) );
  INV_X1 U7658 ( .A(n6131), .ZN(n6133) );
  NAND2_X1 U7659 ( .A1(n6133), .A2(n6132), .ZN(n6134) );
  NAND2_X1 U7660 ( .A1(n9020), .A2(n6134), .ZN(n6152) );
  NAND2_X1 U7661 ( .A1(n6995), .A2(n7936), .ZN(n6138) );
  NAND2_X1 U7662 ( .A1(n6135), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6136) );
  XNOR2_X1 U7663 ( .A(n6136), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9950) );
  AOI22_X1 U7664 ( .A1(n9950), .A2(n6157), .B1(n6456), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7665 ( .A1(n9378), .A2(n4508), .ZN(n6148) );
  NAND2_X1 U7666 ( .A1(n6198), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6146) );
  INV_X1 U7667 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9380) );
  OR2_X1 U7668 ( .A1(n5805), .A2(n9380), .ZN(n6145) );
  INV_X1 U7669 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7670 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7671 ( .A1(n6162), .A2(n6142), .ZN(n9379) );
  OR2_X1 U7672 ( .A1(n5804), .A2(n9379), .ZN(n6144) );
  INV_X1 U7673 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9479) );
  OR2_X1 U7674 ( .A1(n6080), .A2(n9479), .ZN(n6143) );
  OR2_X1 U7675 ( .A1(n9404), .A2(n6326), .ZN(n6147) );
  NAND2_X1 U7676 ( .A1(n6148), .A2(n6147), .ZN(n6149) );
  XNOR2_X1 U7677 ( .A(n6149), .B(n7030), .ZN(n6153) );
  NAND2_X1 U7678 ( .A1(n6152), .A2(n6153), .ZN(n9066) );
  NAND2_X1 U7679 ( .A1(n9378), .A2(n6307), .ZN(n6151) );
  OR2_X1 U7680 ( .A1(n9404), .A2(n5773), .ZN(n6150) );
  NAND2_X1 U7681 ( .A1(n6151), .A2(n6150), .ZN(n9069) );
  NAND2_X1 U7682 ( .A1(n9066), .A2(n9069), .ZN(n6156) );
  INV_X1 U7683 ( .A(n6152), .ZN(n6155) );
  INV_X1 U7684 ( .A(n6153), .ZN(n6154) );
  NAND2_X1 U7685 ( .A1(n6155), .A2(n6154), .ZN(n9067) );
  NAND2_X1 U7686 ( .A1(n7176), .A2(n7936), .ZN(n6159) );
  AOI22_X1 U7687 ( .A1(n5811), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9184), .B2(
        n6157), .ZN(n6158) );
  NAND2_X1 U7688 ( .A1(n9473), .A2(n4508), .ZN(n6169) );
  NAND2_X1 U7689 ( .A1(n6198), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6167) );
  INV_X1 U7690 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7691 ( .A1(n6162), .A2(n6161), .ZN(n6163) );
  NAND2_X1 U7692 ( .A1(n6177), .A2(n6163), .ZN(n9358) );
  OR2_X1 U7693 ( .A1(n9358), .A2(n5804), .ZN(n6166) );
  INV_X1 U7694 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9359) );
  OR2_X1 U7695 ( .A1(n5805), .A2(n9359), .ZN(n6165) );
  INV_X1 U7696 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9176) );
  OR2_X1 U7697 ( .A1(n6080), .A2(n9176), .ZN(n6164) );
  NAND4_X1 U7698 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n9347)
         );
  NAND2_X1 U7699 ( .A1(n9347), .A2(n5997), .ZN(n6168) );
  NAND2_X1 U7700 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  XNOR2_X1 U7701 ( .A(n6170), .B(n7030), .ZN(n6173) );
  AND2_X1 U7702 ( .A1(n9347), .A2(n6306), .ZN(n6171) );
  AOI21_X1 U7703 ( .B1(n9473), .B2(n5997), .A(n6171), .ZN(n6172) );
  XNOR2_X1 U7704 ( .A(n6173), .B(n6172), .ZN(n8986) );
  NAND2_X1 U7705 ( .A1(n6173), .A2(n6172), .ZN(n6174) );
  NAND2_X1 U7706 ( .A1(n7372), .A2(n7936), .ZN(n6176) );
  NAND2_X1 U7707 ( .A1(n6456), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7708 ( .A1(n9467), .A2(n4508), .ZN(n6186) );
  INV_X1 U7709 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9043) );
  NAND2_X1 U7710 ( .A1(n6177), .A2(n9043), .ZN(n6178) );
  NAND2_X1 U7711 ( .A1(n6196), .A2(n6178), .ZN(n9338) );
  NOR2_X1 U7712 ( .A1(n9338), .A2(n5804), .ZN(n6184) );
  INV_X1 U7713 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7714 ( .A1(n6462), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6179) );
  OAI21_X1 U7715 ( .B1(n6639), .B2(n6180), .A(n6179), .ZN(n6183) );
  INV_X1 U7716 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n6181) );
  NOR2_X1 U7717 ( .A1(n6080), .A2(n6181), .ZN(n6182) );
  NAND2_X1 U7718 ( .A1(n9321), .A2(n5997), .ZN(n6185) );
  NAND2_X1 U7719 ( .A1(n6186), .A2(n6185), .ZN(n6187) );
  XNOR2_X1 U7720 ( .A(n6187), .B(n5751), .ZN(n6190) );
  NAND2_X1 U7721 ( .A1(n9467), .A2(n5997), .ZN(n6189) );
  NAND2_X1 U7722 ( .A1(n9321), .A2(n6306), .ZN(n6188) );
  NAND2_X1 U7723 ( .A1(n6189), .A2(n6188), .ZN(n6191) );
  NAND2_X1 U7724 ( .A1(n6190), .A2(n6191), .ZN(n9039) );
  INV_X1 U7725 ( .A(n6190), .ZN(n6193) );
  INV_X1 U7726 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7727 ( .A1(n6193), .A2(n6192), .ZN(n9040) );
  NAND2_X1 U7728 ( .A1(n7386), .A2(n7936), .ZN(n6195) );
  NAND2_X1 U7729 ( .A1(n6456), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7730 ( .A1(n9328), .A2(n4508), .ZN(n6203) );
  INV_X1 U7731 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8994) );
  NAND2_X1 U7732 ( .A1(n6196), .A2(n8994), .ZN(n6197) );
  AND2_X1 U7733 ( .A1(n6214), .A2(n6197), .ZN(n9329) );
  NAND2_X1 U7734 ( .A1(n9329), .A2(n6299), .ZN(n6201) );
  AOI22_X1 U7735 ( .A1(n6462), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n5878), .B2(
        P1_REG1_REG_21__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7736 ( .A1(n6198), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6199) );
  INV_X1 U7737 ( .A(n9306), .ZN(n9349) );
  NAND2_X1 U7738 ( .A1(n9349), .A2(n6307), .ZN(n6202) );
  NAND2_X1 U7739 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  XNOR2_X1 U7740 ( .A(n6204), .B(n5751), .ZN(n6206) );
  NOR2_X1 U7741 ( .A1(n9306), .A2(n5773), .ZN(n6205) );
  AOI21_X1 U7742 ( .B1(n9328), .B2(n5997), .A(n6205), .ZN(n6207) );
  XNOR2_X1 U7743 ( .A(n6206), .B(n6207), .ZN(n8993) );
  NAND2_X1 U7744 ( .A1(n8991), .A2(n8993), .ZN(n6210) );
  INV_X1 U7745 ( .A(n6206), .ZN(n6208) );
  NAND2_X1 U7746 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7747 ( .A1(n7492), .A2(n7936), .ZN(n6212) );
  NAND2_X1 U7748 ( .A1(n6456), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6211) );
  INV_X1 U7749 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U7750 ( .A1(n6214), .A2(n9052), .ZN(n6215) );
  NAND2_X1 U7751 ( .A1(n6230), .A2(n6215), .ZN(n9310) );
  OR2_X1 U7752 ( .A1(n9310), .A2(n5804), .ZN(n6221) );
  INV_X1 U7753 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n6218) );
  NAND2_X1 U7754 ( .A1(n6462), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7755 ( .A1(n5878), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6216) );
  OAI211_X1 U7756 ( .C1(n6639), .C2(n6218), .A(n6217), .B(n6216), .ZN(n6219)
         );
  INV_X1 U7757 ( .A(n6219), .ZN(n6220) );
  NAND2_X1 U7758 ( .A1(n6221), .A2(n6220), .ZN(n9322) );
  AND2_X1 U7759 ( .A1(n9322), .A2(n6306), .ZN(n6222) );
  AOI21_X1 U7760 ( .B1(n9458), .B2(n6307), .A(n6222), .ZN(n6226) );
  NAND2_X1 U7761 ( .A1(n9458), .A2(n4508), .ZN(n6224) );
  NAND2_X1 U7762 ( .A1(n9322), .A2(n5997), .ZN(n6223) );
  NAND2_X1 U7763 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  XNOR2_X1 U7764 ( .A(n6225), .B(n7030), .ZN(n9050) );
  NAND2_X1 U7765 ( .A1(n7632), .A2(n7936), .ZN(n6228) );
  NAND2_X1 U7766 ( .A1(n6456), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7767 ( .A1(n9453), .A2(n4508), .ZN(n6239) );
  INV_X1 U7768 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8980) );
  NAND2_X1 U7769 ( .A1(n6230), .A2(n8980), .ZN(n6231) );
  NAND2_X1 U7770 ( .A1(n6245), .A2(n6231), .ZN(n9296) );
  OR2_X1 U7771 ( .A1(n9296), .A2(n5804), .ZN(n6237) );
  INV_X1 U7772 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6234) );
  NAND2_X1 U7773 ( .A1(n5878), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U7774 ( .A1(n6462), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6232) );
  OAI211_X1 U7775 ( .C1(n6639), .C2(n6234), .A(n6233), .B(n6232), .ZN(n6235)
         );
  INV_X1 U7776 ( .A(n6235), .ZN(n6236) );
  NAND2_X1 U7777 ( .A1(n6237), .A2(n6236), .ZN(n9110) );
  NAND2_X1 U7778 ( .A1(n9110), .A2(n5997), .ZN(n6238) );
  NAND2_X1 U7779 ( .A1(n6239), .A2(n6238), .ZN(n6240) );
  AND2_X1 U7780 ( .A1(n9110), .A2(n6306), .ZN(n6241) );
  AOI21_X1 U7781 ( .B1(n9453), .B2(n5997), .A(n6241), .ZN(n8976) );
  NAND2_X1 U7782 ( .A1(n8977), .A2(n8976), .ZN(n9031) );
  NAND2_X2 U7783 ( .A1(n6242), .A2(n4359), .ZN(n9030) );
  NAND2_X1 U7784 ( .A1(n7700), .A2(n7936), .ZN(n6244) );
  NAND2_X1 U7785 ( .A1(n6456), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7786 ( .A1(n9282), .A2(n4508), .ZN(n6253) );
  INV_X1 U7787 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9034) );
  NAND2_X1 U7788 ( .A1(n6245), .A2(n9034), .ZN(n6246) );
  AND2_X1 U7789 ( .A1(n6267), .A2(n6246), .ZN(n9283) );
  NAND2_X1 U7790 ( .A1(n9283), .A2(n6299), .ZN(n6251) );
  INV_X1 U7791 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9510) );
  NAND2_X1 U7792 ( .A1(n5878), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7793 ( .A1(n6462), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6247) );
  OAI211_X1 U7794 ( .C1(n6639), .C2(n9510), .A(n6248), .B(n6247), .ZN(n6249)
         );
  INV_X1 U7795 ( .A(n6249), .ZN(n6250) );
  NAND2_X1 U7796 ( .A1(n6251), .A2(n6250), .ZN(n9260) );
  NAND2_X1 U7797 ( .A1(n9260), .A2(n5997), .ZN(n6252) );
  NAND2_X1 U7798 ( .A1(n6253), .A2(n6252), .ZN(n6254) );
  XNOR2_X1 U7799 ( .A(n6254), .B(n7030), .ZN(n6256) );
  AND2_X1 U7800 ( .A1(n9260), .A2(n5772), .ZN(n6255) );
  AOI21_X1 U7801 ( .B1(n9282), .B2(n5997), .A(n6255), .ZN(n6257) );
  NAND2_X1 U7802 ( .A1(n6256), .A2(n6257), .ZN(n6261) );
  INV_X1 U7803 ( .A(n6256), .ZN(n6259) );
  INV_X1 U7804 ( .A(n6257), .ZN(n6258) );
  NAND2_X1 U7805 ( .A1(n6259), .A2(n6258), .ZN(n6260) );
  NAND2_X1 U7806 ( .A1(n6261), .A2(n6260), .ZN(n9029) );
  INV_X1 U7807 ( .A(n6261), .ZN(n6262) );
  NAND2_X1 U7808 ( .A1(n7745), .A2(n7936), .ZN(n6264) );
  NAND2_X1 U7809 ( .A1(n6456), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U7810 ( .A1(n9267), .A2(n4508), .ZN(n6275) );
  INV_X1 U7811 ( .A(n6267), .ZN(n6265) );
  INV_X1 U7812 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7813 ( .A1(n6267), .A2(n6266), .ZN(n6268) );
  NAND2_X1 U7814 ( .A1(n6282), .A2(n6268), .ZN(n9002) );
  OR2_X1 U7815 ( .A1(n9002), .A2(n5804), .ZN(n6273) );
  INV_X1 U7816 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9506) );
  NAND2_X1 U7817 ( .A1(n6462), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7818 ( .A1(n5878), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7819 ( .C1(n6639), .C2(n9506), .A(n6270), .B(n6269), .ZN(n6271)
         );
  INV_X1 U7820 ( .A(n6271), .ZN(n6272) );
  INV_X1 U7821 ( .A(n9280), .ZN(n9109) );
  NAND2_X1 U7822 ( .A1(n9109), .A2(n5997), .ZN(n6274) );
  NAND2_X1 U7823 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  XNOR2_X1 U7824 ( .A(n6276), .B(n5751), .ZN(n6278) );
  OAI22_X1 U7825 ( .A1(n9508), .A2(n6326), .B1(n9280), .B2(n5773), .ZN(n6277)
         );
  XNOR2_X1 U7826 ( .A(n6278), .B(n6277), .ZN(n9000) );
  NOR2_X1 U7827 ( .A1(n6278), .A2(n6277), .ZN(n9077) );
  NAND2_X1 U7828 ( .A1(n7802), .A2(n7936), .ZN(n6280) );
  NAND2_X1 U7829 ( .A1(n6456), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U7830 ( .A1(n9248), .A2(n4508), .ZN(n6290) );
  INV_X1 U7831 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U7832 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U7833 ( .A1(n9249), .A2(n6299), .ZN(n6288) );
  INV_X1 U7834 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U7835 ( .A1(n6462), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7836 ( .A1(n5878), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U7837 ( .C1(n9502), .C2(n6639), .A(n6285), .B(n6284), .ZN(n6286)
         );
  INV_X1 U7838 ( .A(n6286), .ZN(n6287) );
  NAND2_X1 U7839 ( .A1(n9261), .A2(n5997), .ZN(n6289) );
  NAND2_X1 U7840 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  XNOR2_X1 U7841 ( .A(n6291), .B(n7030), .ZN(n6293) );
  AND2_X1 U7842 ( .A1(n9261), .A2(n5772), .ZN(n6292) );
  AOI21_X1 U7843 ( .B1(n9248), .B2(n5997), .A(n6292), .ZN(n6294) );
  XNOR2_X1 U7844 ( .A(n6293), .B(n6294), .ZN(n9076) );
  INV_X1 U7845 ( .A(n6293), .ZN(n6296) );
  INV_X1 U7846 ( .A(n6294), .ZN(n6295) );
  NAND2_X1 U7847 ( .A1(n7807), .A2(n7936), .ZN(n6298) );
  NAND2_X1 U7848 ( .A1(n6456), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n6297) );
  XNOR2_X1 U7849 ( .A(n6313), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9230) );
  NAND2_X1 U7850 ( .A1(n9230), .A2(n6299), .ZN(n6304) );
  INV_X1 U7851 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U7852 ( .A1(n6462), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7853 ( .A1(n5878), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6300) );
  OAI211_X1 U7854 ( .C1(n9499), .C2(n6639), .A(n6301), .B(n6300), .ZN(n6302)
         );
  INV_X1 U7855 ( .A(n6302), .ZN(n6303) );
  AOI22_X1 U7856 ( .A1(n6479), .A2(n4508), .B1(n5997), .B2(n9108), .ZN(n6305)
         );
  XNOR2_X1 U7857 ( .A(n6305), .B(n5751), .ZN(n6309) );
  AOI22_X1 U7858 ( .A1(n6479), .A2(n6307), .B1(n6306), .B2(n9108), .ZN(n6308)
         );
  NAND2_X1 U7859 ( .A1(n6309), .A2(n6308), .ZN(n6370) );
  OAI21_X1 U7860 ( .B1(n6309), .B2(n6308), .A(n6370), .ZN(n6473) );
  NAND2_X1 U7861 ( .A1(n8966), .A2(n7936), .ZN(n6311) );
  NAND2_X1 U7862 ( .A1(n6456), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7863 ( .A1(n6455), .A2(n6307), .ZN(n6323) );
  INV_X1 U7864 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6476) );
  INV_X1 U7865 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6312) );
  OAI21_X1 U7866 ( .B1(n6313), .B2(n6476), .A(n6312), .ZN(n6316) );
  INV_X1 U7867 ( .A(n6313), .ZN(n6315) );
  AND2_X1 U7868 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n6314) );
  NAND2_X1 U7869 ( .A1(n6315), .A2(n6314), .ZN(n9202) );
  NAND2_X1 U7870 ( .A1(n6316), .A2(n9202), .ZN(n6364) );
  OR2_X1 U7871 ( .A1(n6364), .A2(n5804), .ZN(n6321) );
  INV_X1 U7872 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7873 ( .A1(n6462), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U7874 ( .A1(n5878), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6317) );
  OAI211_X1 U7875 ( .C1(n6639), .C2(n6450), .A(n6318), .B(n6317), .ZN(n6319)
         );
  INV_X1 U7876 ( .A(n6319), .ZN(n6320) );
  NAND2_X1 U7877 ( .A1(n9107), .A2(n6306), .ZN(n6322) );
  NAND2_X1 U7878 ( .A1(n6323), .A2(n6322), .ZN(n6324) );
  XNOR2_X1 U7879 ( .A(n6324), .B(n7030), .ZN(n6328) );
  NAND2_X1 U7880 ( .A1(n6455), .A2(n4508), .ZN(n6325) );
  OAI21_X1 U7881 ( .B1(n9222), .B2(n6326), .A(n6325), .ZN(n6327) );
  XNOR2_X1 U7882 ( .A(n6328), .B(n6327), .ZN(n6353) );
  INV_X1 U7883 ( .A(n6353), .ZN(n6371) );
  NAND3_X1 U7884 ( .A1(n7749), .A2(P1_B_REG_SCAN_IN), .A3(n7705), .ZN(n6329)
         );
  OAI211_X1 U7885 ( .C1(P1_B_REG_SCAN_IN), .C2(n7705), .A(n6329), .B(n6330), 
        .ZN(n9965) );
  OR2_X1 U7886 ( .A1(n9965), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7887 ( .A1(n6331), .A2(n7749), .ZN(n6332) );
  NAND2_X1 U7888 ( .A1(n6333), .A2(n6332), .ZN(n6520) );
  OR2_X1 U7889 ( .A1(n9965), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U7890 ( .A1(n6331), .A2(n7705), .ZN(n6334) );
  NOR4_X1 U7891 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6344) );
  NOR4_X1 U7892 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6343) );
  NOR4_X1 U7893 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6339) );
  NOR4_X1 U7894 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6338) );
  NOR4_X1 U7895 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6337) );
  NOR4_X1 U7896 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6336) );
  NAND4_X1 U7897 ( .A1(n6339), .A2(n6338), .A3(n6337), .A4(n6336), .ZN(n6340)
         );
  NOR4_X1 U7898 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6341), .A4(n6340), .ZN(n6342) );
  AND3_X1 U7899 ( .A1(n6344), .A2(n6343), .A3(n6342), .ZN(n6345) );
  OR3_X1 U7900 ( .A1(n6520), .A2(n6507), .A3(n6484), .ZN(n6366) );
  NAND2_X1 U7901 ( .A1(n6346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6347) );
  XNOR2_X1 U7902 ( .A(n6347), .B(n4807), .ZN(n7628) );
  AND2_X1 U7903 ( .A1(n7628), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6348) );
  INV_X1 U7904 ( .A(n9966), .ZN(n6521) );
  NAND2_X1 U7905 ( .A1(n5753), .A2(n6350), .ZN(n6493) );
  AND2_X1 U7906 ( .A1(n9982), .A2(n6493), .ZN(n6351) );
  NAND3_X1 U7907 ( .A1(n6371), .A2(n9080), .A3(n6370), .ZN(n6352) );
  NAND3_X1 U7908 ( .A1(n6475), .A2(n6353), .A3(n9080), .ZN(n6375) );
  NOR2_X1 U7909 ( .A1(n6917), .A2(n8122), .ZN(n6916) );
  NAND2_X1 U7910 ( .A1(n6362), .A2(n6916), .ZN(n6355) );
  INV_X1 U7911 ( .A(n8122), .ZN(n6438) );
  NAND2_X1 U7912 ( .A1(n9966), .A2(n9184), .ZN(n6354) );
  OR2_X1 U7913 ( .A1(n9202), .A2(n5804), .ZN(n6360) );
  INV_X1 U7914 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U7915 ( .A1(n6462), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U7916 ( .A1(n6198), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6356) );
  OAI211_X1 U7917 ( .C1(n6487), .C2(n6080), .A(n6357), .B(n6356), .ZN(n6358)
         );
  INV_X1 U7918 ( .A(n6358), .ZN(n6359) );
  AND2_X1 U7919 ( .A1(n6362), .A2(n4378), .ZN(n6363) );
  NAND2_X1 U7920 ( .A1(n6363), .A2(n9891), .ZN(n9070) );
  INV_X1 U7921 ( .A(n9891), .ZN(n9861) );
  NAND2_X1 U7922 ( .A1(n9108), .A2(n9062), .ZN(n6369) );
  INV_X1 U7923 ( .A(n6364), .ZN(n9213) );
  NAND2_X1 U7924 ( .A1(n6366), .A2(n9982), .ZN(n6615) );
  NAND4_X1 U7925 ( .A1(n6615), .A2(n6913), .A3(n6492), .A4(n7628), .ZN(n6365)
         );
  NAND2_X1 U7926 ( .A1(n6365), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6367) );
  NAND3_X1 U7927 ( .A1(n6916), .A2(n9966), .A3(n6366), .ZN(n6616) );
  NAND2_X1 U7928 ( .A1(n6367), .A2(n6616), .ZN(n9082) );
  AOI22_X1 U7929 ( .A1(n9213), .A2(n9082), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6368) );
  OAI211_X1 U7930 ( .C1(n7944), .C2(n9070), .A(n6369), .B(n6368), .ZN(n6373)
         );
  NOR3_X1 U7931 ( .A1(n6371), .A2(n9103), .A3(n6370), .ZN(n6372) );
  AOI211_X1 U7932 ( .C1(n6455), .C2(n6480), .A(n6373), .B(n6372), .ZN(n6374)
         );
  NAND3_X1 U7933 ( .A1(n4900), .A2(n6375), .A3(n6374), .ZN(P1_U3218) );
  AND2_X1 U7934 ( .A1(n6376), .A2(n6920), .ZN(n6706) );
  NAND2_X1 U7935 ( .A1(n5771), .A2(n5774), .ZN(n6377) );
  NAND2_X1 U7936 ( .A1(n9127), .A2(n6839), .ZN(n8084) );
  OR2_X1 U7937 ( .A1(n9127), .A2(n4839), .ZN(n6378) );
  NAND2_X1 U7938 ( .A1(n6675), .A2(n6378), .ZN(n7333) );
  NAND2_X1 U7939 ( .A1(n9126), .A2(n9969), .ZN(n8023) );
  NAND2_X1 U7940 ( .A1(n7333), .A2(n7961), .ZN(n7332) );
  INV_X1 U7941 ( .A(n9969), .ZN(n7338) );
  OR2_X1 U7942 ( .A1(n9126), .A2(n7338), .ZN(n6379) );
  NAND2_X1 U7943 ( .A1(n7332), .A2(n6379), .ZN(n6888) );
  OR2_X1 U7944 ( .A1(n9125), .A2(n7089), .ZN(n8026) );
  NAND2_X1 U7945 ( .A1(n9125), .A2(n7089), .ZN(n8024) );
  NAND2_X1 U7946 ( .A1(n8026), .A2(n8024), .ZN(n6890) );
  INV_X1 U7947 ( .A(n7089), .ZN(n6889) );
  OR2_X1 U7948 ( .A1(n9125), .A2(n6889), .ZN(n6380) );
  OR2_X1 U7949 ( .A1(n9124), .A2(n9976), .ZN(n7828) );
  NAND2_X1 U7950 ( .A1(n9124), .A2(n9976), .ZN(n7830) );
  NAND2_X1 U7951 ( .A1(n7828), .A2(n7830), .ZN(n7217) );
  INV_X1 U7952 ( .A(n7217), .ZN(n7222) );
  NAND2_X1 U7953 ( .A1(n9124), .A2(n4509), .ZN(n6381) );
  OR2_X1 U7954 ( .A1(n9123), .A2(n7008), .ZN(n8091) );
  NAND2_X1 U7955 ( .A1(n9123), .A2(n7008), .ZN(n7826) );
  NAND2_X1 U7956 ( .A1(n8091), .A2(n7826), .ZN(n7824) );
  OR2_X1 U7957 ( .A1(n9123), .A2(n9413), .ZN(n6382) );
  NAND2_X1 U7958 ( .A1(n9122), .A2(n7352), .ZN(n7833) );
  NAND2_X1 U7959 ( .A1(n8017), .A2(n7833), .ZN(n7968) );
  INV_X1 U7960 ( .A(n9122), .ZN(n7004) );
  NAND2_X1 U7961 ( .A1(n7004), .A2(n7352), .ZN(n6383) );
  OR2_X1 U7962 ( .A1(n9121), .A2(n7308), .ZN(n8016) );
  NAND2_X1 U7963 ( .A1(n9121), .A2(n7308), .ZN(n7841) );
  NAND2_X1 U7964 ( .A1(n8016), .A2(n7841), .ZN(n7969) );
  INV_X1 U7965 ( .A(n7969), .ZN(n7244) );
  INV_X1 U7966 ( .A(n7308), .ZN(n7270) );
  NAND2_X1 U7967 ( .A1(n9121), .A2(n7270), .ZN(n6384) );
  NAND2_X1 U7968 ( .A1(n7235), .A2(n6384), .ZN(n7312) );
  AND2_X1 U7969 ( .A1(n7320), .A2(n9120), .ZN(n6385) );
  OAI22_X1 U7970 ( .A1(n7312), .A2(n6385), .B1(n9120), .B2(n7320), .ZN(n7391)
         );
  OR2_X1 U7971 ( .A1(n7398), .A2(n7442), .ZN(n8033) );
  NAND2_X1 U7972 ( .A1(n7398), .A2(n7442), .ZN(n7848) );
  NAND2_X1 U7973 ( .A1(n8033), .A2(n7848), .ZN(n7392) );
  NAND2_X1 U7974 ( .A1(n7391), .A2(n7392), .ZN(n6387) );
  INV_X1 U7975 ( .A(n7442), .ZN(n9119) );
  OR2_X1 U7976 ( .A1(n7398), .A2(n9119), .ZN(n6386) );
  NAND2_X1 U7977 ( .A1(n6387), .A2(n6386), .ZN(n7440) );
  NOR2_X1 U7978 ( .A1(n9844), .A2(n9118), .ZN(n6389) );
  NAND2_X1 U7979 ( .A1(n9844), .A2(n9118), .ZN(n6388) );
  OR2_X1 U7980 ( .A1(n7646), .A2(n7757), .ZN(n7859) );
  NAND2_X1 U7981 ( .A1(n7646), .A2(n7757), .ZN(n7858) );
  NAND2_X1 U7982 ( .A1(n7859), .A2(n7858), .ZN(n7976) );
  NAND2_X1 U7983 ( .A1(n7615), .A2(n7976), .ZN(n6391) );
  INV_X1 U7984 ( .A(n7757), .ZN(n9117) );
  NAND2_X1 U7985 ( .A1(n7646), .A2(n9117), .ZN(n6390) );
  NAND2_X1 U7986 ( .A1(n6391), .A2(n6390), .ZN(n7752) );
  OR2_X1 U7987 ( .A1(n9830), .A2(n9116), .ZN(n6392) );
  NAND2_X1 U7988 ( .A1(n7752), .A2(n6392), .ZN(n6394) );
  NAND2_X1 U7989 ( .A1(n9830), .A2(n9116), .ZN(n6393) );
  NAND2_X1 U7990 ( .A1(n6394), .A2(n6393), .ZN(n7727) );
  OR2_X1 U7991 ( .A1(n7797), .A2(n9115), .ZN(n6395) );
  NOR2_X1 U7992 ( .A1(n9100), .A2(n9114), .ZN(n6396) );
  OR2_X1 U7993 ( .A1(n9017), .A2(n9402), .ZN(n8047) );
  NAND2_X1 U7994 ( .A1(n9017), .A2(n9402), .ZN(n8011) );
  NAND2_X1 U7995 ( .A1(n8047), .A2(n8011), .ZN(n7810) );
  INV_X1 U7996 ( .A(n9402), .ZN(n9113) );
  OR2_X1 U7997 ( .A1(n9483), .A2(n9112), .ZN(n6397) );
  NAND2_X1 U7998 ( .A1(n9386), .A2(n6397), .ZN(n6399) );
  NAND2_X1 U7999 ( .A1(n9483), .A2(n9112), .ZN(n6398) );
  NAND2_X1 U8000 ( .A1(n6399), .A2(n6398), .ZN(n9374) );
  OR2_X1 U8001 ( .A1(n9378), .A2(n9404), .ZN(n7882) );
  NAND2_X1 U8002 ( .A1(n9378), .A2(n9404), .ZN(n8013) );
  NAND2_X1 U8003 ( .A1(n7882), .A2(n8013), .ZN(n9375) );
  INV_X1 U8004 ( .A(n9404), .ZN(n9111) );
  NAND2_X1 U8005 ( .A1(n9378), .A2(n9111), .ZN(n6400) );
  OR2_X1 U8006 ( .A1(n9473), .A2(n9347), .ZN(n6401) );
  NOR2_X1 U8007 ( .A1(n9467), .A2(n9321), .ZN(n6402) );
  INV_X1 U8008 ( .A(n9467), .ZN(n9342) );
  NAND2_X1 U8009 ( .A1(n9328), .A2(n9306), .ZN(n7896) );
  NAND2_X1 U8010 ( .A1(n7998), .A2(n7896), .ZN(n6432) );
  NAND2_X1 U8011 ( .A1(n9317), .A2(n6432), .ZN(n6404) );
  NAND2_X1 U8012 ( .A1(n9328), .A2(n9349), .ZN(n6403) );
  NOR2_X1 U8013 ( .A1(n9453), .A2(n9110), .ZN(n6405) );
  NAND2_X1 U8014 ( .A1(n9453), .A2(n9110), .ZN(n7905) );
  OR2_X1 U8015 ( .A1(n9282), .A2(n9260), .ZN(n6406) );
  NAND2_X1 U8016 ( .A1(n6407), .A2(n6406), .ZN(n9255) );
  NAND2_X1 U8017 ( .A1(n9267), .A2(n9280), .ZN(n7917) );
  NAND2_X1 U8018 ( .A1(n9237), .A2(n7917), .ZN(n9257) );
  OR2_X1 U8019 ( .A1(n9267), .A2(n9109), .ZN(n6408) );
  NOR2_X1 U8020 ( .A1(n9248), .A2(n9261), .ZN(n7985) );
  NAND2_X1 U8021 ( .A1(n6479), .A2(n9243), .ZN(n8058) );
  OR2_X1 U8022 ( .A1(n6479), .A2(n9108), .ZN(n6409) );
  NAND2_X1 U8023 ( .A1(n6455), .A2(n9222), .ZN(n8059) );
  OR2_X1 U8024 ( .A1(n6412), .A2(n7071), .ZN(n6415) );
  OR2_X1 U8025 ( .A1(n6413), .A2(n8066), .ZN(n6414) );
  NAND2_X1 U8026 ( .A1(n6415), .A2(n6414), .ZN(n9824) );
  INV_X1 U8027 ( .A(n6920), .ZN(n6624) );
  NAND3_X1 U8028 ( .A1(n8079), .A2(n6839), .A3(n6624), .ZN(n7334) );
  OR2_X1 U8029 ( .A1(n7334), .A2(n7338), .ZN(n7335) );
  INV_X1 U8030 ( .A(n7320), .ZN(n9983) );
  NAND2_X1 U8031 ( .A1(n7317), .A2(n9983), .ZN(n7394) );
  INV_X1 U8032 ( .A(n7646), .ZN(n7712) );
  INV_X1 U8033 ( .A(n9483), .ZN(n9393) );
  NAND2_X1 U8034 ( .A1(n9387), .A2(n9393), .ZN(n9388) );
  INV_X1 U8035 ( .A(n9328), .ZN(n9518) );
  NAND2_X1 U8036 ( .A1(n9281), .A2(n9508), .ZN(n9264) );
  NAND2_X1 U8037 ( .A1(n9229), .A2(n6455), .ZN(n6416) );
  NAND2_X1 U8038 ( .A1(n6416), .A2(n9228), .ZN(n6417) );
  NOR2_X1 U8039 ( .A1(n6468), .A2(n6417), .ZN(n9212) );
  NOR2_X1 U8040 ( .A1(n6376), .A2(n6624), .ZN(n6711) );
  INV_X1 U8041 ( .A(n5771), .ZN(n6619) );
  NAND2_X1 U8042 ( .A1(n6619), .A2(n5774), .ZN(n6418) );
  NAND2_X1 U8043 ( .A1(n8086), .A2(n7964), .ZN(n6679) );
  NAND2_X1 U8044 ( .A1(n6679), .A2(n8082), .ZN(n8025) );
  INV_X1 U8045 ( .A(n7961), .ZN(n6419) );
  INV_X1 U8046 ( .A(n8026), .ZN(n6420) );
  NAND2_X1 U8047 ( .A1(n8091), .A2(n7828), .ZN(n8027) );
  INV_X1 U8048 ( .A(n8027), .ZN(n6421) );
  NAND2_X1 U8049 ( .A1(n7218), .A2(n6421), .ZN(n6424) );
  INV_X1 U8050 ( .A(n7830), .ZN(n6422) );
  NAND2_X1 U8051 ( .A1(n6422), .A2(n8091), .ZN(n8094) );
  AND2_X1 U8052 ( .A1(n8094), .A2(n7826), .ZN(n6423) );
  INV_X1 U8053 ( .A(n8017), .ZN(n6425) );
  NOR2_X1 U8054 ( .A1(n6425), .A2(n7969), .ZN(n6426) );
  INV_X1 U8055 ( .A(n9120), .ZN(n7266) );
  OR2_X1 U8056 ( .A1(n7320), .A2(n7266), .ZN(n7842) );
  NAND2_X1 U8057 ( .A1(n7320), .A2(n7266), .ZN(n7845) );
  NAND2_X1 U8058 ( .A1(n7314), .A2(n7972), .ZN(n7313) );
  NAND2_X1 U8059 ( .A1(n7313), .A2(n7842), .ZN(n7389) );
  INV_X1 U8060 ( .A(n7392), .ZN(n7973) );
  NAND2_X1 U8061 ( .A1(n7389), .A2(n7973), .ZN(n6427) );
  INV_X1 U8062 ( .A(n9118), .ZN(n7642) );
  NAND2_X1 U8063 ( .A1(n9844), .A2(n7642), .ZN(n7857) );
  OR2_X1 U8064 ( .A1(n9844), .A2(n7642), .ZN(n7621) );
  AND2_X1 U8065 ( .A1(n7859), .A2(n7621), .ZN(n7853) );
  XNOR2_X1 U8066 ( .A(n9830), .B(n9116), .ZN(n7979) );
  NAND2_X1 U8067 ( .A1(n7755), .A2(n7979), .ZN(n6428) );
  INV_X1 U8068 ( .A(n9116), .ZN(n7854) );
  NAND2_X1 U8069 ( .A1(n9830), .A2(n7854), .ZN(n7856) );
  INV_X1 U8070 ( .A(n9115), .ZN(n9093) );
  NAND2_X1 U8071 ( .A1(n7797), .A2(n9093), .ZN(n7867) );
  NAND2_X1 U8072 ( .A1(n7869), .A2(n7867), .ZN(n7978) );
  INV_X1 U8073 ( .A(n9114), .ZN(n9013) );
  OR2_X1 U8074 ( .A1(n9100), .A2(n9013), .ZN(n8046) );
  NAND2_X1 U8075 ( .A1(n9100), .A2(n9013), .ZN(n8043) );
  NAND2_X1 U8076 ( .A1(n8046), .A2(n8043), .ZN(n7865) );
  INV_X1 U8077 ( .A(n7869), .ZN(n8042) );
  INV_X1 U8078 ( .A(n7810), .ZN(n7981) );
  INV_X1 U8079 ( .A(n9112), .ZN(n9372) );
  AND2_X1 U8080 ( .A1(n9483), .A2(n9372), .ZN(n8012) );
  OR2_X1 U8081 ( .A1(n9483), .A2(n9372), .ZN(n9368) );
  AND2_X1 U8082 ( .A1(n7882), .A2(n9368), .ZN(n8000) );
  INV_X1 U8083 ( .A(n9347), .ZN(n9373) );
  OR2_X1 U8084 ( .A1(n9473), .A2(n9373), .ZN(n7883) );
  NAND2_X1 U8085 ( .A1(n9473), .A2(n9373), .ZN(n8008) );
  NAND2_X1 U8086 ( .A1(n9363), .A2(n7959), .ZN(n6431) );
  NAND2_X1 U8087 ( .A1(n6431), .A2(n8008), .ZN(n9344) );
  OR2_X1 U8088 ( .A1(n9467), .A2(n9365), .ZN(n7895) );
  NAND2_X1 U8089 ( .A1(n9467), .A2(n9365), .ZN(n7889) );
  NAND2_X1 U8090 ( .A1(n9344), .A2(n9345), .ZN(n9343) );
  INV_X1 U8091 ( .A(n9322), .ZN(n9293) );
  OR2_X1 U8092 ( .A1(n9458), .A2(n9293), .ZN(n8002) );
  NAND2_X1 U8093 ( .A1(n9458), .A2(n9293), .ZN(n7900) );
  AND2_X1 U8094 ( .A1(n9453), .A2(n9307), .ZN(n7958) );
  OR2_X1 U8095 ( .A1(n9453), .A2(n9307), .ZN(n8003) );
  INV_X1 U8096 ( .A(n9260), .ZN(n9294) );
  OR2_X1 U8097 ( .A1(n9282), .A2(n9294), .ZN(n8006) );
  NAND2_X1 U8098 ( .A1(n9282), .A2(n9294), .ZN(n9256) );
  AND2_X1 U8099 ( .A1(n7917), .A2(n9256), .ZN(n8107) );
  NAND2_X1 U8100 ( .A1(n9275), .A2(n8107), .ZN(n9238) );
  INV_X1 U8101 ( .A(n9261), .ZN(n9221) );
  OR2_X1 U8102 ( .A1(n9248), .A2(n9221), .ZN(n6434) );
  AND2_X1 U8103 ( .A1(n6434), .A2(n9237), .ZN(n8109) );
  NAND2_X1 U8104 ( .A1(n9238), .A2(n8109), .ZN(n6435) );
  NAND2_X1 U8105 ( .A1(n9248), .A2(n9221), .ZN(n8055) );
  NAND2_X1 U8106 ( .A1(n6435), .A2(n8055), .ZN(n9220) );
  INV_X1 U8107 ( .A(n9225), .ZN(n7915) );
  INV_X1 U8108 ( .A(n7987), .ZN(n6436) );
  NAND3_X1 U8109 ( .A1(n6437), .A2(n6436), .A3(n8060), .ZN(n6441) );
  NAND2_X1 U8110 ( .A1(n5753), .A2(n9184), .ZN(n6440) );
  NAND2_X1 U8111 ( .A1(n6350), .A2(n6438), .ZN(n6439) );
  NAND2_X1 U8112 ( .A1(n6441), .A2(n9351), .ZN(n6442) );
  OR2_X1 U8113 ( .A1(n6460), .A2(n6442), .ZN(n6445) );
  INV_X1 U8114 ( .A(n6493), .ZN(n7953) );
  OAI22_X1 U8115 ( .A1(n9243), .A2(n9403), .B1(n7944), .B2(n9405), .ZN(n6443)
         );
  INV_X1 U8116 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8117 ( .A1(n6445), .A2(n6444), .ZN(n9217) );
  AND2_X1 U8118 ( .A1(n6520), .A2(n9966), .ZN(n6446) );
  AND2_X1 U8119 ( .A1(n6913), .A2(n6446), .ZN(n6448) );
  OR2_X1 U8120 ( .A1(n9390), .A2(n8070), .ZN(n6447) );
  INV_X1 U8121 ( .A(n6484), .ZN(n6449) );
  AND2_X1 U8122 ( .A1(n6449), .A2(n6507), .ZN(n6915) );
  INV_X1 U8123 ( .A(n9529), .ZN(n6451) );
  NAND2_X1 U8124 ( .A1(n6455), .A2(n6451), .ZN(n6452) );
  NAND2_X1 U8125 ( .A1(n6453), .A2(n6452), .ZN(P1_U3519) );
  AOI21_X1 U8126 ( .B1(n6455), .B2(n9107), .A(n6454), .ZN(n6459) );
  NAND2_X1 U8127 ( .A1(n8132), .A2(n7936), .ZN(n6458) );
  NAND2_X1 U8128 ( .A1(n6456), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6457) );
  OR2_X1 U8129 ( .A1(n6470), .A2(n7944), .ZN(n8063) );
  NAND2_X1 U8130 ( .A1(n6470), .A2(n7944), .ZN(n8113) );
  NAND2_X1 U8131 ( .A1(n8063), .A2(n8113), .ZN(n7989) );
  XNOR2_X1 U8132 ( .A(n6459), .B(n7989), .ZN(n9200) );
  INV_X1 U8133 ( .A(n9886), .ZN(n9858) );
  AND2_X1 U8134 ( .A1(n9858), .A2(P1_B_REG_SCAN_IN), .ZN(n6461) );
  NOR2_X1 U8135 ( .A1(n9405), .A2(n6461), .ZN(n9191) );
  INV_X1 U8136 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n6465) );
  NAND2_X1 U8137 ( .A1(n6462), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U8138 ( .A1(n5878), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6463) );
  OAI211_X1 U8139 ( .C1(n6639), .C2(n6465), .A(n6464), .B(n6463), .ZN(n9105)
         );
  AOI22_X1 U8140 ( .A1(n9107), .A2(n9346), .B1(n9191), .B2(n9105), .ZN(n6466)
         );
  OAI21_X1 U8141 ( .B1(n6467), .B2(n9400), .A(n6466), .ZN(n9208) );
  INV_X1 U8142 ( .A(n6468), .ZN(n6469) );
  AOI211_X1 U8143 ( .C1(n6470), .C2(n6469), .A(n9390), .B(n9195), .ZN(n9201)
         );
  OAI21_X1 U8144 ( .B1(n6475), .B2(n4346), .A(n9080), .ZN(n6483) );
  OAI22_X1 U8145 ( .A1(n9221), .A2(n9094), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6476), .ZN(n6478) );
  NOR2_X1 U8146 ( .A1(n9222), .A2(n9070), .ZN(n6477) );
  AOI211_X1 U8147 ( .C1(n9230), .C2(n9082), .A(n6478), .B(n6477), .ZN(n6482)
         );
  NAND3_X1 U8148 ( .A1(n6483), .A2(n6482), .A3(n6481), .ZN(P1_U3212) );
  NOR2_X1 U8149 ( .A1(n6484), .A2(n6507), .ZN(n6485) );
  INV_X1 U8150 ( .A(n6488), .ZN(n6489) );
  OAI21_X1 U8151 ( .B1(n6490), .B2(n9992), .A(n6489), .ZN(P1_U3552) );
  INV_X1 U8152 ( .A(n7628), .ZN(n6491) );
  AND2_X2 U8153 ( .A1(n9890), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND2_X1 U8154 ( .A1(n6493), .A2(n6492), .ZN(n6494) );
  NAND2_X1 U8155 ( .A1(n6494), .A2(n7628), .ZN(n9179) );
  NAND2_X1 U8156 ( .A1(n9179), .A2(n5814), .ZN(n9859) );
  NAND2_X1 U8157 ( .A1(n9859), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8158 ( .A(n6878), .ZN(n6796) );
  XNOR2_X1 U8159 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U8160 ( .A1(n6496), .A2(P2_U3152), .ZN(n8968) );
  INV_X2 U8161 ( .A(n8968), .ZN(n8963) );
  NAND2_X1 U8162 ( .A1(n6495), .A2(P2_U3152), .ZN(n8973) );
  OAI222_X1 U8163 ( .A1(n8963), .A2(n4976), .B1(n8973), .B2(n6512), .C1(
        P2_U3152), .C2(n8248), .ZN(P2_U3357) );
  OR2_X1 U8164 ( .A1(n6496), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8339) );
  INV_X1 U8165 ( .A(n8339), .ZN(n9535) );
  AOI22_X1 U8166 ( .A1(n9918), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9535), .ZN(n6497) );
  OAI21_X1 U8167 ( .B1(n6505), .B2(n9537), .A(n6497), .ZN(P1_U3348) );
  INV_X1 U8168 ( .A(n6550), .ZN(n9909) );
  INV_X1 U8169 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6498) );
  OAI222_X1 U8170 ( .A1(P1_U3084), .A2(n9909), .B1(n9537), .B2(n6501), .C1(
        n6498), .C2(n8339), .ZN(P1_U3349) );
  AOI22_X1 U8171 ( .A1(n9129), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9535), .ZN(n6499) );
  OAI21_X1 U8172 ( .B1(n6503), .B2(n9537), .A(n6499), .ZN(P1_U3347) );
  INV_X1 U8173 ( .A(n8973), .ZN(n7631) );
  OAI222_X1 U8174 ( .A1(n8963), .A2(n6500), .B1(n8970), .B2(n6516), .C1(
        P2_U3152), .C2(n8237), .ZN(P2_U3355) );
  OAI222_X1 U8175 ( .A1(n8963), .A2(n4565), .B1(n8970), .B2(n6501), .C1(
        P2_U3152), .C2(n8226), .ZN(P2_U3354) );
  OAI222_X1 U8176 ( .A1(n8963), .A2(n6502), .B1(n8970), .B2(n6514), .C1(
        P2_U3152), .C2(n6810), .ZN(P2_U3356) );
  OAI222_X1 U8177 ( .A1(n8963), .A2(n6504), .B1(n8970), .B2(n6503), .C1(
        P2_U3152), .C2(n8204), .ZN(P2_U3352) );
  OAI222_X1 U8178 ( .A1(n8963), .A2(n6506), .B1(n8970), .B2(n6505), .C1(
        P2_U3152), .C2(n8215), .ZN(P2_U3353) );
  INV_X1 U8179 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6510) );
  INV_X1 U8180 ( .A(n6507), .ZN(n6508) );
  NAND2_X1 U8181 ( .A1(n6508), .A2(n9966), .ZN(n6509) );
  OAI21_X1 U8182 ( .B1(n9966), .B2(n6510), .A(n6509), .ZN(P1_U3440) );
  INV_X1 U8183 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6511) );
  OAI222_X1 U8184 ( .A1(P1_U3084), .A2(n5764), .B1(n9537), .B2(n6512), .C1(
        n6511), .C2(n8339), .ZN(P1_U3352) );
  INV_X1 U8185 ( .A(n6548), .ZN(n9897) );
  INV_X1 U8186 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6513) );
  OAI222_X1 U8187 ( .A1(P1_U3084), .A2(n9897), .B1(n9537), .B2(n6514), .C1(
        n6513), .C2(n8339), .ZN(P1_U3351) );
  INV_X1 U8188 ( .A(n6549), .ZN(n9762) );
  INV_X1 U8189 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6515) );
  OAI222_X1 U8190 ( .A1(P1_U3084), .A2(n9762), .B1(n9537), .B2(n6516), .C1(
        n6515), .C2(n8339), .ZN(P1_U3350) );
  OAI222_X1 U8191 ( .A1(n8963), .A2(n6517), .B1(n8970), .B2(n6518), .C1(
        P2_U3152), .C2(n8193), .ZN(P2_U3351) );
  INV_X1 U8192 ( .A(n6572), .ZN(n6566) );
  OAI222_X1 U8193 ( .A1(n8339), .A2(n6519), .B1(n9537), .B2(n6518), .C1(
        P1_U3084), .C2(n6566), .ZN(P1_U3346) );
  INV_X1 U8194 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6523) );
  NOR2_X1 U8195 ( .A1(n6521), .A2(n6520), .ZN(n6914) );
  INV_X1 U8196 ( .A(n6914), .ZN(n6522) );
  OAI21_X1 U8197 ( .B1(n9966), .B2(n6523), .A(n6522), .ZN(P1_U3441) );
  INV_X1 U8198 ( .A(n6524), .ZN(n6526) );
  INV_X1 U8199 ( .A(n6821), .ZN(n8182) );
  OAI222_X1 U8200 ( .A1(n8963), .A2(n6525), .B1(n8970), .B2(n6526), .C1(
        P2_U3152), .C2(n8182), .ZN(P2_U3350) );
  INV_X1 U8201 ( .A(n6593), .ZN(n6564) );
  OAI222_X1 U8202 ( .A1(n8339), .A2(n6527), .B1(n9537), .B2(n6526), .C1(
        P1_U3084), .C2(n6564), .ZN(P1_U3345) );
  INV_X1 U8203 ( .A(n6528), .ZN(n6530) );
  INV_X1 U8204 ( .A(n6597), .ZN(n9942) );
  OAI222_X1 U8205 ( .A1(n8339), .A2(n6529), .B1(n9537), .B2(n6530), .C1(n9942), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8206 ( .A(n6823), .ZN(n8171) );
  OAI222_X1 U8207 ( .A1(n8963), .A2(n6531), .B1(n8970), .B2(n6530), .C1(n8171), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  AOI22_X1 U8208 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6566), .B1(n6572), .B2(
        n7040), .ZN(n6540) );
  NAND2_X1 U8209 ( .A1(n9129), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6538) );
  MUX2_X1 U8210 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6532), .S(n6549), .Z(n9770)
         );
  MUX2_X1 U8211 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6534), .S(n6546), .Z(n9877)
         );
  NAND3_X1 U8212 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .A3(n9877), .ZN(n9876) );
  OAI21_X1 U8213 ( .B1(n5764), .B2(n6534), .A(n9876), .ZN(n9895) );
  OAI21_X1 U8214 ( .B1(n9897), .B2(n6533), .A(n9893), .ZN(n9771) );
  NAND2_X1 U8215 ( .A1(n9770), .A2(n9771), .ZN(n9769) );
  OAI21_X1 U8216 ( .B1(n6532), .B2(n9762), .A(n9769), .ZN(n9908) );
  AOI22_X1 U8217 ( .A1(n6550), .A2(n5832), .B1(P1_REG2_REG_4__SCAN_IN), .B2(
        n9909), .ZN(n9907) );
  NOR2_X1 U8218 ( .A1(n6550), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6535) );
  MUX2_X1 U8219 ( .A(n6536), .B(P1_REG2_REG_5__SCAN_IN), .S(n9918), .Z(n9926)
         );
  MUX2_X1 U8220 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6537), .S(n9129), .Z(n9131)
         );
  NAND2_X1 U8221 ( .A1(n9132), .A2(n9131), .ZN(n9130) );
  NAND2_X1 U8222 ( .A1(n6538), .A2(n9130), .ZN(n6539) );
  NOR2_X1 U8223 ( .A1(n6540), .A2(n6539), .ZN(n6565) );
  AOI21_X1 U8224 ( .B1(n6540), .B2(n6539), .A(n6565), .ZN(n6559) );
  NAND2_X1 U8225 ( .A1(n9861), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9864) );
  NOR2_X1 U8226 ( .A1(n9864), .A2(n9886), .ZN(n6541) );
  AND2_X1 U8227 ( .A1(n9179), .A2(n6541), .ZN(n9960) );
  OR2_X1 U8228 ( .A1(n9886), .A2(P1_U3084), .ZN(n9180) );
  INV_X1 U8229 ( .A(n9180), .ZN(n7808) );
  AND2_X1 U8230 ( .A1(n9891), .A2(n7808), .ZN(n6542) );
  NAND2_X1 U8231 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6959) );
  OAI21_X1 U8232 ( .B1(n9943), .B2(n6566), .A(n6959), .ZN(n6543) );
  AOI21_X1 U8233 ( .B1(n9866), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6543), .ZN(
        n6558) );
  AOI22_X1 U8234 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6572), .B1(n6566), .B2(
        n5909), .ZN(n6554) );
  NAND2_X1 U8235 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n9918), .ZN(n6544) );
  OAI21_X1 U8236 ( .B1(n9918), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6544), .ZN(
        n9920) );
  AOI22_X1 U8237 ( .A1(n6550), .A2(P1_REG1_REG_4__SCAN_IN), .B1(n5833), .B2(
        n9909), .ZN(n9904) );
  INV_X1 U8238 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9867) );
  INV_X1 U8239 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6545) );
  MUX2_X1 U8240 ( .A(n6545), .B(P1_REG1_REG_1__SCAN_IN), .S(n6546), .Z(n9871)
         );
  NOR3_X1 U8241 ( .A1(n9862), .A2(n9867), .A3(n9871), .ZN(n9870) );
  AOI21_X1 U8242 ( .B1(n6546), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9870), .ZN(
        n9885) );
  INV_X1 U8243 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6547) );
  MUX2_X1 U8244 ( .A(n6547), .B(P1_REG1_REG_2__SCAN_IN), .S(n6548), .Z(n9884)
         );
  NOR2_X1 U8245 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  AOI21_X1 U8246 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6548), .A(n9883), .ZN(
        n9766) );
  AOI22_X1 U8247 ( .A1(n6549), .A2(n5806), .B1(P1_REG1_REG_3__SCAN_IN), .B2(
        n9762), .ZN(n9767) );
  NOR2_X1 U8248 ( .A1(n9766), .A2(n9767), .ZN(n9765) );
  AOI21_X1 U8249 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6549), .A(n9765), .ZN(
        n9903) );
  NAND2_X1 U8250 ( .A1(n9904), .A2(n9903), .ZN(n9902) );
  OR2_X1 U8251 ( .A1(n6550), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U8252 ( .A1(n9902), .A2(n6551), .ZN(n9921) );
  NOR2_X1 U8253 ( .A1(n9920), .A2(n9921), .ZN(n9919) );
  AOI21_X1 U8254 ( .B1(n9918), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9919), .ZN(
        n9134) );
  NOR2_X1 U8255 ( .A1(n9129), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6552) );
  AOI21_X1 U8256 ( .B1(n9129), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6552), .ZN(
        n9135) );
  NAND2_X1 U8257 ( .A1(n9134), .A2(n9135), .ZN(n9133) );
  OAI21_X1 U8258 ( .B1(n9129), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9133), .ZN(
        n6553) );
  NAND2_X1 U8259 ( .A1(n6554), .A2(n6553), .ZN(n6571) );
  OAI21_X1 U8260 ( .B1(n6554), .B2(n6553), .A(n6571), .ZN(n6556) );
  NOR2_X1 U8261 ( .A1(n9864), .A2(n9858), .ZN(n6555) );
  NAND2_X1 U8262 ( .A1(n6556), .A2(n9959), .ZN(n6557) );
  OAI211_X1 U8263 ( .C1(n6559), .C2(n9935), .A(n6558), .B(n6557), .ZN(P1_U3248) );
  INV_X1 U8264 ( .A(n6560), .ZN(n6562) );
  INV_X1 U8265 ( .A(n6825), .ZN(n8160) );
  OAI222_X1 U8266 ( .A1(n8963), .A2(n6561), .B1(n8970), .B2(n6562), .C1(n8160), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8267 ( .A(n6651), .ZN(n6588) );
  OAI222_X1 U8268 ( .A1(n8339), .A2(n6563), .B1(n9537), .B2(n6562), .C1(n6588), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  NOR2_X1 U8269 ( .A1(n6564), .A2(n7240), .ZN(n6594) );
  AOI21_X1 U8270 ( .B1(n6564), .B2(n7240), .A(n6594), .ZN(n6567) );
  AOI21_X1 U8271 ( .B1(n7040), .B2(n6566), .A(n6565), .ZN(n6595) );
  XOR2_X1 U8272 ( .A(n6567), .B(n6595), .Z(n6578) );
  INV_X1 U8273 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n6570) );
  NOR2_X1 U8274 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6568), .ZN(n7269) );
  AOI21_X1 U8275 ( .B1(n9951), .B2(n6593), .A(n7269), .ZN(n6569) );
  OAI21_X1 U8276 ( .B1(n9964), .B2(n6570), .A(n6569), .ZN(n6577) );
  OAI21_X1 U8277 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6572), .A(n6571), .ZN(
        n6575) );
  MUX2_X1 U8278 ( .A(n6573), .B(P1_REG1_REG_8__SCAN_IN), .S(n6593), .Z(n6574)
         );
  NOR2_X1 U8279 ( .A1(n6574), .A2(n6575), .ZN(n6587) );
  INV_X1 U8280 ( .A(n9959), .ZN(n9882) );
  AOI211_X1 U8281 ( .C1(n6575), .C2(n6574), .A(n6587), .B(n9882), .ZN(n6576)
         );
  AOI211_X1 U8282 ( .C1(n6578), .C2(n9960), .A(n6577), .B(n6576), .ZN(n6579)
         );
  INV_X1 U8283 ( .A(n6579), .ZN(P1_U3249) );
  INV_X1 U8284 ( .A(n6983), .ZN(n6831) );
  INV_X1 U8285 ( .A(n6580), .ZN(n6582) );
  INV_X1 U8286 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6581) );
  OAI222_X1 U8287 ( .A1(P2_U3152), .A2(n6831), .B1(n8970), .B2(n6582), .C1(
        n6581), .C2(n8963), .ZN(P2_U3347) );
  INV_X1 U8288 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6583) );
  INV_X1 U8289 ( .A(n6652), .ZN(n9145) );
  OAI222_X1 U8290 ( .A1(n8339), .A2(n6583), .B1(n9537), .B2(n6582), .C1(n9145), 
        .C2(P1_U3084), .ZN(P1_U3342) );
  NAND2_X1 U8291 ( .A1(n10008), .A2(n6753), .ZN(n6584) );
  NAND2_X1 U8292 ( .A1(n6584), .A2(n6804), .ZN(n6586) );
  OR2_X1 U8293 ( .A1(n10008), .A2(n5684), .ZN(n6585) );
  NAND2_X1 U8294 ( .A1(n6586), .A2(n6585), .ZN(n8587) );
  NOR2_X1 U8295 ( .A1(n10002), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8296 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6604) );
  AOI21_X1 U8297 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n6593), .A(n6587), .ZN(
        n9934) );
  AOI22_X1 U8298 ( .A1(n6597), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n5951), .B2(
        n9942), .ZN(n9933) );
  NAND2_X1 U8299 ( .A1(n9934), .A2(n9933), .ZN(n9932) );
  OAI21_X1 U8300 ( .B1(n6597), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9932), .ZN(
        n6590) );
  AOI22_X1 U8301 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6651), .B1(n6588), .B2(
        n5970), .ZN(n6589) );
  NAND2_X1 U8302 ( .A1(n6589), .A2(n6590), .ZN(n6643) );
  OAI21_X1 U8303 ( .B1(n6590), .B2(n6589), .A(n6643), .ZN(n6591) );
  NAND2_X1 U8304 ( .A1(n6591), .A2(n9959), .ZN(n6603) );
  NOR2_X1 U8305 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6592), .ZN(n7410) );
  OAI22_X1 U8306 ( .A1(n6595), .A2(n6594), .B1(n6593), .B2(
        P1_REG2_REG_8__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U8307 ( .A1(n6597), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6596) );
  OAI21_X1 U8308 ( .B1(n6597), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6596), .ZN(
        n9937) );
  NOR2_X1 U8309 ( .A1(n9938), .A2(n9937), .ZN(n9936) );
  AOI21_X1 U8310 ( .B1(n6597), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9936), .ZN(
        n6600) );
  NAND2_X1 U8311 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6651), .ZN(n6598) );
  OAI21_X1 U8312 ( .B1(n6651), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6598), .ZN(
        n6599) );
  NOR2_X1 U8313 ( .A1(n6600), .A2(n6599), .ZN(n6650) );
  AOI211_X1 U8314 ( .C1(n6600), .C2(n6599), .A(n6650), .B(n9935), .ZN(n6601)
         );
  AOI211_X1 U8315 ( .C1(n9951), .C2(n6651), .A(n7410), .B(n6601), .ZN(n6602)
         );
  OAI211_X1 U8316 ( .C1(n9964), .C2(n6604), .A(n6603), .B(n6602), .ZN(P1_U3251) );
  INV_X1 U8317 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U8318 ( .A1(P2_U3966), .A2(n6763), .ZN(n6605) );
  OAI21_X1 U8319 ( .B1(P2_U3966), .B2(n6606), .A(n6605), .ZN(P2_U3552) );
  INV_X1 U8320 ( .A(n6607), .ZN(n6609) );
  INV_X1 U8321 ( .A(n6697), .ZN(n6648) );
  OAI222_X1 U8322 ( .A1(n8339), .A2(n6608), .B1(n9537), .B2(n6609), .C1(
        P1_U3084), .C2(n6648), .ZN(P1_U3341) );
  INV_X1 U8323 ( .A(n6985), .ZN(n8149) );
  OAI222_X1 U8324 ( .A1(n8963), .A2(n6610), .B1(n8970), .B2(n6609), .C1(
        P2_U3152), .C2(n8149), .ZN(P2_U3346) );
  OAI21_X1 U8326 ( .B1(n6614), .B2(n6611), .A(n6612), .ZN(n9887) );
  NAND2_X1 U8327 ( .A1(n9887), .A2(n9080), .ZN(n6618) );
  NAND4_X1 U8328 ( .A1(n6616), .A2(n9966), .A3(n6913), .A4(n6615), .ZN(n9061)
         );
  AOI22_X1 U8329 ( .A1(n6480), .A2(n6920), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9061), .ZN(n6617) );
  OAI211_X1 U8330 ( .C1(n6619), .C2(n9070), .A(n6618), .B(n6617), .ZN(P1_U3230) );
  INV_X1 U8331 ( .A(n6620), .ZN(n6641) );
  AOI22_X1 U8332 ( .A1(n6969), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9535), .ZN(n6621) );
  OAI21_X1 U8333 ( .B1(n6641), .B2(n9537), .A(n6621), .ZN(P1_U3340) );
  INV_X1 U8334 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6626) );
  INV_X1 U8335 ( .A(n9405), .ZN(n9348) );
  AND2_X1 U8336 ( .A1(n6376), .A2(n6624), .ZN(n8078) );
  NOR2_X1 U8337 ( .A1(n6711), .A2(n8078), .ZN(n7965) );
  INV_X1 U8338 ( .A(n6917), .ZN(n6622) );
  NOR3_X1 U8339 ( .A1(n7965), .A2(n6622), .A3(n4378), .ZN(n6623) );
  AOI21_X1 U8340 ( .B1(n9348), .B2(n5771), .A(n6623), .ZN(n6923) );
  OAI21_X1 U8341 ( .B1(n6624), .B2(n6917), .A(n6923), .ZN(n6664) );
  NAND2_X1 U8342 ( .A1(n6664), .A2(n9989), .ZN(n6625) );
  OAI21_X1 U8343 ( .B1(n9989), .B2(n6626), .A(n6625), .ZN(P1_U3454) );
  XNOR2_X1 U8344 ( .A(n6628), .B(n6629), .ZN(n6630) );
  XNOR2_X1 U8345 ( .A(n6631), .B(n6630), .ZN(n6634) );
  AOI22_X1 U8346 ( .A1(n6480), .A2(n5774), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n9061), .ZN(n6633) );
  AOI22_X1 U8347 ( .A1(n9062), .A2(n6376), .B1(n9099), .B2(n9127), .ZN(n6632)
         );
  OAI211_X1 U8348 ( .C1(n6634), .C2(n9103), .A(n6633), .B(n6632), .ZN(P1_U3220) );
  INV_X1 U8349 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n6638) );
  INV_X1 U8350 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6635) );
  OR2_X1 U8351 ( .A1(n5805), .A2(n6635), .ZN(n6637) );
  NAND2_X1 U8352 ( .A1(n5878), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6636) );
  OAI211_X1 U8353 ( .C1(n6639), .C2(n6638), .A(n6637), .B(n6636), .ZN(n9192)
         );
  NAND2_X1 U8354 ( .A1(n9192), .A2(P1_U4006), .ZN(n6640) );
  OAI21_X1 U8355 ( .B1(P1_U4006), .B2(n5504), .A(n6640), .ZN(P1_U3586) );
  INV_X1 U8356 ( .A(n7208), .ZN(n7203) );
  OAI222_X1 U8357 ( .A1(n8963), .A2(n6642), .B1(n8973), .B2(n6641), .C1(n7203), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  AOI22_X1 U8358 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6652), .B1(n9145), .B2(
        n5988), .ZN(n9143) );
  OAI21_X1 U8359 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n6651), .A(n6643), .ZN(
        n9142) );
  NAND2_X1 U8360 ( .A1(n9143), .A2(n9142), .ZN(n9141) );
  OAI21_X1 U8361 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6652), .A(n9141), .ZN(
        n6646) );
  MUX2_X1 U8362 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6644), .S(n6697), .Z(n6645)
         );
  NAND2_X1 U8363 ( .A1(n6645), .A2(n6646), .ZN(n6693) );
  OAI21_X1 U8364 ( .B1(n6646), .B2(n6645), .A(n6693), .ZN(n6658) );
  NAND2_X1 U8365 ( .A1(n9866), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6647) );
  NAND2_X1 U8366 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7641) );
  OAI211_X1 U8367 ( .C1(n9943), .C2(n6648), .A(n6647), .B(n7641), .ZN(n6657)
         );
  NOR2_X1 U8368 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6652), .ZN(n6649) );
  AOI21_X1 U8369 ( .B1(n6652), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6649), .ZN(
        n9150) );
  AOI21_X1 U8370 ( .B1(n6651), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6650), .ZN(
        n9149) );
  NAND2_X1 U8371 ( .A1(n9150), .A2(n9149), .ZN(n9148) );
  OAI21_X1 U8372 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6652), .A(n9148), .ZN(
        n6655) );
  NAND2_X1 U8373 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6697), .ZN(n6653) );
  OAI21_X1 U8374 ( .B1(n6697), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6653), .ZN(
        n6654) );
  NOR2_X1 U8375 ( .A1(n6654), .A2(n6655), .ZN(n6696) );
  AOI211_X1 U8376 ( .C1(n6655), .C2(n6654), .A(n6696), .B(n9935), .ZN(n6656)
         );
  AOI211_X1 U8377 ( .C1(n6658), .C2(n9959), .A(n6657), .B(n6656), .ZN(n6659)
         );
  INV_X1 U8378 ( .A(n6659), .ZN(P1_U3253) );
  INV_X1 U8379 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6661) );
  INV_X1 U8380 ( .A(n6660), .ZN(n6662) );
  INV_X1 U8381 ( .A(n8508), .ZN(n7206) );
  OAI222_X1 U8382 ( .A1(n8963), .A2(n6661), .B1(n8973), .B2(n6662), .C1(n7206), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8383 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6663) );
  INV_X1 U8384 ( .A(n7380), .ZN(n7374) );
  OAI222_X1 U8385 ( .A1(n8339), .A2(n6663), .B1(n9537), .B2(n6662), .C1(n7374), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  NAND2_X1 U8386 ( .A1(n6664), .A2(n9994), .ZN(n6665) );
  OAI21_X1 U8387 ( .B1(n9994), .B2(n9867), .A(n6665), .ZN(P1_U3523) );
  NAND2_X1 U8388 ( .A1(n6668), .A2(n6667), .ZN(n6669) );
  XOR2_X1 U8389 ( .A(n6666), .B(n6669), .Z(n6674) );
  AOI22_X1 U8390 ( .A1(n9062), .A2(n9127), .B1(n9099), .B2(n9125), .ZN(n6673)
         );
  INV_X1 U8391 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7337) );
  NAND2_X1 U8392 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9774) );
  INV_X1 U8393 ( .A(n9774), .ZN(n6671) );
  NOR2_X1 U8394 ( .A1(n9087), .A2(n9969), .ZN(n6670) );
  AOI211_X1 U8395 ( .C1(n7337), .C2(n9082), .A(n6671), .B(n6670), .ZN(n6672)
         );
  OAI211_X1 U8396 ( .C1(n6674), .C2(n9103), .A(n6673), .B(n6672), .ZN(P1_U3216) );
  NAND2_X1 U8397 ( .A1(n6676), .A2(n7964), .ZN(n6677) );
  NAND2_X1 U8398 ( .A1(n6675), .A2(n6677), .ZN(n7330) );
  OAI21_X1 U8399 ( .B1(n5774), .B2(n6920), .A(n4839), .ZN(n6678) );
  NAND3_X1 U8400 ( .A1(n6678), .A2(n9228), .A3(n7334), .ZN(n7326) );
  INV_X1 U8401 ( .A(n7326), .ZN(n6684) );
  NAND2_X1 U8402 ( .A1(n7330), .A2(n9824), .ZN(n6683) );
  OAI21_X1 U8403 ( .B1(n7964), .B2(n8086), .A(n6679), .ZN(n6680) );
  NAND2_X1 U8404 ( .A1(n6680), .A2(n9351), .ZN(n6682) );
  AOI22_X1 U8405 ( .A1(n9346), .A2(n5771), .B1(n9126), .B2(n9348), .ZN(n6681)
         );
  NAND3_X1 U8406 ( .A1(n6683), .A2(n6682), .A3(n6681), .ZN(n7327) );
  AOI211_X1 U8407 ( .C1(n9973), .C2(n7330), .A(n6684), .B(n7327), .ZN(n6842)
         );
  INV_X1 U8408 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6685) );
  OAI22_X1 U8409 ( .A1(n9529), .A2(n6839), .B1(n9989), .B2(n6685), .ZN(n6686)
         );
  INV_X1 U8410 ( .A(n6686), .ZN(n6687) );
  OAI21_X1 U8411 ( .B1(n6842), .B2(n9988), .A(n6687), .ZN(P1_U3460) );
  INV_X1 U8412 ( .A(n6688), .ZN(n6690) );
  OAI222_X1 U8413 ( .A1(n8339), .A2(n6689), .B1(n9537), .B2(n6690), .C1(
        P1_U3084), .C2(n7501), .ZN(P1_U3338) );
  INV_X1 U8414 ( .A(n8526), .ZN(n8520) );
  OAI222_X1 U8415 ( .A1(n8963), .A2(n6691), .B1(n8973), .B2(n6690), .C1(
        P2_U3152), .C2(n8520), .ZN(P2_U3343) );
  INV_X1 U8416 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8417 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6692), .S(n6969), .Z(n6695)
         );
  OAI21_X1 U8418 ( .B1(n6697), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6693), .ZN(
        n6694) );
  NAND2_X1 U8419 ( .A1(n6695), .A2(n6694), .ZN(n6965) );
  OAI21_X1 U8420 ( .B1(n6695), .B2(n6694), .A(n6965), .ZN(n6702) );
  MUX2_X1 U8421 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n9822), .S(n6969), .Z(n6698)
         );
  INV_X1 U8422 ( .A(n6698), .ZN(n6699) );
  AOI211_X1 U8423 ( .C1(n6700), .C2(n6699), .A(n6968), .B(n9935), .ZN(n6701)
         );
  AOI21_X1 U8424 ( .B1(n9959), .B2(n6702), .A(n6701), .ZN(n6704) );
  AND2_X1 U8425 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7678) );
  AOI21_X1 U8426 ( .B1(n9951), .B2(n6969), .A(n7678), .ZN(n6703) );
  OAI211_X1 U8427 ( .C1(n9964), .C2(n6705), .A(n6704), .B(n6703), .ZN(P1_U3254) );
  OR2_X1 U8428 ( .A1(n6707), .A2(n6706), .ZN(n6708) );
  NAND2_X1 U8429 ( .A1(n6709), .A2(n6708), .ZN(n7080) );
  INV_X1 U8430 ( .A(n9973), .ZN(n6718) );
  OAI21_X1 U8431 ( .B1(n7967), .B2(n6711), .A(n6710), .ZN(n6716) );
  INV_X1 U8432 ( .A(n6376), .ZN(n6712) );
  OAI22_X1 U8433 ( .A1(n6712), .A2(n9403), .B1(n4748), .B2(n9405), .ZN(n6715)
         );
  INV_X1 U8434 ( .A(n9824), .ZN(n6713) );
  NOR2_X1 U8435 ( .A1(n7080), .A2(n6713), .ZN(n6714) );
  AOI211_X1 U8436 ( .C1(n9351), .C2(n6716), .A(n6715), .B(n6714), .ZN(n7083)
         );
  XNOR2_X1 U8437 ( .A(n8079), .B(n6920), .ZN(n6717) );
  NAND2_X1 U8438 ( .A1(n6717), .A2(n9228), .ZN(n7075) );
  OAI211_X1 U8439 ( .C1(n7080), .C2(n6718), .A(n7083), .B(n7075), .ZN(n6844)
         );
  INV_X1 U8440 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6719) );
  OAI22_X1 U8441 ( .A1(n9529), .A2(n8079), .B1(n9989), .B2(n6719), .ZN(n6720)
         );
  AOI21_X1 U8442 ( .B1(n6844), .B2(n9989), .A(n6720), .ZN(n6721) );
  INV_X1 U8443 ( .A(n6721), .ZN(P1_U3457) );
  OAI211_X1 U8444 ( .C1(n6724), .C2(n6723), .A(n6769), .B(n9080), .ZN(n6729)
         );
  INV_X1 U8445 ( .A(n6725), .ZN(n7086) );
  NAND2_X1 U8446 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n9905) );
  OAI21_X1 U8447 ( .B1(n9087), .B2(n7089), .A(n9905), .ZN(n6727) );
  INV_X1 U8448 ( .A(n9126), .ZN(n6892) );
  INV_X1 U8449 ( .A(n9124), .ZN(n7003) );
  OAI22_X1 U8450 ( .A1(n6892), .A2(n9094), .B1(n9070), .B2(n7003), .ZN(n6726)
         );
  AOI211_X1 U8451 ( .C1(n7086), .C2(n9082), .A(n6727), .B(n6726), .ZN(n6728)
         );
  NAND2_X1 U8452 ( .A1(n6729), .A2(n6728), .ZN(P1_U3228) );
  NAND2_X1 U8453 ( .A1(n6730), .A2(n8295), .ZN(n6732) );
  NAND2_X1 U8454 ( .A1(n6731), .A2(n8257), .ZN(n6933) );
  NAND2_X1 U8455 ( .A1(n6732), .A2(n6733), .ZN(n6857) );
  NAND2_X1 U8456 ( .A1(n6857), .A2(n6734), .ZN(n6737) );
  NAND2_X1 U8457 ( .A1(n6763), .A2(n7158), .ZN(n7046) );
  INV_X1 U8458 ( .A(n6858), .ZN(n6735) );
  AOI21_X1 U8459 ( .B1(n6737), .B2(n6736), .A(n6735), .ZN(n6767) );
  INV_X1 U8460 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10009) );
  NOR2_X1 U8461 ( .A1(n6739), .A2(n7801), .ZN(n10010) );
  NOR4_X1 U8462 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6743) );
  NOR4_X1 U8463 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6742) );
  NOR4_X1 U8464 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6741) );
  NOR4_X1 U8465 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n6740) );
  NAND4_X1 U8466 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6749)
         );
  NOR2_X1 U8467 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n6747) );
  NOR4_X1 U8468 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n6746) );
  NOR4_X1 U8469 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6745) );
  NOR4_X1 U8470 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6744) );
  NAND4_X1 U8471 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6748)
         );
  INV_X1 U8472 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10012) );
  NOR2_X1 U8473 ( .A1(n7746), .A2(n7801), .ZN(n10014) );
  INV_X1 U8474 ( .A(n10008), .ZN(n6751) );
  INV_X1 U8475 ( .A(n6760), .ZN(n6752) );
  NOR2_X1 U8476 ( .A1(n10088), .A2(n6753), .ZN(n6754) );
  NOR2_X1 U8477 ( .A1(n10016), .A2(n8257), .ZN(n6946) );
  AND2_X1 U8478 ( .A1(n10008), .A2(n6946), .ZN(n6755) );
  NAND2_X1 U8479 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  INV_X1 U8480 ( .A(n7180), .ZN(n6758) );
  NAND2_X1 U8481 ( .A1(n6759), .A2(n6758), .ZN(n6880) );
  INV_X1 U8482 ( .A(n7181), .ZN(n6930) );
  NAND2_X1 U8483 ( .A1(n6880), .A2(n6930), .ZN(n6926) );
  AOI22_X1 U8484 ( .A1(n7054), .A2(n8459), .B1(n6926), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U8485 ( .A1(n6763), .A2(n8804), .ZN(n6764) );
  OAI21_X1 U8486 ( .B1(n8256), .B2(n8838), .A(n6764), .ZN(n7047) );
  NAND2_X1 U8487 ( .A1(n8335), .A2(n7047), .ZN(n6765) );
  OAI211_X1 U8488 ( .C1(n6767), .C2(n8477), .A(n6766), .B(n6765), .ZN(P2_U3224) );
  NAND2_X1 U8489 ( .A1(n6769), .A2(n6768), .ZN(n6773) );
  XNOR2_X1 U8490 ( .A(n6771), .B(n6770), .ZN(n6772) );
  XNOR2_X1 U8491 ( .A(n6773), .B(n6772), .ZN(n6777) );
  AOI22_X1 U8492 ( .A1(n9062), .A2(n9125), .B1(n9099), .B2(n9123), .ZN(n6776)
         );
  AND2_X1 U8493 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9917) );
  NOR2_X1 U8494 ( .A1(n9096), .A2(n7228), .ZN(n6774) );
  AOI211_X1 U8495 ( .C1(n4509), .C2(n6480), .A(n9917), .B(n6774), .ZN(n6775)
         );
  OAI211_X1 U8496 ( .C1(n6777), .C2(n9103), .A(n6776), .B(n6775), .ZN(P1_U3225) );
  INV_X1 U8497 ( .A(n6778), .ZN(n6855) );
  AOI22_X1 U8498 ( .A1(n9175), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9535), .ZN(n6779) );
  OAI21_X1 U8499 ( .B1(n6855), .B2(n9537), .A(n6779), .ZN(P1_U3336) );
  NAND2_X1 U8500 ( .A1(n6825), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6792) );
  MUX2_X1 U8501 ( .A(n5130), .B(P2_REG2_REG_10__SCAN_IN), .S(n6825), .Z(n6780)
         );
  INV_X1 U8502 ( .A(n6780), .ZN(n8156) );
  NAND2_X1 U8503 ( .A1(n6823), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6791) );
  MUX2_X1 U8504 ( .A(n5111), .B(P2_REG2_REG_9__SCAN_IN), .S(n6823), .Z(n6781)
         );
  INV_X1 U8505 ( .A(n6781), .ZN(n8168) );
  MUX2_X1 U8506 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6782), .S(n6821), .Z(n8178)
         );
  MUX2_X1 U8507 ( .A(n7170), .B(P2_REG2_REG_7__SCAN_IN), .S(n8193), .Z(n8189)
         );
  NAND2_X1 U8508 ( .A1(n6818), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6790) );
  MUX2_X1 U8509 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6783), .S(n6818), .Z(n8200)
         );
  NAND2_X1 U8510 ( .A1(n6816), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6789) );
  MUX2_X1 U8511 ( .A(n7134), .B(P2_REG2_REG_5__SCAN_IN), .S(n6816), .Z(n6784)
         );
  INV_X1 U8512 ( .A(n6784), .ZN(n8212) );
  MUX2_X1 U8513 ( .A(n6785), .B(P2_REG2_REG_4__SCAN_IN), .S(n8226), .Z(n8222)
         );
  MUX2_X1 U8514 ( .A(n6786), .B(P2_REG2_REG_3__SCAN_IN), .S(n8237), .Z(n8233)
         );
  INV_X1 U8515 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6788) );
  INV_X1 U8516 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7052) );
  MUX2_X1 U8517 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7052), .S(n8248), .Z(n6787)
         );
  INV_X1 U8518 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10005) );
  OR3_X1 U8519 ( .A1(n6787), .A2(n9996), .A3(n10005), .ZN(n8243) );
  OAI21_X1 U8520 ( .B1(n7052), .B2(n8248), .A(n8243), .ZN(n9784) );
  MUX2_X1 U8521 ( .A(n6788), .B(P2_REG2_REG_2__SCAN_IN), .S(n6810), .Z(n9783)
         );
  NAND2_X1 U8522 ( .A1(n9784), .A2(n9783), .ZN(n9782) );
  OAI21_X1 U8523 ( .B1(n6788), .B2(n6810), .A(n9782), .ZN(n8234) );
  NAND2_X1 U8524 ( .A1(n8233), .A2(n8234), .ZN(n8232) );
  OAI21_X1 U8525 ( .B1(n8237), .B2(n6786), .A(n8232), .ZN(n8223) );
  NAND2_X1 U8526 ( .A1(n8222), .A2(n8223), .ZN(n8221) );
  OAI21_X1 U8527 ( .B1(n8226), .B2(n6785), .A(n8221), .ZN(n8211) );
  NAND2_X1 U8528 ( .A1(n8212), .A2(n8211), .ZN(n8210) );
  NAND2_X1 U8529 ( .A1(n6789), .A2(n8210), .ZN(n8201) );
  NAND2_X1 U8530 ( .A1(n8200), .A2(n8201), .ZN(n8199) );
  NAND2_X1 U8531 ( .A1(n6790), .A2(n8199), .ZN(n8190) );
  NAND2_X1 U8532 ( .A1(n8189), .A2(n8190), .ZN(n8188) );
  OAI21_X1 U8533 ( .B1(n8193), .B2(n7170), .A(n8188), .ZN(n8179) );
  NAND2_X1 U8534 ( .A1(n8178), .A2(n8179), .ZN(n8177) );
  OAI21_X1 U8535 ( .B1(n8182), .B2(n6782), .A(n8177), .ZN(n8167) );
  NAND2_X1 U8536 ( .A1(n8168), .A2(n8167), .ZN(n8166) );
  NAND2_X1 U8537 ( .A1(n6791), .A2(n8166), .ZN(n8157) );
  NAND2_X1 U8538 ( .A1(n8156), .A2(n8157), .ZN(n8155) );
  NAND2_X1 U8539 ( .A1(n6792), .A2(n8155), .ZN(n6795) );
  MUX2_X1 U8540 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n5148), .S(n6983), .Z(n6793)
         );
  INV_X1 U8541 ( .A(n6793), .ZN(n6794) );
  NOR2_X1 U8542 ( .A1(n6795), .A2(n6794), .ZN(n6977) );
  AOI21_X1 U8543 ( .B1(n6795), .B2(n6794), .A(n6977), .ZN(n6834) );
  NOR2_X1 U8544 ( .A1(n6803), .A2(P2_U3152), .ZN(n8967) );
  AOI21_X1 U8545 ( .B1(n6796), .B2(n8967), .A(n5684), .ZN(n6799) );
  NAND2_X1 U8546 ( .A1(n10008), .A2(n6797), .ZN(n6798) );
  NAND2_X1 U8547 ( .A1(n6799), .A2(n6798), .ZN(n6806) );
  NAND2_X1 U8548 ( .A1(n6806), .A2(n6804), .ZN(n6800) );
  NAND2_X1 U8549 ( .A1(n6800), .A2(n8492), .ZN(n6802) );
  NOR2_X1 U8550 ( .A1(n6803), .A2(n8971), .ZN(n6801) );
  NOR2_X1 U8551 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5145), .ZN(n8458) );
  AOI21_X1 U8552 ( .B1(n10002), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8458), .ZN(
        n6830) );
  AND2_X1 U8553 ( .A1(n6804), .A2(n8971), .ZN(n6805) );
  INV_X1 U8554 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6807) );
  MUX2_X1 U8555 ( .A(n6807), .B(P2_REG1_REG_11__SCAN_IN), .S(n6983), .Z(n6827)
         );
  INV_X1 U8556 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6819) );
  INV_X1 U8557 ( .A(n8237), .ZN(n6813) );
  INV_X1 U8558 ( .A(n6810), .ZN(n9780) );
  INV_X1 U8559 ( .A(n8248), .ZN(n6809) );
  INV_X1 U8560 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6808) );
  INV_X1 U8561 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10105) );
  INV_X1 U8562 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6811) );
  MUX2_X1 U8563 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6811), .S(n6810), .Z(n9777)
         );
  NOR2_X1 U8564 ( .A1(n9778), .A2(n9777), .ZN(n9776) );
  AOI21_X1 U8565 ( .B1(P2_REG1_REG_2__SCAN_IN), .B2(n9780), .A(n9776), .ZN(
        n8229) );
  INV_X1 U8566 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6812) );
  MUX2_X1 U8567 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6812), .S(n8237), .Z(n8228)
         );
  INV_X1 U8568 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6814) );
  MUX2_X1 U8569 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6814), .S(n8226), .Z(n8217)
         );
  NAND2_X1 U8570 ( .A1(n6816), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6815) );
  OAI21_X1 U8571 ( .B1(n6816), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6815), .ZN(
        n8206) );
  NOR2_X1 U8572 ( .A1(n8207), .A2(n8206), .ZN(n8205) );
  AOI21_X1 U8573 ( .B1(n6816), .B2(P2_REG1_REG_5__SCAN_IN), .A(n8205), .ZN(
        n8196) );
  NAND2_X1 U8574 ( .A1(n6818), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6817) );
  OAI21_X1 U8575 ( .B1(n6818), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6817), .ZN(
        n8195) );
  NOR2_X1 U8576 ( .A1(n8196), .A2(n8195), .ZN(n8194) );
  MUX2_X1 U8577 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6819), .S(n8193), .Z(n8184)
         );
  INV_X1 U8578 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6820) );
  MUX2_X1 U8579 ( .A(n6820), .B(P2_REG1_REG_8__SCAN_IN), .S(n6821), .Z(n8173)
         );
  INV_X1 U8580 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6822) );
  MUX2_X1 U8581 ( .A(n6822), .B(P2_REG1_REG_9__SCAN_IN), .S(n6823), .Z(n8162)
         );
  NOR2_X1 U8582 ( .A1(n8163), .A2(n8162), .ZN(n8161) );
  AOI21_X1 U8583 ( .B1(n6823), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8161), .ZN(
        n8152) );
  INV_X1 U8584 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6824) );
  MUX2_X1 U8585 ( .A(n6824), .B(P2_REG1_REG_10__SCAN_IN), .S(n6825), .Z(n8151)
         );
  AOI21_X1 U8586 ( .B1(n6827), .B2(n6826), .A(n6982), .ZN(n6828) );
  NAND2_X1 U8587 ( .A1(n9995), .A2(n6828), .ZN(n6829) );
  OAI211_X1 U8588 ( .C1(n9998), .C2(n6831), .A(n6830), .B(n6829), .ZN(n6832)
         );
  INV_X1 U8589 ( .A(n6832), .ZN(n6833) );
  OAI21_X1 U8590 ( .B1(n6834), .B2(n8578), .A(n6833), .ZN(P2_U3256) );
  INV_X1 U8591 ( .A(n6835), .ZN(n6838) );
  OAI222_X1 U8592 ( .A1(P2_U3152), .A2(n8545), .B1(n8973), .B2(n6838), .C1(
        n6836), .C2(n8963), .ZN(P2_U3342) );
  INV_X1 U8593 ( .A(n9160), .ZN(n7509) );
  OAI222_X1 U8594 ( .A1(P1_U3084), .A2(n7509), .B1(n9537), .B2(n6838), .C1(
        n6837), .C2(n8339), .ZN(P1_U3337) );
  OAI22_X1 U8595 ( .A1(n9491), .A2(n6839), .B1(n9994), .B2(n6547), .ZN(n6840)
         );
  INV_X1 U8596 ( .A(n6840), .ZN(n6841) );
  OAI21_X1 U8597 ( .B1(n6842), .B2(n9992), .A(n6841), .ZN(P1_U3525) );
  OAI22_X1 U8598 ( .A1(n9491), .A2(n8079), .B1(n9994), .B2(n6545), .ZN(n6843)
         );
  AOI21_X1 U8599 ( .B1(n6844), .B2(n9994), .A(n6843), .ZN(n6845) );
  INV_X1 U8600 ( .A(n6845), .ZN(P1_U3524) );
  XOR2_X1 U8601 ( .A(n6848), .B(n6847), .Z(n6849) );
  XNOR2_X1 U8602 ( .A(n6846), .B(n6849), .ZN(n6854) );
  AOI22_X1 U8603 ( .A1(n9099), .A2(n9122), .B1(n6480), .B2(n9413), .ZN(n6853)
         );
  NOR2_X1 U8604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6850), .ZN(n9128) );
  NOR2_X1 U8605 ( .A1(n9096), .A2(n9411), .ZN(n6851) );
  AOI211_X1 U8606 ( .C1(n9062), .C2(n9124), .A(n9128), .B(n6851), .ZN(n6852)
         );
  OAI211_X1 U8607 ( .C1(n6854), .C2(n9103), .A(n6853), .B(n6852), .ZN(P1_U3237) );
  INV_X1 U8608 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6856) );
  INV_X1 U8609 ( .A(n8559), .ZN(n8556) );
  OAI222_X1 U8610 ( .A1(n8963), .A2(n6856), .B1(n8973), .B2(n6855), .C1(n8556), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  NAND2_X1 U8611 ( .A1(n8505), .A2(n8309), .ZN(n6860) );
  XNOR2_X1 U8612 ( .A(n7069), .B(n8308), .ZN(n6861) );
  XNOR2_X1 U8613 ( .A(n6860), .B(n6861), .ZN(n6899) );
  INV_X1 U8614 ( .A(n6860), .ZN(n6863) );
  INV_X1 U8615 ( .A(n6861), .ZN(n6862) );
  NAND2_X1 U8616 ( .A1(n6863), .A2(n6862), .ZN(n6864) );
  NAND2_X1 U8617 ( .A1(n8504), .A2(n8295), .ZN(n6865) );
  XNOR2_X1 U8618 ( .A(n4996), .B(n8318), .ZN(n6866) );
  XNOR2_X1 U8619 ( .A(n6865), .B(n6866), .ZN(n8249) );
  INV_X1 U8620 ( .A(n6865), .ZN(n6867) );
  AND2_X1 U8621 ( .A1(n6867), .A2(n6866), .ZN(n6868) );
  NAND2_X1 U8622 ( .A1(n8503), .A2(n8309), .ZN(n6869) );
  XNOR2_X1 U8623 ( .A(n5033), .B(n8308), .ZN(n6870) );
  NAND2_X1 U8624 ( .A1(n6869), .A2(n6870), .ZN(n6874) );
  INV_X1 U8625 ( .A(n6869), .ZN(n6872) );
  INV_X1 U8626 ( .A(n6870), .ZN(n6871) );
  NAND2_X1 U8627 ( .A1(n6872), .A2(n6871), .ZN(n6873) );
  AND2_X1 U8628 ( .A1(n6874), .A2(n6873), .ZN(n6906) );
  XNOR2_X1 U8629 ( .A(n7148), .B(n8318), .ZN(n7021) );
  NAND2_X1 U8630 ( .A1(n8502), .A2(n8309), .ZN(n7020) );
  XNOR2_X1 U8631 ( .A(n7021), .B(n7020), .ZN(n7018) );
  XNOR2_X1 U8632 ( .A(n7019), .B(n7018), .ZN(n6886) );
  INV_X1 U8633 ( .A(n7123), .ZN(n6884) );
  INV_X1 U8634 ( .A(n6875), .ZN(n6877) );
  AND3_X1 U8635 ( .A1(n6878), .A2(n6877), .A3(n6876), .ZN(n6879) );
  NAND2_X1 U8636 ( .A1(n6880), .A2(n6879), .ZN(n6881) );
  INV_X1 U8637 ( .A(n8335), .ZN(n8406) );
  AOI22_X1 U8638 ( .A1(n8804), .A2(n8503), .B1(n8501), .B2(n8806), .ZN(n7132)
         );
  AOI22_X1 U8639 ( .A1(n8459), .A2(n7189), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6882) );
  OAI21_X1 U8640 ( .B1(n8406), .B2(n7132), .A(n6882), .ZN(n6883) );
  AOI21_X1 U8641 ( .B1(n6884), .B2(n8472), .A(n6883), .ZN(n6885) );
  OAI21_X1 U8642 ( .B1(n6886), .B2(n8477), .A(n6885), .ZN(P2_U3229) );
  OAI21_X1 U8643 ( .B1(n6888), .B2(n6890), .A(n6887), .ZN(n7091) );
  AOI211_X1 U8644 ( .C1(n6889), .C2(n7335), .A(n9390), .B(n7227), .ZN(n7085)
         );
  XNOR2_X1 U8645 ( .A(n7822), .B(n6890), .ZN(n6891) );
  OAI222_X1 U8646 ( .A1(n9405), .A2(n7003), .B1(n9403), .B2(n6892), .C1(n6891), 
        .C2(n9400), .ZN(n7084) );
  AOI211_X1 U8647 ( .C1(n9986), .C2(n7091), .A(n7085), .B(n7084), .ZN(n6898)
         );
  INV_X1 U8648 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6893) );
  OAI22_X1 U8649 ( .A1(n9529), .A2(n7089), .B1(n9989), .B2(n6893), .ZN(n6894)
         );
  INV_X1 U8650 ( .A(n6894), .ZN(n6895) );
  OAI21_X1 U8651 ( .B1(n6898), .B2(n9988), .A(n6895), .ZN(P1_U3466) );
  OAI22_X1 U8652 ( .A1(n9491), .A2(n7089), .B1(n9994), .B2(n5833), .ZN(n6896)
         );
  INV_X1 U8653 ( .A(n6896), .ZN(n6897) );
  OAI21_X1 U8654 ( .B1(n6898), .B2(n9992), .A(n6897), .ZN(P1_U3527) );
  XNOR2_X1 U8655 ( .A(n6900), .B(n6899), .ZN(n6903) );
  AOI22_X1 U8656 ( .A1(n8461), .A2(n6730), .B1(n8460), .B2(n8504), .ZN(n6902)
         );
  AOI22_X1 U8657 ( .A1(n7069), .A2(n8459), .B1(n6926), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6901) );
  OAI211_X1 U8658 ( .C1(n6903), .C2(n8477), .A(n6902), .B(n6901), .ZN(P2_U3239) );
  OAI21_X1 U8659 ( .B1(n6906), .B2(n6905), .A(n6904), .ZN(n6909) );
  INV_X1 U8660 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n9671) );
  NOR2_X1 U8661 ( .A1(n9671), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8220) );
  INV_X1 U8662 ( .A(n8220), .ZN(n6907) );
  OAI21_X1 U8663 ( .B1(n8490), .B2(n10044), .A(n6907), .ZN(n6908) );
  AOI21_X1 U8664 ( .B1(n8441), .B2(n6909), .A(n6908), .ZN(n6912) );
  INV_X1 U8665 ( .A(n6910), .ZN(n6948) );
  AOI22_X1 U8666 ( .A1(n8460), .A2(n8502), .B1(n8472), .B2(n6948), .ZN(n6911)
         );
  OAI211_X1 U8667 ( .C1(n7063), .C2(n8485), .A(n6912), .B(n6911), .ZN(P2_U3232) );
  NAND3_X1 U8668 ( .A1(n6915), .A2(n6914), .A3(n6913), .ZN(n7038) );
  INV_X1 U8669 ( .A(n9397), .ZN(n7231) );
  OAI21_X1 U8670 ( .B1(n7231), .B2(n6917), .A(n9392), .ZN(n6921) );
  OAI22_X1 U8671 ( .A1(n9409), .A2(n5717), .B1(n6918), .B2(n9820), .ZN(n6919)
         );
  AOI21_X1 U8672 ( .B1(n6921), .B2(n6920), .A(n6919), .ZN(n6922) );
  OAI21_X1 U8673 ( .B1(n6923), .B2(n9826), .A(n6922), .ZN(P1_U3291) );
  INV_X1 U8674 ( .A(n5519), .ZN(n6924) );
  AOI21_X1 U8675 ( .B1(n7158), .B2(n8319), .A(n6924), .ZN(n6929) );
  INV_X1 U8676 ( .A(n8475), .ZN(n8439) );
  AOI22_X1 U8677 ( .A1(n6925), .A2(n8439), .B1(n8460), .B2(n6730), .ZN(n6928)
         );
  AOI22_X1 U8678 ( .A1(n7158), .A2(n8459), .B1(n6926), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n6927) );
  OAI211_X1 U8679 ( .C1(n6929), .C2(n8477), .A(n6928), .B(n6927), .ZN(P2_U3234) );
  INV_X1 U8680 ( .A(n7196), .ZN(n6931) );
  NAND4_X1 U8681 ( .A1(n6931), .A2(n7194), .A3(n7183), .A4(n6930), .ZN(n7057)
         );
  NOR2_X1 U8682 ( .A1(n6933), .A2(n8828), .ZN(n6932) );
  XNOR2_X1 U8683 ( .A(n6934), .B(n6933), .ZN(n8821) );
  NAND2_X1 U8684 ( .A1(n8821), .A2(n8828), .ZN(n8845) );
  INV_X1 U8685 ( .A(n8845), .ZN(n7664) );
  NAND2_X1 U8686 ( .A1(n8831), .A2(n7664), .ZN(n6935) );
  NAND2_X1 U8687 ( .A1(n6936), .A2(n7046), .ZN(n6938) );
  NAND2_X1 U8688 ( .A1(n4316), .A2(n10024), .ZN(n6937) );
  NAND2_X1 U8689 ( .A1(n6938), .A2(n6937), .ZN(n7056) );
  NAND2_X1 U8690 ( .A1(n7056), .A2(n7060), .ZN(n6940) );
  NAND2_X1 U8691 ( .A1(n8256), .A2(n10032), .ZN(n6939) );
  NAND2_X1 U8692 ( .A1(n6940), .A2(n6939), .ZN(n7112) );
  NAND2_X1 U8693 ( .A1(n7112), .A2(n7110), .ZN(n6941) );
  NAND2_X1 U8694 ( .A1(n7063), .A2(n10037), .ZN(n7114) );
  NAND2_X1 U8695 ( .A1(n6941), .A2(n7114), .ZN(n6942) );
  XOR2_X1 U8696 ( .A(n7113), .B(n6942), .Z(n10042) );
  XNOR2_X1 U8697 ( .A(n7127), .B(n7113), .ZN(n6945) );
  OAI222_X1 U8698 ( .A1(n8838), .A2(n7149), .B1(n8840), .B2(n7063), .C1(n6945), 
        .C2(n8817), .ZN(n10046) );
  NOR2_X1 U8699 ( .A1(n8831), .A2(n6785), .ZN(n6951) );
  INV_X1 U8700 ( .A(n7057), .ZN(n6947) );
  NAND2_X1 U8701 ( .A1(n7094), .A2(n10037), .ZN(n7120) );
  XNOR2_X1 U8702 ( .A(n7120), .B(n10044), .ZN(n10043) );
  INV_X1 U8703 ( .A(n8852), .ZN(n8797) );
  AOI22_X1 U8704 ( .A1(n8856), .A2(n10043), .B1(n6948), .B2(n8797), .ZN(n6949)
         );
  OAI21_X1 U8705 ( .B1(n10044), .B2(n8800), .A(n6949), .ZN(n6950) );
  AOI211_X1 U8706 ( .C1(n8831), .C2(n10046), .A(n6951), .B(n6950), .ZN(n6952)
         );
  OAI21_X1 U8707 ( .B1(n8812), .B2(n10042), .A(n6952), .ZN(P2_U3292) );
  NAND2_X1 U8708 ( .A1(n6955), .A2(n6954), .ZN(n6956) );
  XNOR2_X1 U8709 ( .A(n6957), .B(n6956), .ZN(n6958) );
  NAND2_X1 U8710 ( .A1(n6958), .A2(n9080), .ZN(n6963) );
  INV_X1 U8711 ( .A(n6959), .ZN(n6961) );
  INV_X1 U8712 ( .A(n9123), .ZN(n7035) );
  OAI22_X1 U8713 ( .A1(n9096), .A2(n7039), .B1(n9094), .B2(n7035), .ZN(n6960)
         );
  AOI211_X1 U8714 ( .C1(n9099), .C2(n9121), .A(n6961), .B(n6960), .ZN(n6962)
         );
  OAI211_X1 U8715 ( .C1(n7352), .C2(n9087), .A(n6963), .B(n6962), .ZN(P1_U3211) );
  INV_X1 U8716 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6975) );
  MUX2_X1 U8717 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6964), .S(n7380), .Z(n6967)
         );
  OAI21_X1 U8718 ( .B1(n6969), .B2(P1_REG1_REG_13__SCAN_IN), .A(n6965), .ZN(
        n6966) );
  NAND2_X1 U8719 ( .A1(n6967), .A2(n6966), .ZN(n7379) );
  OAI21_X1 U8720 ( .B1(n6967), .B2(n6966), .A(n7379), .ZN(n6972) );
  NOR2_X1 U8721 ( .A1(n7728), .A2(n6970), .ZN(n7376) );
  AOI211_X1 U8722 ( .C1(n6970), .C2(n7728), .A(n7376), .B(n9935), .ZN(n6971)
         );
  AOI21_X1 U8723 ( .B1(n9959), .B2(n6972), .A(n6971), .ZN(n6974) );
  AND2_X1 U8724 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7796) );
  AOI21_X1 U8725 ( .B1(n9951), .B2(n7380), .A(n7796), .ZN(n6973) );
  OAI211_X1 U8726 ( .C1(n9964), .C2(n6975), .A(n6974), .B(n6973), .ZN(P1_U3255) );
  NAND2_X1 U8727 ( .A1(n6985), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6979) );
  MUX2_X1 U8728 ( .A(n7530), .B(P2_REG2_REG_12__SCAN_IN), .S(n6985), .Z(n6976)
         );
  INV_X1 U8729 ( .A(n6976), .ZN(n8138) );
  NOR2_X1 U8730 ( .A1(n6983), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6978) );
  NOR2_X1 U8731 ( .A1(n6978), .A2(n6977), .ZN(n8139) );
  NAND2_X1 U8732 ( .A1(n8138), .A2(n8139), .ZN(n8137) );
  NAND2_X1 U8733 ( .A1(n6979), .A2(n8137), .ZN(n6981) );
  AOI22_X1 U8734 ( .A1(n7208), .A2(n5188), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7203), .ZN(n6980) );
  NOR2_X1 U8735 ( .A1(n6981), .A2(n6980), .ZN(n7202) );
  AOI21_X1 U8736 ( .B1(n6981), .B2(n6980), .A(n7202), .ZN(n6994) );
  AOI22_X1 U8737 ( .A1(n7208), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5185), .B2(
        n7203), .ZN(n6987) );
  MUX2_X1 U8738 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n6984), .S(n6985), .Z(n8142)
         );
  NAND2_X1 U8739 ( .A1(n8141), .A2(n8142), .ZN(n8140) );
  OAI21_X1 U8740 ( .B1(n6987), .B2(n6986), .A(n7207), .ZN(n6988) );
  NAND2_X1 U8741 ( .A1(n6988), .A2(n9995), .ZN(n6993) );
  INV_X1 U8742 ( .A(n9998), .ZN(n9781) );
  INV_X1 U8743 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n6990) );
  OAI22_X1 U8744 ( .A1(n8587), .A2(n6990), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6989), .ZN(n6991) );
  AOI21_X1 U8745 ( .B1(n9781), .B2(n7208), .A(n6991), .ZN(n6992) );
  OAI211_X1 U8746 ( .C1(n6994), .C2(n8578), .A(n6993), .B(n6992), .ZN(P2_U3258) );
  INV_X1 U8747 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6996) );
  INV_X1 U8748 ( .A(n6995), .ZN(n6997) );
  INV_X1 U8749 ( .A(n9950), .ZN(n9173) );
  OAI222_X1 U8750 ( .A1(n8339), .A2(n6996), .B1(n9537), .B2(n6997), .C1(
        P1_U3084), .C2(n9173), .ZN(P1_U3335) );
  INV_X1 U8751 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6998) );
  INV_X1 U8752 ( .A(n8573), .ZN(n8565) );
  OAI222_X1 U8753 ( .A1(n8963), .A2(n6998), .B1(n8973), .B2(n6997), .C1(
        P2_U3152), .C2(n8565), .ZN(P2_U3340) );
  OAI21_X1 U8754 ( .B1(n4377), .B2(n7824), .A(n6999), .ZN(n9415) );
  AOI21_X1 U8755 ( .B1(n7226), .B2(n9413), .A(n9390), .ZN(n7000) );
  AND2_X1 U8756 ( .A1(n7000), .A2(n7036), .ZN(n9416) );
  OAI21_X1 U8757 ( .B1(n7218), .B2(n7217), .A(n7828), .ZN(n7001) );
  XNOR2_X1 U8758 ( .A(n7001), .B(n7824), .ZN(n7002) );
  OAI222_X1 U8759 ( .A1(n9405), .A2(n7004), .B1(n9403), .B2(n7003), .C1(n7002), 
        .C2(n9400), .ZN(n9410) );
  AOI211_X1 U8760 ( .C1(n9986), .C2(n9415), .A(n9416), .B(n9410), .ZN(n7011)
         );
  OAI22_X1 U8761 ( .A1(n9529), .A2(n7008), .B1(n9989), .B2(n5882), .ZN(n7005)
         );
  INV_X1 U8762 ( .A(n7005), .ZN(n7006) );
  OAI21_X1 U8763 ( .B1(n7011), .B2(n9988), .A(n7006), .ZN(P1_U3472) );
  INV_X1 U8764 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7007) );
  OAI22_X1 U8765 ( .A1(n9491), .A2(n7008), .B1(n9994), .B2(n7007), .ZN(n7009)
         );
  INV_X1 U8766 ( .A(n7009), .ZN(n7010) );
  OAI21_X1 U8767 ( .B1(n7011), .B2(n9992), .A(n7010), .ZN(P1_U3529) );
  NOR2_X1 U8768 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9740), .ZN(n8198) );
  AOI22_X1 U8769 ( .A1(n8500), .A2(n8806), .B1(n8804), .B2(n8502), .ZN(n7139)
         );
  NOR2_X1 U8770 ( .A1(n8406), .A2(n7139), .ZN(n7012) );
  AOI211_X1 U8771 ( .C1(n10049), .C2(n8459), .A(n8198), .B(n7012), .ZN(n7027)
         );
  NAND2_X1 U8772 ( .A1(n8501), .A2(n8295), .ZN(n7013) );
  XNOR2_X1 U8773 ( .A(n10049), .B(n8308), .ZN(n7014) );
  NAND2_X1 U8774 ( .A1(n7013), .A2(n7014), .ZN(n7281) );
  INV_X1 U8775 ( .A(n7013), .ZN(n7016) );
  INV_X1 U8776 ( .A(n7014), .ZN(n7015) );
  NAND2_X1 U8777 ( .A1(n7016), .A2(n7015), .ZN(n7017) );
  AND2_X1 U8778 ( .A1(n7281), .A2(n7017), .ZN(n7278) );
  INV_X1 U8779 ( .A(n7020), .ZN(n7023) );
  INV_X1 U8780 ( .A(n7021), .ZN(n7022) );
  NAND2_X1 U8781 ( .A1(n7023), .A2(n7022), .ZN(n7024) );
  NAND2_X1 U8782 ( .A1(n7286), .A2(n7278), .ZN(n7253) );
  OAI21_X1 U8783 ( .B1(n7278), .B2(n7286), .A(n7253), .ZN(n7025) );
  NAND2_X1 U8784 ( .A1(n7025), .A2(n8441), .ZN(n7026) );
  OAI211_X1 U8785 ( .C1(n8483), .C2(n7145), .A(n7027), .B(n7026), .ZN(P2_U3241) );
  OAI21_X1 U8786 ( .B1(n7029), .B2(n7968), .A(n7028), .ZN(n7348) );
  INV_X1 U8787 ( .A(n7348), .ZN(n7045) );
  NOR2_X1 U8788 ( .A1(n4378), .A2(n7030), .ZN(n7031) );
  INV_X1 U8789 ( .A(n9121), .ZN(n7367) );
  INV_X1 U8790 ( .A(n7245), .ZN(n7032) );
  AOI21_X1 U8791 ( .B1(n7968), .B2(n7033), .A(n7032), .ZN(n7034) );
  OAI222_X1 U8792 ( .A1(n9405), .A2(n7367), .B1(n9403), .B2(n7035), .C1(n9400), 
        .C2(n7034), .ZN(n7346) );
  INV_X2 U8793 ( .A(n9826), .ZN(n9409) );
  NAND2_X1 U8794 ( .A1(n7346), .A2(n9409), .ZN(n7044) );
  AOI211_X1 U8795 ( .C1(n7037), .C2(n7036), .A(n9390), .B(n7238), .ZN(n7347)
         );
  OR2_X1 U8796 ( .A1(n7038), .A2(n9184), .ZN(n9199) );
  NOR2_X1 U8797 ( .A1(n9392), .A2(n7352), .ZN(n7042) );
  OAI22_X1 U8798 ( .A1(n9409), .A2(n7040), .B1(n7039), .B2(n9820), .ZN(n7041)
         );
  AOI211_X1 U8799 ( .C1(n7347), .C2(n9818), .A(n7042), .B(n7041), .ZN(n7043)
         );
  OAI211_X1 U8800 ( .C1(n7045), .C2(n9408), .A(n7044), .B(n7043), .ZN(P1_U3284) );
  XOR2_X1 U8801 ( .A(n6936), .B(n7046), .Z(n10020) );
  INV_X1 U8802 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9699) );
  XNOR2_X1 U8803 ( .A(n5519), .B(n6936), .ZN(n7048) );
  AOI21_X1 U8804 ( .B1(n7048), .B2(n8848), .A(n7047), .ZN(n10025) );
  OAI21_X1 U8805 ( .B1(n9699), .B2(n8852), .A(n10025), .ZN(n7049) );
  NAND2_X1 U8806 ( .A1(n8831), .A2(n7049), .ZN(n7051) );
  NAND2_X1 U8807 ( .A1(n7054), .A2(n7158), .ZN(n10021) );
  NAND3_X1 U8808 ( .A1(n8856), .A2(n10022), .A3(n10021), .ZN(n7050) );
  OAI211_X1 U8809 ( .C1(n8831), .C2(n7052), .A(n7051), .B(n7050), .ZN(n7053)
         );
  AOI21_X1 U8810 ( .B1(n8854), .B2(n7054), .A(n7053), .ZN(n7055) );
  OAI21_X1 U8811 ( .B1(n8812), .B2(n10020), .A(n7055), .ZN(P2_U3295) );
  XOR2_X1 U8812 ( .A(n7056), .B(n7060), .Z(n10029) );
  OR2_X1 U8813 ( .A1(n7057), .A2(n8583), .ZN(n7172) );
  NAND2_X1 U8814 ( .A1(n10022), .A2(n7069), .ZN(n7058) );
  NAND2_X1 U8815 ( .A1(n7058), .A2(n10089), .ZN(n7059) );
  OR2_X1 U8816 ( .A1(n7059), .A2(n7094), .ZN(n10030) );
  OAI22_X1 U8817 ( .A1(n7172), .A2(n10030), .B1(n9625), .B2(n8852), .ZN(n7068)
         );
  NAND2_X1 U8818 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  NAND2_X1 U8819 ( .A1(n7099), .A2(n7062), .ZN(n7065) );
  OAI22_X1 U8820 ( .A1(n4316), .A2(n8840), .B1(n7063), .B2(n8838), .ZN(n7064)
         );
  AOI21_X1 U8821 ( .B1(n7065), .B2(n8848), .A(n7064), .ZN(n10031) );
  NAND2_X1 U8822 ( .A1(n4314), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7066) );
  OAI21_X1 U8823 ( .B1(n4314), .B2(n10031), .A(n7066), .ZN(n7067) );
  AOI211_X1 U8824 ( .C1(n8854), .C2(n7069), .A(n7068), .B(n7067), .ZN(n7070)
         );
  OAI21_X1 U8825 ( .B1(n8812), .B2(n10029), .A(n7070), .ZN(P2_U3294) );
  AND2_X1 U8826 ( .A1(n7071), .A2(n9184), .ZN(n7072) );
  AND2_X1 U8827 ( .A1(n9409), .A2(n7072), .ZN(n9819) );
  INV_X1 U8828 ( .A(n9819), .ZN(n7079) );
  OAI22_X1 U8829 ( .A1(n9409), .A2(n6534), .B1(n7073), .B2(n9820), .ZN(n7074)
         );
  AOI21_X1 U8830 ( .B1(n9831), .B2(n5774), .A(n7074), .ZN(n7078) );
  INV_X1 U8831 ( .A(n7075), .ZN(n7076) );
  NAND2_X1 U8832 ( .A1(n7076), .A2(n9397), .ZN(n7077) );
  OAI211_X1 U8833 ( .C1(n7080), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7081)
         );
  INV_X1 U8834 ( .A(n7081), .ZN(n7082) );
  OAI21_X1 U8835 ( .B1(n7083), .B2(n9826), .A(n7082), .ZN(P1_U3290) );
  INV_X1 U8836 ( .A(n7084), .ZN(n7093) );
  NAND2_X1 U8837 ( .A1(n7085), .A2(n9818), .ZN(n7088) );
  INV_X1 U8838 ( .A(n9820), .ZN(n9339) );
  AOI22_X1 U8839 ( .A1(n9826), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7086), .B2(
        n9339), .ZN(n7087) );
  OAI211_X1 U8840 ( .C1(n7089), .C2(n9392), .A(n7088), .B(n7087), .ZN(n7090)
         );
  AOI21_X1 U8841 ( .B1(n9414), .B2(n7091), .A(n7090), .ZN(n7092) );
  OAI21_X1 U8842 ( .B1(n7093), .B2(n9826), .A(n7092), .ZN(P1_U3287) );
  XNOR2_X1 U8843 ( .A(n7110), .B(n7112), .ZN(n10039) );
  INV_X1 U8844 ( .A(n10039), .ZN(n7108) );
  OR2_X1 U8845 ( .A1(n7094), .A2(n10037), .ZN(n7095) );
  AND2_X1 U8846 ( .A1(n7120), .A2(n7095), .ZN(n10035) );
  NAND2_X1 U8847 ( .A1(n8856), .A2(n10035), .ZN(n7096) );
  OAI21_X1 U8848 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n8852), .A(n7096), .ZN(
        n7097) );
  AOI21_X1 U8849 ( .B1(n8854), .B2(n4996), .A(n7097), .ZN(n7107) );
  NAND2_X1 U8850 ( .A1(n10039), .A2(n7664), .ZN(n7105) );
  NAND3_X1 U8851 ( .A1(n7099), .A2(n7110), .A3(n7098), .ZN(n7100) );
  NAND2_X1 U8852 ( .A1(n7101), .A2(n7100), .ZN(n7103) );
  OAI22_X1 U8853 ( .A1(n8256), .A2(n8840), .B1(n7118), .B2(n8838), .ZN(n7102)
         );
  AOI21_X1 U8854 ( .B1(n7103), .B2(n8848), .A(n7102), .ZN(n7104) );
  AND2_X1 U8855 ( .A1(n7105), .A2(n7104), .ZN(n10041) );
  MUX2_X1 U8856 ( .A(n10041), .B(n6786), .S(n4314), .Z(n7106) );
  OAI211_X1 U8857 ( .C1(n7108), .C2(n8859), .A(n7107), .B(n7106), .ZN(P2_U3293) );
  NAND2_X1 U8858 ( .A1(n7109), .A2(n7152), .ZN(n7130) );
  NAND2_X1 U8859 ( .A1(n7112), .A2(n7111), .ZN(n7117) );
  INV_X1 U8860 ( .A(n7113), .ZN(n7115) );
  OR2_X1 U8861 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  NAND2_X1 U8862 ( .A1(n7118), .A2(n10044), .ZN(n7151) );
  XOR2_X1 U8863 ( .A(n7130), .B(n7119), .Z(n7191) );
  INV_X1 U8864 ( .A(n7172), .ZN(n8793) );
  OAI21_X1 U8865 ( .B1(n7120), .B2(n5033), .A(n7189), .ZN(n7121) );
  AND3_X1 U8866 ( .A1(n7121), .A2(n10089), .A3(n7142), .ZN(n7188) );
  NAND2_X1 U8867 ( .A1(n8793), .A2(n7188), .ZN(n7122) );
  OAI21_X1 U8868 ( .B1(n8852), .B2(n7123), .A(n7122), .ZN(n7124) );
  AOI21_X1 U8869 ( .B1(n8854), .B2(n7189), .A(n7124), .ZN(n7137) );
  INV_X1 U8870 ( .A(n7125), .ZN(n7126) );
  OR2_X1 U8871 ( .A1(n7127), .A2(n7126), .ZN(n7129) );
  NAND2_X1 U8872 ( .A1(n7129), .A2(n7128), .ZN(n7131) );
  XOR2_X1 U8873 ( .A(n7131), .B(n7130), .Z(n7133) );
  OAI21_X1 U8874 ( .B1(n7133), .B2(n8817), .A(n7132), .ZN(n7187) );
  INV_X1 U8875 ( .A(n7187), .ZN(n7135) );
  MUX2_X1 U8876 ( .A(n7135), .B(n7134), .S(n4314), .Z(n7136) );
  OAI211_X1 U8877 ( .C1(n8812), .C2(n7191), .A(n7137), .B(n7136), .ZN(P2_U3291) );
  XNOR2_X1 U8878 ( .A(n7138), .B(n7154), .ZN(n7141) );
  INV_X1 U8879 ( .A(n7139), .ZN(n7140) );
  AOI21_X1 U8880 ( .B1(n7141), .B2(n8848), .A(n7140), .ZN(n10056) );
  INV_X1 U8881 ( .A(n7171), .ZN(n7144) );
  AOI21_X1 U8882 ( .B1(n7142), .B2(n10049), .A(n10096), .ZN(n7143) );
  NAND2_X1 U8883 ( .A1(n7144), .A2(n7143), .ZN(n10051) );
  OAI22_X1 U8884 ( .A1(n7172), .A2(n10051), .B1(n7145), .B2(n8852), .ZN(n7147)
         );
  NOR2_X1 U8885 ( .A1(n8831), .A2(n6783), .ZN(n7146) );
  AOI211_X1 U8886 ( .C1(n8854), .C2(n10049), .A(n7147), .B(n7146), .ZN(n7157)
         );
  INV_X1 U8887 ( .A(n8812), .ZN(n8769) );
  NAND2_X1 U8888 ( .A1(n7149), .A2(n7148), .ZN(n7150) );
  AND2_X1 U8889 ( .A1(n7151), .A2(n7150), .ZN(n7153) );
  NAND2_X1 U8890 ( .A1(n7155), .A2(n7154), .ZN(n10052) );
  NAND3_X1 U8891 ( .A1(n8769), .A2(n10053), .A3(n10052), .ZN(n7156) );
  OAI211_X1 U8892 ( .C1(n4314), .C2(n10056), .A(n7157), .B(n7156), .ZN(
        P2_U3290) );
  OAI21_X1 U8893 ( .B1(n8854), .B2(n8856), .A(n7158), .ZN(n7161) );
  OAI22_X1 U8894 ( .A1(n10017), .A2(n8817), .B1(n4316), .B2(n8838), .ZN(n10019) );
  AOI21_X1 U8895 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n8797), .A(n10019), .ZN(
        n7159) );
  MUX2_X1 U8896 ( .A(n7159), .B(n9996), .S(n4314), .Z(n7160) );
  OAI211_X1 U8897 ( .C1(n10017), .C2(n8812), .A(n7161), .B(n7160), .ZN(
        P2_U3296) );
  NAND2_X1 U8898 ( .A1(n8501), .A2(n10049), .ZN(n7162) );
  INV_X1 U8899 ( .A(n7415), .ZN(n7163) );
  AOI21_X1 U8900 ( .B1(n7166), .B2(n7164), .A(n7163), .ZN(n10057) );
  XOR2_X1 U8901 ( .A(n7165), .B(n7166), .Z(n7169) );
  OAI22_X1 U8902 ( .A1(n7168), .A2(n8838), .B1(n7167), .B2(n8840), .ZN(n7257)
         );
  AOI21_X1 U8903 ( .B1(n7169), .B2(n8848), .A(n7257), .ZN(n10060) );
  MUX2_X1 U8904 ( .A(n10060), .B(n7170), .S(n4314), .Z(n7175) );
  OAI211_X1 U8905 ( .C1(n7171), .C2(n10059), .A(n7425), .B(n10089), .ZN(n10058) );
  OAI22_X1 U8906 ( .A1(n7172), .A2(n10058), .B1(n7260), .B2(n8852), .ZN(n7173)
         );
  AOI21_X1 U8907 ( .B1(n8854), .B2(n7252), .A(n7173), .ZN(n7174) );
  OAI211_X1 U8908 ( .C1(n10057), .C2(n8812), .A(n7175), .B(n7174), .ZN(
        P2_U3289) );
  INV_X1 U8909 ( .A(n7176), .ZN(n7178) );
  OAI222_X1 U8910 ( .A1(n8339), .A2(n7177), .B1(n9537), .B2(n7178), .C1(n8070), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8911 ( .A1(n8963), .A2(n7179), .B1(n8973), .B2(n7178), .C1(
        P2_U3152), .C2(n8828), .ZN(P2_U3339) );
  OR2_X1 U8912 ( .A1(n7181), .A2(n7180), .ZN(n7182) );
  INV_X1 U8913 ( .A(n7198), .ZN(n7185) );
  INV_X1 U8914 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7193) );
  AND2_X1 U8915 ( .A1(n8257), .A2(n8583), .ZN(n7186) );
  NAND2_X1 U8916 ( .A1(n8342), .A2(n7186), .ZN(n9806) );
  AOI211_X1 U8917 ( .C1(n10088), .C2(n7189), .A(n7188), .B(n7187), .ZN(n7190)
         );
  OAI21_X1 U8918 ( .B1(n10085), .B2(n7191), .A(n7190), .ZN(n7199) );
  NAND2_X1 U8919 ( .A1(n7199), .A2(n10120), .ZN(n7192) );
  OAI21_X1 U8920 ( .B1(n10120), .B2(n7193), .A(n7192), .ZN(P2_U3525) );
  INV_X1 U8921 ( .A(n7194), .ZN(n7195) );
  OR2_X1 U8922 ( .A1(n7196), .A2(n7195), .ZN(n7197) );
  INV_X1 U8923 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7201) );
  NAND2_X1 U8924 ( .A1(n7199), .A2(n10104), .ZN(n7200) );
  OAI21_X1 U8925 ( .B1(n10104), .B2(n7201), .A(n7200), .ZN(P2_U3466) );
  AOI21_X1 U8926 ( .B1(n7203), .B2(n5188), .A(n7202), .ZN(n7205) );
  AOI22_X1 U8927 ( .A1(n8508), .A2(n7694), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7206), .ZN(n7204) );
  NOR2_X1 U8928 ( .A1(n7205), .A2(n7204), .ZN(n8509) );
  AOI21_X1 U8929 ( .B1(n7205), .B2(n7204), .A(n8509), .ZN(n7216) );
  AOI22_X1 U8930 ( .A1(n8508), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n5207), .B2(
        n7206), .ZN(n7210) );
  OAI21_X1 U8931 ( .B1(n7210), .B2(n7209), .A(n8506), .ZN(n7211) );
  NAND2_X1 U8932 ( .A1(n7211), .A2(n9995), .ZN(n7215) );
  INV_X1 U8933 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7212) );
  NAND2_X1 U8934 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7591) );
  OAI21_X1 U8935 ( .B1(n8587), .B2(n7212), .A(n7591), .ZN(n7213) );
  AOI21_X1 U8936 ( .B1(n9781), .B2(n8508), .A(n7213), .ZN(n7214) );
  OAI211_X1 U8937 ( .C1(n7216), .C2(n8578), .A(n7215), .B(n7214), .ZN(P2_U3259) );
  XNOR2_X1 U8938 ( .A(n7218), .B(n7217), .ZN(n7219) );
  NAND2_X1 U8939 ( .A1(n7219), .A2(n9351), .ZN(n7221) );
  AOI22_X1 U8940 ( .A1(n9346), .A2(n9125), .B1(n9123), .B2(n9348), .ZN(n7220)
         );
  NAND2_X1 U8941 ( .A1(n7221), .A2(n7220), .ZN(n9977) );
  INV_X1 U8942 ( .A(n9977), .ZN(n7234) );
  NAND2_X1 U8943 ( .A1(n7223), .A2(n7222), .ZN(n7224) );
  AND2_X1 U8944 ( .A1(n7225), .A2(n7224), .ZN(n9979) );
  OAI211_X1 U8945 ( .C1(n7227), .C2(n9976), .A(n9228), .B(n7226), .ZN(n9975)
         );
  OAI22_X1 U8946 ( .A1(n9409), .A2(n6536), .B1(n7228), .B2(n9820), .ZN(n7229)
         );
  AOI21_X1 U8947 ( .B1(n9831), .B2(n4509), .A(n7229), .ZN(n7230) );
  OAI21_X1 U8948 ( .B1(n9975), .B2(n7231), .A(n7230), .ZN(n7232) );
  AOI21_X1 U8949 ( .B1(n9979), .B2(n9414), .A(n7232), .ZN(n7233) );
  OAI21_X1 U8950 ( .B1(n7234), .B2(n9826), .A(n7233), .ZN(P1_U3286) );
  INV_X1 U8951 ( .A(n7235), .ZN(n7236) );
  AOI21_X1 U8952 ( .B1(n7244), .B2(n7237), .A(n7236), .ZN(n7304) );
  INV_X1 U8953 ( .A(n7304), .ZN(n7251) );
  INV_X1 U8954 ( .A(n7238), .ZN(n7239) );
  AOI211_X1 U8955 ( .C1(n7270), .C2(n7239), .A(n9390), .B(n7317), .ZN(n7303)
         );
  NOR2_X1 U8956 ( .A1(n9392), .A2(n7308), .ZN(n7242) );
  OAI22_X1 U8957 ( .A1(n9409), .A2(n7240), .B1(n7267), .B2(n9820), .ZN(n7241)
         );
  AOI211_X1 U8958 ( .C1(n7303), .C2(n9818), .A(n7242), .B(n7241), .ZN(n7250)
         );
  NAND2_X1 U8959 ( .A1(n7243), .A2(n9351), .ZN(n7248) );
  AOI21_X1 U8960 ( .B1(n7245), .B2(n8017), .A(n7244), .ZN(n7247) );
  AOI22_X1 U8961 ( .A1(n9346), .A2(n9122), .B1(n9120), .B2(n9348), .ZN(n7246)
         );
  OAI21_X1 U8962 ( .B1(n7248), .B2(n7247), .A(n7246), .ZN(n7302) );
  NAND2_X1 U8963 ( .A1(n7302), .A2(n9409), .ZN(n7249) );
  OAI211_X1 U8964 ( .C1(n7251), .C2(n9408), .A(n7250), .B(n7249), .ZN(P1_U3283) );
  NAND2_X1 U8965 ( .A1(n8500), .A2(n8295), .ZN(n7274) );
  XNOR2_X1 U8966 ( .A(n7252), .B(n8308), .ZN(n7275) );
  XNOR2_X1 U8967 ( .A(n7274), .B(n7275), .ZN(n7280) );
  NAND2_X1 U8968 ( .A1(n7253), .A2(n7281), .ZN(n7254) );
  XOR2_X1 U8969 ( .A(n7280), .B(n7254), .Z(n7255) );
  NAND2_X1 U8970 ( .A1(n7255), .A2(n8441), .ZN(n7259) );
  NOR2_X1 U8971 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5055), .ZN(n8187) );
  NOR2_X1 U8972 ( .A1(n8490), .A2(n10059), .ZN(n7256) );
  AOI211_X1 U8973 ( .C1(n8335), .C2(n7257), .A(n8187), .B(n7256), .ZN(n7258)
         );
  OAI211_X1 U8974 ( .C1(n8483), .C2(n7260), .A(n7259), .B(n7258), .ZN(P2_U3215) );
  CLKBUF_X1 U8975 ( .A(n7261), .Z(n7262) );
  NAND2_X1 U8976 ( .A1(n7263), .A2(n7262), .ZN(n7265) );
  XNOR2_X1 U8977 ( .A(n7265), .B(n7264), .ZN(n7273) );
  OAI22_X1 U8978 ( .A1(n9096), .A2(n7267), .B1(n9070), .B2(n7266), .ZN(n7268)
         );
  AOI211_X1 U8979 ( .C1(n9062), .C2(n9122), .A(n7269), .B(n7268), .ZN(n7272)
         );
  NAND2_X1 U8980 ( .A1(n6480), .A2(n7270), .ZN(n7271) );
  OAI211_X1 U8981 ( .C1(n7273), .C2(n9103), .A(n7272), .B(n7271), .ZN(P1_U3219) );
  INV_X1 U8982 ( .A(n7274), .ZN(n7277) );
  INV_X1 U8983 ( .A(n7275), .ZN(n7276) );
  NAND2_X1 U8984 ( .A1(n7277), .A2(n7276), .ZN(n7279) );
  AND2_X1 U8985 ( .A1(n7278), .A2(n7279), .ZN(n7285) );
  INV_X1 U8986 ( .A(n7279), .ZN(n7284) );
  INV_X1 U8987 ( .A(n7280), .ZN(n7282) );
  AND2_X1 U8988 ( .A1(n7282), .A2(n7281), .ZN(n7283) );
  XNOR2_X1 U8989 ( .A(n10064), .B(n8318), .ZN(n7289) );
  NAND2_X1 U8990 ( .A1(n8499), .A2(n8309), .ZN(n7287) );
  XNOR2_X1 U8991 ( .A(n7289), .B(n7287), .ZN(n7357) );
  INV_X1 U8992 ( .A(n7287), .ZN(n7288) );
  AND2_X1 U8993 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  XNOR2_X1 U8994 ( .A(n10072), .B(n8308), .ZN(n7294) );
  INV_X1 U8995 ( .A(n7294), .ZN(n7292) );
  AND2_X1 U8996 ( .A1(n8498), .A2(n8295), .ZN(n7293) );
  INV_X1 U8997 ( .A(n7293), .ZN(n7291) );
  NAND2_X1 U8998 ( .A1(n7292), .A2(n7291), .ZN(n7573) );
  NAND2_X1 U8999 ( .A1(n7294), .A2(n7293), .ZN(n7456) );
  NAND2_X1 U9000 ( .A1(n7573), .A2(n7456), .ZN(n7295) );
  XNOR2_X1 U9001 ( .A(n7457), .B(n7295), .ZN(n7301) );
  NOR2_X1 U9002 ( .A1(n5108), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8165) );
  INV_X1 U9003 ( .A(n8165), .ZN(n7297) );
  NAND2_X1 U9004 ( .A1(n8459), .A2(n7554), .ZN(n7296) );
  OAI211_X1 U9005 ( .C1(n8483), .C2(n7550), .A(n7297), .B(n7296), .ZN(n7298)
         );
  INV_X1 U9006 ( .A(n7298), .ZN(n7300) );
  INV_X1 U9007 ( .A(n8451), .ZN(n8497) );
  AOI22_X1 U9008 ( .A1(n8461), .A2(n8499), .B1(n8460), .B2(n8497), .ZN(n7299)
         );
  OAI211_X1 U9009 ( .C1(n7301), .C2(n8477), .A(n7300), .B(n7299), .ZN(P2_U3233) );
  AOI211_X1 U9010 ( .C1(n7304), .C2(n9986), .A(n7303), .B(n7302), .ZN(n7311)
         );
  OAI22_X1 U9011 ( .A1(n9491), .A2(n7308), .B1(n9994), .B2(n6573), .ZN(n7305)
         );
  INV_X1 U9012 ( .A(n7305), .ZN(n7306) );
  OAI21_X1 U9013 ( .B1(n7311), .B2(n9992), .A(n7306), .ZN(P1_U3531) );
  INV_X1 U9014 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7307) );
  OAI22_X1 U9015 ( .A1(n9529), .A2(n7308), .B1(n9989), .B2(n7307), .ZN(n7309)
         );
  INV_X1 U9016 ( .A(n7309), .ZN(n7310) );
  OAI21_X1 U9017 ( .B1(n7311), .B2(n9988), .A(n7310), .ZN(P1_U3478) );
  XNOR2_X1 U9018 ( .A(n7312), .B(n7972), .ZN(n9987) );
  INV_X1 U9019 ( .A(n9987), .ZN(n7324) );
  OAI211_X1 U9020 ( .C1(n7314), .C2(n7972), .A(n7313), .B(n9351), .ZN(n7316)
         );
  AOI22_X1 U9021 ( .A1(n9119), .A2(n9348), .B1(n9346), .B2(n9121), .ZN(n7315)
         );
  NAND2_X1 U9022 ( .A1(n7316), .A2(n7315), .ZN(n9985) );
  OAI211_X1 U9023 ( .C1(n7317), .C2(n9983), .A(n9228), .B(n7394), .ZN(n9981)
         );
  INV_X1 U9024 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7318) );
  OAI22_X1 U9025 ( .A1(n9409), .A2(n7318), .B1(n7368), .B2(n9820), .ZN(n7319)
         );
  AOI21_X1 U9026 ( .B1(n9831), .B2(n7320), .A(n7319), .ZN(n7321) );
  OAI21_X1 U9027 ( .B1(n9981), .B2(n9199), .A(n7321), .ZN(n7322) );
  AOI21_X1 U9028 ( .B1(n9985), .B2(n9409), .A(n7322), .ZN(n7323) );
  OAI21_X1 U9029 ( .B1(n7324), .B2(n9408), .A(n7323), .ZN(P1_U3282) );
  AOI22_X1 U9030 ( .A1(n9831), .A2(n4839), .B1(n9339), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7325) );
  OAI21_X1 U9031 ( .B1(n9199), .B2(n7326), .A(n7325), .ZN(n7329) );
  MUX2_X1 U9032 ( .A(n7327), .B(P1_REG2_REG_2__SCAN_IN), .S(n9826), .Z(n7328)
         );
  AOI211_X1 U9033 ( .C1(n9819), .C2(n7330), .A(n7329), .B(n7328), .ZN(n7331)
         );
  INV_X1 U9034 ( .A(n7331), .ZN(P1_U3289) );
  OAI21_X1 U9035 ( .B1(n7333), .B2(n7961), .A(n7332), .ZN(n9972) );
  INV_X1 U9036 ( .A(n7334), .ZN(n7336) );
  OAI211_X1 U9037 ( .C1(n7336), .C2(n9969), .A(n9228), .B(n7335), .ZN(n9968)
         );
  AOI22_X1 U9038 ( .A1(n9831), .A2(n7338), .B1(n9339), .B2(n7337), .ZN(n7339)
         );
  OAI21_X1 U9039 ( .B1(n9968), .B2(n9199), .A(n7339), .ZN(n7344) );
  XNOR2_X1 U9040 ( .A(n7961), .B(n8025), .ZN(n7342) );
  NAND2_X1 U9041 ( .A1(n9972), .A2(n9824), .ZN(n7341) );
  AOI22_X1 U9042 ( .A1(n9346), .A2(n9127), .B1(n9125), .B2(n9348), .ZN(n7340)
         );
  OAI211_X1 U9043 ( .C1(n9400), .C2(n7342), .A(n7341), .B(n7340), .ZN(n9970)
         );
  MUX2_X1 U9044 ( .A(n9970), .B(P1_REG2_REG_3__SCAN_IN), .S(n9826), .Z(n7343)
         );
  AOI211_X1 U9045 ( .C1(n9819), .C2(n9972), .A(n7344), .B(n7343), .ZN(n7345)
         );
  INV_X1 U9046 ( .A(n7345), .ZN(P1_U3288) );
  AOI211_X1 U9047 ( .C1(n9986), .C2(n7348), .A(n7347), .B(n7346), .ZN(n7355)
         );
  OAI22_X1 U9048 ( .A1(n9491), .A2(n7352), .B1(n9994), .B2(n5909), .ZN(n7349)
         );
  INV_X1 U9049 ( .A(n7349), .ZN(n7350) );
  OAI21_X1 U9050 ( .B1(n7355), .B2(n9992), .A(n7350), .ZN(P1_U3530) );
  INV_X1 U9051 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7351) );
  OAI22_X1 U9052 ( .A1(n9529), .A2(n7352), .B1(n9989), .B2(n7351), .ZN(n7353)
         );
  INV_X1 U9053 ( .A(n7353), .ZN(n7354) );
  OAI21_X1 U9054 ( .B1(n7355), .B2(n9988), .A(n7354), .ZN(P1_U3475) );
  XOR2_X1 U9055 ( .A(n7357), .B(n7356), .Z(n7361) );
  AOI22_X1 U9056 ( .A1(n8461), .A2(n8500), .B1(n8460), .B2(n8498), .ZN(n7359)
         );
  AOI22_X1 U9057 ( .A1(n8459), .A2(n10064), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n7358) );
  OAI211_X1 U9058 ( .C1(n7427), .C2(n8483), .A(n7359), .B(n7358), .ZN(n7360)
         );
  AOI21_X1 U9059 ( .B1(n7361), .B2(n8441), .A(n7360), .ZN(n7362) );
  INV_X1 U9060 ( .A(n7362), .ZN(P2_U3223) );
  XNOR2_X1 U9061 ( .A(n7364), .B(n7365), .ZN(n7366) );
  NAND2_X1 U9062 ( .A1(n7366), .A2(n9080), .ZN(n7371) );
  AND2_X1 U9063 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9940) );
  OAI22_X1 U9064 ( .A1(n9096), .A2(n7368), .B1(n9094), .B2(n7367), .ZN(n7369)
         );
  AOI211_X1 U9065 ( .C1(n9099), .C2(n9119), .A(n9940), .B(n7369), .ZN(n7370)
         );
  OAI211_X1 U9066 ( .C1(n9983), .C2(n9087), .A(n7371), .B(n7370), .ZN(P1_U3229) );
  INV_X1 U9067 ( .A(n7372), .ZN(n8258) );
  OAI222_X1 U9068 ( .A1(n8339), .A2(n7373), .B1(P1_U3084), .B2(n8122), .C1(
        n9537), .C2(n8258), .ZN(P1_U3333) );
  NOR2_X1 U9069 ( .A1(n7375), .A2(n7374), .ZN(n7377) );
  NOR2_X1 U9070 ( .A1(n7377), .A2(n7376), .ZN(n7494) );
  XNOR2_X1 U9071 ( .A(n7494), .B(n7501), .ZN(n7378) );
  NOR2_X1 U9072 ( .A1(n7738), .A2(n7378), .ZN(n7495) );
  AOI211_X1 U9073 ( .C1(n7378), .C2(n7738), .A(n7495), .B(n9935), .ZN(n7385)
         );
  OAI21_X1 U9074 ( .B1(n7380), .B2(P1_REG1_REG_14__SCAN_IN), .A(n7379), .ZN(
        n7500) );
  XNOR2_X1 U9075 ( .A(n7501), .B(n7500), .ZN(n7381) );
  NOR2_X1 U9076 ( .A1(n6079), .A2(n7381), .ZN(n7502) );
  AOI211_X1 U9077 ( .C1(n7381), .C2(n6079), .A(n7502), .B(n9882), .ZN(n7384)
         );
  NAND2_X1 U9078 ( .A1(n9866), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7382) );
  NAND2_X1 U9079 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9092) );
  OAI211_X1 U9080 ( .C1(n9943), .C2(n7501), .A(n7382), .B(n9092), .ZN(n7383)
         );
  OR3_X1 U9081 ( .A1(n7385), .A2(n7384), .A3(n7383), .ZN(P1_U3256) );
  INV_X1 U9082 ( .A(n7386), .ZN(n7401) );
  OAI222_X1 U9083 ( .A1(n8963), .A2(n7388), .B1(n8973), .B2(n7401), .C1(n7387), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  XNOR2_X1 U9084 ( .A(n7389), .B(n7392), .ZN(n7390) );
  AOI222_X1 U9085 ( .A1(n9351), .A2(n7390), .B1(n9118), .B2(n9348), .C1(n9120), 
        .C2(n9346), .ZN(n9789) );
  XNOR2_X1 U9086 ( .A(n7391), .B(n7392), .ZN(n9792) );
  NAND2_X1 U9087 ( .A1(n9792), .A2(n9414), .ZN(n7400) );
  OAI22_X1 U9088 ( .A1(n9409), .A2(n7393), .B1(n7408), .B2(n9820), .ZN(n7397)
         );
  INV_X1 U9089 ( .A(n7394), .ZN(n7395) );
  INV_X1 U9090 ( .A(n7398), .ZN(n9790) );
  OAI211_X1 U9091 ( .C1(n7395), .C2(n9790), .A(n9228), .B(n7447), .ZN(n9788)
         );
  NOR2_X1 U9092 ( .A1(n9788), .A2(n9199), .ZN(n7396) );
  AOI211_X1 U9093 ( .C1(n9831), .C2(n7398), .A(n7397), .B(n7396), .ZN(n7399)
         );
  OAI211_X1 U9094 ( .C1(n9826), .C2(n9789), .A(n7400), .B(n7399), .ZN(P1_U3281) );
  OAI222_X1 U9095 ( .A1(n8339), .A2(n7402), .B1(P1_U3084), .B2(n8066), .C1(
        n9537), .C2(n7401), .ZN(P1_U3332) );
  XNOR2_X1 U9096 ( .A(n7404), .B(n7403), .ZN(n7405) );
  XNOR2_X1 U9097 ( .A(n7406), .B(n7405), .ZN(n7407) );
  NAND2_X1 U9098 ( .A1(n7407), .A2(n9080), .ZN(n7412) );
  OAI22_X1 U9099 ( .A1(n9096), .A2(n7408), .B1(n9070), .B2(n7642), .ZN(n7409)
         );
  AOI211_X1 U9100 ( .C1(n9062), .C2(n9120), .A(n7410), .B(n7409), .ZN(n7411)
         );
  OAI211_X1 U9101 ( .C1(n9790), .C2(n9087), .A(n7412), .B(n7411), .ZN(P1_U3215) );
  NAND2_X1 U9102 ( .A1(n7413), .A2(n10059), .ZN(n7414) );
  NAND2_X1 U9103 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  INV_X1 U9104 ( .A(n10069), .ZN(n7433) );
  INV_X1 U9105 ( .A(n7420), .ZN(n7421) );
  AOI21_X1 U9106 ( .B1(n4885), .B2(n7419), .A(n7421), .ZN(n7424) );
  AOI22_X1 U9107 ( .A1(n8500), .A2(n8804), .B1(n8806), .B2(n8498), .ZN(n7423)
         );
  NAND2_X1 U9108 ( .A1(n10069), .A2(n7664), .ZN(n7422) );
  OAI211_X1 U9109 ( .C1(n7424), .C2(n8817), .A(n7423), .B(n7422), .ZN(n10067)
         );
  NAND2_X1 U9110 ( .A1(n10067), .A2(n8831), .ZN(n7432) );
  INV_X1 U9111 ( .A(n8856), .ZN(n8601) );
  NAND2_X1 U9112 ( .A1(n7425), .A2(n10064), .ZN(n7426) );
  NAND2_X1 U9113 ( .A1(n7548), .A2(n7426), .ZN(n10066) );
  NOR2_X1 U9114 ( .A1(n8852), .A2(n7427), .ZN(n7428) );
  AOI21_X1 U9115 ( .B1(n4314), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7428), .ZN(
        n7429) );
  OAI21_X1 U9116 ( .B1(n8601), .B2(n10066), .A(n7429), .ZN(n7430) );
  AOI21_X1 U9117 ( .B1(n8854), .B2(n10064), .A(n7430), .ZN(n7431) );
  OAI211_X1 U9118 ( .C1(n7433), .C2(n8859), .A(n7432), .B(n7431), .ZN(P2_U3288) );
  XNOR2_X1 U9119 ( .A(n7435), .B(n7434), .ZN(n7439) );
  AND2_X1 U9120 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9147) );
  OAI22_X1 U9121 ( .A1(n9096), .A2(n7450), .B1(n9070), .B2(n7757), .ZN(n7436)
         );
  AOI211_X1 U9122 ( .C1(n9062), .C2(n9119), .A(n9147), .B(n7436), .ZN(n7438)
         );
  NAND2_X1 U9123 ( .A1(n9844), .A2(n6480), .ZN(n7437) );
  OAI211_X1 U9124 ( .C1(n7439), .C2(n9103), .A(n7438), .B(n7437), .ZN(P1_U3234) );
  XNOR2_X1 U9125 ( .A(n9844), .B(n9118), .ZN(n7849) );
  INV_X1 U9126 ( .A(n7849), .ZN(n7977) );
  XNOR2_X1 U9127 ( .A(n7440), .B(n7977), .ZN(n9848) );
  XNOR2_X1 U9128 ( .A(n7441), .B(n7849), .ZN(n7445) );
  OAI22_X1 U9129 ( .A1(n7442), .A2(n9403), .B1(n7757), .B2(n9405), .ZN(n7443)
         );
  INV_X1 U9130 ( .A(n7443), .ZN(n7444) );
  OAI21_X1 U9131 ( .B1(n7445), .B2(n9400), .A(n7444), .ZN(n7446) );
  AOI21_X1 U9132 ( .B1(n9848), .B2(n9824), .A(n7446), .ZN(n9850) );
  NAND2_X1 U9133 ( .A1(n7447), .A2(n9844), .ZN(n7448) );
  NAND2_X1 U9134 ( .A1(n7448), .A2(n9228), .ZN(n7449) );
  OR2_X1 U9135 ( .A1(n7616), .A2(n7449), .ZN(n9846) );
  OAI22_X1 U9136 ( .A1(n9409), .A2(n7451), .B1(n7450), .B2(n9820), .ZN(n7452)
         );
  AOI21_X1 U9137 ( .B1(n9844), .B2(n9831), .A(n7452), .ZN(n7453) );
  OAI21_X1 U9138 ( .B1(n9846), .B2(n9199), .A(n7453), .ZN(n7454) );
  AOI21_X1 U9139 ( .B1(n9848), .B2(n9819), .A(n7454), .ZN(n7455) );
  OAI21_X1 U9140 ( .B1(n9850), .B2(n9826), .A(n7455), .ZN(P1_U3280) );
  NAND2_X1 U9141 ( .A1(n7457), .A2(n7456), .ZN(n7574) );
  XNOR2_X1 U9142 ( .A(n7578), .B(n8318), .ZN(n7458) );
  NOR2_X1 U9143 ( .A1(n8451), .A2(n8319), .ZN(n7459) );
  NAND2_X1 U9144 ( .A1(n7458), .A2(n7459), .ZN(n7470) );
  INV_X1 U9145 ( .A(n7458), .ZN(n8452) );
  INV_X1 U9146 ( .A(n7459), .ZN(n7460) );
  NAND2_X1 U9147 ( .A1(n8452), .A2(n7460), .ZN(n7461) );
  NAND2_X1 U9148 ( .A1(n7470), .A2(n7461), .ZN(n7577) );
  INV_X1 U9149 ( .A(n7577), .ZN(n7462) );
  AND2_X1 U9150 ( .A1(n7573), .A2(n7462), .ZN(n7467) );
  XNOR2_X1 U9151 ( .A(n10087), .B(n8318), .ZN(n7463) );
  NOR2_X1 U9152 ( .A1(n8390), .A2(n8319), .ZN(n7464) );
  NAND2_X1 U9153 ( .A1(n7463), .A2(n7464), .ZN(n7471) );
  INV_X1 U9154 ( .A(n7463), .ZN(n8391) );
  INV_X1 U9155 ( .A(n7464), .ZN(n7465) );
  NAND2_X1 U9156 ( .A1(n8391), .A2(n7465), .ZN(n7466) );
  AND2_X1 U9157 ( .A1(n7471), .A2(n7466), .ZN(n7469) );
  AND2_X1 U9158 ( .A1(n7467), .A2(n7469), .ZN(n7468) );
  NAND2_X1 U9159 ( .A1(n7574), .A2(n7468), .ZN(n8387) );
  INV_X1 U9160 ( .A(n7469), .ZN(n8449) );
  OR2_X1 U9161 ( .A1(n8449), .A2(n7470), .ZN(n8386) );
  AND2_X1 U9162 ( .A1(n7471), .A2(n8386), .ZN(n7472) );
  NAND2_X1 U9163 ( .A1(n8387), .A2(n7472), .ZN(n7477) );
  XNOR2_X1 U9164 ( .A(n8398), .B(n8318), .ZN(n7473) );
  NOR2_X1 U9165 ( .A1(n7660), .A2(n8319), .ZN(n7474) );
  NAND2_X1 U9166 ( .A1(n7473), .A2(n7474), .ZN(n7483) );
  INV_X1 U9167 ( .A(n7473), .ZN(n7482) );
  INV_X1 U9168 ( .A(n7474), .ZN(n7475) );
  NAND2_X1 U9169 ( .A1(n7482), .A2(n7475), .ZN(n7476) );
  AND2_X1 U9170 ( .A1(n7483), .A2(n7476), .ZN(n8388) );
  NAND2_X2 U9171 ( .A1(n7477), .A2(n8388), .ZN(n8392) );
  XNOR2_X1 U9172 ( .A(n7681), .B(n8318), .ZN(n7478) );
  NOR2_X1 U9173 ( .A1(n7590), .A2(n8319), .ZN(n7479) );
  NAND2_X1 U9174 ( .A1(n7478), .A2(n7479), .ZN(n7587) );
  INV_X1 U9175 ( .A(n7478), .ZN(n7584) );
  INV_X1 U9176 ( .A(n7479), .ZN(n7480) );
  NAND2_X1 U9177 ( .A1(n7584), .A2(n7480), .ZN(n7481) );
  AND2_X1 U9178 ( .A1(n7587), .A2(n7481), .ZN(n7484) );
  AOI21_X1 U9179 ( .B1(n8392), .B2(n4725), .A(n8477), .ZN(n7487) );
  NOR3_X1 U9180 ( .A1(n8475), .A2(n7482), .A3(n7660), .ZN(n7486) );
  OAI21_X1 U9181 ( .B1(n7487), .B2(n7486), .A(n7589), .ZN(n7491) );
  INV_X1 U9182 ( .A(n7660), .ZN(n8495) );
  OAI22_X1 U9183 ( .A1(n8483), .A2(n7667), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6989), .ZN(n7489) );
  INV_X1 U9184 ( .A(n7781), .ZN(n8493) );
  AND2_X1 U9185 ( .A1(n8460), .A2(n8493), .ZN(n7488) );
  AOI211_X1 U9186 ( .C1(n8461), .C2(n8495), .A(n7489), .B(n7488), .ZN(n7490)
         );
  OAI211_X1 U9187 ( .C1(n4578), .C2(n8490), .A(n7491), .B(n7490), .ZN(P2_U3236) );
  INV_X1 U9188 ( .A(n7492), .ZN(n8343) );
  OAI222_X1 U9189 ( .A1(n8339), .A2(n7493), .B1(n9537), .B2(n8343), .C1(n6349), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  NOR2_X1 U9190 ( .A1(n7494), .A2(n7501), .ZN(n7496) );
  NAND2_X1 U9191 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9160), .ZN(n7497) );
  OAI21_X1 U9192 ( .B1(n9160), .B2(P1_REG2_REG_16__SCAN_IN), .A(n7497), .ZN(
        n7498) );
  AOI211_X1 U9193 ( .C1(n7499), .C2(n7498), .A(n9155), .B(n9935), .ZN(n7512)
         );
  NOR2_X1 U9194 ( .A1(n7501), .A2(n7500), .ZN(n7503) );
  NOR2_X1 U9195 ( .A1(n7503), .A2(n7502), .ZN(n7506) );
  MUX2_X1 U9196 ( .A(n7504), .B(P1_REG1_REG_16__SCAN_IN), .S(n9160), .Z(n7505)
         );
  NOR2_X1 U9197 ( .A1(n7506), .A2(n7505), .ZN(n9159) );
  AOI211_X1 U9198 ( .C1(n7506), .C2(n7505), .A(n9159), .B(n9882), .ZN(n7511)
         );
  NAND2_X1 U9199 ( .A1(n9866), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7508) );
  NAND2_X1 U9200 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n7507) );
  OAI211_X1 U9201 ( .C1(n9943), .C2(n7509), .A(n7508), .B(n7507), .ZN(n7510)
         );
  OR3_X1 U9202 ( .A1(n7512), .A2(n7511), .A3(n7510), .ZN(P1_U3257) );
  NAND2_X1 U9203 ( .A1(n7514), .A2(n7513), .ZN(n7526) );
  INV_X1 U9204 ( .A(n7526), .ZN(n7515) );
  XNOR2_X1 U9205 ( .A(n7516), .B(n7515), .ZN(n7517) );
  NAND2_X1 U9206 ( .A1(n7517), .A2(n8848), .ZN(n7520) );
  OAI22_X1 U9207 ( .A1(n7590), .A2(n8838), .B1(n8390), .B2(n8840), .ZN(n7518)
         );
  INV_X1 U9208 ( .A(n7518), .ZN(n7519) );
  NAND2_X1 U9209 ( .A1(n7520), .A2(n7519), .ZN(n10098) );
  INV_X1 U9210 ( .A(n10098), .ZN(n7535) );
  AND2_X1 U9211 ( .A1(n7543), .A2(n7537), .ZN(n7536) );
  NAND2_X1 U9212 ( .A1(n7578), .A2(n8497), .ZN(n7522) );
  AND2_X1 U9213 ( .A1(n7536), .A2(n7522), .ZN(n7521) );
  NAND2_X1 U9214 ( .A1(n7538), .A2(n7521), .ZN(n7608) );
  NAND2_X1 U9215 ( .A1(n10072), .A2(n7562), .ZN(n7557) );
  AND2_X1 U9216 ( .A1(n7610), .A2(n7607), .ZN(n7524) );
  NAND2_X1 U9217 ( .A1(n7608), .A2(n7524), .ZN(n7609) );
  INV_X1 U9218 ( .A(n8390), .ZN(n8496) );
  NAND2_X1 U9219 ( .A1(n10087), .A2(n8496), .ZN(n7525) );
  NAND2_X1 U9220 ( .A1(n7527), .A2(n7526), .ZN(n7651) );
  OAI21_X1 U9221 ( .B1(n7527), .B2(n7526), .A(n7651), .ZN(n10100) );
  INV_X1 U9222 ( .A(n7578), .ZN(n10079) );
  INV_X1 U9223 ( .A(n10087), .ZN(n7606) );
  NAND2_X1 U9224 ( .A1(n7603), .A2(n7606), .ZN(n7528) );
  INV_X1 U9225 ( .A(n7528), .ZN(n7529) );
  INV_X1 U9226 ( .A(n8398), .ZN(n10095) );
  OAI21_X1 U9227 ( .B1(n7529), .B2(n10095), .A(n7665), .ZN(n10097) );
  OAI22_X1 U9228 ( .A1(n8831), .A2(n7530), .B1(n8395), .B2(n8852), .ZN(n7531)
         );
  AOI21_X1 U9229 ( .B1(n8854), .B2(n8398), .A(n7531), .ZN(n7532) );
  OAI21_X1 U9230 ( .B1(n8601), .B2(n10097), .A(n7532), .ZN(n7533) );
  AOI21_X1 U9231 ( .B1(n10100), .B2(n8769), .A(n7533), .ZN(n7534) );
  OAI21_X1 U9232 ( .B1(n4314), .B2(n7535), .A(n7534), .ZN(P2_U3284) );
  NAND2_X1 U9233 ( .A1(n7538), .A2(n7536), .ZN(n7558) );
  INV_X1 U9234 ( .A(n7558), .ZN(n7540) );
  AOI21_X1 U9235 ( .B1(n7538), .B2(n7537), .A(n7543), .ZN(n7539) );
  NOR2_X1 U9236 ( .A1(n7540), .A2(n7539), .ZN(n10071) );
  AOI22_X1 U9237 ( .A1(n8497), .A2(n8806), .B1(n8804), .B2(n8499), .ZN(n7547)
         );
  INV_X1 U9238 ( .A(n7541), .ZN(n7545) );
  AND3_X1 U9239 ( .A1(n7420), .A2(n7543), .A3(n7542), .ZN(n7544) );
  OAI21_X1 U9240 ( .B1(n7545), .B2(n7544), .A(n8848), .ZN(n7546) );
  OAI211_X1 U9241 ( .C1(n10071), .C2(n8845), .A(n7547), .B(n7546), .ZN(n10074)
         );
  NAND2_X1 U9242 ( .A1(n10074), .A2(n8831), .ZN(n7556) );
  AND2_X1 U9243 ( .A1(n7548), .A2(n7554), .ZN(n7549) );
  OR2_X1 U9244 ( .A1(n7549), .A2(n7566), .ZN(n10073) );
  NOR2_X1 U9245 ( .A1(n8852), .A2(n7550), .ZN(n7551) );
  AOI21_X1 U9246 ( .B1(n4314), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7551), .ZN(
        n7552) );
  OAI21_X1 U9247 ( .B1(n8601), .B2(n10073), .A(n7552), .ZN(n7553) );
  AOI21_X1 U9248 ( .B1(n8854), .B2(n7554), .A(n7553), .ZN(n7555) );
  OAI211_X1 U9249 ( .C1(n10071), .C2(n8859), .A(n7556), .B(n7555), .ZN(
        P2_U3287) );
  NAND2_X1 U9250 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  XNOR2_X1 U9251 ( .A(n7559), .B(n7560), .ZN(n10078) );
  XNOR2_X1 U9252 ( .A(n7561), .B(n7560), .ZN(n7564) );
  OAI22_X1 U9253 ( .A1(n7562), .A2(n8840), .B1(n8390), .B2(n8838), .ZN(n7563)
         );
  AOI21_X1 U9254 ( .B1(n7564), .B2(n8848), .A(n7563), .ZN(n7565) );
  OAI21_X1 U9255 ( .B1(n10078), .B2(n8845), .A(n7565), .ZN(n10081) );
  NAND2_X1 U9256 ( .A1(n10081), .A2(n8831), .ZN(n7572) );
  NOR2_X1 U9257 ( .A1(n7566), .A2(n10079), .ZN(n7567) );
  OR2_X1 U9258 ( .A1(n7603), .A2(n7567), .ZN(n10080) );
  NOR2_X1 U9259 ( .A1(n8852), .A2(n7581), .ZN(n7568) );
  AOI21_X1 U9260 ( .B1(n4314), .B2(P2_REG2_REG_10__SCAN_IN), .A(n7568), .ZN(
        n7569) );
  OAI21_X1 U9261 ( .B1(n8601), .B2(n10080), .A(n7569), .ZN(n7570) );
  AOI21_X1 U9262 ( .B1(n8854), .B2(n7578), .A(n7570), .ZN(n7571) );
  OAI211_X1 U9263 ( .C1(n10078), .C2(n8859), .A(n7572), .B(n7571), .ZN(
        P2_U3286) );
  NAND2_X1 U9264 ( .A1(n7574), .A2(n7573), .ZN(n7576) );
  OR2_X1 U9265 ( .A1(n7576), .A2(n7577), .ZN(n8450) );
  INV_X1 U9266 ( .A(n8450), .ZN(n7575) );
  AOI211_X1 U9267 ( .C1(n7577), .C2(n7576), .A(n8477), .B(n7575), .ZN(n7583)
         );
  AOI22_X1 U9268 ( .A1(n8461), .A2(n8498), .B1(n8460), .B2(n8496), .ZN(n7580)
         );
  AOI22_X1 U9269 ( .A1(n8459), .A2(n7578), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7579) );
  OAI211_X1 U9270 ( .C1(n7581), .C2(n8483), .A(n7580), .B(n7579), .ZN(n7582)
         );
  OR2_X1 U9271 ( .A1(n7583), .A2(n7582), .ZN(P2_U3219) );
  INV_X1 U9272 ( .A(n7589), .ZN(n7586) );
  NOR3_X1 U9273 ( .A1(n8475), .A2(n7584), .A3(n7590), .ZN(n7585) );
  AOI21_X1 U9274 ( .B1(n7586), .B2(n8441), .A(n7585), .ZN(n7598) );
  XNOR2_X1 U9275 ( .A(n7775), .B(n8318), .ZN(n7713) );
  NAND2_X1 U9276 ( .A1(n8493), .A2(n8309), .ZN(n7714) );
  XNOR2_X1 U9277 ( .A(n7713), .B(n7714), .ZN(n7597) );
  INV_X1 U9278 ( .A(n7775), .ZN(n9801) );
  INV_X1 U9279 ( .A(n8841), .ZN(n8602) );
  INV_X1 U9280 ( .A(n7590), .ZN(n8494) );
  AOI22_X1 U9281 ( .A1(n8460), .A2(n8602), .B1(n8461), .B2(n8494), .ZN(n7594)
         );
  OAI21_X1 U9282 ( .B1(n8483), .B2(n7693), .A(n7591), .ZN(n7592) );
  INV_X1 U9283 ( .A(n7592), .ZN(n7593) );
  OAI211_X1 U9284 ( .C1(n9801), .C2(n8490), .A(n7594), .B(n7593), .ZN(n7595)
         );
  AOI21_X1 U9285 ( .B1(n4373), .B2(n8441), .A(n7595), .ZN(n7596) );
  OAI21_X1 U9286 ( .B1(n7598), .B2(n7597), .A(n7596), .ZN(P2_U3217) );
  XNOR2_X1 U9287 ( .A(n7599), .B(n7600), .ZN(n7602) );
  OAI22_X1 U9288 ( .A1(n8451), .A2(n8840), .B1(n7660), .B2(n8838), .ZN(n7601)
         );
  AOI21_X1 U9289 ( .B1(n7602), .B2(n8848), .A(n7601), .ZN(n10092) );
  XNOR2_X1 U9290 ( .A(n7603), .B(n10087), .ZN(n10090) );
  INV_X1 U9291 ( .A(n8456), .ZN(n7604) );
  AOI22_X1 U9292 ( .A1(n4314), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7604), .B2(
        n8797), .ZN(n7605) );
  OAI21_X1 U9293 ( .B1(n7606), .B2(n8800), .A(n7605), .ZN(n7613) );
  AND2_X1 U9294 ( .A1(n7608), .A2(n7607), .ZN(n7611) );
  OAI21_X1 U9295 ( .B1(n7611), .B2(n7610), .A(n7609), .ZN(n10086) );
  NOR2_X1 U9296 ( .A1(n10086), .A2(n8812), .ZN(n7612) );
  AOI211_X1 U9297 ( .C1(n8856), .C2(n10090), .A(n7613), .B(n7612), .ZN(n7614)
         );
  OAI21_X1 U9298 ( .B1(n4314), .B2(n10092), .A(n7614), .ZN(P2_U3285) );
  XOR2_X1 U9299 ( .A(n7615), .B(n7976), .Z(n7708) );
  INV_X1 U9300 ( .A(n7708), .ZN(n7627) );
  INV_X1 U9301 ( .A(n7616), .ZN(n7617) );
  AOI211_X1 U9302 ( .C1(n7646), .C2(n7617), .A(n9390), .B(n7753), .ZN(n7707)
         );
  NOR2_X1 U9303 ( .A1(n7712), .A2(n9392), .ZN(n7620) );
  INV_X1 U9304 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7618) );
  OAI22_X1 U9305 ( .A1(n9409), .A2(n7618), .B1(n7643), .B2(n9820), .ZN(n7619)
         );
  AOI211_X1 U9306 ( .C1(n7707), .C2(n9818), .A(n7620), .B(n7619), .ZN(n7626)
         );
  NAND2_X1 U9307 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  XOR2_X1 U9308 ( .A(n7976), .B(n7623), .Z(n7624) );
  OAI222_X1 U9309 ( .A1(n9403), .A2(n7642), .B1(n9405), .B2(n7854), .C1(n9400), 
        .C2(n7624), .ZN(n7706) );
  NAND2_X1 U9310 ( .A1(n7706), .A2(n9409), .ZN(n7625) );
  OAI211_X1 U9311 ( .C1(n7627), .C2(n9408), .A(n7626), .B(n7625), .ZN(P1_U3279) );
  INV_X1 U9312 ( .A(n7632), .ZN(n7630) );
  NOR2_X1 U9313 ( .A1(n7628), .A2(P1_U3084), .ZN(n8126) );
  AOI21_X1 U9314 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9535), .A(n8126), .ZN(
        n7629) );
  OAI21_X1 U9315 ( .B1(n7630), .B2(n9537), .A(n7629), .ZN(P1_U3330) );
  NAND2_X1 U9316 ( .A1(n7632), .A2(n7631), .ZN(n7634) );
  OAI211_X1 U9317 ( .C1(n7635), .C2(n8963), .A(n7634), .B(n7633), .ZN(P2_U3335) );
  INV_X1 U9318 ( .A(n7637), .ZN(n7638) );
  AOI21_X1 U9319 ( .B1(n7640), .B2(n7639), .A(n7638), .ZN(n7649) );
  INV_X1 U9320 ( .A(n7641), .ZN(n7645) );
  OAI22_X1 U9321 ( .A1(n9096), .A2(n7643), .B1(n9094), .B2(n7642), .ZN(n7644)
         );
  AOI211_X1 U9322 ( .C1(n9099), .C2(n9116), .A(n7645), .B(n7644), .ZN(n7648)
         );
  NAND2_X1 U9323 ( .A1(n7646), .A2(n6480), .ZN(n7647) );
  OAI211_X1 U9324 ( .C1(n7649), .C2(n9103), .A(n7648), .B(n7647), .ZN(P1_U3222) );
  OR2_X1 U9325 ( .A1(n8398), .A2(n8495), .ZN(n7650) );
  NAND2_X1 U9326 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  INV_X1 U9327 ( .A(n7682), .ZN(n7655) );
  NAND2_X1 U9328 ( .A1(n7652), .A2(n7653), .ZN(n7654) );
  NAND2_X1 U9329 ( .A1(n7658), .A2(n7657), .ZN(n7659) );
  AOI21_X1 U9330 ( .B1(n7656), .B2(n7659), .A(n8817), .ZN(n7662) );
  OAI22_X1 U9331 ( .A1(n7781), .A2(n8838), .B1(n7660), .B2(n8840), .ZN(n7661)
         );
  OR2_X1 U9332 ( .A1(n7662), .A2(n7661), .ZN(n7663) );
  AOI21_X1 U9333 ( .B1(n9809), .B2(n7664), .A(n7663), .ZN(n9811) );
  INV_X1 U9334 ( .A(n8859), .ZN(n7671) );
  AND2_X1 U9335 ( .A1(n7665), .A2(n7681), .ZN(n7666) );
  OR2_X1 U9336 ( .A1(n7666), .A2(n7692), .ZN(n9807) );
  OAI22_X1 U9337 ( .A1(n8831), .A2(n5188), .B1(n7667), .B2(n8852), .ZN(n7668)
         );
  AOI21_X1 U9338 ( .B1(n8854), .B2(n7681), .A(n7668), .ZN(n7669) );
  OAI21_X1 U9339 ( .B1(n9807), .B2(n8601), .A(n7669), .ZN(n7670) );
  AOI21_X1 U9340 ( .B1(n9809), .B2(n7671), .A(n7670), .ZN(n7672) );
  OAI21_X1 U9341 ( .B1(n9811), .B2(n4314), .A(n7672), .ZN(P2_U3283) );
  NOR2_X1 U9342 ( .A1(n4372), .A2(n7673), .ZN(n7674) );
  XNOR2_X1 U9343 ( .A(n7675), .B(n7674), .ZN(n7676) );
  NAND2_X1 U9344 ( .A1(n7676), .A2(n9080), .ZN(n7680) );
  OAI22_X1 U9345 ( .A1(n9096), .A2(n9821), .B1(n9094), .B2(n7757), .ZN(n7677)
         );
  AOI211_X1 U9346 ( .C1(n9099), .C2(n9115), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI211_X1 U9347 ( .C1(n7762), .C2(n9087), .A(n7680), .B(n7679), .ZN(P1_U3232) );
  OAI21_X1 U9348 ( .B1(n7684), .B2(n7683), .A(n7777), .ZN(n9805) );
  INV_X1 U9349 ( .A(n9805), .ZN(n7699) );
  NAND2_X1 U9350 ( .A1(n7685), .A2(n8848), .ZN(n7690) );
  AOI21_X1 U9351 ( .B1(n7656), .B2(n7687), .A(n7686), .ZN(n7689) );
  AOI22_X1 U9352 ( .A1(n8806), .A2(n8602), .B1(n8494), .B2(n8804), .ZN(n7688)
         );
  OAI21_X1 U9353 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(n9803) );
  INV_X1 U9354 ( .A(n7782), .ZN(n7691) );
  OAI21_X1 U9355 ( .B1(n9801), .B2(n7692), .A(n7691), .ZN(n9802) );
  OAI22_X1 U9356 ( .A1(n8831), .A2(n7694), .B1(n7693), .B2(n8852), .ZN(n7695)
         );
  AOI21_X1 U9357 ( .B1(n8854), .B2(n7775), .A(n7695), .ZN(n7696) );
  OAI21_X1 U9358 ( .B1(n9802), .B2(n8601), .A(n7696), .ZN(n7697) );
  AOI21_X1 U9359 ( .B1(n9803), .B2(n8831), .A(n7697), .ZN(n7698) );
  OAI21_X1 U9360 ( .B1(n7699), .B2(n8812), .A(n7698), .ZN(P2_U3282) );
  INV_X1 U9361 ( .A(n7700), .ZN(n7704) );
  OAI222_X1 U9362 ( .A1(P2_U3152), .A2(n7702), .B1(n8973), .B2(n7704), .C1(
        n7701), .C2(n8963), .ZN(P2_U3334) );
  OAI222_X1 U9363 ( .A1(P1_U3084), .A2(n7705), .B1(n9537), .B2(n7704), .C1(
        n7703), .C2(n8339), .ZN(P1_U3329) );
  AOI211_X1 U9364 ( .C1(n7708), .C2(n9986), .A(n7707), .B(n7706), .ZN(n7710)
         );
  MUX2_X1 U9365 ( .A(n6014), .B(n7710), .S(n9989), .Z(n7709) );
  OAI21_X1 U9366 ( .B1(n7712), .B2(n9529), .A(n7709), .ZN(P1_U3490) );
  MUX2_X1 U9367 ( .A(n6644), .B(n7710), .S(n9994), .Z(n7711) );
  OAI21_X1 U9368 ( .B1(n7712), .B2(n9491), .A(n7711), .ZN(P1_U3535) );
  NOR2_X1 U9369 ( .A1(n8841), .A2(n8319), .ZN(n7763) );
  INV_X1 U9370 ( .A(n7713), .ZN(n7715) );
  XNOR2_X1 U9371 ( .A(n8603), .B(n8308), .ZN(n7716) );
  NAND2_X1 U9372 ( .A1(n7764), .A2(n7766), .ZN(n7718) );
  XOR2_X1 U9373 ( .A(n7763), .B(n7718), .Z(n7722) );
  INV_X1 U9374 ( .A(n8820), .ZN(n8606) );
  AOI22_X1 U9375 ( .A1(n8461), .A2(n8493), .B1(n8460), .B2(n8606), .ZN(n7719)
         );
  NAND2_X1 U9376 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8513) );
  OAI211_X1 U9377 ( .C1(n7783), .C2(n8483), .A(n7719), .B(n8513), .ZN(n7720)
         );
  AOI21_X1 U9378 ( .B1(n8603), .B2(n8459), .A(n7720), .ZN(n7721) );
  OAI21_X1 U9379 ( .B1(n7722), .B2(n8477), .A(n7721), .ZN(P2_U3243) );
  INV_X1 U9380 ( .A(n7723), .ZN(n7733) );
  AOI211_X1 U9381 ( .C1(n7724), .C2(n7978), .A(n9400), .B(n7733), .ZN(n7726)
         );
  OAI22_X1 U9382 ( .A1(n7854), .A2(n9403), .B1(n9013), .B2(n9405), .ZN(n7725)
         );
  NOR2_X1 U9383 ( .A1(n7726), .A2(n7725), .ZN(n9840) );
  XOR2_X1 U9384 ( .A(n7727), .B(n7978), .Z(n9842) );
  NAND2_X1 U9385 ( .A1(n9842), .A2(n9414), .ZN(n7732) );
  OAI22_X1 U9386 ( .A1(n9409), .A2(n7728), .B1(n7794), .B2(n9820), .ZN(n7730)
         );
  OAI211_X1 U9387 ( .C1(n4370), .C2(n4676), .A(n9228), .B(n7739), .ZN(n9839)
         );
  NOR2_X1 U9388 ( .A1(n9839), .A2(n9199), .ZN(n7729) );
  AOI211_X1 U9389 ( .C1(n9831), .C2(n7797), .A(n7730), .B(n7729), .ZN(n7731)
         );
  OAI211_X1 U9390 ( .C1(n9826), .C2(n9840), .A(n7732), .B(n7731), .ZN(P1_U3277) );
  OAI21_X1 U9391 ( .B1(n7733), .B2(n8042), .A(n7865), .ZN(n7735) );
  NAND2_X1 U9392 ( .A1(n7735), .A2(n7734), .ZN(n7736) );
  AOI222_X1 U9393 ( .A1(n9351), .A2(n7736), .B1(n9113), .B2(n9348), .C1(n9115), 
        .C2(n9346), .ZN(n9835) );
  XNOR2_X1 U9394 ( .A(n7737), .B(n7865), .ZN(n9838) );
  NAND2_X1 U9395 ( .A1(n9838), .A2(n9414), .ZN(n7744) );
  OAI22_X1 U9396 ( .A1(n9409), .A2(n7738), .B1(n9095), .B2(n9820), .ZN(n7742)
         );
  INV_X1 U9397 ( .A(n7739), .ZN(n7740) );
  INV_X1 U9398 ( .A(n9100), .ZN(n9836) );
  OAI211_X1 U9399 ( .C1(n7740), .C2(n9836), .A(n9228), .B(n7814), .ZN(n9834)
         );
  NOR2_X1 U9400 ( .A1(n9834), .A2(n9199), .ZN(n7741) );
  AOI211_X1 U9401 ( .C1(n9831), .C2(n9100), .A(n7742), .B(n7741), .ZN(n7743)
         );
  OAI211_X1 U9402 ( .C1(n9826), .C2(n9835), .A(n7744), .B(n7743), .ZN(P1_U3276) );
  INV_X1 U9403 ( .A(n7745), .ZN(n7750) );
  INV_X1 U9404 ( .A(n7746), .ZN(n7747) );
  OAI222_X1 U9405 ( .A1(n8963), .A2(n7748), .B1(n8970), .B2(n7750), .C1(
        P2_U3152), .C2(n7747), .ZN(P2_U3333) );
  OAI222_X1 U9406 ( .A1(n8339), .A2(n7751), .B1(n9537), .B2(n7750), .C1(
        P1_U3084), .C2(n7749), .ZN(P1_U3328) );
  INV_X1 U9407 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7758) );
  XNOR2_X1 U9408 ( .A(n7752), .B(n7979), .ZN(n9825) );
  INV_X1 U9409 ( .A(n7753), .ZN(n7754) );
  AOI211_X1 U9410 ( .C1(n9830), .C2(n7754), .A(n9390), .B(n4370), .ZN(n9817)
         );
  XOR2_X1 U9411 ( .A(n7979), .B(n7755), .Z(n7756) );
  OAI222_X1 U9412 ( .A1(n9405), .A2(n9093), .B1(n9403), .B2(n7757), .C1(n9400), 
        .C2(n7756), .ZN(n9823) );
  AOI211_X1 U9413 ( .C1(n9986), .C2(n9825), .A(n9817), .B(n9823), .ZN(n7760)
         );
  MUX2_X1 U9414 ( .A(n7758), .B(n7760), .S(n9989), .Z(n7759) );
  OAI21_X1 U9415 ( .B1(n7762), .B2(n9529), .A(n7759), .ZN(P1_U3493) );
  MUX2_X1 U9416 ( .A(n6692), .B(n7760), .S(n9994), .Z(n7761) );
  OAI21_X1 U9417 ( .B1(n7762), .B2(n9491), .A(n7761), .ZN(P1_U3536) );
  XNOR2_X1 U9418 ( .A(n8938), .B(n8318), .ZN(n8262) );
  NOR2_X1 U9419 ( .A1(n8820), .A2(n8319), .ZN(n8263) );
  XNOR2_X1 U9420 ( .A(n8262), .B(n8263), .ZN(n7769) );
  NAND2_X1 U9421 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  NAND2_X1 U9422 ( .A1(n7766), .A2(n7765), .ZN(n7768) );
  INV_X1 U9423 ( .A(n8267), .ZN(n7767) );
  AOI21_X1 U9424 ( .B1(n7769), .B2(n7768), .A(n7767), .ZN(n7774) );
  INV_X1 U9425 ( .A(n8839), .ZN(n8805) );
  AOI22_X1 U9426 ( .A1(n8461), .A2(n8602), .B1(n8460), .B2(n8805), .ZN(n7771)
         );
  NOR2_X1 U9427 ( .A1(n9735), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8532) );
  INV_X1 U9428 ( .A(n8532), .ZN(n7770) );
  OAI211_X1 U9429 ( .C1(n8851), .C2(n8483), .A(n7771), .B(n7770), .ZN(n7772)
         );
  AOI21_X1 U9430 ( .B1(n8938), .B2(n8459), .A(n7772), .ZN(n7773) );
  OAI21_X1 U9431 ( .B1(n7774), .B2(n8477), .A(n7773), .ZN(P2_U3228) );
  OR2_X1 U9432 ( .A1(n7775), .A2(n8493), .ZN(n7776) );
  XNOR2_X1 U9433 ( .A(n8605), .B(n8604), .ZN(n9799) );
  INV_X1 U9434 ( .A(n9799), .ZN(n7789) );
  XNOR2_X1 U9435 ( .A(n7779), .B(n7778), .ZN(n7780) );
  OAI222_X1 U9436 ( .A1(n8838), .A2(n8820), .B1(n8840), .B2(n7781), .C1(n8817), 
        .C2(n7780), .ZN(n9797) );
  INV_X1 U9437 ( .A(n8603), .ZN(n9795) );
  OAI21_X1 U9438 ( .B1(n7782), .B2(n9795), .A(n8855), .ZN(n9796) );
  OAI22_X1 U9439 ( .A1(n8831), .A2(n7784), .B1(n7783), .B2(n8852), .ZN(n7785)
         );
  AOI21_X1 U9440 ( .B1(n8854), .B2(n8603), .A(n7785), .ZN(n7786) );
  OAI21_X1 U9441 ( .B1(n9796), .B2(n8601), .A(n7786), .ZN(n7787) );
  AOI21_X1 U9442 ( .B1(n9797), .B2(n8831), .A(n7787), .ZN(n7788) );
  OAI21_X1 U9443 ( .B1(n8812), .B2(n7789), .A(n7788), .ZN(P2_U3281) );
  NAND2_X1 U9444 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  XOR2_X1 U9445 ( .A(n7793), .B(n7792), .Z(n7800) );
  OAI22_X1 U9446 ( .A1(n9096), .A2(n7794), .B1(n9094), .B2(n7854), .ZN(n7795)
         );
  AOI211_X1 U9447 ( .C1(n9099), .C2(n9114), .A(n7796), .B(n7795), .ZN(n7799)
         );
  NAND2_X1 U9448 ( .A1(n7797), .A2(n6480), .ZN(n7798) );
  OAI211_X1 U9449 ( .C1(n7800), .C2(n9103), .A(n7799), .B(n7798), .ZN(P1_U3213) );
  INV_X1 U9450 ( .A(n7801), .ZN(n7804) );
  INV_X1 U9451 ( .A(n7802), .ZN(n7806) );
  OAI222_X1 U9452 ( .A1(P2_U3152), .A2(n7804), .B1(n8970), .B2(n7806), .C1(
        n7803), .C2(n8963), .ZN(P2_U3332) );
  OAI222_X1 U9453 ( .A1(P1_U3084), .A2(n6331), .B1(n9537), .B2(n7806), .C1(
        n7805), .C2(n8339), .ZN(P1_U3327) );
  INV_X1 U9454 ( .A(n7807), .ZN(n8972) );
  AOI21_X1 U9455 ( .B1(n9535), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7808), .ZN(
        n7809) );
  OAI21_X1 U9456 ( .B1(n8972), .B2(n9537), .A(n7809), .ZN(P1_U3326) );
  XNOR2_X1 U9457 ( .A(n7811), .B(n7810), .ZN(n7812) );
  OAI222_X1 U9458 ( .A1(n9403), .A2(n9013), .B1(n9405), .B2(n9372), .C1(n7812), 
        .C2(n9400), .ZN(n9487) );
  INV_X1 U9459 ( .A(n9487), .ZN(n7820) );
  XNOR2_X1 U9460 ( .A(n7813), .B(n7981), .ZN(n9489) );
  NAND2_X1 U9461 ( .A1(n9489), .A2(n9414), .ZN(n7819) );
  AOI211_X1 U9462 ( .C1(n9017), .C2(n7814), .A(n9390), .B(n9387), .ZN(n9488)
         );
  INV_X1 U9463 ( .A(n9017), .ZN(n9530) );
  NOR2_X1 U9464 ( .A1(n9530), .A2(n9392), .ZN(n7817) );
  OAI22_X1 U9465 ( .A1(n9409), .A2(n7815), .B1(n9014), .B2(n9820), .ZN(n7816)
         );
  AOI211_X1 U9466 ( .C1(n9488), .C2(n9818), .A(n7817), .B(n7816), .ZN(n7818)
         );
  OAI211_X1 U9467 ( .C1(n9826), .C2(n7820), .A(n7819), .B(n7818), .ZN(P1_U3275) );
  MUX2_X1 U9468 ( .A(n9453), .B(n9110), .S(n7948), .Z(n7821) );
  AND2_X1 U9469 ( .A1(n7859), .A2(n8033), .ZN(n7840) );
  INV_X1 U9470 ( .A(n7948), .ZN(n7929) );
  NAND2_X1 U9471 ( .A1(n8024), .A2(n7929), .ZN(n7823) );
  AND2_X1 U9472 ( .A1(n7830), .A2(n8024), .ZN(n8029) );
  INV_X1 U9473 ( .A(n7824), .ZN(n7966) );
  NAND2_X1 U9474 ( .A1(n7966), .A2(n7828), .ZN(n7825) );
  AOI21_X1 U9475 ( .B1(n7829), .B2(n8029), .A(n7825), .ZN(n7827) );
  NAND2_X1 U9476 ( .A1(n7833), .A2(n7826), .ZN(n8093) );
  OAI21_X1 U9477 ( .B1(n7827), .B2(n8093), .A(n8017), .ZN(n7836) );
  NAND2_X1 U9478 ( .A1(n7828), .A2(n8026), .ZN(n7962) );
  INV_X1 U9479 ( .A(n7962), .ZN(n8092) );
  NAND2_X1 U9480 ( .A1(n7829), .A2(n8092), .ZN(n7831) );
  NAND3_X1 U9481 ( .A1(n7831), .A2(n7966), .A3(n7830), .ZN(n7832) );
  NAND3_X1 U9482 ( .A1(n7832), .A2(n8017), .A3(n8091), .ZN(n7834) );
  NAND2_X1 U9483 ( .A1(n7834), .A2(n7833), .ZN(n7835) );
  INV_X1 U9484 ( .A(n7841), .ZN(n7837) );
  OAI211_X1 U9485 ( .C1(n7844), .C2(n7837), .A(n7845), .B(n8016), .ZN(n7838)
         );
  NAND3_X1 U9486 ( .A1(n7838), .A2(n8033), .A3(n7842), .ZN(n7839) );
  MUX2_X1 U9487 ( .A(n7840), .B(n7839), .S(n7929), .Z(n7851) );
  INV_X1 U9488 ( .A(n8016), .ZN(n7843) );
  AND2_X1 U9489 ( .A1(n7842), .A2(n7841), .ZN(n8032) );
  OAI21_X1 U9490 ( .B1(n7844), .B2(n7843), .A(n8032), .ZN(n7846) );
  AND2_X1 U9491 ( .A1(n7848), .A2(n7845), .ZN(n8035) );
  NAND2_X1 U9492 ( .A1(n7846), .A2(n8035), .ZN(n7847) );
  MUX2_X1 U9493 ( .A(n7848), .B(n7847), .S(n7948), .Z(n7850) );
  NAND4_X1 U9494 ( .A1(n7851), .A2(n7850), .A3(n7858), .A4(n7849), .ZN(n7864)
         );
  INV_X1 U9495 ( .A(n7858), .ZN(n7852) );
  OR2_X1 U9496 ( .A1(n7853), .A2(n7852), .ZN(n7855) );
  OR2_X1 U9497 ( .A1(n9830), .A2(n7854), .ZN(n7866) );
  AND2_X1 U9498 ( .A1(n7855), .A2(n7866), .ZN(n8038) );
  AND2_X1 U9499 ( .A1(n8038), .A2(n7869), .ZN(n7862) );
  NAND2_X1 U9500 ( .A1(n7867), .A2(n7856), .ZN(n8015) );
  NAND2_X1 U9501 ( .A1(n7858), .A2(n7857), .ZN(n8037) );
  AND2_X1 U9502 ( .A1(n8037), .A2(n7859), .ZN(n7860) );
  NOR2_X1 U9503 ( .A1(n8015), .A2(n7860), .ZN(n7861) );
  MUX2_X1 U9504 ( .A(n7862), .B(n7861), .S(n7948), .Z(n7863) );
  NAND2_X1 U9505 ( .A1(n7864), .A2(n7863), .ZN(n7873) );
  NAND2_X1 U9506 ( .A1(n7869), .A2(n7866), .ZN(n7868) );
  NAND2_X1 U9507 ( .A1(n7868), .A2(n7867), .ZN(n7871) );
  NAND2_X1 U9508 ( .A1(n8015), .A2(n7869), .ZN(n7870) );
  MUX2_X1 U9509 ( .A(n7871), .B(n7870), .S(n7929), .Z(n7872) );
  NAND3_X1 U9510 ( .A1(n7873), .A2(n4433), .A3(n7872), .ZN(n7875) );
  MUX2_X1 U9511 ( .A(n8046), .B(n8043), .S(n7948), .Z(n7874) );
  NAND3_X1 U9512 ( .A1(n7875), .A2(n7981), .A3(n7874), .ZN(n7877) );
  INV_X1 U9513 ( .A(n8012), .ZN(n7878) );
  MUX2_X1 U9514 ( .A(n8047), .B(n8011), .S(n7929), .Z(n7876) );
  NAND3_X1 U9515 ( .A1(n7877), .A2(n7960), .A3(n7876), .ZN(n7881) );
  AND2_X1 U9516 ( .A1(n8013), .A2(n7878), .ZN(n7879) );
  MUX2_X1 U9517 ( .A(n8000), .B(n7879), .S(n7948), .Z(n7880) );
  NAND2_X1 U9518 ( .A1(n7881), .A2(n7880), .ZN(n7886) );
  AND2_X1 U9519 ( .A1(n8008), .A2(n8013), .ZN(n7995) );
  NAND2_X1 U9520 ( .A1(n7895), .A2(n7883), .ZN(n7996) );
  AOI21_X1 U9521 ( .B1(n7886), .B2(n7995), .A(n7996), .ZN(n7888) );
  AND2_X1 U9522 ( .A1(n7883), .A2(n7882), .ZN(n7885) );
  NAND2_X1 U9523 ( .A1(n7889), .A2(n8008), .ZN(n7884) );
  AOI21_X1 U9524 ( .B1(n7886), .B2(n7885), .A(n7884), .ZN(n7887) );
  MUX2_X1 U9525 ( .A(n7888), .B(n7887), .S(n7948), .Z(n7898) );
  NAND2_X1 U9526 ( .A1(n7898), .A2(n7998), .ZN(n7893) );
  INV_X1 U9527 ( .A(n7889), .ZN(n7890) );
  NAND2_X1 U9528 ( .A1(n7998), .A2(n7890), .ZN(n7891) );
  AND2_X1 U9529 ( .A1(n7891), .A2(n7896), .ZN(n7892) );
  AND2_X1 U9530 ( .A1(n7892), .A2(n7900), .ZN(n7994) );
  NAND2_X1 U9531 ( .A1(n7893), .A2(n7994), .ZN(n7894) );
  NAND2_X1 U9532 ( .A1(n7894), .A2(n8002), .ZN(n7903) );
  INV_X1 U9533 ( .A(n7895), .ZN(n7897) );
  OAI21_X1 U9534 ( .B1(n7898), .B2(n7897), .A(n7896), .ZN(n7899) );
  NAND2_X1 U9535 ( .A1(n7901), .A2(n7900), .ZN(n7902) );
  OAI21_X1 U9536 ( .B1(n9277), .B2(n7905), .A(n7904), .ZN(n7906) );
  NAND2_X1 U9537 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  NAND2_X1 U9538 ( .A1(n7909), .A2(n7908), .ZN(n7923) );
  NAND2_X1 U9539 ( .A1(n7917), .A2(n9261), .ZN(n7910) );
  NAND2_X1 U9540 ( .A1(n8060), .A2(n7910), .ZN(n7913) );
  NAND2_X1 U9541 ( .A1(n9248), .A2(n9237), .ZN(n7911) );
  NAND2_X1 U9542 ( .A1(n8058), .A2(n7911), .ZN(n7912) );
  MUX2_X1 U9543 ( .A(n7913), .B(n7912), .S(n7948), .Z(n7914) );
  INV_X1 U9544 ( .A(n7985), .ZN(n7922) );
  NAND2_X1 U9545 ( .A1(n9237), .A2(n9221), .ZN(n7916) );
  NAND2_X1 U9546 ( .A1(n8055), .A2(n7916), .ZN(n7920) );
  NOR2_X1 U9547 ( .A1(n7917), .A2(n9261), .ZN(n7918) );
  NOR2_X1 U9548 ( .A1(n7918), .A2(n9248), .ZN(n7919) );
  MUX2_X1 U9549 ( .A(n7920), .B(n7919), .S(n7929), .Z(n7921) );
  OAI21_X1 U9550 ( .B1(n7923), .B2(n7922), .A(n7921), .ZN(n7924) );
  NAND2_X1 U9551 ( .A1(n7925), .A2(n7924), .ZN(n7928) );
  MUX2_X1 U9552 ( .A(n8058), .B(n8060), .S(n7948), .Z(n7926) );
  AND2_X1 U9553 ( .A1(n7987), .A2(n7926), .ZN(n7927) );
  NAND2_X1 U9554 ( .A1(n7928), .A2(n7927), .ZN(n7931) );
  MUX2_X1 U9555 ( .A(n8059), .B(n8062), .S(n7929), .Z(n7930) );
  INV_X1 U9556 ( .A(n7944), .ZN(n9106) );
  NOR2_X1 U9557 ( .A1(n7932), .A2(n9106), .ZN(n7933) );
  MUX2_X1 U9558 ( .A(n7948), .B(n7933), .S(n9206), .Z(n7952) );
  NAND2_X1 U9559 ( .A1(n8959), .A2(n7936), .ZN(n7935) );
  NAND2_X1 U9560 ( .A1(n6456), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7934) );
  NAND2_X1 U9561 ( .A1(n8134), .A2(n7936), .ZN(n7938) );
  NAND2_X1 U9562 ( .A1(n6456), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7937) );
  INV_X1 U9563 ( .A(n9105), .ZN(n7940) );
  OR2_X1 U9564 ( .A1(n9188), .A2(n7940), .ZN(n7991) );
  NAND2_X1 U9565 ( .A1(n7991), .A2(n9192), .ZN(n7939) );
  AND2_X1 U9566 ( .A1(n9189), .A2(n7939), .ZN(n7946) );
  INV_X1 U9567 ( .A(n7946), .ZN(n8068) );
  NAND2_X1 U9568 ( .A1(n9188), .A2(n7940), .ZN(n8112) );
  INV_X1 U9569 ( .A(n9192), .ZN(n7942) );
  NAND2_X1 U9570 ( .A1(n9188), .A2(n7942), .ZN(n7941) );
  NAND2_X1 U9571 ( .A1(n8112), .A2(n7941), .ZN(n7945) );
  INV_X1 U9572 ( .A(n7945), .ZN(n8064) );
  OAI211_X1 U9573 ( .C1(n7948), .C2(n7944), .A(n8068), .B(n8064), .ZN(n7951)
         );
  NAND2_X1 U9574 ( .A1(n9189), .A2(n7942), .ZN(n7992) );
  OAI21_X1 U9575 ( .B1(n7943), .B2(n7945), .A(n7992), .ZN(n7950) );
  NOR2_X1 U9576 ( .A1(n7947), .A2(n7946), .ZN(n7949) );
  NAND2_X1 U9577 ( .A1(n6349), .A2(n6350), .ZN(n7954) );
  INV_X1 U9578 ( .A(n8112), .ZN(n7990) );
  INV_X1 U9579 ( .A(n7958), .ZN(n8100) );
  NAND2_X1 U9580 ( .A1(n8100), .A2(n8003), .ZN(n9290) );
  NOR2_X1 U9581 ( .A1(n7962), .A2(n7961), .ZN(n7963) );
  NAND4_X1 U9582 ( .A1(n7965), .A2(n7964), .A3(n7963), .A4(n8029), .ZN(n7971)
         );
  NAND2_X1 U9583 ( .A1(n7967), .A2(n7966), .ZN(n7970) );
  NOR4_X1 U9584 ( .A1(n7971), .A2(n7970), .A3(n7969), .A4(n7968), .ZN(n7974)
         );
  NAND3_X1 U9585 ( .A1(n7974), .A2(n7973), .A3(n7972), .ZN(n7975) );
  NOR4_X1 U9586 ( .A1(n7978), .A2(n7977), .A3(n7976), .A4(n7975), .ZN(n7980)
         );
  NAND4_X1 U9587 ( .A1(n7981), .A2(n4433), .A3(n7980), .A4(n7979), .ZN(n7982)
         );
  NOR4_X1 U9588 ( .A1(n9362), .A2(n9375), .A3(n9398), .A4(n7982), .ZN(n7983)
         );
  NAND4_X1 U9589 ( .A1(n9304), .A2(n9318), .A3(n9345), .A4(n7983), .ZN(n7984)
         );
  NOR4_X1 U9590 ( .A1(n9257), .A2(n9277), .A3(n9290), .A4(n7984), .ZN(n7986)
         );
  OR2_X1 U9591 ( .A1(n7985), .A2(n4326), .ZN(n9239) );
  NAND4_X1 U9592 ( .A1(n7987), .A2(n9225), .A3(n7986), .A4(n9239), .ZN(n7988)
         );
  NOR4_X1 U9593 ( .A1(n8119), .A2(n7990), .A3(n7989), .A4(n7988), .ZN(n7993)
         );
  AND2_X1 U9594 ( .A1(n7992), .A2(n7991), .ZN(n8075) );
  AOI21_X1 U9595 ( .B1(n7993), .B2(n8075), .A(n6350), .ZN(n8072) );
  INV_X1 U9596 ( .A(n7994), .ZN(n8010) );
  INV_X1 U9597 ( .A(n7995), .ZN(n7999) );
  INV_X1 U9598 ( .A(n7996), .ZN(n7997) );
  OAI211_X1 U9599 ( .C1(n8000), .C2(n7999), .A(n7998), .B(n7997), .ZN(n8001)
         );
  INV_X1 U9600 ( .A(n8001), .ZN(n8004) );
  OAI211_X1 U9601 ( .C1(n8010), .C2(n8004), .A(n8003), .B(n8002), .ZN(n8005)
         );
  NAND2_X1 U9602 ( .A1(n8100), .A2(n8005), .ZN(n8007) );
  AND2_X1 U9603 ( .A1(n8007), .A2(n8006), .ZN(n8105) );
  INV_X1 U9604 ( .A(n8008), .ZN(n8009) );
  NOR2_X1 U9605 ( .A1(n8010), .A2(n8009), .ZN(n8101) );
  NOR2_X1 U9606 ( .A1(n8012), .A2(n4798), .ZN(n8014) );
  NAND2_X1 U9607 ( .A1(n8014), .A2(n8013), .ZN(n8049) );
  INV_X1 U9608 ( .A(n8015), .ZN(n8039) );
  INV_X1 U9609 ( .A(n8037), .ZN(n8021) );
  INV_X1 U9610 ( .A(n8035), .ZN(n8019) );
  NAND2_X1 U9611 ( .A1(n8017), .A2(n8016), .ZN(n8018) );
  NOR2_X1 U9612 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND4_X1 U9613 ( .A1(n8043), .A2(n8039), .A3(n8021), .A4(n8020), .ZN(n8022)
         );
  OR2_X1 U9614 ( .A1(n8049), .A2(n8022), .ZN(n8077) );
  AND2_X1 U9615 ( .A1(n8024), .A2(n8023), .ZN(n8087) );
  NAND3_X1 U9616 ( .A1(n8025), .A2(n8087), .A3(n8094), .ZN(n8031) );
  NAND2_X1 U9617 ( .A1(n8026), .A2(n8089), .ZN(n8028) );
  AOI21_X1 U9618 ( .B1(n8029), .B2(n8028), .A(n8027), .ZN(n8030) );
  AOI21_X1 U9619 ( .B1(n8031), .B2(n8030), .A(n8093), .ZN(n8050) );
  INV_X1 U9620 ( .A(n8032), .ZN(n8034) );
  AOI21_X1 U9621 ( .B1(n8035), .B2(n8034), .A(n4786), .ZN(n8036) );
  NOR2_X1 U9622 ( .A1(n8037), .A2(n8036), .ZN(n8041) );
  INV_X1 U9623 ( .A(n8038), .ZN(n8040) );
  OAI211_X1 U9624 ( .C1(n8041), .C2(n8040), .A(n8043), .B(n8039), .ZN(n8045)
         );
  NAND2_X1 U9625 ( .A1(n8043), .A2(n8042), .ZN(n8044) );
  AND4_X1 U9626 ( .A1(n8047), .A2(n8046), .A3(n8045), .A4(n8044), .ZN(n8048)
         );
  OR2_X1 U9627 ( .A1(n8049), .A2(n8048), .ZN(n8076) );
  OAI21_X1 U9628 ( .B1(n8077), .B2(n8050), .A(n8076), .ZN(n8051) );
  NAND3_X1 U9629 ( .A1(n8100), .A2(n8101), .A3(n8051), .ZN(n8052) );
  NAND2_X1 U9630 ( .A1(n8105), .A2(n8052), .ZN(n8053) );
  NAND2_X1 U9631 ( .A1(n8107), .A2(n8053), .ZN(n8054) );
  AND2_X1 U9632 ( .A1(n8109), .A2(n8054), .ZN(n8061) );
  INV_X1 U9633 ( .A(n8055), .ZN(n8056) );
  NAND2_X1 U9634 ( .A1(n8060), .A2(n8056), .ZN(n8057) );
  NAND3_X1 U9635 ( .A1(n8059), .A2(n8058), .A3(n8057), .ZN(n8110) );
  AOI21_X1 U9636 ( .B1(n8061), .B2(n8060), .A(n8110), .ZN(n8065) );
  NAND2_X1 U9637 ( .A1(n8063), .A2(n8062), .ZN(n8114) );
  OAI211_X1 U9638 ( .C1(n8065), .C2(n8114), .A(n8064), .B(n8113), .ZN(n8067)
         );
  NOR2_X1 U9639 ( .A1(n8072), .A2(n8069), .ZN(n8071) );
  MUX2_X1 U9640 ( .A(n8072), .B(n8071), .S(n8070), .Z(n8073) );
  INV_X1 U9641 ( .A(n8075), .ZN(n8118) );
  INV_X1 U9642 ( .A(n8076), .ZN(n8103) );
  INV_X1 U9643 ( .A(n8077), .ZN(n8099) );
  INV_X1 U9644 ( .A(n8078), .ZN(n8081) );
  NAND2_X1 U9645 ( .A1(n5771), .A2(n8079), .ZN(n8080) );
  NAND3_X1 U9646 ( .A1(n8081), .A2(n6350), .A3(n8080), .ZN(n8083) );
  NAND2_X1 U9647 ( .A1(n8083), .A2(n8082), .ZN(n8085) );
  OAI21_X1 U9648 ( .B1(n8086), .B2(n8085), .A(n8084), .ZN(n8090) );
  INV_X1 U9649 ( .A(n8087), .ZN(n8088) );
  AOI21_X1 U9650 ( .B1(n8090), .B2(n8089), .A(n8088), .ZN(n8097) );
  NAND2_X1 U9651 ( .A1(n8092), .A2(n8091), .ZN(n8096) );
  INV_X1 U9652 ( .A(n8093), .ZN(n8095) );
  OAI211_X1 U9653 ( .C1(n8097), .C2(n8096), .A(n8095), .B(n8094), .ZN(n8098)
         );
  AND2_X1 U9654 ( .A1(n8099), .A2(n8098), .ZN(n8102) );
  OAI211_X1 U9655 ( .C1(n8103), .C2(n8102), .A(n8101), .B(n8100), .ZN(n8104)
         );
  NAND2_X1 U9656 ( .A1(n8105), .A2(n8104), .ZN(n8106) );
  NAND2_X1 U9657 ( .A1(n8107), .A2(n8106), .ZN(n8108) );
  AND3_X1 U9658 ( .A1(n9225), .A2(n8109), .A3(n8108), .ZN(n8111) );
  NOR2_X1 U9659 ( .A1(n8111), .A2(n8110), .ZN(n8115) );
  OAI211_X1 U9660 ( .C1(n8115), .C2(n8114), .A(n8113), .B(n8112), .ZN(n8116)
         );
  INV_X1 U9661 ( .A(n8116), .ZN(n8117) );
  OR2_X1 U9662 ( .A1(n8118), .A2(n8117), .ZN(n8120) );
  NAND2_X1 U9663 ( .A1(n8120), .A2(n7956), .ZN(n8125) );
  INV_X1 U9664 ( .A(n8121), .ZN(n8124) );
  NAND3_X1 U9665 ( .A1(n8125), .A2(n9184), .A3(n8122), .ZN(n8123) );
  OAI211_X1 U9666 ( .C1(n8125), .C2(n8124), .A(n8123), .B(n8126), .ZN(n8130)
         );
  INV_X1 U9667 ( .A(n8126), .ZN(n8128) );
  NAND4_X1 U9668 ( .A1(n4378), .A2(n9861), .A3(n9858), .A4(n9966), .ZN(n8127)
         );
  OAI211_X1 U9669 ( .C1(n5753), .C2(n8128), .A(n8127), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8129) );
  INV_X1 U9670 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8133) );
  INV_X1 U9671 ( .A(n8132), .ZN(n8965) );
  OAI222_X1 U9672 ( .A1(n8339), .A2(n8133), .B1(P1_U3084), .B2(n8131), .C1(
        n9537), .C2(n8965), .ZN(P1_U3324) );
  INV_X1 U9673 ( .A(n8134), .ZN(n8341) );
  OAI222_X1 U9674 ( .A1(n8970), .A2(n8341), .B1(P2_U3152), .B2(n8136), .C1(
        n8135), .C2(n8963), .ZN(P2_U3328) );
  OAI211_X1 U9675 ( .C1(n8139), .C2(n8138), .A(n9997), .B(n8137), .ZN(n8148)
         );
  OAI21_X1 U9676 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8146) );
  NOR2_X1 U9677 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8143), .ZN(n8397) );
  INV_X1 U9678 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8144) );
  NOR2_X1 U9679 ( .A1(n8587), .A2(n8144), .ZN(n8145) );
  AOI211_X1 U9680 ( .C1(n9995), .C2(n8146), .A(n8397), .B(n8145), .ZN(n8147)
         );
  OAI211_X1 U9681 ( .C1(n9998), .C2(n8149), .A(n8148), .B(n8147), .ZN(P2_U3257) );
  NOR2_X1 U9682 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9725), .ZN(n8154) );
  AOI211_X1 U9683 ( .C1(n8152), .C2(n8151), .A(n8150), .B(n10000), .ZN(n8153)
         );
  AOI211_X1 U9684 ( .C1(n10002), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n8154), .B(
        n8153), .ZN(n8159) );
  OAI211_X1 U9685 ( .C1(n8157), .C2(n8156), .A(n9997), .B(n8155), .ZN(n8158)
         );
  OAI211_X1 U9686 ( .C1(n9998), .C2(n8160), .A(n8159), .B(n8158), .ZN(P2_U3255) );
  AOI211_X1 U9687 ( .C1(n8163), .C2(n8162), .A(n8161), .B(n10000), .ZN(n8164)
         );
  AOI211_X1 U9688 ( .C1(n10002), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n8165), .B(
        n8164), .ZN(n8170) );
  OAI211_X1 U9689 ( .C1(n8168), .C2(n8167), .A(n9997), .B(n8166), .ZN(n8169)
         );
  OAI211_X1 U9690 ( .C1(n9998), .C2(n8171), .A(n8170), .B(n8169), .ZN(P2_U3254) );
  NOR2_X1 U9691 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9719), .ZN(n8176) );
  AOI211_X1 U9692 ( .C1(n8174), .C2(n8173), .A(n8172), .B(n10000), .ZN(n8175)
         );
  AOI211_X1 U9693 ( .C1(n10002), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n8176), .B(
        n8175), .ZN(n8181) );
  OAI211_X1 U9694 ( .C1(n8179), .C2(n8178), .A(n9997), .B(n8177), .ZN(n8180)
         );
  OAI211_X1 U9695 ( .C1(n9998), .C2(n8182), .A(n8181), .B(n8180), .ZN(P2_U3253) );
  AOI211_X1 U9696 ( .C1(n8185), .C2(n8184), .A(n8183), .B(n10000), .ZN(n8186)
         );
  AOI211_X1 U9697 ( .C1(n10002), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n8187), .B(
        n8186), .ZN(n8192) );
  OAI211_X1 U9698 ( .C1(n8190), .C2(n8189), .A(n9997), .B(n8188), .ZN(n8191)
         );
  OAI211_X1 U9699 ( .C1(n9998), .C2(n8193), .A(n8192), .B(n8191), .ZN(P2_U3252) );
  AOI211_X1 U9700 ( .C1(n8196), .C2(n8195), .A(n8194), .B(n10000), .ZN(n8197)
         );
  AOI211_X1 U9701 ( .C1(n10002), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n8198), .B(
        n8197), .ZN(n8203) );
  OAI211_X1 U9702 ( .C1(n8201), .C2(n8200), .A(n9997), .B(n8199), .ZN(n8202)
         );
  OAI211_X1 U9703 ( .C1(n9998), .C2(n8204), .A(n8203), .B(n8202), .ZN(P2_U3251) );
  NOR2_X1 U9704 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5016), .ZN(n8209) );
  AOI211_X1 U9705 ( .C1(n8207), .C2(n8206), .A(n8205), .B(n10000), .ZN(n8208)
         );
  AOI211_X1 U9706 ( .C1(n10002), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n8209), .B(
        n8208), .ZN(n8214) );
  OAI211_X1 U9707 ( .C1(n8212), .C2(n8211), .A(n9997), .B(n8210), .ZN(n8213)
         );
  OAI211_X1 U9708 ( .C1(n9998), .C2(n8215), .A(n8214), .B(n8213), .ZN(P2_U3250) );
  AOI211_X1 U9709 ( .C1(n8218), .C2(n8217), .A(n8216), .B(n10000), .ZN(n8219)
         );
  AOI211_X1 U9710 ( .C1(n10002), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n8220), .B(
        n8219), .ZN(n8225) );
  OAI211_X1 U9711 ( .C1(n8223), .C2(n8222), .A(n9997), .B(n8221), .ZN(n8224)
         );
  OAI211_X1 U9712 ( .C1(n9998), .C2(n8226), .A(n8225), .B(n8224), .ZN(P2_U3249) );
  INV_X1 U9713 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9706) );
  NOR2_X1 U9714 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9706), .ZN(n8231) );
  AOI211_X1 U9715 ( .C1(n8229), .C2(n8228), .A(n8227), .B(n10000), .ZN(n8230)
         );
  AOI211_X1 U9716 ( .C1(n10002), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n8231), .B(
        n8230), .ZN(n8236) );
  OAI211_X1 U9717 ( .C1(n8234), .C2(n8233), .A(n9997), .B(n8232), .ZN(n8235)
         );
  OAI211_X1 U9718 ( .C1(n9998), .C2(n8237), .A(n8236), .B(n8235), .ZN(P2_U3248) );
  NAND2_X1 U9719 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n8240) );
  AOI211_X1 U9720 ( .C1(n8240), .C2(n8239), .A(n8238), .B(n10000), .ZN(n8242)
         );
  INV_X1 U9721 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10125) );
  OAI22_X1 U9722 ( .A1(n8587), .A2(n10125), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9699), .ZN(n8241) );
  NOR2_X1 U9723 ( .A1(n8242), .A2(n8241), .ZN(n8247) );
  NOR2_X1 U9724 ( .A1(n10005), .A2(n9996), .ZN(n8245) );
  MUX2_X1 U9725 ( .A(n7052), .B(P2_REG2_REG_1__SCAN_IN), .S(n8248), .Z(n8244)
         );
  OAI211_X1 U9726 ( .C1(n8245), .C2(n8244), .A(n9997), .B(n8243), .ZN(n8246)
         );
  OAI211_X1 U9727 ( .C1(n9998), .C2(n8248), .A(n8247), .B(n8246), .ZN(P2_U3246) );
  XNOR2_X1 U9728 ( .A(n8250), .B(n8249), .ZN(n8252) );
  NAND2_X1 U9729 ( .A1(n8459), .A2(n4996), .ZN(n8251) );
  OAI21_X1 U9730 ( .B1(n8477), .B2(n8252), .A(n8251), .ZN(n8253) );
  AOI21_X1 U9731 ( .B1(n8460), .B2(n8503), .A(n8253), .ZN(n8255) );
  MUX2_X1 U9732 ( .A(n8483), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n8254) );
  OAI211_X1 U9733 ( .C1(n8256), .C2(n8485), .A(n8255), .B(n8254), .ZN(P2_U3220) );
  OAI222_X1 U9734 ( .A1(n8963), .A2(n8259), .B1(n8973), .B2(n8258), .C1(n8257), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  NOR2_X1 U9735 ( .A1(n8632), .A2(n8319), .ZN(n8260) );
  XNOR2_X1 U9736 ( .A(n8260), .B(n8318), .ZN(n8326) );
  INV_X1 U9737 ( .A(n8326), .ZN(n8327) );
  NOR3_X1 U9738 ( .A1(n8620), .A2(n8459), .A3(n8327), .ZN(n8261) );
  AOI21_X1 U9739 ( .B1(n8620), .B2(n8327), .A(n8261), .ZN(n8333) );
  INV_X1 U9740 ( .A(n8262), .ZN(n8265) );
  INV_X1 U9741 ( .A(n8263), .ZN(n8264) );
  NAND2_X1 U9742 ( .A1(n8265), .A2(n8264), .ZN(n8266) );
  XNOR2_X1 U9743 ( .A(n8934), .B(n8318), .ZN(n8268) );
  NOR2_X1 U9744 ( .A1(n8839), .A2(n8319), .ZN(n8269) );
  NAND2_X1 U9745 ( .A1(n8268), .A2(n8269), .ZN(n8272) );
  INV_X1 U9746 ( .A(n8268), .ZN(n8468) );
  INV_X1 U9747 ( .A(n8269), .ZN(n8270) );
  NAND2_X1 U9748 ( .A1(n8468), .A2(n8270), .ZN(n8271) );
  NAND2_X1 U9749 ( .A1(n8272), .A2(n8271), .ZN(n8413) );
  NAND2_X1 U9750 ( .A1(n8467), .A2(n8272), .ZN(n8277) );
  XNOR2_X1 U9751 ( .A(n8929), .B(n8318), .ZN(n8273) );
  AND2_X1 U9752 ( .A1(n8788), .A2(n8295), .ZN(n8274) );
  NAND2_X1 U9753 ( .A1(n8273), .A2(n8274), .ZN(n8278) );
  INV_X1 U9754 ( .A(n8273), .ZN(n8366) );
  INV_X1 U9755 ( .A(n8274), .ZN(n8275) );
  NAND2_X1 U9756 ( .A1(n8366), .A2(n8275), .ZN(n8276) );
  AND2_X1 U9757 ( .A1(n8278), .A2(n8276), .ZN(n8465) );
  XNOR2_X1 U9758 ( .A(n8925), .B(n8318), .ZN(n8280) );
  NAND2_X1 U9759 ( .A1(n8807), .A2(n8309), .ZN(n8281) );
  XNOR2_X1 U9760 ( .A(n8280), .B(n8281), .ZN(n8367) );
  AND2_X1 U9761 ( .A1(n8367), .A2(n8278), .ZN(n8279) );
  INV_X1 U9762 ( .A(n8280), .ZN(n8282) );
  NAND2_X1 U9763 ( .A1(n8282), .A2(n8281), .ZN(n8283) );
  XNOR2_X1 U9764 ( .A(n8919), .B(n8318), .ZN(n8284) );
  NOR2_X1 U9765 ( .A1(n8610), .A2(n8319), .ZN(n8285) );
  NAND2_X1 U9766 ( .A1(n8284), .A2(n8285), .ZN(n8289) );
  INV_X1 U9767 ( .A(n8284), .ZN(n8378) );
  INV_X1 U9768 ( .A(n8285), .ZN(n8286) );
  NAND2_X1 U9769 ( .A1(n8378), .A2(n8286), .ZN(n8287) );
  NAND2_X1 U9770 ( .A1(n8289), .A2(n8287), .ZN(n8434) );
  XNOR2_X1 U9771 ( .A(n8755), .B(n8318), .ZN(n8291) );
  NOR2_X1 U9772 ( .A1(n8611), .A2(n8319), .ZN(n8292) );
  XNOR2_X1 U9773 ( .A(n8291), .B(n8292), .ZN(n8376) );
  INV_X1 U9774 ( .A(n8291), .ZN(n8293) );
  NAND2_X1 U9775 ( .A1(n8293), .A2(n8292), .ZN(n8294) );
  NAND2_X1 U9776 ( .A1(n8379), .A2(n8294), .ZN(n8296) );
  XNOR2_X1 U9777 ( .A(n8907), .B(n8308), .ZN(n8297) );
  XNOR2_X1 U9778 ( .A(n8296), .B(n8297), .ZN(n8442) );
  NAND2_X1 U9779 ( .A1(n8758), .A2(n8295), .ZN(n8440) );
  NAND2_X1 U9780 ( .A1(n8442), .A2(n8440), .ZN(n8300) );
  INV_X1 U9781 ( .A(n8296), .ZN(n8298) );
  NAND2_X1 U9782 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  XNOR2_X1 U9783 ( .A(n8902), .B(n8318), .ZN(n8305) );
  XNOR2_X1 U9784 ( .A(n8897), .B(n8318), .ZN(n8421) );
  NOR2_X1 U9785 ( .A1(n8713), .A2(n8319), .ZN(n8356) );
  INV_X1 U9786 ( .A(n8301), .ZN(n8303) );
  INV_X1 U9787 ( .A(n8421), .ZN(n8302) );
  NOR2_X1 U9788 ( .A1(n8423), .A2(n8319), .ZN(n8306) );
  INV_X1 U9789 ( .A(n8306), .ZN(n8425) );
  OAI21_X1 U9790 ( .B1(n8306), .B2(n8421), .A(n8418), .ZN(n8307) );
  XNOR2_X1 U9791 ( .A(n8893), .B(n8308), .ZN(n8476) );
  NAND2_X1 U9792 ( .A1(n8614), .A2(n8309), .ZN(n8310) );
  NOR2_X1 U9793 ( .A1(n8476), .A2(n8310), .ZN(n8311) );
  AOI21_X1 U9794 ( .B1(n8476), .B2(n8310), .A(n8311), .ZN(n8402) );
  INV_X1 U9795 ( .A(n8311), .ZN(n8316) );
  XNOR2_X1 U9796 ( .A(n8888), .B(n8318), .ZN(n8312) );
  NOR2_X1 U9797 ( .A1(n8404), .A2(n8319), .ZN(n8313) );
  NAND2_X1 U9798 ( .A1(n8312), .A2(n8313), .ZN(n8317) );
  INV_X1 U9799 ( .A(n8312), .ZN(n8348) );
  INV_X1 U9800 ( .A(n8313), .ZN(n8314) );
  NAND2_X1 U9801 ( .A1(n8348), .A2(n8314), .ZN(n8315) );
  NAND2_X1 U9802 ( .A1(n8317), .A2(n8315), .ZN(n8478) );
  XNOR2_X1 U9803 ( .A(n8881), .B(n8318), .ZN(n8320) );
  NOR2_X1 U9804 ( .A1(n8681), .A2(n8319), .ZN(n8321) );
  NAND2_X1 U9805 ( .A1(n8320), .A2(n8321), .ZN(n8325) );
  INV_X1 U9806 ( .A(n8320), .ZN(n8323) );
  INV_X1 U9807 ( .A(n8321), .ZN(n8322) );
  NAND2_X1 U9808 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  AND2_X1 U9809 ( .A1(n8325), .A2(n8324), .ZN(n8346) );
  NOR3_X1 U9810 ( .A1(n8620), .A2(n8326), .A3(n8459), .ZN(n8329) );
  NOR2_X1 U9811 ( .A1(n8876), .A2(n8327), .ZN(n8328) );
  OAI21_X1 U9812 ( .B1(n8620), .B2(n8490), .A(n8477), .ZN(n8330) );
  OAI211_X1 U9813 ( .C1(n8333), .C2(n8332), .A(n8331), .B(n8330), .ZN(n8337)
         );
  NAND2_X1 U9814 ( .A1(n8491), .A2(n8806), .ZN(n8334) );
  OAI21_X1 U9815 ( .B1(n8681), .B2(n8840), .A(n8334), .ZN(n8638) );
  AOI22_X1 U9816 ( .A1(n8335), .A2(n8638), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8336) );
  OAI211_X1 U9817 ( .C1(n8645), .C2(n8483), .A(n8337), .B(n8336), .ZN(P2_U3222) );
  INV_X1 U9818 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8340) );
  OAI222_X1 U9819 ( .A1(n9537), .A2(n8341), .B1(P1_U3084), .B2(n8338), .C1(
        n8340), .C2(n8339), .ZN(P1_U3323) );
  OAI222_X1 U9820 ( .A1(n8963), .A2(n8344), .B1(n8973), .B2(n8343), .C1(
        P2_U3152), .C2(n8342), .ZN(P2_U3336) );
  INV_X1 U9821 ( .A(n8345), .ZN(n8480) );
  INV_X1 U9822 ( .A(n8346), .ZN(n8347) );
  NOR3_X1 U9823 ( .A1(n8348), .A2(n8404), .A3(n8475), .ZN(n8350) );
  OAI21_X1 U9824 ( .B1(n8351), .B2(n8350), .A(n8349), .ZN(n8355) );
  AOI22_X1 U9825 ( .A1(n8472), .A2(n8656), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8354) );
  AOI22_X1 U9826 ( .A1(n8460), .A2(n8660), .B1(n8461), .B2(n8661), .ZN(n8353)
         );
  NAND2_X1 U9827 ( .A1(n8881), .A2(n8459), .ZN(n8352) );
  NAND4_X1 U9828 ( .A1(n8355), .A2(n8354), .A3(n8353), .A4(n8352), .ZN(
        P2_U3216) );
  INV_X1 U9829 ( .A(n8713), .ZN(n8744) );
  AOI22_X1 U9830 ( .A1(n8357), .A2(n8441), .B1(n8439), .B2(n8744), .ZN(n8363)
         );
  NAND2_X1 U9831 ( .A1(n8357), .A2(n8356), .ZN(n8420) );
  INV_X1 U9832 ( .A(n8420), .ZN(n8362) );
  INV_X1 U9833 ( .A(n8724), .ZN(n8358) );
  OAI22_X1 U9834 ( .A1(n8483), .A2(n8358), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9724), .ZN(n8360) );
  INV_X1 U9835 ( .A(n8460), .ZN(n8484) );
  OAI22_X1 U9836 ( .A1(n8423), .A2(n8484), .B1(n8485), .B2(n8612), .ZN(n8359)
         );
  AOI211_X1 U9837 ( .C1(n8902), .C2(n8459), .A(n8360), .B(n8359), .ZN(n8361)
         );
  OAI21_X1 U9838 ( .B1(n8363), .B2(n8362), .A(n8361), .ZN(P2_U3218) );
  OAI21_X1 U9839 ( .B1(n8367), .B2(n8364), .A(n8365), .ZN(n8374) );
  NOR3_X1 U9840 ( .A1(n8367), .A2(n8366), .A3(n8475), .ZN(n8368) );
  OAI21_X1 U9841 ( .B1(n8368), .B2(n8461), .A(n8788), .ZN(n8372) );
  INV_X1 U9842 ( .A(n8610), .ZN(n8789) );
  NAND2_X1 U9843 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8585) );
  OAI21_X1 U9844 ( .B1(n8483), .B2(n8369), .A(n8585), .ZN(n8370) );
  AOI21_X1 U9845 ( .B1(n8460), .B2(n8789), .A(n8370), .ZN(n8371) );
  OAI211_X1 U9846 ( .C1(n8784), .C2(n8490), .A(n8372), .B(n8371), .ZN(n8373)
         );
  AOI21_X1 U9847 ( .B1(n8374), .B2(n8441), .A(n8373), .ZN(n8375) );
  INV_X1 U9848 ( .A(n8375), .ZN(P2_U3221) );
  INV_X1 U9849 ( .A(n8376), .ZN(n8377) );
  AOI21_X1 U9850 ( .B1(n8431), .B2(n8377), .A(n8477), .ZN(n8381) );
  NOR3_X1 U9851 ( .A1(n8378), .A2(n8610), .A3(n8475), .ZN(n8380) );
  OAI21_X1 U9852 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8385) );
  AOI22_X1 U9853 ( .A1(n8472), .A2(n8753), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8384) );
  AOI22_X1 U9854 ( .A1(n8461), .A2(n8789), .B1(n8460), .B2(n8758), .ZN(n8383)
         );
  NAND2_X1 U9855 ( .A1(n8912), .A2(n8459), .ZN(n8382) );
  NAND4_X1 U9856 ( .A1(n8385), .A2(n8384), .A3(n8383), .A4(n8382), .ZN(
        P2_U3225) );
  AND2_X1 U9857 ( .A1(n8387), .A2(n8386), .ZN(n8453) );
  INV_X1 U9858 ( .A(n8388), .ZN(n8389) );
  AOI21_X1 U9859 ( .B1(n8453), .B2(n8389), .A(n8477), .ZN(n8394) );
  NOR3_X1 U9860 ( .A1(n8475), .A2(n8391), .A3(n8390), .ZN(n8393) );
  OAI21_X1 U9861 ( .B1(n8394), .B2(n8393), .A(n8392), .ZN(n8401) );
  NOR2_X1 U9862 ( .A1(n8483), .A2(n8395), .ZN(n8396) );
  AOI211_X1 U9863 ( .C1(n8398), .C2(n8459), .A(n8397), .B(n8396), .ZN(n8400)
         );
  AOI22_X1 U9864 ( .A1(n8460), .A2(n8494), .B1(n8461), .B2(n8496), .ZN(n8399)
         );
  NAND3_X1 U9865 ( .A1(n8401), .A2(n8400), .A3(n8399), .ZN(P2_U3226) );
  INV_X1 U9866 ( .A(n8893), .ZN(n8696) );
  OAI211_X1 U9867 ( .C1(n8403), .C2(n8402), .A(n8479), .B(n8441), .ZN(n8409)
         );
  OAI22_X1 U9868 ( .A1(n8404), .A2(n8838), .B1(n8423), .B2(n8840), .ZN(n8688)
         );
  INV_X1 U9869 ( .A(n8688), .ZN(n8405) );
  OAI22_X1 U9870 ( .A1(n8406), .A2(n8405), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9712), .ZN(n8407) );
  AOI21_X1 U9871 ( .B1(n8693), .B2(n8472), .A(n8407), .ZN(n8408) );
  OAI211_X1 U9872 ( .C1(n8696), .C2(n8490), .A(n8409), .B(n8408), .ZN(P2_U3227) );
  AOI22_X1 U9873 ( .A1(n8460), .A2(n8788), .B1(n8461), .B2(n8606), .ZN(n8411)
         );
  NOR2_X1 U9874 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9691), .ZN(n8543) );
  INV_X1 U9875 ( .A(n8543), .ZN(n8410) );
  OAI211_X1 U9876 ( .C1(n8483), .C2(n8829), .A(n8411), .B(n8410), .ZN(n8416)
         );
  INV_X1 U9877 ( .A(n8467), .ZN(n8412) );
  AOI211_X1 U9878 ( .C1(n8414), .C2(n8413), .A(n8477), .B(n8412), .ZN(n8415)
         );
  AOI211_X1 U9879 ( .C1(n8934), .C2(n8459), .A(n8416), .B(n8415), .ZN(n8417)
         );
  INV_X1 U9880 ( .A(n8417), .ZN(P2_U3230) );
  INV_X1 U9881 ( .A(n8897), .ZN(n8706) );
  INV_X1 U9882 ( .A(n8418), .ZN(n8419) );
  NAND2_X1 U9883 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  XNOR2_X1 U9884 ( .A(n8422), .B(n8421), .ZN(n8426) );
  OAI22_X1 U9885 ( .A1(n8426), .A2(n8477), .B1(n8423), .B2(n8475), .ZN(n8424)
         );
  OAI21_X1 U9886 ( .B1(n8426), .B2(n8425), .A(n8424), .ZN(n8430) );
  OAI22_X1 U9887 ( .A1(n8483), .A2(n8703), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9705), .ZN(n8428) );
  NOR2_X1 U9888 ( .A1(n8485), .A2(n8713), .ZN(n8427) );
  AOI211_X1 U9889 ( .C1(n8460), .C2(n8614), .A(n8428), .B(n8427), .ZN(n8429)
         );
  OAI211_X1 U9890 ( .C1(n8706), .C2(n8490), .A(n8430), .B(n8429), .ZN(P2_U3231) );
  INV_X1 U9891 ( .A(n8431), .ZN(n8432) );
  AOI211_X1 U9892 ( .C1(n8434), .C2(n8433), .A(n8477), .B(n8432), .ZN(n8438)
         );
  AOI22_X1 U9893 ( .A1(n8472), .A2(n8773), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8436) );
  INV_X1 U9894 ( .A(n8611), .ZN(n8765) );
  AOI22_X1 U9895 ( .A1(n8460), .A2(n8765), .B1(n8461), .B2(n8807), .ZN(n8435)
         );
  OAI211_X1 U9896 ( .C1(n8770), .C2(n8490), .A(n8436), .B(n8435), .ZN(n8437)
         );
  OR2_X1 U9897 ( .A1(n8438), .A2(n8437), .ZN(P2_U3235) );
  NAND2_X1 U9898 ( .A1(n8439), .A2(n8758), .ZN(n8444) );
  NAND2_X1 U9899 ( .A1(n8441), .A2(n8440), .ZN(n8443) );
  MUX2_X1 U9900 ( .A(n8444), .B(n8443), .S(n8442), .Z(n8448) );
  NOR2_X1 U9901 ( .A1(n8483), .A2(n8736), .ZN(n8446) );
  OAI22_X1 U9902 ( .A1(n8713), .A2(n8484), .B1(n8485), .B2(n8611), .ZN(n8445)
         );
  AOI211_X1 U9903 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8446), 
        .B(n8445), .ZN(n8447) );
  OAI211_X1 U9904 ( .C1(n8739), .C2(n8490), .A(n8448), .B(n8447), .ZN(P2_U3237) );
  AOI21_X1 U9905 ( .B1(n8450), .B2(n8449), .A(n8477), .ZN(n8455) );
  NOR3_X1 U9906 ( .A1(n8475), .A2(n8452), .A3(n8451), .ZN(n8454) );
  OAI21_X1 U9907 ( .B1(n8455), .B2(n8454), .A(n8453), .ZN(n8464) );
  NOR2_X1 U9908 ( .A1(n8483), .A2(n8456), .ZN(n8457) );
  AOI211_X1 U9909 ( .C1(n10087), .C2(n8459), .A(n8458), .B(n8457), .ZN(n8463)
         );
  AOI22_X1 U9910 ( .A1(n8461), .A2(n8497), .B1(n8460), .B2(n8495), .ZN(n8462)
         );
  NAND3_X1 U9911 ( .A1(n8464), .A2(n8463), .A3(n8462), .ZN(P2_U3238) );
  INV_X1 U9912 ( .A(n8929), .ZN(n8801) );
  INV_X1 U9913 ( .A(n8465), .ZN(n8466) );
  AOI21_X1 U9914 ( .B1(n8467), .B2(n8466), .A(n8477), .ZN(n8470) );
  NOR3_X1 U9915 ( .A1(n8468), .A2(n8839), .A3(n8475), .ZN(n8469) );
  OAI21_X1 U9916 ( .B1(n8470), .B2(n8469), .A(n8364), .ZN(n8474) );
  NOR2_X1 U9917 ( .A1(n9650), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8563) );
  OAI22_X1 U9918 ( .A1(n8839), .A2(n8485), .B1(n8484), .B2(n8609), .ZN(n8471)
         );
  AOI211_X1 U9919 ( .C1(n8472), .C2(n8798), .A(n8563), .B(n8471), .ZN(n8473)
         );
  OAI211_X1 U9920 ( .C1(n8801), .C2(n8490), .A(n8474), .B(n8473), .ZN(P2_U3240) );
  INV_X1 U9921 ( .A(n8888), .ZN(n8671) );
  NOR3_X1 U9922 ( .A1(n8476), .A2(n8714), .A3(n8475), .ZN(n8482) );
  AOI21_X1 U9923 ( .B1(n8479), .B2(n8478), .A(n8477), .ZN(n8481) );
  OAI21_X1 U9924 ( .B1(n8482), .B2(n8481), .A(n8480), .ZN(n8489) );
  NOR2_X1 U9925 ( .A1(n8483), .A2(n8672), .ZN(n8487) );
  OAI22_X1 U9926 ( .A1(n8714), .A2(n8485), .B1(n8484), .B2(n8681), .ZN(n8486)
         );
  AOI211_X1 U9927 ( .C1(P2_REG3_REG_26__SCAN_IN), .C2(P2_U3152), .A(n8487), 
        .B(n8486), .ZN(n8488) );
  OAI211_X1 U9928 ( .C1(n8671), .C2(n8490), .A(n8489), .B(n8488), .ZN(P2_U3242) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8592), .S(P2_U3966), .Z(
        P2_U3583) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8629), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9931 ( .A(n8491), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8492), .Z(
        P2_U3581) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8660), .S(P2_U3966), .Z(
        P2_U3580) );
  INV_X1 U9933 ( .A(n8681), .ZN(n8617) );
  MUX2_X1 U9934 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8617), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9935 ( .A(n8661), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8492), .Z(
        P2_U3578) );
  MUX2_X1 U9936 ( .A(n8614), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8492), .Z(
        P2_U3577) );
  MUX2_X1 U9937 ( .A(n8729), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8492), .Z(
        P2_U3576) );
  MUX2_X1 U9938 ( .A(n8744), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8492), .Z(
        P2_U3575) );
  MUX2_X1 U9939 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8758), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8765), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8789), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8807), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9943 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8788), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U9944 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8805), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8606), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8602), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9947 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8493), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9948 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8494), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8495), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8496), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8497), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U9952 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8498), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U9953 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8499), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8500), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8501), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U9956 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8502), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U9957 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8503), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U9958 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8504), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U9959 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8505), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U9960 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n6730), .S(P2_U3966), .Z(
        P2_U3553) );
  XNOR2_X1 U9961 ( .A(n8519), .B(n8520), .ZN(n8507) );
  INV_X1 U9962 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U9963 ( .A1(n9800), .A2(n8507), .ZN(n8521) );
  AOI211_X1 U9964 ( .C1(n8507), .C2(n9800), .A(n8521), .B(n10000), .ZN(n8518)
         );
  NOR2_X1 U9965 ( .A1(n8508), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8510) );
  NOR2_X1 U9966 ( .A1(n8510), .A2(n8509), .ZN(n8525) );
  XNOR2_X1 U9967 ( .A(n8525), .B(n8526), .ZN(n8511) );
  NOR2_X1 U9968 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8511), .ZN(n8527) );
  AOI21_X1 U9969 ( .B1(n8511), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8527), .ZN(
        n8512) );
  NOR2_X1 U9970 ( .A1(n8512), .A2(n8578), .ZN(n8517) );
  INV_X1 U9971 ( .A(n8513), .ZN(n8514) );
  AOI21_X1 U9972 ( .B1(n10002), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8514), .ZN(
        n8515) );
  OAI21_X1 U9973 ( .B1(n9998), .B2(n8520), .A(n8515), .ZN(n8516) );
  OR3_X1 U9974 ( .A1(n8518), .A2(n8517), .A3(n8516), .ZN(P2_U3260) );
  NOR2_X1 U9975 ( .A1(n8520), .A2(n8519), .ZN(n8522) );
  XNOR2_X1 U9976 ( .A(n8545), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8523) );
  OAI21_X1 U9977 ( .B1(n8524), .B2(n8523), .A(n8546), .ZN(n8536) );
  NOR2_X1 U9978 ( .A1(n8526), .A2(n8525), .ZN(n8528) );
  NOR2_X1 U9979 ( .A1(n8528), .A2(n8527), .ZN(n8531) );
  MUX2_X1 U9980 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n5251), .S(n8545), .Z(n8529)
         );
  INV_X1 U9981 ( .A(n8529), .ZN(n8530) );
  NAND2_X1 U9982 ( .A1(n8530), .A2(n8531), .ZN(n8539) );
  OAI211_X1 U9983 ( .C1(n8531), .C2(n8530), .A(n9997), .B(n8539), .ZN(n8534)
         );
  AOI21_X1 U9984 ( .B1(n10002), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8532), .ZN(
        n8533) );
  OAI211_X1 U9985 ( .C1(n9998), .C2(n8545), .A(n8534), .B(n8533), .ZN(n8535)
         );
  AOI21_X1 U9986 ( .B1(n8536), .B2(n9995), .A(n8535), .ZN(n8537) );
  INV_X1 U9987 ( .A(n8537), .ZN(P2_U3261) );
  NAND2_X1 U9988 ( .A1(n8538), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U9989 ( .A1(n8540), .A2(n8539), .ZN(n8542) );
  XNOR2_X1 U9990 ( .A(n8559), .B(n8830), .ZN(n8541) );
  NAND2_X1 U9991 ( .A1(n8541), .A2(n8542), .ZN(n8555) );
  OAI211_X1 U9992 ( .C1(n8542), .C2(n8541), .A(n9997), .B(n8555), .ZN(n8554)
         );
  AOI21_X1 U9993 ( .B1(n10002), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8543), .ZN(
        n8553) );
  OR2_X1 U9994 ( .A1(n9998), .A2(n8556), .ZN(n8552) );
  XNOR2_X1 U9995 ( .A(n8559), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8549) );
  NAND2_X1 U9996 ( .A1(n8545), .A2(n8544), .ZN(n8547) );
  AOI21_X1 U9997 ( .B1(n8549), .B2(n8548), .A(n8558), .ZN(n8550) );
  NAND2_X1 U9998 ( .A1(n9995), .A2(n8550), .ZN(n8551) );
  NAND4_X1 U9999 ( .A1(n8554), .A2(n8553), .A3(n8552), .A4(n8551), .ZN(
        P2_U3262) );
  OAI21_X1 U10000 ( .B1(n8830), .B2(n8556), .A(n8555), .ZN(n8572) );
  XNOR2_X1 U10001 ( .A(n8573), .B(n8572), .ZN(n8557) );
  NOR2_X1 U10002 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8557), .ZN(n8574) );
  AOI21_X1 U10003 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n8557), .A(n8574), .ZN(
        n8569) );
  INV_X1 U10004 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8560) );
  AOI22_X1 U10005 ( .A1(n8573), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n8560), .B2(
        n8565), .ZN(n8561) );
  NAND2_X1 U10006 ( .A1(n8562), .A2(n8561), .ZN(n8570) );
  OAI21_X1 U10007 ( .B1(n8562), .B2(n8561), .A(n8570), .ZN(n8567) );
  AOI21_X1 U10008 ( .B1(n10002), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8563), .ZN(
        n8564) );
  OAI21_X1 U10009 ( .B1(n9998), .B2(n8565), .A(n8564), .ZN(n8566) );
  AOI21_X1 U10010 ( .B1(n8567), .B2(n9995), .A(n8566), .ZN(n8568) );
  OAI21_X1 U10011 ( .B1(n8569), .B2(n8578), .A(n8568), .ZN(P2_U3263) );
  OAI21_X1 U10012 ( .B1(n8573), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8570), .ZN(
        n8571) );
  XOR2_X1 U10013 ( .A(n8571), .B(P2_REG1_REG_19__SCAN_IN), .Z(n8580) );
  NOR2_X1 U10014 ( .A1(n8573), .A2(n8572), .ZN(n8575) );
  NOR2_X1 U10015 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  XOR2_X1 U10016 ( .A(n8577), .B(n8576), .Z(n8579) );
  OAI22_X1 U10017 ( .A1(n8580), .A2(n10000), .B1(n8579), .B2(n8578), .ZN(n8584) );
  NAND2_X1 U10018 ( .A1(n8579), .A2(n9997), .ZN(n8582) );
  NAND2_X1 U10019 ( .A1(n8580), .A2(n9995), .ZN(n8581) );
  INV_X1 U10020 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8586) );
  OAI21_X1 U10021 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8588) );
  NAND2_X1 U10022 ( .A1(n8701), .A2(n8696), .ZN(n8690) );
  NAND2_X1 U10023 ( .A1(n8596), .A2(n8621), .ZN(n8595) );
  XNOR2_X1 U10024 ( .A(n8862), .B(n8595), .ZN(n8864) );
  NOR2_X1 U10025 ( .A1(n8831), .A2(n8589), .ZN(n8593) );
  INV_X1 U10026 ( .A(n8971), .ZN(n8590) );
  AND2_X1 U10027 ( .A1(n8590), .A2(P2_B_REG_SCAN_IN), .ZN(n8591) );
  NOR2_X1 U10028 ( .A1(n8838), .A2(n8591), .ZN(n8630) );
  NAND2_X1 U10029 ( .A1(n8592), .A2(n8630), .ZN(n8867) );
  NOR2_X1 U10030 ( .A1(n4314), .A2(n8867), .ZN(n8598) );
  AOI211_X1 U10031 ( .C1(n8862), .C2(n8854), .A(n8593), .B(n8598), .ZN(n8594)
         );
  OAI21_X1 U10032 ( .B1(n8864), .B2(n8601), .A(n8594), .ZN(P2_U3265) );
  OAI21_X1 U10033 ( .B1(n8596), .B2(n8621), .A(n8595), .ZN(n8868) );
  NOR2_X1 U10034 ( .A1(n8831), .A2(n8597), .ZN(n8599) );
  AOI211_X1 U10035 ( .C1(n8865), .C2(n8854), .A(n8599), .B(n8598), .ZN(n8600)
         );
  OAI21_X1 U10036 ( .B1(n8868), .B2(n8601), .A(n8600), .ZN(P2_U3266) );
  INV_X1 U10037 ( .A(n8902), .ZN(n8726) );
  NAND2_X1 U10038 ( .A1(n8938), .A2(n8606), .ZN(n8607) );
  OAI21_X1 U10039 ( .B1(n8805), .B2(n8934), .A(n8813), .ZN(n8795) );
  NOR2_X1 U10040 ( .A1(n8929), .A2(n8788), .ZN(n8608) );
  INV_X1 U10041 ( .A(n8643), .ZN(n8622) );
  AOI21_X1 U10042 ( .B1(n8869), .B2(n8622), .A(n8621), .ZN(n8870) );
  AOI22_X1 U10043 ( .A1(n4314), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n8797), .B2(
        n8623), .ZN(n8624) );
  OAI21_X1 U10044 ( .B1(n8625), .B2(n8800), .A(n8624), .ZN(n8635) );
  INV_X1 U10045 ( .A(n8626), .ZN(n8628) );
  INV_X1 U10046 ( .A(n8630), .ZN(n8631) );
  INV_X1 U10047 ( .A(n8633), .ZN(n8872) );
  OAI21_X1 U10048 ( .B1(n8874), .B2(n8812), .A(n8636), .ZN(P2_U3267) );
  XNOR2_X1 U10049 ( .A(n8637), .B(n8641), .ZN(n8639) );
  AOI21_X1 U10050 ( .B1(n8639), .B2(n8848), .A(n8638), .ZN(n8879) );
  OAI21_X1 U10051 ( .B1(n8642), .B2(n8641), .A(n8640), .ZN(n8875) );
  NAND2_X1 U10052 ( .A1(n8875), .A2(n8769), .ZN(n8650) );
  INV_X1 U10053 ( .A(n8655), .ZN(n8644) );
  AOI21_X1 U10054 ( .B1(n8876), .B2(n8644), .A(n8643), .ZN(n8877) );
  NOR2_X1 U10055 ( .A1(n8620), .A2(n8800), .ZN(n8648) );
  OAI22_X1 U10056 ( .A1(n8831), .A2(n8646), .B1(n8852), .B2(n8645), .ZN(n8647)
         );
  AOI211_X1 U10057 ( .C1(n8877), .C2(n8856), .A(n8648), .B(n8647), .ZN(n8649)
         );
  OAI211_X1 U10058 ( .C1(n4314), .C2(n8879), .A(n8650), .B(n8649), .ZN(
        P2_U3268) );
  OAI21_X1 U10059 ( .B1(n8653), .B2(n8652), .A(n8651), .ZN(n8654) );
  INV_X1 U10060 ( .A(n8654), .ZN(n8885) );
  AOI21_X1 U10061 ( .B1(n8881), .B2(n8669), .A(n8655), .ZN(n8882) );
  AOI22_X1 U10062 ( .A1(n4314), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8656), .B2(
        n8797), .ZN(n8657) );
  OAI21_X1 U10063 ( .B1(n8618), .B2(n8800), .A(n8657), .ZN(n8664) );
  XNOR2_X1 U10064 ( .A(n8659), .B(n8658), .ZN(n8662) );
  AOI222_X1 U10065 ( .A1(n8848), .A2(n8662), .B1(n8661), .B2(n8804), .C1(n8660), .C2(n8806), .ZN(n8884) );
  NOR2_X1 U10066 ( .A1(n8884), .A2(n4314), .ZN(n8663) );
  OAI21_X1 U10067 ( .B1(n8885), .B2(n8812), .A(n8665), .ZN(P2_U3269) );
  OAI21_X1 U10068 ( .B1(n8667), .B2(n8679), .A(n8666), .ZN(n8668) );
  INV_X1 U10069 ( .A(n8668), .ZN(n8890) );
  INV_X1 U10070 ( .A(n8669), .ZN(n8670) );
  AOI211_X1 U10071 ( .C1(n8888), .C2(n8690), .A(n10096), .B(n8670), .ZN(n8887)
         );
  NOR2_X1 U10072 ( .A1(n8671), .A2(n8800), .ZN(n8675) );
  OAI22_X1 U10073 ( .A1(n8831), .A2(n8673), .B1(n8672), .B2(n8852), .ZN(n8674)
         );
  AOI211_X1 U10074 ( .C1(n8887), .C2(n8793), .A(n8675), .B(n8674), .ZN(n8683)
         );
  INV_X1 U10075 ( .A(n8676), .ZN(n8677) );
  OAI222_X1 U10076 ( .A1(n8838), .A2(n8681), .B1(n8840), .B2(n8714), .C1(n8817), .C2(n8680), .ZN(n8886) );
  NAND2_X1 U10077 ( .A1(n8886), .A2(n8831), .ZN(n8682) );
  OAI211_X1 U10078 ( .C1(n8890), .C2(n8812), .A(n8683), .B(n8682), .ZN(
        P2_U3270) );
  OAI21_X1 U10079 ( .B1(n8685), .B2(n8686), .A(n8684), .ZN(n8891) );
  XNOR2_X1 U10080 ( .A(n8687), .B(n8686), .ZN(n8689) );
  AOI21_X1 U10081 ( .B1(n8689), .B2(n8848), .A(n8688), .ZN(n8895) );
  INV_X1 U10082 ( .A(n8701), .ZN(n8692) );
  INV_X1 U10083 ( .A(n8690), .ZN(n8691) );
  AOI211_X1 U10084 ( .C1(n8893), .C2(n8692), .A(n10096), .B(n8691), .ZN(n8892)
         );
  AOI22_X1 U10085 ( .A1(n8892), .A2(n8828), .B1(n8797), .B2(n8693), .ZN(n8694)
         );
  AOI21_X1 U10086 ( .B1(n8895), .B2(n8694), .A(n4314), .ZN(n8698) );
  OAI22_X1 U10087 ( .A1(n8696), .A2(n8800), .B1(n8831), .B2(n8695), .ZN(n8697)
         );
  AOI211_X1 U10088 ( .C1(n8891), .C2(n8769), .A(n8698), .B(n8697), .ZN(n8699)
         );
  INV_X1 U10089 ( .A(n8699), .ZN(P2_U3271) );
  XNOR2_X1 U10090 ( .A(n8700), .B(n8708), .ZN(n8901) );
  INV_X1 U10091 ( .A(n8723), .ZN(n8702) );
  AOI21_X1 U10092 ( .B1(n8897), .B2(n8702), .A(n8701), .ZN(n8898) );
  INV_X1 U10093 ( .A(n8703), .ZN(n8704) );
  AOI22_X1 U10094 ( .A1(n4314), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8704), .B2(
        n8797), .ZN(n8705) );
  OAI21_X1 U10095 ( .B1(n8706), .B2(n8800), .A(n8705), .ZN(n8718) );
  INV_X1 U10096 ( .A(n8707), .ZN(n8710) );
  OAI21_X1 U10097 ( .B1(n8710), .B2(n8709), .A(n8708), .ZN(n8712) );
  AND3_X1 U10098 ( .A1(n8711), .A2(n8848), .A3(n8712), .ZN(n8716) );
  OAI22_X1 U10099 ( .A1(n8714), .A2(n8838), .B1(n8713), .B2(n8840), .ZN(n8715)
         );
  NOR2_X1 U10100 ( .A1(n8716), .A2(n8715), .ZN(n8900) );
  NOR2_X1 U10101 ( .A1(n8900), .A2(n4314), .ZN(n8717) );
  AOI211_X1 U10102 ( .C1(n8898), .C2(n8856), .A(n8718), .B(n8717), .ZN(n8719)
         );
  OAI21_X1 U10103 ( .B1(n8901), .B2(n8812), .A(n8719), .ZN(P2_U3272) );
  OAI21_X1 U10104 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(n8906) );
  AOI21_X1 U10105 ( .B1(n8902), .B2(n8734), .A(n8723), .ZN(n8903) );
  AOI22_X1 U10106 ( .A1(n4314), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8724), .B2(
        n8797), .ZN(n8725) );
  OAI21_X1 U10107 ( .B1(n8726), .B2(n8800), .A(n8725), .ZN(n8732) );
  OAI21_X1 U10108 ( .B1(n8728), .B2(n8727), .A(n8707), .ZN(n8730) );
  AOI222_X1 U10109 ( .A1(n8848), .A2(n8730), .B1(n8758), .B2(n8804), .C1(n8729), .C2(n8806), .ZN(n8905) );
  NOR2_X1 U10110 ( .A1(n8905), .A2(n4314), .ZN(n8731) );
  AOI211_X1 U10111 ( .C1(n8903), .C2(n8856), .A(n8732), .B(n8731), .ZN(n8733)
         );
  OAI21_X1 U10112 ( .B1(n8906), .B2(n8812), .A(n8733), .ZN(P2_U3273) );
  XOR2_X1 U10113 ( .A(n8743), .B(n4349), .Z(n8911) );
  INV_X1 U10114 ( .A(n8734), .ZN(n8735) );
  AOI21_X1 U10115 ( .B1(n8907), .B2(n8750), .A(n8735), .ZN(n8908) );
  INV_X1 U10116 ( .A(n8736), .ZN(n8737) );
  AOI22_X1 U10117 ( .A1(n4314), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8737), .B2(
        n8797), .ZN(n8738) );
  OAI21_X1 U10118 ( .B1(n8739), .B2(n8800), .A(n8738), .ZN(n8747) );
  NAND2_X1 U10119 ( .A1(n8740), .A2(n8741), .ZN(n8742) );
  XOR2_X1 U10120 ( .A(n8743), .B(n8742), .Z(n8745) );
  AOI222_X1 U10121 ( .A1(n8848), .A2(n8745), .B1(n8765), .B2(n8804), .C1(n8744), .C2(n8806), .ZN(n8910) );
  NOR2_X1 U10122 ( .A1(n8910), .A2(n4314), .ZN(n8746) );
  AOI211_X1 U10123 ( .C1(n8908), .C2(n8856), .A(n8747), .B(n8746), .ZN(n8748)
         );
  OAI21_X1 U10124 ( .B1(n8911), .B2(n8812), .A(n8748), .ZN(P2_U3274) );
  XNOR2_X1 U10125 ( .A(n8749), .B(n8756), .ZN(n8916) );
  INV_X1 U10126 ( .A(n8772), .ZN(n8752) );
  INV_X1 U10127 ( .A(n8750), .ZN(n8751) );
  AOI21_X1 U10128 ( .B1(n8912), .B2(n8752), .A(n8751), .ZN(n8913) );
  AOI22_X1 U10129 ( .A1(n4314), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8753), .B2(
        n8797), .ZN(n8754) );
  OAI21_X1 U10130 ( .B1(n8755), .B2(n8800), .A(n8754), .ZN(n8761) );
  OAI21_X1 U10131 ( .B1(n8757), .B2(n5337), .A(n8740), .ZN(n8759) );
  AOI222_X1 U10132 ( .A1(n8848), .A2(n8759), .B1(n8758), .B2(n8806), .C1(n8789), .C2(n8804), .ZN(n8915) );
  NOR2_X1 U10133 ( .A1(n8915), .A2(n4314), .ZN(n8760) );
  AOI211_X1 U10134 ( .C1(n8913), .C2(n8856), .A(n8761), .B(n8760), .ZN(n8762)
         );
  OAI21_X1 U10135 ( .B1(n8916), .B2(n8812), .A(n8762), .ZN(P2_U3275) );
  NAND2_X1 U10136 ( .A1(n8785), .A2(n8763), .ZN(n8764) );
  XOR2_X1 U10137 ( .A(n8767), .B(n8764), .Z(n8766) );
  AOI222_X1 U10138 ( .A1(n8848), .A2(n8766), .B1(n8807), .B2(n8804), .C1(n8765), .C2(n8806), .ZN(n8922) );
  OR2_X1 U10139 ( .A1(n8768), .A2(n8767), .ZN(n8918) );
  NAND3_X1 U10140 ( .A1(n8918), .A2(n8917), .A3(n8769), .ZN(n8778) );
  NOR2_X1 U10141 ( .A1(n8780), .A2(n8770), .ZN(n8771) );
  NOR2_X1 U10142 ( .A1(n8772), .A2(n8771), .ZN(n8920) );
  NAND2_X1 U10143 ( .A1(n8919), .A2(n8854), .ZN(n8775) );
  AOI22_X1 U10144 ( .A1(n4314), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8773), .B2(
        n8797), .ZN(n8774) );
  NAND2_X1 U10145 ( .A1(n8775), .A2(n8774), .ZN(n8776) );
  AOI21_X1 U10146 ( .B1(n8920), .B2(n8856), .A(n8776), .ZN(n8777) );
  OAI211_X1 U10147 ( .C1(n4314), .C2(n8922), .A(n8778), .B(n8777), .ZN(
        P2_U3276) );
  XOR2_X1 U10148 ( .A(n8779), .B(n8787), .Z(n8928) );
  INV_X1 U10149 ( .A(n8796), .ZN(n8781) );
  AOI211_X1 U10150 ( .C1(n8925), .C2(n8781), .A(n10096), .B(n8780), .ZN(n8924)
         );
  AOI22_X1 U10151 ( .A1(n4314), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8782), .B2(
        n8797), .ZN(n8783) );
  OAI21_X1 U10152 ( .B1(n8784), .B2(n8800), .A(n8783), .ZN(n8792) );
  OAI21_X1 U10153 ( .B1(n8787), .B2(n8786), .A(n8785), .ZN(n8790) );
  AOI222_X1 U10154 ( .A1(n8848), .A2(n8790), .B1(n8789), .B2(n8806), .C1(n8788), .C2(n8804), .ZN(n8927) );
  NOR2_X1 U10155 ( .A1(n8927), .A2(n4314), .ZN(n8791) );
  AOI211_X1 U10156 ( .C1(n8924), .C2(n8793), .A(n8792), .B(n8791), .ZN(n8794)
         );
  OAI21_X1 U10157 ( .B1(n8812), .B2(n8928), .A(n8794), .ZN(P2_U3277) );
  XNOR2_X1 U10158 ( .A(n8795), .B(n4317), .ZN(n8933) );
  AOI21_X1 U10159 ( .B1(n8929), .B2(n8823), .A(n8796), .ZN(n8930) );
  AOI22_X1 U10160 ( .A1(n4314), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8798), .B2(
        n8797), .ZN(n8799) );
  OAI21_X1 U10161 ( .B1(n8801), .B2(n8800), .A(n8799), .ZN(n8810) );
  OAI21_X1 U10162 ( .B1(n8803), .B2(n4317), .A(n8802), .ZN(n8808) );
  AOI222_X1 U10163 ( .A1(n8848), .A2(n8808), .B1(n8807), .B2(n8806), .C1(n8805), .C2(n8804), .ZN(n8932) );
  NOR2_X1 U10164 ( .A1(n8932), .A2(n4314), .ZN(n8809) );
  AOI211_X1 U10165 ( .C1(n8930), .C2(n8856), .A(n8810), .B(n8809), .ZN(n8811)
         );
  OAI21_X1 U10166 ( .B1(n8812), .B2(n8933), .A(n8811), .ZN(P2_U3278) );
  OAI21_X1 U10167 ( .B1(n8814), .B2(n8815), .A(n8813), .ZN(n8935) );
  INV_X1 U10168 ( .A(n8935), .ZN(n8835) );
  XNOR2_X1 U10169 ( .A(n8816), .B(n8815), .ZN(n8818) );
  OAI222_X1 U10170 ( .A1(n8840), .A2(n8820), .B1(n8838), .B2(n8819), .C1(n8818), .C2(n8817), .ZN(n8827) );
  INV_X1 U10171 ( .A(n8821), .ZN(n8825) );
  AOI21_X1 U10172 ( .B1(n8822), .B2(n8934), .A(n10096), .ZN(n8824) );
  AOI21_X1 U10173 ( .B1(n8824), .B2(n8823), .A(n8827), .ZN(n8936) );
  OAI21_X1 U10174 ( .B1(n8835), .B2(n8825), .A(n8936), .ZN(n8826) );
  OAI211_X1 U10175 ( .C1(n8828), .C2(n8827), .A(n8826), .B(n8831), .ZN(n8834)
         );
  OAI22_X1 U10176 ( .A1(n8831), .A2(n8830), .B1(n8829), .B2(n8852), .ZN(n8832)
         );
  AOI21_X1 U10177 ( .B1(n8934), .B2(n8854), .A(n8832), .ZN(n8833) );
  OAI211_X1 U10178 ( .C1(n8835), .C2(n8859), .A(n8834), .B(n8833), .ZN(
        P2_U3279) );
  XNOR2_X1 U10179 ( .A(n8836), .B(n8837), .ZN(n8849) );
  OAI22_X1 U10180 ( .A1(n8841), .A2(n8840), .B1(n8839), .B2(n8838), .ZN(n8847)
         );
  NOR2_X1 U10181 ( .A1(n8843), .A2(n8842), .ZN(n8844) );
  NOR2_X1 U10182 ( .A1(n8942), .A2(n8845), .ZN(n8846) );
  AOI211_X1 U10183 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8941)
         );
  NAND2_X1 U10184 ( .A1(n4314), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8850) );
  OAI21_X1 U10185 ( .B1(n8852), .B2(n8851), .A(n8850), .ZN(n8853) );
  AOI21_X1 U10186 ( .B1(n8854), .B2(n8938), .A(n8853), .ZN(n8858) );
  XNOR2_X1 U10187 ( .A(n8855), .B(n4582), .ZN(n8939) );
  NAND2_X1 U10188 ( .A1(n8939), .A2(n8856), .ZN(n8857) );
  OAI211_X1 U10189 ( .C1(n8942), .C2(n8859), .A(n8858), .B(n8857), .ZN(n8860)
         );
  INV_X1 U10190 ( .A(n8860), .ZN(n8861) );
  OAI21_X1 U10191 ( .B1(n8941), .B2(n4314), .A(n8861), .ZN(P2_U3280) );
  NAND2_X1 U10192 ( .A1(n8862), .A2(n10088), .ZN(n8863) );
  OAI211_X1 U10193 ( .C1(n8864), .C2(n10096), .A(n8867), .B(n8863), .ZN(n8943)
         );
  MUX2_X1 U10194 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8943), .S(n10120), .Z(
        P2_U3551) );
  NAND2_X1 U10195 ( .A1(n8865), .A2(n10088), .ZN(n8866) );
  OAI211_X1 U10196 ( .C1(n8868), .C2(n10096), .A(n8867), .B(n8866), .ZN(n8944)
         );
  MUX2_X1 U10197 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8944), .S(n10120), .Z(
        P2_U3550) );
  AOI22_X1 U10198 ( .A1(n8870), .A2(n10089), .B1(n10088), .B2(n8869), .ZN(
        n8871) );
  MUX2_X1 U10199 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8945), .S(n10120), .Z(
        P2_U3549) );
  INV_X1 U10200 ( .A(n8875), .ZN(n8880) );
  AOI22_X1 U10201 ( .A1(n8877), .A2(n10089), .B1(n10088), .B2(n8876), .ZN(
        n8878) );
  OAI211_X1 U10202 ( .C1(n8880), .C2(n10085), .A(n8879), .B(n8878), .ZN(n8946)
         );
  MUX2_X1 U10203 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8946), .S(n10120), .Z(
        P2_U3548) );
  AOI22_X1 U10204 ( .A1(n8882), .A2(n10089), .B1(n10088), .B2(n8881), .ZN(
        n8883) );
  OAI211_X1 U10205 ( .C1(n8885), .C2(n10085), .A(n8884), .B(n8883), .ZN(n8947)
         );
  MUX2_X1 U10206 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8947), .S(n10120), .Z(
        P2_U3547) );
  OAI21_X1 U10207 ( .B1(n8890), .B2(n10085), .A(n8889), .ZN(n8948) );
  MUX2_X1 U10208 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8948), .S(n10120), .Z(
        P2_U3546) );
  INV_X1 U10209 ( .A(n8891), .ZN(n8896) );
  AOI21_X1 U10210 ( .B1(n10088), .B2(n8893), .A(n8892), .ZN(n8894) );
  OAI211_X1 U10211 ( .C1(n8896), .C2(n10085), .A(n8895), .B(n8894), .ZN(n8949)
         );
  MUX2_X1 U10212 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8949), .S(n10120), .Z(
        P2_U3545) );
  AOI22_X1 U10213 ( .A1(n8898), .A2(n10089), .B1(n10088), .B2(n8897), .ZN(
        n8899) );
  OAI211_X1 U10214 ( .C1(n8901), .C2(n10085), .A(n8900), .B(n8899), .ZN(n8950)
         );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8950), .S(n10120), .Z(
        P2_U3544) );
  AOI22_X1 U10216 ( .A1(n8903), .A2(n10089), .B1(n10088), .B2(n8902), .ZN(
        n8904) );
  OAI211_X1 U10217 ( .C1(n8906), .C2(n10085), .A(n8905), .B(n8904), .ZN(n8951)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8951), .S(n10120), .Z(
        P2_U3543) );
  AOI22_X1 U10219 ( .A1(n8908), .A2(n10089), .B1(n10088), .B2(n8907), .ZN(
        n8909) );
  OAI211_X1 U10220 ( .C1(n8911), .C2(n10085), .A(n8910), .B(n8909), .ZN(n8952)
         );
  MUX2_X1 U10221 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8952), .S(n10120), .Z(
        P2_U3542) );
  AOI22_X1 U10222 ( .A1(n8913), .A2(n10089), .B1(n10088), .B2(n8912), .ZN(
        n8914) );
  OAI211_X1 U10223 ( .C1(n8916), .C2(n10085), .A(n8915), .B(n8914), .ZN(n8953)
         );
  MUX2_X1 U10224 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8953), .S(n10120), .Z(
        P2_U3541) );
  NAND3_X1 U10225 ( .A1(n8918), .A2(n8917), .A3(n10101), .ZN(n8923) );
  AOI22_X1 U10226 ( .A1(n8920), .A2(n10089), .B1(n10088), .B2(n8919), .ZN(
        n8921) );
  NAND3_X1 U10227 ( .A1(n8923), .A2(n8922), .A3(n8921), .ZN(n8954) );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8954), .S(n10120), .Z(
        P2_U3540) );
  AOI21_X1 U10229 ( .B1(n10088), .B2(n8925), .A(n8924), .ZN(n8926) );
  OAI211_X1 U10230 ( .C1(n8928), .C2(n10085), .A(n8927), .B(n8926), .ZN(n8955)
         );
  MUX2_X1 U10231 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8955), .S(n10120), .Z(
        P2_U3539) );
  AOI22_X1 U10232 ( .A1(n8930), .A2(n10089), .B1(n10088), .B2(n8929), .ZN(
        n8931) );
  OAI211_X1 U10233 ( .C1(n8933), .C2(n10085), .A(n8932), .B(n8931), .ZN(n8956)
         );
  MUX2_X1 U10234 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8956), .S(n10120), .Z(
        P2_U3538) );
  AOI22_X1 U10235 ( .A1(n8935), .A2(n10101), .B1(n10088), .B2(n8934), .ZN(
        n8937) );
  NAND2_X1 U10236 ( .A1(n8937), .A2(n8936), .ZN(n8957) );
  MUX2_X1 U10237 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8957), .S(n10120), .Z(
        P2_U3537) );
  AOI22_X1 U10238 ( .A1(n8939), .A2(n10089), .B1(n10088), .B2(n8938), .ZN(
        n8940) );
  OAI211_X1 U10239 ( .C1(n9806), .C2(n8942), .A(n8941), .B(n8940), .ZN(n8958)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8958), .S(n10120), .Z(
        P2_U3536) );
  MUX2_X1 U10241 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8943), .S(n10104), .Z(
        P2_U3519) );
  MUX2_X1 U10242 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8944), .S(n10104), .Z(
        P2_U3518) );
  MUX2_X1 U10243 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8945), .S(n10104), .Z(
        P2_U3517) );
  MUX2_X1 U10244 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8946), .S(n10104), .Z(
        P2_U3516) );
  MUX2_X1 U10245 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8947), .S(n10104), .Z(
        P2_U3515) );
  MUX2_X1 U10246 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8948), .S(n10104), .Z(
        P2_U3514) );
  MUX2_X1 U10247 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8949), .S(n10104), .Z(
        P2_U3513) );
  MUX2_X1 U10248 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8950), .S(n10104), .Z(
        P2_U3512) );
  MUX2_X1 U10249 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8951), .S(n10104), .Z(
        P2_U3511) );
  MUX2_X1 U10250 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8952), .S(n10104), .Z(
        P2_U3510) );
  MUX2_X1 U10251 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8953), .S(n10104), .Z(
        P2_U3509) );
  MUX2_X1 U10252 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8954), .S(n10104), .Z(
        P2_U3508) );
  MUX2_X1 U10253 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8955), .S(n10104), .Z(
        P2_U3507) );
  MUX2_X1 U10254 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8956), .S(n10104), .Z(
        P2_U3505) );
  MUX2_X1 U10255 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8957), .S(n10104), .Z(
        P2_U3502) );
  MUX2_X1 U10256 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8958), .S(n10104), .Z(
        P2_U3499) );
  INV_X1 U10257 ( .A(n8959), .ZN(n9534) );
  NOR4_X1 U10258 ( .A1(n8960), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4919), .A4(
        P2_U3152), .ZN(n8961) );
  AOI21_X1 U10259 ( .B1(n8968), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8961), .ZN(
        n8962) );
  OAI21_X1 U10260 ( .B1(n9534), .B2(n8970), .A(n8962), .ZN(P2_U3327) );
  OAI222_X1 U10261 ( .A1(n4923), .A2(P2_U3152), .B1(n8973), .B2(n8965), .C1(
        n8964), .C2(n8963), .ZN(P2_U3329) );
  INV_X1 U10262 ( .A(n8966), .ZN(n9538) );
  AOI21_X1 U10263 ( .B1(n8968), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8967), .ZN(
        n8969) );
  OAI21_X1 U10264 ( .B1(n9538), .B2(n8970), .A(n8969), .ZN(P2_U3330) );
  OAI222_X1 U10265 ( .A1(n8963), .A2(n8974), .B1(n8973), .B2(n8972), .C1(n8971), .C2(P2_U3152), .ZN(P2_U3331) );
  MUX2_X1 U10266 ( .A(n8975), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10267 ( .A(n9031), .ZN(n8979) );
  AOI21_X1 U10268 ( .B1(n8977), .B2(n9030), .A(n8976), .ZN(n8978) );
  AOI21_X1 U10269 ( .B1(n8979), .B2(n9030), .A(n8978), .ZN(n8984) );
  OAI22_X1 U10270 ( .A1(n9293), .A2(n9094), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8980), .ZN(n8982) );
  OAI22_X1 U10271 ( .A1(n9294), .A2(n9070), .B1(n9096), .B2(n9296), .ZN(n8981)
         );
  AOI211_X1 U10272 ( .C1(n9453), .C2(n6480), .A(n8982), .B(n8981), .ZN(n8983)
         );
  OAI21_X1 U10273 ( .B1(n8984), .B2(n9103), .A(n8983), .ZN(P1_U3214) );
  XOR2_X1 U10274 ( .A(n8986), .B(n8985), .Z(n8990) );
  NAND2_X1 U10275 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9186) );
  OAI21_X1 U10276 ( .B1(n9365), .B2(n9070), .A(n9186), .ZN(n8988) );
  OAI22_X1 U10277 ( .A1(n9096), .A2(n9358), .B1(n9094), .B2(n9404), .ZN(n8987)
         );
  AOI211_X1 U10278 ( .C1(n9473), .C2(n6480), .A(n8988), .B(n8987), .ZN(n8989)
         );
  OAI21_X1 U10279 ( .B1(n8990), .B2(n9103), .A(n8989), .ZN(P1_U3217) );
  XOR2_X1 U10280 ( .A(n8992), .B(n8993), .Z(n8999) );
  OAI22_X1 U10281 ( .A1(n9293), .A2(n9070), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8994), .ZN(n8997) );
  INV_X1 U10282 ( .A(n9329), .ZN(n8995) );
  OAI22_X1 U10283 ( .A1(n9096), .A2(n8995), .B1(n9365), .B2(n9094), .ZN(n8996)
         );
  AOI211_X1 U10284 ( .C1(n9328), .C2(n6480), .A(n8997), .B(n8996), .ZN(n8998)
         );
  OAI21_X1 U10285 ( .B1(n8999), .B2(n9103), .A(n8998), .ZN(P1_U3221) );
  AOI21_X1 U10286 ( .B1(n9001), .B2(n9000), .A(n9078), .ZN(n9007) );
  NAND2_X1 U10287 ( .A1(n9261), .A2(n9099), .ZN(n9004) );
  INV_X1 U10288 ( .A(n9002), .ZN(n9268) );
  AOI22_X1 U10289 ( .A1(n9268), .A2(n9082), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9003) );
  OAI211_X1 U10290 ( .C1(n9294), .C2(n9094), .A(n9004), .B(n9003), .ZN(n9005)
         );
  AOI21_X1 U10291 ( .B1(n9267), .B2(n6480), .A(n9005), .ZN(n9006) );
  OAI21_X1 U10292 ( .B1(n9007), .B2(n9103), .A(n9006), .ZN(P1_U3223) );
  INV_X1 U10293 ( .A(n9009), .ZN(n9010) );
  AOI21_X1 U10294 ( .B1(n9011), .B2(n9008), .A(n9010), .ZN(n9019) );
  OAI22_X1 U10295 ( .A1(n9094), .A2(n9013), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9012), .ZN(n9016) );
  OAI22_X1 U10296 ( .A1(n9096), .A2(n9014), .B1(n9070), .B2(n9372), .ZN(n9015)
         );
  AOI211_X1 U10297 ( .C1(n9017), .C2(n6480), .A(n9016), .B(n9015), .ZN(n9018)
         );
  OAI21_X1 U10298 ( .B1(n9019), .B2(n9103), .A(n9018), .ZN(P1_U3224) );
  OAI21_X1 U10299 ( .B1(n9022), .B2(n9021), .A(n9020), .ZN(n9023) );
  NAND2_X1 U10300 ( .A1(n9023), .A2(n9080), .ZN(n9028) );
  OAI22_X1 U10301 ( .A1(n9070), .A2(n9404), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9024), .ZN(n9026) );
  OAI22_X1 U10302 ( .A1(n9096), .A2(n9394), .B1(n9094), .B2(n9402), .ZN(n9025)
         );
  AOI211_X1 U10303 ( .C1(n9483), .C2(n6480), .A(n9026), .B(n9025), .ZN(n9027)
         );
  NAND2_X1 U10304 ( .A1(n9028), .A2(n9027), .ZN(P1_U3226) );
  AND3_X1 U10305 ( .A1(n9031), .A2(n9030), .A3(n9029), .ZN(n9032) );
  OAI21_X1 U10306 ( .B1(n9033), .B2(n9032), .A(n9080), .ZN(n9038) );
  OAI22_X1 U10307 ( .A1(n9307), .A2(n9094), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9034), .ZN(n9036) );
  NOR2_X1 U10308 ( .A1(n9280), .A2(n9070), .ZN(n9035) );
  AOI211_X1 U10309 ( .C1(n9283), .C2(n9082), .A(n9036), .B(n9035), .ZN(n9037)
         );
  OAI211_X1 U10310 ( .C1(n9512), .C2(n9087), .A(n9038), .B(n9037), .ZN(
        P1_U3227) );
  NAND2_X1 U10311 ( .A1(n9040), .A2(n9039), .ZN(n9041) );
  XNOR2_X1 U10312 ( .A(n9042), .B(n9041), .ZN(n9047) );
  OAI22_X1 U10313 ( .A1(n9306), .A2(n9070), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9043), .ZN(n9045) );
  OAI22_X1 U10314 ( .A1(n9096), .A2(n9338), .B1(n9094), .B2(n9373), .ZN(n9044)
         );
  AOI211_X1 U10315 ( .C1(n9467), .C2(n6480), .A(n9045), .B(n9044), .ZN(n9046)
         );
  OAI21_X1 U10316 ( .B1(n9047), .B2(n9103), .A(n9046), .ZN(P1_U3231) );
  NAND2_X1 U10317 ( .A1(n9049), .A2(n9048), .ZN(n9051) );
  XNOR2_X1 U10318 ( .A(n9051), .B(n9050), .ZN(n9056) );
  OAI22_X1 U10319 ( .A1(n9307), .A2(n9070), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9052), .ZN(n9054) );
  OAI22_X1 U10320 ( .A1(n9306), .A2(n9094), .B1(n9096), .B2(n9310), .ZN(n9053)
         );
  AOI211_X1 U10321 ( .C1(n9458), .C2(n6480), .A(n9054), .B(n9053), .ZN(n9055)
         );
  OAI21_X1 U10322 ( .B1(n9056), .B2(n9103), .A(n9055), .ZN(P1_U3233) );
  OAI21_X1 U10323 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9060) );
  NAND2_X1 U10324 ( .A1(n9060), .A2(n9080), .ZN(n9065) );
  AOI22_X1 U10325 ( .A1(n6480), .A2(n4839), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        n9061), .ZN(n9064) );
  AOI22_X1 U10326 ( .A1(n9062), .A2(n5771), .B1(n9099), .B2(n9126), .ZN(n9063)
         );
  NAND3_X1 U10327 ( .A1(n9065), .A2(n9064), .A3(n9063), .ZN(P1_U3235) );
  NAND2_X1 U10328 ( .A1(n9067), .A2(n9066), .ZN(n9068) );
  XOR2_X1 U10329 ( .A(n9069), .B(n9068), .Z(n9074) );
  NAND2_X1 U10330 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9948) );
  OAI21_X1 U10331 ( .B1(n9070), .B2(n9373), .A(n9948), .ZN(n9072) );
  OAI22_X1 U10332 ( .A1(n9096), .A2(n9379), .B1(n9094), .B2(n9372), .ZN(n9071)
         );
  AOI211_X1 U10333 ( .C1(n9378), .C2(n6480), .A(n9072), .B(n9071), .ZN(n9073)
         );
  OAI21_X1 U10334 ( .B1(n9074), .B2(n9103), .A(n9073), .ZN(P1_U3236) );
  INV_X1 U10335 ( .A(n9075), .ZN(n9081) );
  OAI21_X1 U10336 ( .B1(n9078), .B2(n9077), .A(n9076), .ZN(n9079) );
  NAND3_X1 U10337 ( .A1(n9081), .A2(n9080), .A3(n9079), .ZN(n9086) );
  AOI22_X1 U10338 ( .A1(n9249), .A2(n9082), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9083) );
  OAI21_X1 U10339 ( .B1(n9280), .B2(n9094), .A(n9083), .ZN(n9084) );
  AOI21_X1 U10340 ( .B1(n9108), .B2(n9099), .A(n9084), .ZN(n9085) );
  OAI211_X1 U10341 ( .C1(n9504), .C2(n9087), .A(n9086), .B(n9085), .ZN(
        P1_U3238) );
  NAND2_X1 U10342 ( .A1(n9088), .A2(n9089), .ZN(n9090) );
  XOR2_X1 U10343 ( .A(n9091), .B(n9090), .Z(n9104) );
  INV_X1 U10344 ( .A(n9092), .ZN(n9098) );
  OAI22_X1 U10345 ( .A1(n9096), .A2(n9095), .B1(n9094), .B2(n9093), .ZN(n9097)
         );
  AOI211_X1 U10346 ( .C1(n9099), .C2(n9113), .A(n9098), .B(n9097), .ZN(n9102)
         );
  NAND2_X1 U10347 ( .A1(n9100), .A2(n6480), .ZN(n9101) );
  OAI211_X1 U10348 ( .C1(n9104), .C2(n9103), .A(n9102), .B(n9101), .ZN(
        P1_U3239) );
  MUX2_X1 U10349 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9105), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10350 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9106), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10351 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9107), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10352 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9108), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10353 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9261), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10354 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9109), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10355 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9260), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10356 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9110), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10357 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9322), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10358 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9349), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10359 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9321), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10360 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9347), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10361 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9111), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10362 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9112), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10363 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9113), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10364 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9114), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10365 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9115), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10366 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9116), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10367 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9117), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10368 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9118), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10369 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9119), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10370 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9120), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10371 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9121), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10372 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9122), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10373 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9123), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10374 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9124), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10375 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9125), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10376 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9126), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9127), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5771), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6376), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10380 ( .A1(n9866), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9140) );
  AOI21_X1 U10381 ( .B1(n9951), .B2(n9129), .A(n9128), .ZN(n9139) );
  OAI211_X1 U10382 ( .C1(n9132), .C2(n9131), .A(n9960), .B(n9130), .ZN(n9138)
         );
  OAI21_X1 U10383 ( .B1(n9135), .B2(n9134), .A(n9133), .ZN(n9136) );
  NAND2_X1 U10384 ( .A1(n9959), .A2(n9136), .ZN(n9137) );
  NAND4_X1 U10385 ( .A1(n9140), .A2(n9139), .A3(n9138), .A4(n9137), .ZN(
        P1_U3247) );
  OAI21_X1 U10386 ( .B1(n9143), .B2(n9142), .A(n9141), .ZN(n9144) );
  NAND2_X1 U10387 ( .A1(n9144), .A2(n9959), .ZN(n9154) );
  NOR2_X1 U10388 ( .A1(n9943), .A2(n9145), .ZN(n9146) );
  AOI211_X1 U10389 ( .C1(n9866), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9147), .B(
        n9146), .ZN(n9153) );
  OAI21_X1 U10390 ( .B1(n9150), .B2(n9149), .A(n9148), .ZN(n9151) );
  NAND2_X1 U10391 ( .A1(n9151), .A2(n9960), .ZN(n9152) );
  NAND3_X1 U10392 ( .A1(n9154), .A2(n9153), .A3(n9152), .ZN(P1_U3252) );
  INV_X1 U10393 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9169) );
  MUX2_X1 U10394 ( .A(n9156), .B(P1_REG2_REG_17__SCAN_IN), .S(n9175), .Z(n9157) );
  AOI211_X1 U10395 ( .C1(n9158), .C2(n9157), .A(n9170), .B(n9935), .ZN(n9167)
         );
  AOI21_X1 U10396 ( .B1(n9160), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9159), .ZN(
        n9162) );
  XNOR2_X1 U10397 ( .A(n9175), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9161) );
  NOR2_X1 U10398 ( .A1(n9162), .A2(n9161), .ZN(n9174) );
  AOI211_X1 U10399 ( .C1(n9162), .C2(n9161), .A(n9174), .B(n9882), .ZN(n9166)
         );
  INV_X1 U10400 ( .A(n9175), .ZN(n9164) );
  NAND2_X1 U10401 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9163) );
  OAI21_X1 U10402 ( .B1(n9943), .B2(n9164), .A(n9163), .ZN(n9165) );
  NOR3_X1 U10403 ( .A1(n9167), .A2(n9166), .A3(n9165), .ZN(n9168) );
  OAI21_X1 U10404 ( .B1(n9964), .B2(n9169), .A(n9168), .ZN(P1_U3258) );
  INV_X1 U10405 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9187) );
  AOI21_X1 U10406 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n9175), .A(n9170), .ZN(
        n9954) );
  NAND2_X1 U10407 ( .A1(n9950), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9171) );
  OAI21_X1 U10408 ( .B1(n9950), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9171), .ZN(
        n9953) );
  NOR2_X1 U10409 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  AOI21_X1 U10410 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9950), .A(n9952), .ZN(
        n9172) );
  XNOR2_X1 U10411 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9172), .ZN(n9182) );
  AOI22_X1 U10412 ( .A1(n9950), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9479), .B2(
        n9173), .ZN(n9957) );
  AOI21_X1 U10413 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9175), .A(n9174), .ZN(
        n9956) );
  NAND2_X1 U10414 ( .A1(n9957), .A2(n9956), .ZN(n9955) );
  OAI21_X1 U10415 ( .B1(n9950), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9955), .ZN(
        n9177) );
  XOR2_X1 U10416 ( .A(n9177), .B(n9176), .Z(n9178) );
  AOI22_X1 U10417 ( .A1(n9182), .A2(n9960), .B1(n9959), .B2(n9178), .ZN(n9185)
         );
  INV_X1 U10418 ( .A(n9178), .ZN(n9183) );
  INV_X1 U10419 ( .A(n9179), .ZN(n9181) );
  XNOR2_X1 U10420 ( .A(n9189), .B(n4320), .ZN(n9190) );
  NAND2_X1 U10421 ( .A1(n9422), .A2(n9818), .ZN(n9194) );
  AND2_X1 U10422 ( .A1(n9192), .A2(n9191), .ZN(n9421) );
  INV_X1 U10423 ( .A(n9421), .ZN(n9425) );
  NOR2_X1 U10424 ( .A1(n9425), .A2(n9826), .ZN(n9197) );
  AOI21_X1 U10425 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(n9826), .A(n9197), .ZN(
        n9193) );
  OAI211_X1 U10426 ( .C1(n9494), .C2(n9392), .A(n9194), .B(n9193), .ZN(
        P1_U3261) );
  OAI211_X1 U10427 ( .C1(n9497), .C2(n9195), .A(n9228), .B(n4320), .ZN(n9426)
         );
  NOR2_X1 U10428 ( .A1(n9497), .A2(n9392), .ZN(n9196) );
  AOI211_X1 U10429 ( .C1(n9826), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9197), .B(
        n9196), .ZN(n9198) );
  OAI21_X1 U10430 ( .B1(n9199), .B2(n9426), .A(n9198), .ZN(P1_U3262) );
  INV_X1 U10431 ( .A(n9200), .ZN(n9210) );
  NAND2_X1 U10432 ( .A1(n9201), .A2(n9397), .ZN(n9205) );
  INV_X1 U10433 ( .A(n9202), .ZN(n9203) );
  AOI22_X1 U10434 ( .A1(n9203), .A2(n9339), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9826), .ZN(n9204) );
  OAI211_X1 U10435 ( .C1(n9206), .C2(n9392), .A(n9205), .B(n9204), .ZN(n9207)
         );
  AOI21_X1 U10436 ( .B1(n9208), .B2(n9409), .A(n9207), .ZN(n9209) );
  OAI21_X1 U10437 ( .B1(n9210), .B2(n9408), .A(n9209), .ZN(P1_U3355) );
  INV_X1 U10438 ( .A(n9211), .ZN(n9219) );
  NAND2_X1 U10439 ( .A1(n9212), .A2(n9397), .ZN(n9215) );
  AOI22_X1 U10440 ( .A1(n9213), .A2(n9339), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9826), .ZN(n9214) );
  OAI211_X1 U10441 ( .C1(n4667), .C2(n9392), .A(n9215), .B(n9214), .ZN(n9216)
         );
  AOI21_X1 U10442 ( .B1(n9217), .B2(n9409), .A(n9216), .ZN(n9218) );
  OAI21_X1 U10443 ( .B1(n9219), .B2(n9408), .A(n9218), .ZN(P1_U3263) );
  XNOR2_X1 U10444 ( .A(n9220), .B(n9225), .ZN(n9224) );
  OAI22_X1 U10445 ( .A1(n9222), .A2(n9405), .B1(n9221), .B2(n9403), .ZN(n9223)
         );
  AOI21_X1 U10446 ( .B1(n9224), .B2(n9351), .A(n9223), .ZN(n9431) );
  XNOR2_X1 U10447 ( .A(n9226), .B(n9225), .ZN(n9433) );
  NAND2_X1 U10448 ( .A1(n9433), .A2(n9414), .ZN(n9235) );
  INV_X1 U10449 ( .A(n9227), .ZN(n9247) );
  OAI211_X1 U10450 ( .C1(n4666), .C2(n9247), .A(n9229), .B(n9228), .ZN(n9430)
         );
  INV_X1 U10451 ( .A(n9430), .ZN(n9233) );
  AOI22_X1 U10452 ( .A1(n9230), .A2(n9339), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9826), .ZN(n9231) );
  OAI21_X1 U10453 ( .B1(n4666), .B2(n9392), .A(n9231), .ZN(n9232) );
  AOI21_X1 U10454 ( .B1(n9233), .B2(n9397), .A(n9232), .ZN(n9234) );
  OAI211_X1 U10455 ( .C1(n9431), .C2(n9826), .A(n9235), .B(n9234), .ZN(
        P1_U3264) );
  XOR2_X1 U10456 ( .A(n9239), .B(n9236), .Z(n9438) );
  INV_X1 U10457 ( .A(n9438), .ZN(n9254) );
  NAND2_X1 U10458 ( .A1(n9238), .A2(n9237), .ZN(n9241) );
  INV_X1 U10459 ( .A(n9239), .ZN(n9240) );
  XNOR2_X1 U10460 ( .A(n9241), .B(n9240), .ZN(n9242) );
  NAND2_X1 U10461 ( .A1(n9242), .A2(n9351), .ZN(n9246) );
  OAI22_X1 U10462 ( .A1(n9243), .A2(n9405), .B1(n9280), .B2(n9403), .ZN(n9244)
         );
  INV_X1 U10463 ( .A(n9244), .ZN(n9245) );
  NAND2_X1 U10464 ( .A1(n9246), .A2(n9245), .ZN(n9436) );
  AOI211_X1 U10465 ( .C1(n9248), .C2(n9264), .A(n9390), .B(n9247), .ZN(n9437)
         );
  NAND2_X1 U10466 ( .A1(n9437), .A2(n9397), .ZN(n9251) );
  AOI22_X1 U10467 ( .A1(n9249), .A2(n9339), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9826), .ZN(n9250) );
  OAI211_X1 U10468 ( .C1(n9504), .C2(n9392), .A(n9251), .B(n9250), .ZN(n9252)
         );
  AOI21_X1 U10469 ( .B1(n9436), .B2(n9409), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10470 ( .B1(n9254), .B2(n9408), .A(n9253), .ZN(P1_U3265) );
  XNOR2_X1 U10471 ( .A(n9255), .B(n9257), .ZN(n9443) );
  INV_X1 U10472 ( .A(n9443), .ZN(n9273) );
  NAND2_X1 U10473 ( .A1(n9275), .A2(n9256), .ZN(n9258) );
  XNOR2_X1 U10474 ( .A(n9258), .B(n4605), .ZN(n9259) );
  NAND2_X1 U10475 ( .A1(n9259), .A2(n9351), .ZN(n9263) );
  AOI22_X1 U10476 ( .A1(n9261), .A2(n9348), .B1(n9346), .B2(n9260), .ZN(n9262)
         );
  NAND2_X1 U10477 ( .A1(n9263), .A2(n9262), .ZN(n9441) );
  INV_X1 U10478 ( .A(n9281), .ZN(n9266) );
  INV_X1 U10479 ( .A(n9264), .ZN(n9265) );
  AOI211_X1 U10480 ( .C1(n9267), .C2(n9266), .A(n9390), .B(n9265), .ZN(n9442)
         );
  NAND2_X1 U10481 ( .A1(n9442), .A2(n9397), .ZN(n9270) );
  AOI22_X1 U10482 ( .A1(n9268), .A2(n9339), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9826), .ZN(n9269) );
  OAI211_X1 U10483 ( .C1(n9508), .C2(n9392), .A(n9270), .B(n9269), .ZN(n9271)
         );
  AOI21_X1 U10484 ( .B1(n9441), .B2(n9409), .A(n9271), .ZN(n9272) );
  OAI21_X1 U10485 ( .B1(n9273), .B2(n9408), .A(n9272), .ZN(P1_U3266) );
  XOR2_X1 U10486 ( .A(n9277), .B(n9274), .Z(n9448) );
  INV_X1 U10487 ( .A(n9448), .ZN(n9288) );
  INV_X1 U10488 ( .A(n9275), .ZN(n9276) );
  AOI21_X1 U10489 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(n9279) );
  OAI222_X1 U10490 ( .A1(n9405), .A2(n9280), .B1(n9403), .B2(n9307), .C1(n9400), .C2(n9279), .ZN(n9446) );
  AOI211_X1 U10491 ( .C1(n9282), .C2(n4673), .A(n9390), .B(n9281), .ZN(n9447)
         );
  NAND2_X1 U10492 ( .A1(n9447), .A2(n9397), .ZN(n9285) );
  AOI22_X1 U10493 ( .A1(n9283), .A2(n9339), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9826), .ZN(n9284) );
  OAI211_X1 U10494 ( .C1(n9512), .C2(n9392), .A(n9285), .B(n9284), .ZN(n9286)
         );
  AOI21_X1 U10495 ( .B1(n9446), .B2(n9409), .A(n9286), .ZN(n9287) );
  OAI21_X1 U10496 ( .B1(n9288), .B2(n9408), .A(n9287), .ZN(P1_U3267) );
  XOR2_X1 U10497 ( .A(n9290), .B(n9289), .Z(n9455) );
  XNOR2_X1 U10498 ( .A(n9291), .B(n9290), .ZN(n9292) );
  OAI222_X1 U10499 ( .A1(n9405), .A2(n9294), .B1(n9403), .B2(n9293), .C1(n9292), .C2(n9400), .ZN(n9451) );
  AOI211_X1 U10500 ( .C1(n9453), .C2(n9308), .A(n9390), .B(n9295), .ZN(n9452)
         );
  NAND2_X1 U10501 ( .A1(n9452), .A2(n9818), .ZN(n9299) );
  INV_X1 U10502 ( .A(n9296), .ZN(n9297) );
  AOI22_X1 U10503 ( .A1(n9297), .A2(n9339), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9826), .ZN(n9298) );
  OAI211_X1 U10504 ( .C1(n4671), .C2(n9392), .A(n9299), .B(n9298), .ZN(n9300)
         );
  AOI21_X1 U10505 ( .B1(n9451), .B2(n9409), .A(n9300), .ZN(n9301) );
  OAI21_X1 U10506 ( .B1(n9455), .B2(n9408), .A(n9301), .ZN(P1_U3268) );
  XOR2_X1 U10507 ( .A(n9304), .B(n9302), .Z(n9460) );
  XOR2_X1 U10508 ( .A(n9304), .B(n9303), .Z(n9305) );
  OAI222_X1 U10509 ( .A1(n9405), .A2(n9307), .B1(n9403), .B2(n9306), .C1(n9305), .C2(n9400), .ZN(n9456) );
  INV_X1 U10510 ( .A(n9458), .ZN(n9314) );
  INV_X1 U10511 ( .A(n9308), .ZN(n9309) );
  AOI211_X1 U10512 ( .C1(n9458), .C2(n9325), .A(n9390), .B(n9309), .ZN(n9457)
         );
  NAND2_X1 U10513 ( .A1(n9457), .A2(n9397), .ZN(n9313) );
  INV_X1 U10514 ( .A(n9310), .ZN(n9311) );
  AOI22_X1 U10515 ( .A1(n9311), .A2(n9339), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9826), .ZN(n9312) );
  OAI211_X1 U10516 ( .C1(n9314), .C2(n9392), .A(n9313), .B(n9312), .ZN(n9315)
         );
  AOI21_X1 U10517 ( .B1(n9456), .B2(n9409), .A(n9315), .ZN(n9316) );
  OAI21_X1 U10518 ( .B1(n9460), .B2(n9408), .A(n9316), .ZN(P1_U3269) );
  XNOR2_X1 U10519 ( .A(n9317), .B(n9318), .ZN(n9463) );
  INV_X1 U10520 ( .A(n9463), .ZN(n9334) );
  XNOR2_X1 U10521 ( .A(n9319), .B(n9318), .ZN(n9320) );
  NAND2_X1 U10522 ( .A1(n9320), .A2(n9351), .ZN(n9324) );
  AOI22_X1 U10523 ( .A1(n9322), .A2(n9348), .B1(n9346), .B2(n9321), .ZN(n9323)
         );
  NAND2_X1 U10524 ( .A1(n9324), .A2(n9323), .ZN(n9461) );
  INV_X1 U10525 ( .A(n9336), .ZN(n9327) );
  INV_X1 U10526 ( .A(n9325), .ZN(n9326) );
  AOI211_X1 U10527 ( .C1(n9328), .C2(n9327), .A(n9390), .B(n9326), .ZN(n9462)
         );
  NAND2_X1 U10528 ( .A1(n9462), .A2(n9397), .ZN(n9331) );
  AOI22_X1 U10529 ( .A1(n9826), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9329), .B2(
        n9339), .ZN(n9330) );
  OAI211_X1 U10530 ( .C1(n9518), .C2(n9392), .A(n9331), .B(n9330), .ZN(n9332)
         );
  AOI21_X1 U10531 ( .B1(n9461), .B2(n9409), .A(n9332), .ZN(n9333) );
  OAI21_X1 U10532 ( .B1(n9334), .B2(n9408), .A(n9333), .ZN(P1_U3270) );
  XNOR2_X1 U10533 ( .A(n9335), .B(n9345), .ZN(n9470) );
  INV_X1 U10534 ( .A(n9356), .ZN(n9337) );
  AOI211_X1 U10535 ( .C1(n9467), .C2(n9337), .A(n9390), .B(n9336), .ZN(n9466)
         );
  INV_X1 U10536 ( .A(n9338), .ZN(n9340) );
  AOI22_X1 U10537 ( .A1(n9826), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9340), .B2(
        n9339), .ZN(n9341) );
  OAI21_X1 U10538 ( .B1(n9342), .B2(n9392), .A(n9341), .ZN(n9353) );
  OAI21_X1 U10539 ( .B1(n9345), .B2(n9344), .A(n9343), .ZN(n9350) );
  AOI222_X1 U10540 ( .A1(n9351), .A2(n9350), .B1(n9349), .B2(n9348), .C1(n9347), .C2(n9346), .ZN(n9469) );
  NOR2_X1 U10541 ( .A1(n9469), .A2(n9826), .ZN(n9352) );
  AOI211_X1 U10542 ( .C1(n9466), .C2(n9818), .A(n9353), .B(n9352), .ZN(n9354)
         );
  OAI21_X1 U10543 ( .B1(n9470), .B2(n9408), .A(n9354), .ZN(P1_U3271) );
  XNOR2_X1 U10544 ( .A(n9355), .B(n9362), .ZN(n9475) );
  AOI211_X1 U10545 ( .C1(n9473), .C2(n9376), .A(n9390), .B(n9356), .ZN(n9472)
         );
  INV_X1 U10546 ( .A(n9473), .ZN(n9357) );
  NOR2_X1 U10547 ( .A1(n9357), .A2(n9392), .ZN(n9361) );
  OAI22_X1 U10548 ( .A1(n9409), .A2(n9359), .B1(n9358), .B2(n9820), .ZN(n9360)
         );
  AOI211_X1 U10549 ( .C1(n9472), .C2(n9818), .A(n9361), .B(n9360), .ZN(n9367)
         );
  XNOR2_X1 U10550 ( .A(n9363), .B(n9362), .ZN(n9364) );
  OAI222_X1 U10551 ( .A1(n9405), .A2(n9365), .B1(n9403), .B2(n9404), .C1(n9364), .C2(n9400), .ZN(n9471) );
  NAND2_X1 U10552 ( .A1(n9471), .A2(n9409), .ZN(n9366) );
  OAI211_X1 U10553 ( .C1(n9475), .C2(n9408), .A(n9367), .B(n9366), .ZN(
        P1_U3272) );
  NAND2_X1 U10554 ( .A1(n9369), .A2(n9368), .ZN(n9370) );
  XOR2_X1 U10555 ( .A(n9375), .B(n9370), .Z(n9371) );
  OAI222_X1 U10556 ( .A1(n9405), .A2(n9373), .B1(n9403), .B2(n9372), .C1(n9400), .C2(n9371), .ZN(n9476) );
  INV_X1 U10557 ( .A(n9476), .ZN(n9385) );
  XOR2_X1 U10558 ( .A(n9374), .B(n9375), .Z(n9478) );
  NAND2_X1 U10559 ( .A1(n9478), .A2(n9414), .ZN(n9384) );
  INV_X1 U10560 ( .A(n9376), .ZN(n9377) );
  AOI211_X1 U10561 ( .C1(n9378), .C2(n9388), .A(n9390), .B(n9377), .ZN(n9477)
         );
  INV_X1 U10562 ( .A(n9378), .ZN(n9524) );
  NOR2_X1 U10563 ( .A1(n9524), .A2(n9392), .ZN(n9382) );
  OAI22_X1 U10564 ( .A1(n9409), .A2(n9380), .B1(n9379), .B2(n9820), .ZN(n9381)
         );
  AOI211_X1 U10565 ( .C1(n9477), .C2(n9397), .A(n9382), .B(n9381), .ZN(n9383)
         );
  OAI211_X1 U10566 ( .C1(n9826), .C2(n9385), .A(n9384), .B(n9383), .ZN(
        P1_U3273) );
  XNOR2_X1 U10567 ( .A(n9386), .B(n9398), .ZN(n9485) );
  INV_X1 U10568 ( .A(n9387), .ZN(n9391) );
  INV_X1 U10569 ( .A(n9388), .ZN(n9389) );
  AOI211_X1 U10570 ( .C1(n9483), .C2(n9391), .A(n9390), .B(n9389), .ZN(n9482)
         );
  NOR2_X1 U10571 ( .A1(n9393), .A2(n9392), .ZN(n9396) );
  OAI22_X1 U10572 ( .A1(n9409), .A2(n9156), .B1(n9394), .B2(n9820), .ZN(n9395)
         );
  AOI211_X1 U10573 ( .C1(n9482), .C2(n9397), .A(n9396), .B(n9395), .ZN(n9407)
         );
  XNOR2_X1 U10574 ( .A(n9399), .B(n9398), .ZN(n9401) );
  OAI222_X1 U10575 ( .A1(n9405), .A2(n9404), .B1(n9403), .B2(n9402), .C1(n9401), .C2(n9400), .ZN(n9481) );
  NAND2_X1 U10576 ( .A1(n9481), .A2(n9409), .ZN(n9406) );
  OAI211_X1 U10577 ( .C1(n9485), .C2(n9408), .A(n9407), .B(n9406), .ZN(
        P1_U3274) );
  NAND2_X1 U10578 ( .A1(n9410), .A2(n9409), .ZN(n9420) );
  OAI22_X1 U10579 ( .A1(n9409), .A2(n6537), .B1(n9411), .B2(n9820), .ZN(n9412)
         );
  AOI21_X1 U10580 ( .B1(n9831), .B2(n9413), .A(n9412), .ZN(n9419) );
  NAND2_X1 U10581 ( .A1(n9415), .A2(n9414), .ZN(n9418) );
  NAND2_X1 U10582 ( .A1(n9416), .A2(n9818), .ZN(n9417) );
  NAND4_X1 U10583 ( .A1(n9420), .A2(n9419), .A3(n9418), .A4(n9417), .ZN(
        P1_U3285) );
  INV_X1 U10584 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9423) );
  NOR2_X1 U10585 ( .A1(n9422), .A2(n9421), .ZN(n9492) );
  MUX2_X1 U10586 ( .A(n9423), .B(n9492), .S(n9994), .Z(n9424) );
  OAI21_X1 U10587 ( .B1(n9494), .B2(n9491), .A(n9424), .ZN(P1_U3554) );
  INV_X1 U10588 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9427) );
  AND2_X1 U10589 ( .A1(n9426), .A2(n9425), .ZN(n9495) );
  MUX2_X1 U10590 ( .A(n9427), .B(n9495), .S(n9994), .Z(n9428) );
  OAI21_X1 U10591 ( .B1(n9497), .B2(n9491), .A(n9428), .ZN(P1_U3553) );
  INV_X1 U10592 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9429) );
  INV_X1 U10593 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U10594 ( .A1(n9431), .A2(n9430), .ZN(n9432) );
  AOI21_X1 U10595 ( .B1(n9433), .B2(n9986), .A(n9432), .ZN(n9498) );
  MUX2_X1 U10596 ( .A(n9434), .B(n9498), .S(n9994), .Z(n9435) );
  OAI21_X1 U10597 ( .B1(n4666), .B2(n9491), .A(n9435), .ZN(P1_U3550) );
  INV_X1 U10598 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9439) );
  AOI211_X1 U10599 ( .C1(n9438), .C2(n9986), .A(n9437), .B(n9436), .ZN(n9501)
         );
  MUX2_X1 U10600 ( .A(n9439), .B(n9501), .S(n9994), .Z(n9440) );
  OAI21_X1 U10601 ( .B1(n9504), .B2(n9491), .A(n9440), .ZN(P1_U3549) );
  INV_X1 U10602 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9444) );
  AOI211_X1 U10603 ( .C1(n9443), .C2(n9986), .A(n9442), .B(n9441), .ZN(n9505)
         );
  MUX2_X1 U10604 ( .A(n9444), .B(n9505), .S(n9994), .Z(n9445) );
  OAI21_X1 U10605 ( .B1(n9508), .B2(n9491), .A(n9445), .ZN(P1_U3548) );
  INV_X1 U10606 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9449) );
  AOI211_X1 U10607 ( .C1(n9448), .C2(n9986), .A(n9447), .B(n9446), .ZN(n9509)
         );
  MUX2_X1 U10608 ( .A(n9449), .B(n9509), .S(n9994), .Z(n9450) );
  OAI21_X1 U10609 ( .B1(n9512), .B2(n9491), .A(n9450), .ZN(P1_U3547) );
  INV_X1 U10610 ( .A(n9986), .ZN(n9486) );
  AOI211_X1 U10611 ( .C1(n9843), .C2(n9453), .A(n9452), .B(n9451), .ZN(n9454)
         );
  OAI21_X1 U10612 ( .B1(n9455), .B2(n9486), .A(n9454), .ZN(n9513) );
  MUX2_X1 U10613 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9513), .S(n9994), .Z(
        P1_U3546) );
  AOI211_X1 U10614 ( .C1(n9843), .C2(n9458), .A(n9457), .B(n9456), .ZN(n9459)
         );
  OAI21_X1 U10615 ( .B1(n9460), .B2(n9486), .A(n9459), .ZN(n9514) );
  MUX2_X1 U10616 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9514), .S(n9994), .Z(
        P1_U3545) );
  INV_X1 U10617 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9464) );
  AOI211_X1 U10618 ( .C1(n9463), .C2(n9986), .A(n9462), .B(n9461), .ZN(n9515)
         );
  MUX2_X1 U10619 ( .A(n9464), .B(n9515), .S(n9994), .Z(n9465) );
  OAI21_X1 U10620 ( .B1(n9518), .B2(n9491), .A(n9465), .ZN(P1_U3544) );
  AOI21_X1 U10621 ( .B1(n9843), .B2(n9467), .A(n9466), .ZN(n9468) );
  OAI211_X1 U10622 ( .C1(n9470), .C2(n9486), .A(n9469), .B(n9468), .ZN(n9519)
         );
  MUX2_X1 U10623 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9519), .S(n9994), .Z(
        P1_U3543) );
  AOI211_X1 U10624 ( .C1(n9843), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9474)
         );
  OAI21_X1 U10625 ( .B1(n9475), .B2(n9486), .A(n9474), .ZN(n9520) );
  MUX2_X1 U10626 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9520), .S(n9994), .Z(
        P1_U3542) );
  AOI211_X1 U10627 ( .C1(n9478), .C2(n9986), .A(n9477), .B(n9476), .ZN(n9521)
         );
  MUX2_X1 U10628 ( .A(n9479), .B(n9521), .S(n9994), .Z(n9480) );
  OAI21_X1 U10629 ( .B1(n9524), .B2(n9491), .A(n9480), .ZN(P1_U3541) );
  AOI211_X1 U10630 ( .C1(n9843), .C2(n9483), .A(n9482), .B(n9481), .ZN(n9484)
         );
  OAI21_X1 U10631 ( .B1(n9486), .B2(n9485), .A(n9484), .ZN(n9525) );
  MUX2_X1 U10632 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9525), .S(n9994), .Z(
        P1_U3540) );
  AOI211_X1 U10633 ( .C1(n9489), .C2(n9986), .A(n9488), .B(n9487), .ZN(n9526)
         );
  MUX2_X1 U10634 ( .A(n7504), .B(n9526), .S(n9994), .Z(n9490) );
  OAI21_X1 U10635 ( .B1(n9530), .B2(n9491), .A(n9490), .ZN(P1_U3539) );
  MUX2_X1 U10636 ( .A(n6638), .B(n9492), .S(n9989), .Z(n9493) );
  OAI21_X1 U10637 ( .B1(n9494), .B2(n9529), .A(n9493), .ZN(P1_U3522) );
  MUX2_X1 U10638 ( .A(n9495), .B(n6465), .S(n9988), .Z(n9496) );
  OAI21_X1 U10639 ( .B1(n9497), .B2(n9529), .A(n9496), .ZN(P1_U3521) );
  MUX2_X1 U10640 ( .A(n9499), .B(n9498), .S(n9989), .Z(n9500) );
  OAI21_X1 U10641 ( .B1(n4666), .B2(n9529), .A(n9500), .ZN(P1_U3518) );
  MUX2_X1 U10642 ( .A(n9502), .B(n9501), .S(n9989), .Z(n9503) );
  OAI21_X1 U10643 ( .B1(n9504), .B2(n9529), .A(n9503), .ZN(P1_U3517) );
  MUX2_X1 U10644 ( .A(n9506), .B(n9505), .S(n9989), .Z(n9507) );
  OAI21_X1 U10645 ( .B1(n9508), .B2(n9529), .A(n9507), .ZN(P1_U3516) );
  MUX2_X1 U10646 ( .A(n9510), .B(n9509), .S(n9989), .Z(n9511) );
  OAI21_X1 U10647 ( .B1(n9512), .B2(n9529), .A(n9511), .ZN(P1_U3515) );
  MUX2_X1 U10648 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9513), .S(n9989), .Z(
        P1_U3514) );
  MUX2_X1 U10649 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9514), .S(n9989), .Z(
        P1_U3513) );
  INV_X1 U10650 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9516) );
  MUX2_X1 U10651 ( .A(n9516), .B(n9515), .S(n9989), .Z(n9517) );
  OAI21_X1 U10652 ( .B1(n9518), .B2(n9529), .A(n9517), .ZN(P1_U3512) );
  MUX2_X1 U10653 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9519), .S(n9989), .Z(
        P1_U3511) );
  MUX2_X1 U10654 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9520), .S(n9989), .Z(
        P1_U3510) );
  INV_X1 U10655 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9522) );
  MUX2_X1 U10656 ( .A(n9522), .B(n9521), .S(n9989), .Z(n9523) );
  OAI21_X1 U10657 ( .B1(n9524), .B2(n9529), .A(n9523), .ZN(P1_U3508) );
  MUX2_X1 U10658 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9525), .S(n9989), .Z(
        P1_U3505) );
  INV_X1 U10659 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9527) );
  MUX2_X1 U10660 ( .A(n9527), .B(n9526), .S(n9989), .Z(n9528) );
  OAI21_X1 U10661 ( .B1(n9530), .B2(n9529), .A(n9528), .ZN(P1_U3502) );
  NOR4_X1 U10662 ( .A1(n9531), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5899), .A4(
        P1_U3084), .ZN(n9532) );
  AOI21_X1 U10663 ( .B1(n9535), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9532), .ZN(
        n9533) );
  OAI21_X1 U10664 ( .B1(n9534), .B2(n9537), .A(n9533), .ZN(P1_U3322) );
  NAND2_X1 U10665 ( .A1(n9535), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9536) );
  OAI211_X1 U10666 ( .C1(n9538), .C2(n9537), .A(n9864), .B(n9536), .ZN(
        P1_U3325) );
  MUX2_X1 U10667 ( .A(n9539), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U10668 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10157) );
  NOR2_X1 U10669 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9540) );
  AOI21_X1 U10670 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9540), .ZN(n10128) );
  NOR2_X1 U10671 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9541) );
  AOI21_X1 U10672 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9541), .ZN(n10131) );
  NOR2_X1 U10673 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9542) );
  AOI21_X1 U10674 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9542), .ZN(n10134) );
  NOR2_X1 U10675 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9543) );
  AOI21_X1 U10676 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9543), .ZN(n10137) );
  NOR2_X1 U10677 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9544) );
  AOI21_X1 U10678 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9544), .ZN(n10140) );
  INV_X1 U10679 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9931) );
  NOR2_X1 U10680 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9550) );
  XOR2_X1 U10681 ( .A(n9916), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10167) );
  NAND2_X1 U10682 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9548) );
  XOR2_X1 U10683 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10165) );
  NAND2_X1 U10684 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9546) );
  INV_X1 U10685 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9901) );
  XNOR2_X1 U10686 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9901), .ZN(n10153) );
  AOI21_X1 U10687 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10121) );
  NAND3_X1 U10688 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10123) );
  OAI21_X1 U10689 ( .B1(n10121), .B2(n10125), .A(n10123), .ZN(n10152) );
  NAND2_X1 U10690 ( .A1(n10153), .A2(n10152), .ZN(n9545) );
  NAND2_X1 U10691 ( .A1(n9546), .A2(n9545), .ZN(n10164) );
  NAND2_X1 U10692 ( .A1(n10165), .A2(n10164), .ZN(n9547) );
  NAND2_X1 U10693 ( .A1(n9548), .A2(n9547), .ZN(n10166) );
  NAND2_X1 U10694 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10162), .ZN(n9551) );
  NOR2_X1 U10695 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10162), .ZN(n10161) );
  AOI21_X1 U10696 ( .B1(n9931), .B2(n9551), .A(n10161), .ZN(n9552) );
  NAND2_X1 U10697 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n9552), .ZN(n9554) );
  XOR2_X1 U10698 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n9552), .Z(n10160) );
  NAND2_X1 U10699 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10160), .ZN(n9553) );
  NAND2_X1 U10700 ( .A1(n9554), .A2(n9553), .ZN(n9555) );
  NAND2_X1 U10701 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9555), .ZN(n9558) );
  INV_X1 U10702 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9556) );
  XNOR2_X1 U10703 ( .A(n9556), .B(n9555), .ZN(n10159) );
  NAND2_X1 U10704 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10159), .ZN(n9557) );
  NAND2_X1 U10705 ( .A1(n9558), .A2(n9557), .ZN(n9559) );
  NAND2_X1 U10706 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9559), .ZN(n9561) );
  XOR2_X1 U10707 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9559), .Z(n10154) );
  NAND2_X1 U10708 ( .A1(n10154), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U10709 ( .A1(n9561), .A2(n9560), .ZN(n10150) );
  AOI222_X1 U10710 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .B1(P2_ADDR_REG_9__SCAN_IN), .B2(n10150), .C1(P1_ADDR_REG_9__SCAN_IN), 
        .C2(n10150), .ZN(n10149) );
  NAND2_X1 U10711 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9562) );
  OAI21_X1 U10712 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9562), .ZN(n10148) );
  NOR2_X1 U10713 ( .A1(n10149), .A2(n10148), .ZN(n10147) );
  AOI21_X1 U10714 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10147), .ZN(n10146) );
  NAND2_X1 U10715 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9563) );
  OAI21_X1 U10716 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9563), .ZN(n10145) );
  NOR2_X1 U10717 ( .A1(n10146), .A2(n10145), .ZN(n10144) );
  AOI21_X1 U10718 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10144), .ZN(n10143) );
  NOR2_X1 U10719 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9564) );
  AOI21_X1 U10720 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9564), .ZN(n10142) );
  NAND2_X1 U10721 ( .A1(n10143), .A2(n10142), .ZN(n10141) );
  OAI21_X1 U10722 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10141), .ZN(n10139) );
  NAND2_X1 U10723 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  OAI21_X1 U10724 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10138), .ZN(n10136) );
  NAND2_X1 U10725 ( .A1(n10137), .A2(n10136), .ZN(n10135) );
  OAI21_X1 U10726 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10135), .ZN(n10133) );
  NAND2_X1 U10727 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  OAI21_X1 U10728 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10132), .ZN(n10130) );
  NAND2_X1 U10729 ( .A1(n10131), .A2(n10130), .ZN(n10129) );
  OAI21_X1 U10730 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10129), .ZN(n10127) );
  NAND2_X1 U10731 ( .A1(n10128), .A2(n10127), .ZN(n10126) );
  OAI21_X1 U10732 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10126), .ZN(n10156) );
  NOR2_X1 U10733 ( .A1(n10157), .A2(n10156), .ZN(n9565) );
  NAND2_X1 U10734 ( .A1(n10157), .A2(n10156), .ZN(n10155) );
  OAI21_X1 U10735 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n9565), .A(n10155), .ZN(
        n9757) );
  AOI22_X1 U10736 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_f41), .ZN(n9566) );
  OAI221_X1 U10737 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_f41), .A(n9566), .ZN(n9573) );
  AOI22_X1 U10738 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(keyinput_f55), .B1(
        P2_REG3_REG_28__SCAN_IN), .B2(keyinput_f42), .ZN(n9567) );
  OAI221_X1 U10739 ( .B1(P2_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_f42), .A(n9567), .ZN(n9572) );
  AOI22_X1 U10740 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        SI_17_), .B2(keyinput_f15), .ZN(n9568) );
  OAI221_X1 U10741 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        SI_17_), .C2(keyinput_f15), .A(n9568), .ZN(n9571) );
  AOI22_X1 U10742 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(SI_22_), .B2(keyinput_f10), .ZN(n9569) );
  OAI221_X1 U10743 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        SI_22_), .C2(keyinput_f10), .A(n9569), .ZN(n9570) );
  NOR4_X1 U10744 ( .A1(n9573), .A2(n9572), .A3(n9571), .A4(n9570), .ZN(n9602)
         );
  INV_X1 U10745 ( .A(SI_21_), .ZN(n9690) );
  XNOR2_X1 U10746 ( .A(n9690), .B(keyinput_f11), .ZN(n9580) );
  AOI22_X1 U10747 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_2_), .B2(
        keyinput_f30), .ZN(n9574) );
  OAI221_X1 U10748 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_2_), .C2(
        keyinput_f30), .A(n9574), .ZN(n9579) );
  AOI22_X1 U10749 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        SI_25_), .B2(keyinput_f7), .ZN(n9575) );
  OAI221_X1 U10750 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        SI_25_), .C2(keyinput_f7), .A(n9575), .ZN(n9578) );
  AOI22_X1 U10751 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_26_), .B2(
        keyinput_f6), .ZN(n9576) );
  OAI221_X1 U10752 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_26_), .C2(
        keyinput_f6), .A(n9576), .ZN(n9577) );
  NOR4_X1 U10753 ( .A1(n9580), .A2(n9579), .A3(n9578), .A4(n9577), .ZN(n9601)
         );
  AOI22_X1 U10754 ( .A1(n9582), .A2(keyinput_f37), .B1(keyinput_f56), .B2(
        n6989), .ZN(n9581) );
  OAI221_X1 U10755 ( .B1(n9582), .B2(keyinput_f37), .C1(n6989), .C2(
        keyinput_f56), .A(n9581), .ZN(n9590) );
  AOI22_X1 U10756 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput_f47), .B1(
        SI_28_), .B2(keyinput_f4), .ZN(n9583) );
  OAI221_X1 U10757 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .C1(
        SI_28_), .C2(keyinput_f4), .A(n9583), .ZN(n9589) );
  AOI22_X1 U10758 ( .A1(keyinput_f0), .A2(P2_WR_REG_SCAN_IN), .B1(SI_14_), 
        .B2(keyinput_f18), .ZN(n9584) );
  OAI221_X1 U10759 ( .B1(keyinput_f0), .B2(P2_WR_REG_SCAN_IN), .C1(SI_14_), 
        .C2(keyinput_f18), .A(n9584), .ZN(n9588) );
  XNOR2_X1 U10760 ( .A(SI_1_), .B(keyinput_f31), .ZN(n9586) );
  XNOR2_X1 U10761 ( .A(SI_9_), .B(keyinput_f23), .ZN(n9585) );
  NAND2_X1 U10762 ( .A1(n9586), .A2(n9585), .ZN(n9587) );
  NOR4_X1 U10763 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n9600)
         );
  AOI22_X1 U10764 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_f54), .B1(
        P2_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n9591) );
  OAI221_X1 U10765 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_f54), .C1(
        P2_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n9591), .ZN(n9598) );
  AOI22_X1 U10766 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        SI_23_), .B2(keyinput_f9), .ZN(n9592) );
  OAI221_X1 U10767 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_23_), .C2(keyinput_f9), .A(n9592), .ZN(n9597) );
  AOI22_X1 U10768 ( .A1(SI_3_), .A2(keyinput_f29), .B1(SI_11_), .B2(
        keyinput_f21), .ZN(n9593) );
  OAI221_X1 U10769 ( .B1(SI_3_), .B2(keyinput_f29), .C1(SI_11_), .C2(
        keyinput_f21), .A(n9593), .ZN(n9596) );
  AOI22_X1 U10770 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_f62), .B1(
        SI_15_), .B2(keyinput_f17), .ZN(n9594) );
  OAI221_X1 U10771 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .C1(
        SI_15_), .C2(keyinput_f17), .A(n9594), .ZN(n9595) );
  NOR4_X1 U10772 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n9599)
         );
  NAND4_X1 U10773 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n9648)
         );
  INV_X1 U10774 ( .A(SI_24_), .ZN(n9721) );
  AOI22_X1 U10775 ( .A1(n9721), .A2(keyinput_f8), .B1(keyinput_f53), .B2(n5108), .ZN(n9603) );
  OAI221_X1 U10776 ( .B1(n9721), .B2(keyinput_f8), .C1(n5108), .C2(
        keyinput_f53), .A(n9603), .ZN(n9612) );
  AOI22_X1 U10777 ( .A1(n9659), .A2(keyinput_f32), .B1(keyinput_f38), .B2(
        n9724), .ZN(n9604) );
  OAI221_X1 U10778 ( .B1(n9659), .B2(keyinput_f32), .C1(n9724), .C2(
        keyinput_f38), .A(n9604), .ZN(n9611) );
  AOI22_X1 U10779 ( .A1(P2_U3152), .A2(keyinput_f34), .B1(keyinput_f36), .B2(
        n9734), .ZN(n9605) );
  OAI221_X1 U10780 ( .B1(P2_U3152), .B2(keyinput_f34), .C1(n9734), .C2(
        keyinput_f36), .A(n9605), .ZN(n9610) );
  XNOR2_X1 U10781 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_f33), .ZN(n9608) );
  XNOR2_X1 U10782 ( .A(SI_4_), .B(keyinput_f28), .ZN(n9607) );
  NAND2_X1 U10783 ( .A1(n9608), .A2(n9607), .ZN(n9609) );
  NOR4_X1 U10784 ( .A1(n9612), .A2(n9611), .A3(n9610), .A4(n9609), .ZN(n9646)
         );
  AOI22_X1 U10785 ( .A1(n9740), .A2(keyinput_f61), .B1(n9735), .B2(
        keyinput_f48), .ZN(n9613) );
  OAI221_X1 U10786 ( .B1(n9740), .B2(keyinput_f61), .C1(n9735), .C2(
        keyinput_f48), .A(n9613), .ZN(n9620) );
  AOI22_X1 U10787 ( .A1(n9719), .A2(keyinput_f43), .B1(keyinput_f44), .B2(
        n9699), .ZN(n9614) );
  OAI221_X1 U10788 ( .B1(n9719), .B2(keyinput_f43), .C1(n9699), .C2(
        keyinput_f44), .A(n9614), .ZN(n9619) );
  INV_X1 U10789 ( .A(SI_19_), .ZN(n9742) );
  INV_X1 U10790 ( .A(SI_6_), .ZN(n9696) );
  AOI22_X1 U10791 ( .A1(n9742), .A2(keyinput_f13), .B1(keyinput_f26), .B2(
        n9696), .ZN(n9615) );
  OAI221_X1 U10792 ( .B1(n9742), .B2(keyinput_f13), .C1(n9696), .C2(
        keyinput_f26), .A(n9615), .ZN(n9618) );
  AOI22_X1 U10793 ( .A1(n9737), .A2(keyinput_f5), .B1(keyinput_f35), .B2(n5055), .ZN(n9616) );
  OAI221_X1 U10794 ( .B1(n9737), .B2(keyinput_f5), .C1(n5055), .C2(
        keyinput_f35), .A(n9616), .ZN(n9617) );
  NOR4_X1 U10795 ( .A1(n9620), .A2(n9619), .A3(n9618), .A4(n9617), .ZN(n9645)
         );
  AOI22_X1 U10796 ( .A1(n9738), .A2(keyinput_f16), .B1(keyinput_f51), .B2(
        n9705), .ZN(n9621) );
  OAI221_X1 U10797 ( .B1(n9738), .B2(keyinput_f16), .C1(n9705), .C2(
        keyinput_f51), .A(n9621), .ZN(n9630) );
  INV_X1 U10798 ( .A(SI_13_), .ZN(n9623) );
  AOI22_X1 U10799 ( .A1(n9691), .A2(keyinput_f50), .B1(n9623), .B2(
        keyinput_f19), .ZN(n9622) );
  OAI221_X1 U10800 ( .B1(n9691), .B2(keyinput_f50), .C1(n9623), .C2(
        keyinput_f19), .A(n9622), .ZN(n9629) );
  INV_X1 U10801 ( .A(SI_7_), .ZN(n9710) );
  AOI22_X1 U10802 ( .A1(n9710), .A2(keyinput_f25), .B1(keyinput_f59), .B2(
        n9625), .ZN(n9624) );
  OAI221_X1 U10803 ( .B1(n9710), .B2(keyinput_f25), .C1(n9625), .C2(
        keyinput_f59), .A(n9624), .ZN(n9628) );
  INV_X1 U10804 ( .A(SI_31_), .ZN(n9718) );
  AOI22_X1 U10805 ( .A1(n9708), .A2(keyinput_f45), .B1(keyinput_f1), .B2(n9718), .ZN(n9626) );
  OAI221_X1 U10806 ( .B1(n9708), .B2(keyinput_f45), .C1(n9718), .C2(
        keyinput_f1), .A(n9626), .ZN(n9627) );
  NOR4_X1 U10807 ( .A1(n9630), .A2(n9629), .A3(n9628), .A4(n9627), .ZN(n9644)
         );
  AOI22_X1 U10808 ( .A1(n5145), .A2(keyinput_f58), .B1(keyinput_f52), .B2(
        n9671), .ZN(n9631) );
  OAI221_X1 U10809 ( .B1(n5145), .B2(keyinput_f58), .C1(n9671), .C2(
        keyinput_f52), .A(n9631), .ZN(n9642) );
  AOI22_X1 U10810 ( .A1(n9670), .A2(keyinput_f22), .B1(n9633), .B2(
        keyinput_f12), .ZN(n9632) );
  OAI221_X1 U10811 ( .B1(n9670), .B2(keyinput_f22), .C1(n9633), .C2(
        keyinput_f12), .A(n9632), .ZN(n9641) );
  AOI22_X1 U10812 ( .A1(n9636), .A2(keyinput_f27), .B1(keyinput_f3), .B2(n9635), .ZN(n9634) );
  OAI221_X1 U10813 ( .B1(n9636), .B2(keyinput_f27), .C1(n9635), .C2(
        keyinput_f3), .A(n9634), .ZN(n9640) );
  INV_X1 U10814 ( .A(SI_18_), .ZN(n9722) );
  AOI22_X1 U10815 ( .A1(n9638), .A2(keyinput_f24), .B1(n9722), .B2(
        keyinput_f14), .ZN(n9637) );
  OAI221_X1 U10816 ( .B1(n9638), .B2(keyinput_f24), .C1(n9722), .C2(
        keyinput_f14), .A(n9637), .ZN(n9639) );
  NOR4_X1 U10817 ( .A1(n9642), .A2(n9641), .A3(n9640), .A4(n9639), .ZN(n9643)
         );
  NAND4_X1 U10818 ( .A1(n9646), .A2(n9645), .A3(n9644), .A4(n9643), .ZN(n9647)
         );
  OAI22_X1 U10819 ( .A1(keyinput_f60), .A2(n9650), .B1(n9648), .B2(n9647), 
        .ZN(n9649) );
  AOI21_X1 U10820 ( .B1(keyinput_f60), .B2(n9650), .A(n9649), .ZN(n9755) );
  AOI22_X1 U10821 ( .A1(P2_REG3_REG_28__SCAN_IN), .A2(keyinput_g42), .B1(
        SI_15_), .B2(keyinput_g17), .ZN(n9651) );
  OAI221_X1 U10822 ( .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .C1(
        SI_15_), .C2(keyinput_g17), .A(n9651), .ZN(n9658) );
  AOI22_X1 U10823 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_22_), .B2(
        keyinput_g10), .ZN(n9652) );
  OAI221_X1 U10824 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_22_), .C2(
        keyinput_g10), .A(n9652), .ZN(n9657) );
  AOI22_X1 U10825 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(keyinput_g57), .B1(
        SI_13_), .B2(keyinput_g19), .ZN(n9653) );
  OAI221_X1 U10826 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .C1(
        SI_13_), .C2(keyinput_g19), .A(n9653), .ZN(n9656) );
  AOI22_X1 U10827 ( .A1(SI_29_), .A2(keyinput_g3), .B1(SI_5_), .B2(
        keyinput_g27), .ZN(n9654) );
  OAI221_X1 U10828 ( .B1(SI_29_), .B2(keyinput_g3), .C1(SI_5_), .C2(
        keyinput_g27), .A(n9654), .ZN(n9655) );
  NOR4_X1 U10829 ( .A1(n9658), .A2(n9657), .A3(n9656), .A4(n9655), .ZN(n9688)
         );
  XOR2_X1 U10830 ( .A(n9659), .B(keyinput_g32), .Z(n9666) );
  AOI22_X1 U10831 ( .A1(SI_20_), .A2(keyinput_g12), .B1(n5055), .B2(
        keyinput_g35), .ZN(n9660) );
  OAI221_X1 U10832 ( .B1(SI_20_), .B2(keyinput_g12), .C1(n5055), .C2(
        keyinput_g35), .A(n9660), .ZN(n9665) );
  AOI22_X1 U10833 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_g63), .B1(
        P2_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n9661) );
  OAI221_X1 U10834 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .C1(
        P2_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n9661), .ZN(n9664) );
  AOI22_X1 U10835 ( .A1(SI_4_), .A2(keyinput_g28), .B1(SI_9_), .B2(
        keyinput_g23), .ZN(n9662) );
  OAI221_X1 U10836 ( .B1(SI_4_), .B2(keyinput_g28), .C1(SI_9_), .C2(
        keyinput_g23), .A(n9662), .ZN(n9663) );
  NOR4_X1 U10837 ( .A1(n9666), .A2(n9665), .A3(n9664), .A4(n9663), .ZN(n9687)
         );
  AOI22_X1 U10838 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_g62), .B1(
        SI_11_), .B2(keyinput_g21), .ZN(n9667) );
  OAI221_X1 U10839 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .C1(
        SI_11_), .C2(keyinput_g21), .A(n9667), .ZN(n9676) );
  AOI22_X1 U10840 ( .A1(SI_17_), .A2(keyinput_g15), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_g33), .ZN(n9668) );
  OAI221_X1 U10841 ( .B1(SI_17_), .B2(keyinput_g15), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_g33), .A(n9668), .ZN(n9675) );
  AOI22_X1 U10842 ( .A1(n9671), .A2(keyinput_g52), .B1(n9670), .B2(
        keyinput_g22), .ZN(n9669) );
  OAI221_X1 U10843 ( .B1(n9671), .B2(keyinput_g52), .C1(n9670), .C2(
        keyinput_g22), .A(n9669), .ZN(n9674) );
  INV_X1 U10844 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9857) );
  AOI22_X1 U10845 ( .A1(n5016), .A2(keyinput_g49), .B1(keyinput_g0), .B2(n9857), .ZN(n9672) );
  OAI221_X1 U10846 ( .B1(n5016), .B2(keyinput_g49), .C1(n9857), .C2(
        keyinput_g0), .A(n9672), .ZN(n9673) );
  NOR4_X1 U10847 ( .A1(n9676), .A2(n9675), .A3(n9674), .A4(n9673), .ZN(n9686)
         );
  AOI22_X1 U10848 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_2_), 
        .B2(keyinput_g30), .ZN(n9677) );
  OAI221_X1 U10849 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(SI_2_), .C2(keyinput_g30), .A(n9677), .ZN(n9684) );
  AOI22_X1 U10850 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_25_), .B2(
        keyinput_g7), .ZN(n9678) );
  OAI221_X1 U10851 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_25_), .C2(
        keyinput_g7), .A(n9678), .ZN(n9683) );
  AOI22_X1 U10852 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_g37), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n9679) );
  OAI221_X1 U10853 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .C1(
        P2_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n9679), .ZN(n9682) );
  AOI22_X1 U10854 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(SI_8_), .B2(keyinput_g24), .ZN(n9680) );
  OAI221_X1 U10855 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        SI_8_), .C2(keyinput_g24), .A(n9680), .ZN(n9681) );
  NOR4_X1 U10856 ( .A1(n9684), .A2(n9683), .A3(n9682), .A4(n9681), .ZN(n9685)
         );
  NAND4_X1 U10857 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n9753)
         );
  AOI22_X1 U10858 ( .A1(n9691), .A2(keyinput_g50), .B1(n9690), .B2(
        keyinput_g11), .ZN(n9689) );
  OAI221_X1 U10859 ( .B1(n9691), .B2(keyinput_g50), .C1(n9690), .C2(
        keyinput_g11), .A(n9689), .ZN(n9703) );
  INV_X1 U10860 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9693) );
  AOI22_X1 U10861 ( .A1(n9694), .A2(keyinput_g55), .B1(keyinput_g54), .B2(
        n9693), .ZN(n9692) );
  OAI221_X1 U10862 ( .B1(n9694), .B2(keyinput_g55), .C1(n9693), .C2(
        keyinput_g54), .A(n9692), .ZN(n9702) );
  AOI22_X1 U10863 ( .A1(n9696), .A2(keyinput_g26), .B1(keyinput_g4), .B2(n5472), .ZN(n9695) );
  OAI221_X1 U10864 ( .B1(n9696), .B2(keyinput_g26), .C1(n5472), .C2(
        keyinput_g4), .A(n9695), .ZN(n9701) );
  AOI22_X1 U10865 ( .A1(n9699), .A2(keyinput_g44), .B1(n9698), .B2(keyinput_g9), .ZN(n9697) );
  OAI221_X1 U10866 ( .B1(n9699), .B2(keyinput_g44), .C1(n9698), .C2(
        keyinput_g9), .A(n9697), .ZN(n9700) );
  NOR4_X1 U10867 ( .A1(n9703), .A2(n9702), .A3(n9701), .A4(n9700), .ZN(n9751)
         );
  AOI22_X1 U10868 ( .A1(n9706), .A2(keyinput_g40), .B1(n9705), .B2(
        keyinput_g51), .ZN(n9704) );
  OAI221_X1 U10869 ( .B1(n9706), .B2(keyinput_g40), .C1(n9705), .C2(
        keyinput_g51), .A(n9704), .ZN(n9716) );
  AOI22_X1 U10870 ( .A1(n9708), .A2(keyinput_g45), .B1(keyinput_g53), .B2(
        n5108), .ZN(n9707) );
  OAI221_X1 U10871 ( .B1(n9708), .B2(keyinput_g45), .C1(n5108), .C2(
        keyinput_g53), .A(n9707), .ZN(n9715) );
  AOI22_X1 U10872 ( .A1(n5145), .A2(keyinput_g58), .B1(n9710), .B2(
        keyinput_g25), .ZN(n9709) );
  OAI221_X1 U10873 ( .B1(n5145), .B2(keyinput_g58), .C1(n9710), .C2(
        keyinput_g25), .A(n9709), .ZN(n9714) );
  AOI22_X1 U10874 ( .A1(n9712), .A2(keyinput_g47), .B1(keyinput_g56), .B2(
        n6989), .ZN(n9711) );
  OAI221_X1 U10875 ( .B1(n9712), .B2(keyinput_g47), .C1(n6989), .C2(
        keyinput_g56), .A(n9711), .ZN(n9713) );
  NOR4_X1 U10876 ( .A1(n9716), .A2(n9715), .A3(n9714), .A4(n9713), .ZN(n9750)
         );
  AOI22_X1 U10877 ( .A1(n9719), .A2(keyinput_g43), .B1(keyinput_g1), .B2(n9718), .ZN(n9717) );
  OAI221_X1 U10878 ( .B1(n9719), .B2(keyinput_g43), .C1(n9718), .C2(
        keyinput_g1), .A(n9717), .ZN(n9732) );
  AOI22_X1 U10879 ( .A1(n9722), .A2(keyinput_g14), .B1(n9721), .B2(keyinput_g8), .ZN(n9720) );
  OAI221_X1 U10880 ( .B1(n9722), .B2(keyinput_g14), .C1(n9721), .C2(
        keyinput_g8), .A(n9720), .ZN(n9731) );
  AOI22_X1 U10881 ( .A1(n9725), .A2(keyinput_g39), .B1(n9724), .B2(
        keyinput_g38), .ZN(n9723) );
  OAI221_X1 U10882 ( .B1(n9725), .B2(keyinput_g39), .C1(n9724), .C2(
        keyinput_g38), .A(n9723), .ZN(n9730) );
  INV_X1 U10883 ( .A(SI_12_), .ZN(n9726) );
  XOR2_X1 U10884 ( .A(n9726), .B(keyinput_g20), .Z(n9728) );
  XNOR2_X1 U10885 ( .A(SI_1_), .B(keyinput_g31), .ZN(n9727) );
  NAND2_X1 U10886 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  NOR4_X1 U10887 ( .A1(n9732), .A2(n9731), .A3(n9730), .A4(n9729), .ZN(n9749)
         );
  AOI22_X1 U10888 ( .A1(n9735), .A2(keyinput_g48), .B1(n9734), .B2(
        keyinput_g36), .ZN(n9733) );
  OAI221_X1 U10889 ( .B1(n9735), .B2(keyinput_g48), .C1(n9734), .C2(
        keyinput_g36), .A(n9733), .ZN(n9747) );
  AOI22_X1 U10890 ( .A1(n9738), .A2(keyinput_g16), .B1(n9737), .B2(keyinput_g5), .ZN(n9736) );
  OAI221_X1 U10891 ( .B1(n9738), .B2(keyinput_g16), .C1(n9737), .C2(
        keyinput_g5), .A(n9736), .ZN(n9746) );
  AOI22_X1 U10892 ( .A1(n9740), .A2(keyinput_g61), .B1(keyinput_g2), .B2(n5497), .ZN(n9739) );
  OAI221_X1 U10893 ( .B1(n9740), .B2(keyinput_g61), .C1(n5497), .C2(
        keyinput_g2), .A(n9739), .ZN(n9745) );
  AOI22_X1 U10894 ( .A1(n9743), .A2(keyinput_g6), .B1(keyinput_g13), .B2(n9742), .ZN(n9741) );
  OAI221_X1 U10895 ( .B1(n9743), .B2(keyinput_g6), .C1(n9742), .C2(
        keyinput_g13), .A(n9741), .ZN(n9744) );
  NOR4_X1 U10896 ( .A1(n9747), .A2(n9746), .A3(n9745), .A4(n9744), .ZN(n9748)
         );
  NAND4_X1 U10897 ( .A1(n9751), .A2(n9750), .A3(n9749), .A4(n9748), .ZN(n9752)
         );
  OAI22_X1 U10898 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(n9753), .B2(n9752), .ZN(n9754) );
  AOI211_X1 U10899 ( .C1(P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n9755), .B(n9754), .ZN(n9756) );
  XNOR2_X1 U10900 ( .A(n9757), .B(n9756), .ZN(n9761) );
  NOR2_X1 U10901 ( .A1(n9758), .A2(n9759), .ZN(n9760) );
  XOR2_X1 U10902 ( .A(n9761), .B(n9760), .Z(ADD_1071_U4) );
  INV_X1 U10903 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9763) );
  OAI22_X1 U10904 ( .A1(n9964), .A2(n9763), .B1(n9943), .B2(n9762), .ZN(n9764)
         );
  INV_X1 U10905 ( .A(n9764), .ZN(n9775) );
  AOI21_X1 U10906 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9768) );
  NAND2_X1 U10907 ( .A1(n9959), .A2(n9768), .ZN(n9773) );
  OAI211_X1 U10908 ( .C1(n9771), .C2(n9770), .A(n9960), .B(n9769), .ZN(n9772)
         );
  NAND4_X1 U10909 ( .A1(n9775), .A2(n9774), .A3(n9773), .A4(n9772), .ZN(
        P1_U3244) );
  AOI22_X1 U10910 ( .A1(n10002), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9787) );
  AOI211_X1 U10911 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n10000), .ZN(n9779)
         );
  AOI21_X1 U10912 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9786) );
  OAI211_X1 U10913 ( .C1(n9784), .C2(n9783), .A(n9997), .B(n9782), .ZN(n9785)
         );
  NAND3_X1 U10914 ( .A1(n9787), .A2(n9786), .A3(n9785), .ZN(P2_U3247) );
  OAI211_X1 U10915 ( .C1(n9790), .C2(n9982), .A(n9789), .B(n9788), .ZN(n9791)
         );
  AOI21_X1 U10916 ( .B1(n9986), .B2(n9792), .A(n9791), .ZN(n9794) );
  INV_X1 U10917 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9793) );
  AOI22_X1 U10918 ( .A1(n9989), .A2(n9794), .B1(n9793), .B2(n9988), .ZN(
        P1_U3484) );
  AOI22_X1 U10919 ( .A1(n9994), .A2(n9794), .B1(n5970), .B2(n9992), .ZN(
        P1_U3533) );
  INV_X1 U10920 ( .A(n10088), .ZN(n10094) );
  OAI22_X1 U10921 ( .A1(n9796), .A2(n10096), .B1(n9795), .B2(n10094), .ZN(
        n9798) );
  AOI211_X1 U10922 ( .C1(n10101), .C2(n9799), .A(n9798), .B(n9797), .ZN(n9812)
         );
  AOI22_X1 U10923 ( .A1(n10120), .A2(n9812), .B1(n9800), .B2(n10118), .ZN(
        P2_U3535) );
  OAI22_X1 U10924 ( .A1(n9802), .A2(n10096), .B1(n9801), .B2(n10094), .ZN(
        n9804) );
  AOI211_X1 U10925 ( .C1(n9805), .C2(n10101), .A(n9804), .B(n9803), .ZN(n9814)
         );
  AOI22_X1 U10926 ( .A1(n10120), .A2(n9814), .B1(n5207), .B2(n10118), .ZN(
        P2_U3534) );
  INV_X1 U10927 ( .A(n9806), .ZN(n10084) );
  OAI22_X1 U10928 ( .A1(n9807), .A2(n10096), .B1(n4578), .B2(n10094), .ZN(
        n9808) );
  AOI21_X1 U10929 ( .B1(n9809), .B2(n10084), .A(n9808), .ZN(n9810) );
  AND2_X1 U10930 ( .A1(n9811), .A2(n9810), .ZN(n9816) );
  AOI22_X1 U10931 ( .A1(n10120), .A2(n9816), .B1(n5185), .B2(n10118), .ZN(
        P2_U3533) );
  AOI22_X1 U10932 ( .A1(n10104), .A2(n9812), .B1(n5226), .B2(n10102), .ZN(
        P2_U3496) );
  INV_X1 U10933 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9813) );
  AOI22_X1 U10934 ( .A1(n10104), .A2(n9814), .B1(n9813), .B2(n10102), .ZN(
        P2_U3493) );
  INV_X1 U10935 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U10936 ( .A1(n10104), .A2(n9816), .B1(n9815), .B2(n10102), .ZN(
        P2_U3490) );
  AOI22_X1 U10937 ( .A1(n9825), .A2(n9819), .B1(n9818), .B2(n9817), .ZN(n9833)
         );
  OAI22_X1 U10938 ( .A1(n9409), .A2(n9822), .B1(n9821), .B2(n9820), .ZN(n9829)
         );
  AOI21_X1 U10939 ( .B1(n9825), .B2(n9824), .A(n9823), .ZN(n9827) );
  NOR2_X1 U10940 ( .A1(n9827), .A2(n9826), .ZN(n9828) );
  AOI211_X1 U10941 ( .C1(n9831), .C2(n9830), .A(n9829), .B(n9828), .ZN(n9832)
         );
  NAND2_X1 U10942 ( .A1(n9833), .A2(n9832), .ZN(P1_U3278) );
  OAI211_X1 U10943 ( .C1(n9836), .C2(n9982), .A(n9835), .B(n9834), .ZN(n9837)
         );
  AOI21_X1 U10944 ( .B1(n9986), .B2(n9838), .A(n9837), .ZN(n9852) );
  AOI22_X1 U10945 ( .A1(n9994), .A2(n9852), .B1(n6079), .B2(n9992), .ZN(
        P1_U3538) );
  OAI211_X1 U10946 ( .C1(n4676), .C2(n9982), .A(n9840), .B(n9839), .ZN(n9841)
         );
  AOI21_X1 U10947 ( .B1(n9842), .B2(n9986), .A(n9841), .ZN(n9854) );
  AOI22_X1 U10948 ( .A1(n9994), .A2(n9854), .B1(n6964), .B2(n9992), .ZN(
        P1_U3537) );
  NAND2_X1 U10949 ( .A1(n9844), .A2(n9843), .ZN(n9845) );
  NAND2_X1 U10950 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  AOI21_X1 U10951 ( .B1(n9848), .B2(n9973), .A(n9847), .ZN(n9849) );
  AND2_X1 U10952 ( .A1(n9850), .A2(n9849), .ZN(n9856) );
  AOI22_X1 U10953 ( .A1(n9994), .A2(n9856), .B1(n5988), .B2(n9992), .ZN(
        P1_U3534) );
  INV_X1 U10954 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10955 ( .A1(n9989), .A2(n9852), .B1(n9851), .B2(n9988), .ZN(
        P1_U3499) );
  INV_X1 U10956 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9853) );
  AOI22_X1 U10957 ( .A1(n9989), .A2(n9854), .B1(n9853), .B2(n9988), .ZN(
        P1_U3496) );
  INV_X1 U10958 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U10959 ( .A1(n9989), .A2(n9856), .B1(n9855), .B2(n9988), .ZN(
        P1_U3487) );
  XOR2_X1 U10960 ( .A(n9857), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  NOR2_X1 U10961 ( .A1(n9862), .A2(n5717), .ZN(n9878) );
  INV_X1 U10962 ( .A(n9878), .ZN(n9888) );
  AOI22_X1 U10963 ( .A1(n9858), .A2(n9888), .B1(n9862), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9860) );
  AOI21_X1 U10964 ( .B1(n9861), .B2(n9860), .A(n9859), .ZN(n9865) );
  NOR2_X1 U10965 ( .A1(n9886), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9863) );
  OAI22_X1 U10966 ( .A1(n9864), .A2(n9863), .B1(n9862), .B2(P1_U3084), .ZN(
        n9889) );
  AOI22_X1 U10967 ( .A1(n9866), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(n9865), .B2(
        n9889), .ZN(n9869) );
  NAND3_X1 U10968 ( .A1(n9959), .A2(P1_IR_REG_0__SCAN_IN), .A3(n9867), .ZN(
        n9868) );
  OAI211_X1 U10969 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n6918), .A(n9869), .B(
        n9868), .ZN(P1_U3241) );
  NAND2_X1 U10970 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9872) );
  AOI211_X1 U10971 ( .C1(n9872), .C2(n9871), .A(n9870), .B(n9882), .ZN(n9873)
         );
  AOI21_X1 U10972 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(P1_U3084), .A(n9873), 
        .ZN(n9881) );
  INV_X1 U10973 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9874) );
  OAI22_X1 U10974 ( .A1(n9964), .A2(n9874), .B1(n9943), .B2(n5764), .ZN(n9875)
         );
  INV_X1 U10975 ( .A(n9875), .ZN(n9880) );
  OAI211_X1 U10976 ( .C1(n9878), .C2(n9877), .A(n9960), .B(n9876), .ZN(n9879)
         );
  NAND3_X1 U10977 ( .A1(n9881), .A2(n9880), .A3(n9879), .ZN(P1_U3242) );
  AOI211_X1 U10978 ( .C1(n9885), .C2(n9884), .A(n9883), .B(n9882), .ZN(n9899)
         );
  MUX2_X1 U10979 ( .A(n9888), .B(n9887), .S(n9886), .Z(n9892) );
  OAI211_X1 U10980 ( .C1(n9892), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9914)
         );
  OAI211_X1 U10981 ( .C1(n9895), .C2(n9894), .A(n9960), .B(n9893), .ZN(n9896)
         );
  OAI211_X1 U10982 ( .C1(n9943), .C2(n9897), .A(n9914), .B(n9896), .ZN(n9898)
         );
  AOI211_X1 U10983 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(P1_U3084), .A(n9899), 
        .B(n9898), .ZN(n9900) );
  OAI21_X1 U10984 ( .B1(n9964), .B2(n9901), .A(n9900), .ZN(P1_U3243) );
  OAI21_X1 U10985 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9913) );
  INV_X1 U10986 ( .A(n9905), .ZN(n9912) );
  AOI21_X1 U10987 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(n9910) );
  OAI22_X1 U10988 ( .A1(n9910), .A2(n9935), .B1(n9943), .B2(n9909), .ZN(n9911)
         );
  AOI211_X1 U10989 ( .C1(n9959), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9915)
         );
  OAI211_X1 U10990 ( .C1(n9916), .C2(n9964), .A(n9915), .B(n9914), .ZN(
        P1_U3245) );
  AOI21_X1 U10991 ( .B1(n9951), .B2(n9918), .A(n9917), .ZN(n9924) );
  AOI21_X1 U10992 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(n9922) );
  NAND2_X1 U10993 ( .A1(n9959), .A2(n9922), .ZN(n9923) );
  AND2_X1 U10994 ( .A1(n9924), .A2(n9923), .ZN(n9930) );
  AOI21_X1 U10995 ( .B1(n9927), .B2(n9926), .A(n9925), .ZN(n9928) );
  OR2_X1 U10996 ( .A1(n9935), .A2(n9928), .ZN(n9929) );
  OAI211_X1 U10997 ( .C1(n9931), .C2(n9964), .A(n9930), .B(n9929), .ZN(
        P1_U3246) );
  OAI21_X1 U10998 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9941) );
  AOI211_X1 U10999 ( .C1(n9938), .C2(n9937), .A(n9936), .B(n9935), .ZN(n9939)
         );
  AOI211_X1 U11000 ( .C1(n9959), .C2(n9941), .A(n9940), .B(n9939), .ZN(n9947)
         );
  INV_X1 U11001 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9944) );
  OAI22_X1 U11002 ( .A1(n9964), .A2(n9944), .B1(n9943), .B2(n9942), .ZN(n9945)
         );
  INV_X1 U11003 ( .A(n9945), .ZN(n9946) );
  NAND2_X1 U11004 ( .A1(n9947), .A2(n9946), .ZN(P1_U3250) );
  INV_X1 U11005 ( .A(n9948), .ZN(n9949) );
  AOI21_X1 U11006 ( .B1(n9951), .B2(n9950), .A(n9949), .ZN(n9963) );
  AOI21_X1 U11007 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(n9961) );
  OAI21_X1 U11008 ( .B1(n9957), .B2(n9956), .A(n9955), .ZN(n9958) );
  AOI22_X1 U11009 ( .A1(n9961), .A2(n9960), .B1(n9959), .B2(n9958), .ZN(n9962)
         );
  OAI211_X1 U11010 ( .C1(n9964), .C2(n10157), .A(n9963), .B(n9962), .ZN(
        P1_U3259) );
  AND2_X1 U11011 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9967), .ZN(P1_U3292) );
  AND2_X1 U11012 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9967), .ZN(P1_U3293) );
  AND2_X1 U11013 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9967), .ZN(P1_U3294) );
  AND2_X1 U11014 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9967), .ZN(P1_U3295) );
  AND2_X1 U11015 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9967), .ZN(P1_U3296) );
  AND2_X1 U11016 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9967), .ZN(P1_U3297) );
  AND2_X1 U11017 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9967), .ZN(P1_U3298) );
  AND2_X1 U11018 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9967), .ZN(P1_U3299) );
  AND2_X1 U11019 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9967), .ZN(P1_U3300) );
  AND2_X1 U11020 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9967), .ZN(P1_U3301) );
  AND2_X1 U11021 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9967), .ZN(P1_U3302) );
  AND2_X1 U11022 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9967), .ZN(P1_U3303) );
  AND2_X1 U11023 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9967), .ZN(P1_U3304) );
  AND2_X1 U11024 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9967), .ZN(P1_U3305) );
  AND2_X1 U11025 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9967), .ZN(P1_U3306) );
  AND2_X1 U11026 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9967), .ZN(P1_U3307) );
  AND2_X1 U11027 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9967), .ZN(P1_U3308) );
  AND2_X1 U11028 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9967), .ZN(P1_U3309) );
  AND2_X1 U11029 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9967), .ZN(P1_U3310) );
  AND2_X1 U11030 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9967), .ZN(P1_U3311) );
  AND2_X1 U11031 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9967), .ZN(P1_U3312) );
  AND2_X1 U11032 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9967), .ZN(P1_U3313) );
  AND2_X1 U11033 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9967), .ZN(P1_U3314) );
  AND2_X1 U11034 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9967), .ZN(P1_U3315) );
  AND2_X1 U11035 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9967), .ZN(P1_U3316) );
  AND2_X1 U11036 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9967), .ZN(P1_U3317) );
  AND2_X1 U11037 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9967), .ZN(P1_U3318) );
  AND2_X1 U11038 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9967), .ZN(P1_U3319) );
  AND2_X1 U11039 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9967), .ZN(P1_U3320) );
  AND2_X1 U11040 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9967), .ZN(P1_U3321) );
  OAI21_X1 U11041 ( .B1(n9969), .B2(n9982), .A(n9968), .ZN(n9971) );
  AOI211_X1 U11042 ( .C1(n9973), .C2(n9972), .A(n9971), .B(n9970), .ZN(n9990)
         );
  INV_X1 U11043 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11044 ( .A1(n9989), .A2(n9990), .B1(n9974), .B2(n9988), .ZN(
        P1_U3463) );
  OAI21_X1 U11045 ( .B1(n9976), .B2(n9982), .A(n9975), .ZN(n9978) );
  AOI211_X1 U11046 ( .C1(n9979), .C2(n9986), .A(n9978), .B(n9977), .ZN(n9991)
         );
  INV_X1 U11047 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9980) );
  AOI22_X1 U11048 ( .A1(n9989), .A2(n9991), .B1(n9980), .B2(n9988), .ZN(
        P1_U3469) );
  OAI21_X1 U11049 ( .B1(n9983), .B2(n9982), .A(n9981), .ZN(n9984) );
  AOI211_X1 U11050 ( .C1(n9987), .C2(n9986), .A(n9985), .B(n9984), .ZN(n9993)
         );
  AOI22_X1 U11051 ( .A1(n9989), .A2(n9993), .B1(n5952), .B2(n9988), .ZN(
        P1_U3481) );
  AOI22_X1 U11052 ( .A1(n9994), .A2(n9990), .B1(n5806), .B2(n9992), .ZN(
        P1_U3526) );
  AOI22_X1 U11053 ( .A1(n9994), .A2(n9991), .B1(n5855), .B2(n9992), .ZN(
        P1_U3528) );
  AOI22_X1 U11054 ( .A1(n9994), .A2(n9993), .B1(n5951), .B2(n9992), .ZN(
        P1_U3532) );
  AOI22_X1 U11055 ( .A1(n9997), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9995), .ZN(n10006) );
  NAND2_X1 U11056 ( .A1(n9997), .A2(n9996), .ZN(n9999) );
  OAI211_X1 U11057 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n10000), .A(n9999), .B(
        n9998), .ZN(n10001) );
  INV_X1 U11058 ( .A(n10001), .ZN(n10004) );
  AOI22_X1 U11059 ( .A1(n10002), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10003) );
  OAI221_X1 U11060 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n10006), .C1(n10005), .C2(
        n10004), .A(n10003), .ZN(P2_U3245) );
  AND2_X1 U11061 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10011), .ZN(P2_U3297) );
  AND2_X1 U11062 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10011), .ZN(P2_U3298) );
  AND2_X1 U11063 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10011), .ZN(P2_U3299) );
  AND2_X1 U11064 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10011), .ZN(P2_U3300) );
  AND2_X1 U11065 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10011), .ZN(P2_U3301) );
  AND2_X1 U11066 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10011), .ZN(P2_U3302) );
  AND2_X1 U11067 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10011), .ZN(P2_U3303) );
  AND2_X1 U11068 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10011), .ZN(P2_U3304) );
  AND2_X1 U11069 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10011), .ZN(P2_U3305) );
  AND2_X1 U11070 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10011), .ZN(P2_U3306) );
  AND2_X1 U11071 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10011), .ZN(P2_U3307) );
  AND2_X1 U11072 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10011), .ZN(P2_U3308) );
  AND2_X1 U11073 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10011), .ZN(P2_U3309) );
  AND2_X1 U11074 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10011), .ZN(P2_U3310) );
  AND2_X1 U11075 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10011), .ZN(P2_U3311) );
  AND2_X1 U11076 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10011), .ZN(P2_U3312) );
  AND2_X1 U11077 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10011), .ZN(P2_U3313) );
  AND2_X1 U11078 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10011), .ZN(P2_U3314) );
  AND2_X1 U11079 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10011), .ZN(P2_U3315) );
  AND2_X1 U11080 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10011), .ZN(P2_U3316) );
  AND2_X1 U11081 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10011), .ZN(P2_U3317) );
  AND2_X1 U11082 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10011), .ZN(P2_U3318) );
  AND2_X1 U11083 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10011), .ZN(P2_U3319) );
  AND2_X1 U11084 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10011), .ZN(P2_U3320) );
  AND2_X1 U11085 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10011), .ZN(P2_U3321) );
  AND2_X1 U11086 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10011), .ZN(P2_U3322) );
  AND2_X1 U11087 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10011), .ZN(P2_U3323) );
  AND2_X1 U11088 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10011), .ZN(P2_U3324) );
  AND2_X1 U11089 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10011), .ZN(P2_U3325) );
  AND2_X1 U11090 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10011), .ZN(P2_U3326) );
  AOI22_X1 U11091 ( .A1(n10010), .A2(n10013), .B1(n10009), .B2(n10011), .ZN(
        P2_U3437) );
  AOI22_X1 U11092 ( .A1(n10014), .A2(n10013), .B1(n10012), .B2(n10011), .ZN(
        P2_U3438) );
  OAI22_X1 U11093 ( .A1(n10017), .A2(n10085), .B1(n10016), .B2(n10015), .ZN(
        n10018) );
  NOR2_X1 U11094 ( .A1(n10019), .A2(n10018), .ZN(n10106) );
  AOI22_X1 U11095 ( .A1(n10104), .A2(n10106), .B1(n4958), .B2(n10102), .ZN(
        P2_U3451) );
  INV_X1 U11096 ( .A(n10020), .ZN(n10028) );
  NAND3_X1 U11097 ( .A1(n10022), .A2(n10021), .A3(n10089), .ZN(n10023) );
  OAI21_X1 U11098 ( .B1(n10024), .B2(n10094), .A(n10023), .ZN(n10027) );
  INV_X1 U11099 ( .A(n10025), .ZN(n10026) );
  AOI211_X1 U11100 ( .C1(n10101), .C2(n10028), .A(n10027), .B(n10026), .ZN(
        n10107) );
  AOI22_X1 U11101 ( .A1(n10104), .A2(n10107), .B1(n4968), .B2(n10102), .ZN(
        P2_U3454) );
  INV_X1 U11102 ( .A(n10029), .ZN(n10034) );
  OAI211_X1 U11103 ( .C1(n10032), .C2(n10094), .A(n10031), .B(n10030), .ZN(
        n10033) );
  AOI21_X1 U11104 ( .B1(n10034), .B2(n10101), .A(n10033), .ZN(n10108) );
  AOI22_X1 U11105 ( .A1(n10104), .A2(n10108), .B1(n4936), .B2(n10102), .ZN(
        P2_U3457) );
  NAND2_X1 U11106 ( .A1(n10035), .A2(n10089), .ZN(n10036) );
  OAI21_X1 U11107 ( .B1(n10037), .B2(n10094), .A(n10036), .ZN(n10038) );
  AOI21_X1 U11108 ( .B1(n10039), .B2(n10084), .A(n10038), .ZN(n10040) );
  AND2_X1 U11109 ( .A1(n10041), .A2(n10040), .ZN(n10109) );
  AOI22_X1 U11110 ( .A1(n10104), .A2(n10109), .B1(n4981), .B2(n10102), .ZN(
        P2_U3460) );
  INV_X1 U11111 ( .A(n10042), .ZN(n10048) );
  INV_X1 U11112 ( .A(n10043), .ZN(n10045) );
  OAI22_X1 U11113 ( .A1(n10045), .A2(n10096), .B1(n10044), .B2(n10094), .ZN(
        n10047) );
  AOI211_X1 U11114 ( .C1(n10101), .C2(n10048), .A(n10047), .B(n10046), .ZN(
        n10110) );
  AOI22_X1 U11115 ( .A1(n10104), .A2(n10110), .B1(n4999), .B2(n10102), .ZN(
        P2_U3463) );
  NAND2_X1 U11116 ( .A1(n10049), .A2(n10088), .ZN(n10050) );
  AND2_X1 U11117 ( .A1(n10051), .A2(n10050), .ZN(n10055) );
  NAND3_X1 U11118 ( .A1(n10053), .A2(n10052), .A3(n10101), .ZN(n10054) );
  AND3_X1 U11119 ( .A1(n10056), .A2(n10055), .A3(n10054), .ZN(n10112) );
  AOI22_X1 U11120 ( .A1(n10104), .A2(n10112), .B1(n5036), .B2(n10102), .ZN(
        P2_U3469) );
  INV_X1 U11121 ( .A(n10057), .ZN(n10063) );
  OAI21_X1 U11122 ( .B1(n10059), .B2(n10094), .A(n10058), .ZN(n10062) );
  INV_X1 U11123 ( .A(n10060), .ZN(n10061) );
  AOI211_X1 U11124 ( .C1(n10101), .C2(n10063), .A(n10062), .B(n10061), .ZN(
        n10113) );
  AOI22_X1 U11125 ( .A1(n10104), .A2(n10113), .B1(n5054), .B2(n10102), .ZN(
        P2_U3472) );
  INV_X1 U11126 ( .A(n10064), .ZN(n10065) );
  OAI22_X1 U11127 ( .A1(n10066), .A2(n10096), .B1(n10065), .B2(n10094), .ZN(
        n10068) );
  AOI211_X1 U11128 ( .C1(n10084), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        n10114) );
  INV_X1 U11129 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10070) );
  AOI22_X1 U11130 ( .A1(n10104), .A2(n10114), .B1(n10070), .B2(n10102), .ZN(
        P2_U3475) );
  INV_X1 U11131 ( .A(n10071), .ZN(n10076) );
  OAI22_X1 U11132 ( .A1(n10073), .A2(n10096), .B1(n10072), .B2(n10094), .ZN(
        n10075) );
  AOI211_X1 U11133 ( .C1(n10084), .C2(n10076), .A(n10075), .B(n10074), .ZN(
        n10115) );
  INV_X1 U11134 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U11135 ( .A1(n10104), .A2(n10115), .B1(n10077), .B2(n10102), .ZN(
        P2_U3478) );
  INV_X1 U11136 ( .A(n10078), .ZN(n10083) );
  OAI22_X1 U11137 ( .A1(n10080), .A2(n10096), .B1(n10079), .B2(n10094), .ZN(
        n10082) );
  AOI211_X1 U11138 ( .C1(n10084), .C2(n10083), .A(n10082), .B(n10081), .ZN(
        n10116) );
  AOI22_X1 U11139 ( .A1(n10104), .A2(n10116), .B1(n5126), .B2(n10102), .ZN(
        P2_U3481) );
  OR2_X1 U11140 ( .A1(n10086), .A2(n10085), .ZN(n10093) );
  AOI22_X1 U11141 ( .A1(n10090), .A2(n10089), .B1(n10088), .B2(n10087), .ZN(
        n10091) );
  AOI22_X1 U11142 ( .A1(n10104), .A2(n10117), .B1(n5144), .B2(n10102), .ZN(
        P2_U3484) );
  OAI22_X1 U11143 ( .A1(n10097), .A2(n10096), .B1(n10095), .B2(n10094), .ZN(
        n10099) );
  AOI211_X1 U11144 ( .C1(n10101), .C2(n10100), .A(n10099), .B(n10098), .ZN(
        n10119) );
  INV_X1 U11145 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U11146 ( .A1(n10104), .A2(n10119), .B1(n10103), .B2(n10102), .ZN(
        P2_U3487) );
  AOI22_X1 U11147 ( .A1(n10120), .A2(n10106), .B1(n10105), .B2(n10118), .ZN(
        P2_U3520) );
  AOI22_X1 U11148 ( .A1(n10120), .A2(n10107), .B1(n6808), .B2(n10118), .ZN(
        P2_U3521) );
  AOI22_X1 U11149 ( .A1(n10120), .A2(n10108), .B1(n6811), .B2(n10118), .ZN(
        P2_U3522) );
  AOI22_X1 U11150 ( .A1(n10120), .A2(n10109), .B1(n6812), .B2(n10118), .ZN(
        P2_U3523) );
  AOI22_X1 U11151 ( .A1(n10120), .A2(n10110), .B1(n6814), .B2(n10118), .ZN(
        P2_U3524) );
  INV_X1 U11152 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U11153 ( .A1(n10120), .A2(n10112), .B1(n10111), .B2(n10118), .ZN(
        P2_U3526) );
  AOI22_X1 U11154 ( .A1(n10120), .A2(n10113), .B1(n6819), .B2(n10118), .ZN(
        P2_U3527) );
  AOI22_X1 U11155 ( .A1(n10120), .A2(n10114), .B1(n6820), .B2(n10118), .ZN(
        P2_U3528) );
  AOI22_X1 U11156 ( .A1(n10120), .A2(n10115), .B1(n6822), .B2(n10118), .ZN(
        P2_U3529) );
  AOI22_X1 U11157 ( .A1(n10120), .A2(n10116), .B1(n6824), .B2(n10118), .ZN(
        P2_U3530) );
  AOI22_X1 U11158 ( .A1(n10120), .A2(n10117), .B1(n6807), .B2(n10118), .ZN(
        P2_U3531) );
  AOI22_X1 U11159 ( .A1(n10120), .A2(n10119), .B1(n6984), .B2(n10118), .ZN(
        P2_U3532) );
  INV_X1 U11160 ( .A(n10121), .ZN(n10122) );
  NAND2_X1 U11161 ( .A1(n10123), .A2(n10122), .ZN(n10124) );
  XOR2_X1 U11162 ( .A(n10125), .B(n10124), .Z(ADD_1071_U5) );
  XOR2_X1 U11163 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11164 ( .B1(n10128), .B2(n10127), .A(n10126), .ZN(ADD_1071_U56) );
  OAI21_X1 U11165 ( .B1(n10131), .B2(n10130), .A(n10129), .ZN(ADD_1071_U57) );
  OAI21_X1 U11166 ( .B1(n10134), .B2(n10133), .A(n10132), .ZN(ADD_1071_U58) );
  OAI21_X1 U11167 ( .B1(n10137), .B2(n10136), .A(n10135), .ZN(ADD_1071_U59) );
  OAI21_X1 U11168 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(ADD_1071_U60) );
  OAI21_X1 U11169 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(ADD_1071_U61) );
  AOI21_X1 U11170 ( .B1(n10146), .B2(n10145), .A(n10144), .ZN(ADD_1071_U62) );
  AOI21_X1 U11171 ( .B1(n10149), .B2(n10148), .A(n10147), .ZN(ADD_1071_U63) );
  XNOR2_X1 U11172 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10151) );
  XNOR2_X1 U11173 ( .A(n10151), .B(n10150), .ZN(ADD_1071_U47) );
  XOR2_X1 U11174 ( .A(n10153), .B(n10152), .Z(ADD_1071_U54) );
  XOR2_X1 U11175 ( .A(n10154), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  OAI21_X1 U11176 ( .B1(n10157), .B2(n10156), .A(n10155), .ZN(n10158) );
  XNOR2_X1 U11177 ( .A(n10158), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  XOR2_X1 U11178 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10159), .Z(ADD_1071_U49) );
  XOR2_X1 U11179 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10160), .Z(ADD_1071_U50) );
  AOI21_X1 U11180 ( .B1(n10162), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10161), .ZN(
        n10163) );
  XOR2_X1 U11181 ( .A(n10163), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1071_U51) );
  XOR2_X1 U11182 ( .A(n10165), .B(n10164), .Z(ADD_1071_U53) );
  XNOR2_X1 U11183 ( .A(n10167), .B(n10166), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4819 ( .A(n4933), .Z(n4922) );
  CLKBUF_X3 U4913 ( .A(n5001), .Z(n5480) );
endmodule

