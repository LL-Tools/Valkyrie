

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9709, n9710, n9711, n9712, n9714, n9715, n9716, n9717, n9718, n9720,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9736, n9737, n9738, n9739, n9740, n9742, n9743, n9744,
         n9746, n9747, n9748, n9749, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899;

  INV_X2 U11153 ( .A(n20919), .ZN(n20897) );
  INV_X1 U11154 ( .A(n20520), .ZN(n20490) );
  NOR2_X1 U11155 ( .A1(n20536), .A2(n20396), .ZN(n20449) );
  NOR2_X1 U11156 ( .A1(n20536), .A2(n20752), .ZN(n20668) );
  OR2_X1 U11157 ( .A1(n20751), .A2(n20781), .ZN(n20536) );
  NAND2_X1 U11158 ( .A1(n20751), .A2(n16855), .ZN(n20205) );
  OAI21_X1 U11159 ( .B1(n11719), .B2(n11515), .A(n10391), .ZN(n11516) );
  NAND2_X1 U11160 ( .A1(n13900), .A2(n18706), .ZN(n17723) );
  AND2_X1 U11161 ( .A1(n11526), .A2(n13893), .ZN(n20212) );
  AND2_X1 U11162 ( .A1(n11525), .A2(n13893), .ZN(n20148) );
  AND2_X1 U11163 ( .A1(n9991), .A2(n13893), .ZN(n20174) );
  INV_X1 U11164 ( .A(n13047), .ZN(n13339) );
  BUF_X2 U11165 ( .A(n12366), .Z(n12378) );
  NOR2_X2 U11166 ( .A1(n13711), .A2(n13710), .ZN(n13766) );
  CLKBUF_X2 U11168 ( .A(n12091), .Z(n12283) );
  INV_X1 U11169 ( .A(n12090), .ZN(n12282) );
  INV_X1 U11170 ( .A(n13684), .ZN(n9724) );
  INV_X1 U11171 ( .A(n9723), .ZN(n14490) );
  NAND2_X1 U11172 ( .A1(n13634), .A2(n11224), .ZN(n11311) );
  CLKBUF_X2 U11174 ( .A(n11492), .Z(n11982) );
  CLKBUF_X2 U11175 ( .A(n11224), .Z(n9747) );
  CLKBUF_X2 U11176 ( .A(n10825), .Z(n13320) );
  AND2_X4 U11177 ( .A1(n12073), .A2(n20800), .ZN(n12077) );
  INV_X1 U11178 ( .A(n10740), .ZN(n18450) );
  CLKBUF_X2 U11179 ( .A(n11655), .Z(n12290) );
  INV_X1 U11180 ( .A(n18445), .ZN(n18420) );
  INV_X1 U11181 ( .A(n18301), .ZN(n18451) );
  AND2_X2 U11182 ( .A1(n11536), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11641) );
  BUF_X1 U11183 ( .A(n11457), .Z(n20135) );
  CLKBUF_X2 U11184 ( .A(n10937), .Z(n13269) );
  INV_X1 U11185 ( .A(n12035), .ZN(n10037) );
  CLKBUF_X2 U11186 ( .A(n10925), .Z(n13285) );
  NAND2_X1 U11187 ( .A1(n11457), .A2(n9726), .ZN(n11473) );
  NAND2_X1 U11188 ( .A1(n10553), .A2(n9744), .ZN(n11224) );
  NAND2_X2 U11189 ( .A1(n11415), .A2(n11414), .ZN(n20807) );
  AND2_X1 U11190 ( .A1(n12642), .A2(n11537), .ZN(n11560) );
  INV_X1 U11192 ( .A(n10739), .ZN(n18460) );
  INV_X2 U11193 ( .A(n10739), .ZN(n18269) );
  AND4_X1 U11194 ( .A1(n10841), .A2(n10840), .A3(n10839), .A4(n10838), .ZN(
        n10857) );
  BUF_X2 U11195 ( .A(n10811), .Z(n13291) );
  NOR2_X2 U11196 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16805) );
  AND2_X1 U11197 ( .A1(n10554), .A2(n13977), .ZN(n10741) );
  AND2_X1 U11198 ( .A1(n10754), .A2(n10752), .ZN(n10925) );
  AND2_X1 U11199 ( .A1(n10754), .A2(n10554), .ZN(n10825) );
  INV_X1 U11200 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10880) );
  AND2_X1 U11201 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10752) );
  BUF_X1 U11202 ( .A(n13211), .Z(n13328) );
  CLKBUF_X2 U11203 ( .A(n13321), .Z(n13293) );
  NOR2_X1 U11204 ( .A1(n11929), .A2(n16767), .ZN(n10096) );
  AND3_X1 U11205 ( .A1(n11218), .A2(n14306), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11167) );
  AND2_X1 U11206 ( .A1(n11538), .A2(n12642), .ZN(n11574) );
  NAND2_X1 U11207 ( .A1(n10269), .A2(n10268), .ZN(n9726) );
  INV_X2 U11208 ( .A(n20807), .ZN(n11890) );
  INV_X1 U11209 ( .A(n18419), .ZN(n18443) );
  OAI21_X1 U11210 ( .B1(n10544), .B2(n13014), .A(n12825), .ZN(n14104) );
  NOR2_X1 U11211 ( .A1(n15365), .A2(n15363), .ZN(n15351) );
  BUF_X1 U11213 ( .A(n11009), .Z(n12850) );
  NAND2_X1 U11215 ( .A1(n11784), .A2(n11843), .ZN(n11755) );
  NAND2_X1 U11216 ( .A1(n10032), .A2(n9926), .ZN(n11840) );
  OR2_X1 U11217 ( .A1(n12433), .A2(n12434), .ZN(n16298) );
  AND2_X1 U11218 ( .A1(n11655), .A2(n10271), .ZN(n11461) );
  INV_X1 U11219 ( .A(n18459), .ZN(n18402) );
  NAND2_X1 U11220 ( .A1(n18977), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18976) );
  INV_X1 U11221 ( .A(n17027), .ZN(n18330) );
  INV_X1 U11222 ( .A(n13634), .ZN(n11242) );
  CLKBUF_X2 U11223 ( .A(n10741), .Z(n13995) );
  INV_X1 U11224 ( .A(n12386), .ZN(n11683) );
  INV_X1 U11225 ( .A(n15967), .ZN(n10319) );
  NAND2_X1 U11226 ( .A1(n10269), .A2(n10268), .ZN(n9727) );
  INV_X1 U11227 ( .A(n12073), .ZN(n11456) );
  NAND2_X1 U11228 ( .A1(n14600), .A2(n14601), .ZN(n14598) );
  INV_X1 U11229 ( .A(n18707), .ZN(n19943) );
  AOI21_X1 U11230 ( .B1(n14945), .B2(n14936), .A(n9798), .ZN(n15310) );
  NAND2_X1 U11231 ( .A1(n14368), .A2(n14403), .ZN(n14402) );
  INV_X1 U11232 ( .A(n15969), .ZN(n15981) );
  BUF_X1 U11233 ( .A(n12347), .Z(n15967) );
  NAND2_X1 U11234 ( .A1(n15815), .A2(n9829), .ZN(n15732) );
  CLKBUF_X2 U11235 ( .A(n11455), .Z(n16873) );
  NAND2_X1 U11236 ( .A1(n16239), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16509) );
  OAI21_X1 U11237 ( .B1(n20106), .B2(n20105), .A(n20104), .ZN(n20143) );
  NOR2_X1 U11238 ( .A1(n20536), .A2(n20535), .ZN(n20559) );
  INV_X2 U11239 ( .A(n17742), .ZN(n18098) );
  OR2_X1 U11240 ( .A1(n13724), .A2(n13723), .ZN(n18502) );
  NOR2_X1 U11241 ( .A1(n13683), .A2(n13682), .ZN(n9734) );
  OAI21_X1 U11242 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19937), .A(n17710), 
        .ZN(n19045) );
  AND2_X1 U11243 ( .A1(n12052), .A2(n12453), .ZN(n17615) );
  OR2_X1 U11244 ( .A1(n20556), .A2(n20535), .ZN(n20555) );
  INV_X1 U11245 ( .A(n18484), .ZN(n18498) );
  INV_X1 U11246 ( .A(n18946), .ZN(n18966) );
  OR2_X1 U11248 ( .A1(n10258), .A2(n9865), .ZN(n9709) );
  AND3_X1 U11249 ( .A1(n11554), .A2(n11553), .A3(n10471), .ZN(n9710) );
  AND4_X1 U11250 ( .A1(n10623), .A2(n11547), .A3(n11550), .A4(n11548), .ZN(
        n9711) );
  NAND2_X2 U11251 ( .A1(n10245), .A2(n15233), .ZN(n15174) );
  XOR2_X2 U11252 ( .A(n17135), .B(n17134), .Z(n18983) );
  XNOR2_X2 U11253 ( .A(n12712), .B(n12696), .ZN(n16012) );
  NAND4_X2 U11254 ( .A1(n9711), .A2(n9814), .A3(n9763), .A4(n9710), .ZN(n10703) );
  AND2_X4 U11255 ( .A1(n12783), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11909) );
  INV_X1 U11256 ( .A(n18254), .ZN(n10740) );
  NAND2_X4 U11257 ( .A1(n9820), .A2(n9768), .ZN(n10872) );
  AND4_X2 U11258 ( .A1(n10802), .A2(n10801), .A3(n10800), .A4(n10799), .ZN(
        n9820) );
  NAND2_X4 U11259 ( .A1(n13663), .A2(n17415), .ZN(n18445) );
  INV_X4 U11260 ( .A(n13831), .ZN(n14578) );
  BUF_X2 U11261 ( .A(n10722), .Z(n9712) );
  NOR2_X2 U11262 ( .A1(n17420), .A2(n13659), .ZN(n14479) );
  NAND4_X2 U11263 ( .A1(n10621), .A2(n10630), .A3(n10624), .A4(n10628), .ZN(
        n9968) );
  AND2_X2 U11266 ( .A1(n13391), .A2(n14271), .ZN(n14270) );
  OAI21_X2 U11267 ( .B1(n9950), .B2(n9949), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9937) );
  NOR2_X4 U11268 ( .A1(n10227), .A2(n10228), .ZN(n16239) );
  XNOR2_X2 U11269 ( .A(n10151), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14626) );
  BUF_X2 U11271 ( .A(n19045), .Z(n9716) );
  OAI21_X1 U11272 ( .B1(n10138), .B2(n16745), .A(n11931), .ZN(n11932) );
  NAND2_X2 U11273 ( .A1(n10100), .A2(n10099), .ZN(n12432) );
  OAI21_X1 U11274 ( .B1(n11887), .B2(n10731), .A(n11464), .ZN(n12251) );
  XNOR2_X2 U11275 ( .A(n10214), .B(n12098), .ZN(n11929) );
  NAND2_X1 U11276 ( .A1(n11840), .A2(n9765), .ZN(n14600) );
  NAND2_X1 U11277 ( .A1(n9981), .A2(n10393), .ZN(n16377) );
  AND2_X1 U11278 ( .A1(n14795), .A2(n10698), .ZN(n13304) );
  NOR2_X2 U11279 ( .A1(n14809), .A2(n14810), .ZN(n14795) );
  NAND2_X1 U11280 ( .A1(n14863), .A2(n10691), .ZN(n14809) );
  AND2_X1 U11281 ( .A1(n11117), .A2(n15281), .ZN(n11118) );
  NOR3_X1 U11282 ( .A1(n15678), .A2(n9864), .A3(n10001), .ZN(n15616) );
  AND2_X1 U11283 ( .A1(n12232), .A2(n9886), .ZN(n12435) );
  AND2_X1 U11284 ( .A1(n12540), .A2(n12544), .ZN(n13892) );
  AND2_X1 U11285 ( .A1(n10040), .A2(n10597), .ZN(n9801) );
  INV_X1 U11286 ( .A(n17105), .ZN(n10313) );
  NAND2_X1 U11287 ( .A1(n13609), .A2(n13608), .ZN(n20769) );
  OR2_X1 U11288 ( .A1(n13607), .A2(n13606), .ZN(n13609) );
  NAND2_X1 U11289 ( .A1(n18982), .A2(n17136), .ZN(n18969) );
  INV_X1 U11290 ( .A(n16787), .ZN(n15977) );
  AOI21_X1 U11291 ( .B1(n17068), .B2(n18998), .A(n10045), .ZN(n10044) );
  NAND2_X1 U11292 ( .A1(n9985), .A2(n10357), .ZN(n11508) );
  XNOR2_X1 U11293 ( .A(n11513), .B(n11514), .ZN(n16787) );
  CLKBUF_X2 U11294 ( .A(n18501), .Z(n9725) );
  NAND2_X1 U11295 ( .A1(n11477), .A2(n12044), .ZN(n11486) );
  NOR2_X1 U11296 ( .A1(n13011), .A2(n12934), .ZN(n12950) );
  OR2_X1 U11297 ( .A1(n12977), .A2(n12981), .ZN(n13011) );
  NOR2_X2 U11298 ( .A1(n19377), .A2(n19373), .ZN(n13771) );
  AND2_X2 U11299 ( .A1(n9837), .A2(n10047), .ZN(n12366) );
  NAND2_X1 U11300 ( .A1(n11454), .A2(n11461), .ZN(n11464) );
  AND2_X1 U11301 ( .A1(n11461), .A2(n11456), .ZN(n12024) );
  INV_X2 U11302 ( .A(n10915), .ZN(n10866) );
  NAND4_X1 U11303 ( .A1(n20118), .A2(n12035), .A3(n11455), .A4(n12028), .ZN(
        n11463) );
  INV_X1 U11305 ( .A(n12028), .ZN(n20113) );
  AND4_X2 U11306 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n10864) );
  CLKBUF_X2 U11307 ( .A(n13291), .Z(n13319) );
  CLKBUF_X2 U11308 ( .A(n10919), .Z(n13187) );
  AND2_X1 U11309 ( .A1(n12861), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12870) );
  INV_X8 U11310 ( .A(n9799), .ZN(n9717) );
  INV_X2 U11311 ( .A(n18445), .ZN(n18388) );
  CLKBUF_X2 U11312 ( .A(n10924), .Z(n13133) );
  CLKBUF_X2 U11313 ( .A(n13327), .Z(n13132) );
  CLKBUF_X2 U11314 ( .A(n13326), .Z(n13138) );
  BUF_X2 U11315 ( .A(n10773), .Z(n9754) );
  AND2_X1 U11316 ( .A1(n16789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9737) );
  CLKBUF_X1 U11317 ( .A(n9749), .Z(n9718) );
  AND3_X2 U11319 ( .A1(n10277), .A2(n10276), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11430) );
  CLKBUF_X2 U11320 ( .A(n10755), .Z(n14012) );
  NAND2_X2 U11321 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U11322 ( .B1(n10729), .B2(n12812), .A(n9835), .ZN(n10548) );
  AND2_X1 U11323 ( .A1(n9984), .A2(n9982), .ZN(n10681) );
  NAND2_X1 U11324 ( .A1(n10376), .A2(n10375), .ZN(n10011) );
  OR2_X1 U11325 ( .A1(n16332), .A2(n10442), .ZN(n10526) );
  NAND2_X1 U11326 ( .A1(n10640), .A2(n10639), .ZN(n11129) );
  NAND2_X1 U11327 ( .A1(n10385), .A2(n16377), .ZN(n16655) );
  NOR2_X1 U11328 ( .A1(n16363), .A2(n10293), .ZN(n16345) );
  OAI21_X1 U11329 ( .B1(n16575), .B2(n16748), .A(n10264), .ZN(n10263) );
  AND2_X1 U11330 ( .A1(n15216), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10182) );
  CLKBUF_X1 U11331 ( .A(n15174), .Z(n15175) );
  AND2_X1 U11332 ( .A1(n10132), .A2(n16363), .ZN(n16644) );
  INV_X1 U11333 ( .A(n15174), .ZN(n10640) );
  OAI21_X1 U11334 ( .B1(n16575), .B2(n17594), .A(n10279), .ZN(n10278) );
  NAND2_X1 U11335 ( .A1(n10635), .A2(n12491), .ZN(n16226) );
  XNOR2_X1 U11336 ( .A(n14748), .B(n13347), .ZN(n15166) );
  XNOR2_X1 U11337 ( .A(n9929), .B(n9819), .ZN(n16532) );
  NAND2_X1 U11338 ( .A1(n16692), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10386) );
  NOR2_X1 U11339 ( .A1(n17165), .A2(n10305), .ZN(n17316) );
  NAND2_X1 U11340 ( .A1(n16298), .A2(n10265), .ZN(n16575) );
  NAND2_X1 U11341 ( .A1(n10294), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16363) );
  OAI21_X1 U11342 ( .B1(n16617), .B2(n16472), .A(n10399), .ZN(n10398) );
  NOR2_X1 U11343 ( .A1(n16436), .A2(n16722), .ZN(n16435) );
  NAND2_X1 U11344 ( .A1(n10013), .A2(n10012), .ZN(n15312) );
  NOR2_X2 U11345 ( .A1(n16377), .A2(n9914), .ZN(n16322) );
  AOI211_X1 U11346 ( .C1(n16194), .C2(BUF2_REG_29__SCAN_IN), .A(n16097), .B(
        n16096), .ZN(n16098) );
  INV_X1 U11347 ( .A(n16405), .ZN(n16692) );
  NOR2_X1 U11348 ( .A1(n16536), .A2(n9775), .ZN(n9929) );
  NAND2_X1 U11349 ( .A1(n10101), .A2(n10663), .ZN(n16092) );
  AND2_X1 U11350 ( .A1(n16405), .A2(n16674), .ZN(n16672) );
  OR2_X1 U11351 ( .A1(n16410), .A2(n10168), .ZN(n10163) );
  OR2_X1 U11352 ( .A1(n15351), .A2(n15364), .ZN(n10013) );
  XNOR2_X1 U11353 ( .A(n16416), .B(n16417), .ZN(n16436) );
  NAND2_X1 U11354 ( .A1(n9981), .A2(n10392), .ZN(n16405) );
  OAI21_X1 U11355 ( .B1(n10093), .B2(n10171), .A(n16408), .ZN(n16401) );
  NAND2_X1 U11356 ( .A1(n10150), .A2(n10400), .ZN(n16536) );
  INV_X1 U11357 ( .A(n10093), .ZN(n16410) );
  NAND2_X1 U11358 ( .A1(n10411), .A2(n10229), .ZN(n10228) );
  NAND2_X1 U11359 ( .A1(n10094), .A2(n16390), .ZN(n10093) );
  XNOR2_X1 U11360 ( .A(n12810), .B(n12809), .ZN(n15056) );
  NAND2_X1 U11361 ( .A1(n12807), .A2(n12806), .ZN(n12810) );
  AND2_X1 U11362 ( .A1(n10395), .A2(n10394), .ZN(n10393) );
  AND2_X1 U11363 ( .A1(n17324), .A2(n9853), .ZN(n10303) );
  AND2_X1 U11364 ( .A1(n15612), .A2(n14611), .ZN(n16003) );
  AND2_X1 U11365 ( .A1(n12371), .A2(n12021), .ZN(n16009) );
  AND2_X1 U11366 ( .A1(n16389), .A2(n16391), .ZN(n10367) );
  INV_X2 U11367 ( .A(n14862), .ZN(n14863) );
  NAND2_X1 U11368 ( .A1(n10298), .A2(n17519), .ZN(n17513) );
  OAI211_X1 U11369 ( .C1(n20109), .C2(n20101), .A(n20100), .B(n20619), .ZN(
        n20144) );
  NOR2_X1 U11370 ( .A1(n15616), .A2(n15615), .ZN(n16493) );
  XNOR2_X1 U11371 ( .A(n12384), .B(n12383), .ZN(n15993) );
  OAI211_X1 U11372 ( .C1(n10075), .C2(n10051), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n10050), .ZN(n16389) );
  NAND2_X1 U11373 ( .A1(n9946), .A2(n11935), .ZN(n10515) );
  NOR2_X1 U11374 ( .A1(n10110), .A2(n10109), .ZN(n10108) );
  OAI21_X1 U11375 ( .B1(n16388), .B2(n9709), .A(n10082), .ZN(n10085) );
  OAI21_X1 U11376 ( .B1(n16012), .B2(n10732), .A(n12716), .ZN(n10110) );
  AND2_X1 U11377 ( .A1(n18764), .A2(n17086), .ZN(n10300) );
  AND2_X1 U11378 ( .A1(n11931), .A2(n16743), .ZN(n10702) );
  NAND2_X1 U11379 ( .A1(n10049), .A2(n15918), .ZN(n16388) );
  AOI22_X1 U11380 ( .A1(n16861), .A2(n16860), .B1(n16864), .B2(n20489), .ZN(
        n20389) );
  AND3_X2 U11381 ( .A1(n14121), .A2(n10066), .A3(n10064), .ZN(n14368) );
  AND2_X1 U11382 ( .A1(n16858), .A2(n20748), .ZN(n16861) );
  AND2_X1 U11383 ( .A1(n16418), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10192) );
  AND2_X1 U11384 ( .A1(n10387), .A2(n10075), .ZN(n11931) );
  NAND2_X1 U11385 ( .A1(n11731), .A2(n9813), .ZN(n16418) );
  NAND2_X1 U11386 ( .A1(n10075), .A2(n14606), .ZN(n10193) );
  NAND2_X1 U11387 ( .A1(n12011), .A2(n12010), .ZN(n15678) );
  OR2_X1 U11388 ( .A1(n20394), .A2(n16857), .ZN(n16858) );
  NOR2_X1 U11389 ( .A1(n12678), .A2(n12713), .ZN(n16013) );
  INV_X1 U11390 ( .A(n20449), .ZN(n20432) );
  OR2_X1 U11391 ( .A1(n15279), .A2(n11122), .ZN(n11124) );
  INV_X1 U11392 ( .A(n15748), .ZN(n12232) );
  OAI211_X1 U11393 ( .C1(n13047), .C2(n12876), .A(n12875), .B(n12874), .ZN(
        n14335) );
  NAND2_X1 U11394 ( .A1(n11731), .A2(n11930), .ZN(n10075) );
  OR2_X1 U11395 ( .A1(n17526), .A2(n10451), .ZN(n10450) );
  OR2_X1 U11396 ( .A1(n20804), .A2(n20388), .ZN(n16857) );
  OR2_X1 U11397 ( .A1(n11092), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17520) );
  AND2_X1 U11398 ( .A1(n11730), .A2(n11729), .ZN(n11930) );
  NOR2_X2 U11399 ( .A1(n20536), .A2(n20453), .ZN(n20520) );
  AND4_X1 U11400 ( .A1(n14104), .A2(n12860), .A3(n12859), .A4(n14099), .ZN(
        n14105) );
  NOR2_X2 U11401 ( .A1(n20396), .A2(n20205), .ZN(n20201) );
  NOR2_X2 U11402 ( .A1(n20244), .A2(n20752), .ZN(n20362) );
  AOI21_X1 U11403 ( .B1(n18783), .B2(n18830), .A(n10042), .ZN(n10531) );
  NAND2_X1 U11404 ( .A1(n18901), .A2(n17283), .ZN(n18798) );
  NAND2_X1 U11405 ( .A1(n12858), .A2(n12857), .ZN(n14099) );
  OR2_X1 U11406 ( .A1(n11121), .A2(n15524), .ZN(n15313) );
  OAI21_X1 U11407 ( .B1(n11821), .B2(n10476), .A(n16281), .ZN(n10475) );
  OR2_X1 U11408 ( .A1(n20751), .A2(n16855), .ZN(n20556) );
  NAND2_X1 U11409 ( .A1(n10248), .A2(n10996), .ZN(n10009) );
  NAND2_X1 U11410 ( .A1(n20751), .A2(n20781), .ZN(n20244) );
  NOR2_X2 U11411 ( .A1(n15732), .A2(n15734), .ZN(n12440) );
  NAND2_X1 U11412 ( .A1(n18792), .A2(n18831), .ZN(n18873) );
  OAI21_X2 U11413 ( .B1(n13889), .B2(n13892), .A(n13890), .ZN(n20751) );
  AND2_X1 U11414 ( .A1(n10018), .A2(n10017), .ZN(n11726) );
  NAND2_X1 U11415 ( .A1(n9928), .A2(n11625), .ZN(n9941) );
  NAND2_X1 U11416 ( .A1(n18933), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19171) );
  NOR2_X1 U11417 ( .A1(n10625), .A2(n10622), .ZN(n10621) );
  XNOR2_X1 U11418 ( .A(n11107), .B(n11095), .ZN(n12883) );
  OR2_X1 U11419 ( .A1(n18889), .A2(n19140), .ZN(n18831) );
  AND2_X1 U11420 ( .A1(n10629), .A2(n11528), .ZN(n10628) );
  NOR2_X1 U11421 ( .A1(n18888), .A2(n10541), .ZN(n10540) );
  NAND2_X1 U11422 ( .A1(n17339), .A2(n19210), .ZN(n19204) );
  CLKBUF_X1 U11423 ( .A(n14731), .Z(n15142) );
  CLKBUF_X1 U11424 ( .A(n13373), .Z(n15140) );
  AND2_X1 U11425 ( .A1(n16884), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10622) );
  AND2_X1 U11426 ( .A1(n13865), .A2(n13868), .ZN(n20762) );
  AND2_X1 U11427 ( .A1(n10062), .A2(n18830), .ZN(n18888) );
  NAND2_X1 U11428 ( .A1(n10310), .A2(n10313), .ZN(n18889) );
  AND2_X1 U11429 ( .A1(n10015), .A2(n15977), .ZN(n10020) );
  AOI22_X1 U11430 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11604), .B1(
        n20524), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11550) );
  OR2_X1 U11431 ( .A1(n17222), .A2(n9901), .ZN(n10062) );
  OR2_X1 U11432 ( .A1(n13615), .A2(n13616), .ZN(n13617) );
  INV_X1 U11433 ( .A(n10266), .ZN(n10040) );
  AND2_X1 U11434 ( .A1(n17222), .A2(n10311), .ZN(n10310) );
  NAND2_X1 U11435 ( .A1(n10107), .A2(n10105), .ZN(n12540) );
  NOR2_X2 U11436 ( .A1(n11519), .A2(n15977), .ZN(n16884) );
  INV_X1 U11437 ( .A(n18093), .ZN(n18102) );
  OR2_X1 U11438 ( .A1(n21003), .A2(n13882), .ZN(n17547) );
  NAND2_X2 U11439 ( .A1(n15151), .A2(n13858), .ZN(n15160) );
  NAND2_X1 U11440 ( .A1(n14114), .A2(n9841), .ZN(n10160) );
  NAND2_X1 U11441 ( .A1(n10063), .A2(n18976), .ZN(n17222) );
  OAI21_X1 U11442 ( .B1(n10225), .B2(n10106), .A(n10103), .ZN(n12544) );
  AND2_X1 U11443 ( .A1(n9852), .A2(n11518), .ZN(n16862) );
  AND2_X1 U11444 ( .A1(n10225), .A2(n11523), .ZN(n20524) );
  AND2_X1 U11445 ( .A1(n11526), .A2(n10225), .ZN(n11604) );
  AND2_X1 U11446 ( .A1(n10004), .A2(n9858), .ZN(n11036) );
  AND2_X1 U11447 ( .A1(n11354), .A2(n17468), .ZN(n21003) );
  AND2_X1 U11448 ( .A1(n11354), .A2(n11339), .ZN(n13882) );
  NOR2_X1 U11449 ( .A1(n10528), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10063) );
  NAND2_X1 U11450 ( .A1(n11354), .A2(n13553), .ZN(n15533) );
  AND2_X1 U11451 ( .A1(n10183), .A2(n13550), .ZN(n11354) );
  CLKBUF_X1 U11452 ( .A(n13994), .Z(n21167) );
  NOR2_X1 U11453 ( .A1(n11522), .A2(n10383), .ZN(n11523) );
  AND2_X1 U11454 ( .A1(n12846), .A2(n12845), .ZN(n13616) );
  AND2_X1 U11455 ( .A1(n10007), .A2(n9862), .ZN(n12832) );
  NAND2_X1 U11456 ( .A1(n12522), .A2(n12521), .ZN(n12534) );
  OR2_X1 U11457 ( .A1(n12522), .A2(n12521), .ZN(n12523) );
  NOR2_X2 U11458 ( .A1(n19337), .A2(n19121), .ZN(n19183) );
  AND2_X1 U11459 ( .A1(n13869), .A2(n11521), .ZN(n11525) );
  OAI21_X1 U11460 ( .B1(n13869), .B2(n16839), .A(n12519), .ZN(n12522) );
  NAND2_X1 U11461 ( .A1(n11023), .A2(n11022), .ZN(n12840) );
  OAI21_X1 U11462 ( .B1(n18969), .B2(n18968), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17139) );
  AND2_X1 U11463 ( .A1(n10215), .A2(n10204), .ZN(n11520) );
  NAND2_X1 U11464 ( .A1(n10215), .A2(n9815), .ZN(n10224) );
  AND2_X1 U11465 ( .A1(n13869), .A2(n9815), .ZN(n11526) );
  AND2_X1 U11466 ( .A1(n11522), .A2(n10204), .ZN(n11518) );
  NAND2_X1 U11468 ( .A1(n10241), .A2(n10904), .ZN(n14013) );
  NAND2_X1 U11469 ( .A1(n12529), .A2(n12528), .ZN(n12530) );
  NAND2_X1 U11470 ( .A1(n11508), .A2(n10002), .ZN(n10480) );
  AND2_X1 U11471 ( .A1(n11750), .A2(n11749), .ZN(n15877) );
  AND2_X2 U11472 ( .A1(n11193), .A2(n11192), .ZN(n17503) );
  OAI21_X1 U11473 ( .B1(n18999), .B2(n10046), .A(n10044), .ZN(n18985) );
  NAND2_X1 U11474 ( .A1(n10903), .A2(n10902), .ZN(n10904) );
  NAND2_X1 U11475 ( .A1(n10355), .A2(n10353), .ZN(n10455) );
  AND2_X2 U11476 ( .A1(n9960), .A2(n20026), .ZN(n12255) );
  AND2_X1 U11477 ( .A1(n13785), .A2(n13786), .ZN(n13896) );
  AND2_X1 U11478 ( .A1(n11949), .A2(n11953), .ZN(n10579) );
  INV_X1 U11479 ( .A(n10176), .ZN(n10177) );
  NOR2_X1 U11480 ( .A1(n10606), .A2(n15933), .ZN(n10604) );
  OR2_X1 U11481 ( .A1(n11694), .A2(n10650), .ZN(n11746) );
  NAND2_X1 U11482 ( .A1(n10212), .A2(n11511), .ZN(n11514) );
  NAND2_X1 U11483 ( .A1(n11497), .A2(n11496), .ZN(n11509) );
  AND2_X1 U11484 ( .A1(n10883), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10900) );
  OAI21_X1 U11485 ( .B1(n19026), .B2(n10054), .A(n10057), .ZN(n19018) );
  AND2_X1 U11486 ( .A1(n13779), .A2(n10420), .ZN(n13786) );
  NAND2_X1 U11487 ( .A1(n10080), .A2(n10076), .ZN(n10360) );
  OAI21_X1 U11488 ( .B1(n11651), .B2(n11490), .A(n11491), .ZN(n11510) );
  CLKBUF_X3 U11489 ( .A(n11982), .Z(n12377) );
  NAND2_X1 U11490 ( .A1(n11486), .A2(n10077), .ZN(n10080) );
  AND2_X1 U11491 ( .A1(n19015), .A2(n10058), .ZN(n10057) );
  AND2_X1 U11492 ( .A1(n10918), .A2(n10454), .ZN(n10368) );
  NOR2_X1 U11493 ( .A1(n14102), .A2(n10557), .ZN(n10556) );
  INV_X1 U11494 ( .A(n13876), .ZN(n11233) );
  NAND2_X1 U11495 ( .A1(n11486), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11490) );
  AND2_X1 U11496 ( .A1(n11232), .A2(n11231), .ZN(n13876) );
  AND2_X1 U11497 ( .A1(n10887), .A2(n10878), .ZN(n11200) );
  NAND2_X1 U11498 ( .A1(n9964), .A2(n10014), .ZN(n11492) );
  CLKBUF_X1 U11499 ( .A(n12382), .Z(n12376) );
  AND2_X1 U11500 ( .A1(n10875), .A2(n10874), .ZN(n10887) );
  OR2_X1 U11501 ( .A1(n12382), .A2(n11505), .ZN(n10069) );
  NAND2_X1 U11502 ( .A1(n10558), .A2(n11223), .ZN(n10560) );
  AOI21_X1 U11503 ( .B1(n10056), .B2(n17057), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10055) );
  AOI21_X1 U11504 ( .B1(n12022), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10079), 
        .ZN(n10076) );
  OR2_X1 U11505 ( .A1(n17063), .A2(n18635), .ZN(n17069) );
  NAND2_X1 U11506 ( .A1(n10255), .A2(n10254), .ZN(n11209) );
  OR2_X1 U11507 ( .A1(n11227), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n10558) );
  NAND4_X1 U11508 ( .A1(n12023), .A2(n20810), .A3(n12024), .A4(n11460), .ZN(
        n10014) );
  OAI211_X1 U11509 ( .C1(n17492), .C2(n10866), .A(n10870), .B(n10869), .ZN(
        n10892) );
  NOR2_X1 U11510 ( .A1(n11203), .A2(n10860), .ZN(n10876) );
  NAND2_X1 U11511 ( .A1(n10797), .A2(n10798), .ZN(n10295) );
  NAND2_X2 U11512 ( .A1(n11235), .A2(n11333), .ZN(n13629) );
  NOR2_X1 U11513 ( .A1(n11464), .A2(n11890), .ZN(n10262) );
  NAND2_X1 U11514 ( .A1(n10981), .A2(n10980), .ZN(n11186) );
  NAND2_X1 U11515 ( .A1(n10453), .A2(n10452), .ZN(n10877) );
  AND2_X1 U11516 ( .A1(n14239), .A2(n11328), .ZN(n10870) );
  NAND2_X2 U11517 ( .A1(n10866), .A2(n10994), .ZN(n10868) );
  OR2_X1 U11518 ( .A1(n10943), .A2(n10942), .ZN(n11109) );
  OR2_X1 U11519 ( .A1(n16989), .A2(n16988), .ZN(n17114) );
  AND2_X1 U11520 ( .A1(n18707), .A2(n19355), .ZN(n13788) );
  INV_X1 U11521 ( .A(n14481), .ZN(n19369) );
  NAND2_X1 U11522 ( .A1(n10271), .A2(n9727), .ZN(n11466) );
  AND2_X1 U11523 ( .A1(n16873), .A2(n10037), .ZN(n11458) );
  NOR2_X2 U11524 ( .A1(n12331), .A2(n16346), .ZN(n12334) );
  AND2_X2 U11525 ( .A1(n11890), .A2(n11456), .ZN(n11465) );
  BUF_X2 U11526 ( .A(n11456), .Z(n16029) );
  NOR2_X1 U11527 ( .A1(n17733), .A2(n18767), .ZN(n17213) );
  CLKBUF_X1 U11528 ( .A(n10864), .Z(n14157) );
  AND3_X1 U11529 ( .A1(n20113), .A2(n16873), .A3(n11890), .ZN(n10038) );
  INV_X1 U11530 ( .A(n12819), .ZN(n10858) );
  INV_X1 U11531 ( .A(n20118), .ZN(n11470) );
  OR2_X1 U11532 ( .A1(n16969), .A2(n16968), .ZN(n17124) );
  NAND2_X1 U11533 ( .A1(n10864), .A2(n10867), .ZN(n10888) );
  CLKBUF_X1 U11534 ( .A(n10915), .Z(n14306) );
  INV_X1 U11535 ( .A(n10994), .ZN(n11152) );
  INV_X1 U11536 ( .A(n9726), .ZN(n11655) );
  INV_X1 U11537 ( .A(n11457), .ZN(n10271) );
  NOR2_X2 U11538 ( .A1(n13695), .A2(n13694), .ZN(n19365) );
  OR2_X1 U11539 ( .A1(n13739), .A2(n13738), .ZN(n14481) );
  OR2_X1 U11540 ( .A1(n11580), .A2(n11579), .ZN(n12080) );
  INV_X1 U11541 ( .A(n11455), .ZN(n12069) );
  NOR2_X1 U11542 ( .A1(n17655), .A2(n17618), .ZN(n17656) );
  NAND2_X1 U11543 ( .A1(n12819), .A2(n10994), .ZN(n10889) );
  OR2_X1 U11544 ( .A1(n11590), .A2(n11589), .ZN(n11653) );
  NAND2_X1 U11545 ( .A1(n11403), .A2(n11402), .ZN(n12073) );
  INV_X1 U11546 ( .A(n9727), .ZN(n9720) );
  OR3_X1 U11547 ( .A1(n13702), .A2(n13701), .A3(n13700), .ZN(n13711) );
  NAND2_X1 U11548 ( .A1(n10785), .A2(n10784), .ZN(n10865) );
  NAND2_X1 U11549 ( .A1(n10751), .A2(n9757), .ZN(n10915) );
  INV_X2 U11550 ( .A(U214), .ZN(n17655) );
  AND4_X1 U11551 ( .A1(n10777), .A2(n10776), .A3(n10775), .A4(n10774), .ZN(
        n10785) );
  AND4_X1 U11552 ( .A1(n10845), .A2(n10844), .A3(n10843), .A4(n10842), .ZN(
        n10856) );
  AND4_X1 U11553 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10794) );
  AND4_X1 U11554 ( .A1(n10783), .A2(n10782), .A3(n10781), .A4(n10780), .ZN(
        n10784) );
  AND4_X1 U11555 ( .A1(n10833), .A2(n10832), .A3(n10831), .A4(n10830), .ZN(
        n10834) );
  AND4_X1 U11556 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10772) );
  AND4_X1 U11557 ( .A1(n10849), .A2(n10848), .A3(n10847), .A4(n10846), .ZN(
        n10855) );
  AND4_X1 U11558 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10795) );
  AND4_X1 U11559 ( .A1(n10853), .A2(n10852), .A3(n10851), .A4(n10850), .ZN(
        n10854) );
  AND4_X1 U11560 ( .A1(n10819), .A2(n10818), .A3(n10817), .A4(n10816), .ZN(
        n10837) );
  AND4_X1 U11561 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10751) );
  AND2_X1 U11562 ( .A1(n11386), .A2(n11387), .ZN(n9951) );
  AND4_X1 U11563 ( .A1(n10829), .A2(n10828), .A3(n10827), .A4(n10826), .ZN(
        n10835) );
  AND2_X1 U11564 ( .A1(n10779), .A2(n10778), .ZN(n10781) );
  AND4_X1 U11565 ( .A1(n10824), .A2(n10823), .A3(n10822), .A4(n10821), .ZN(
        n10836) );
  AND4_X1 U11566 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10771) );
  INV_X2 U11567 ( .A(n17693), .ZN(U215) );
  AND3_X1 U11568 ( .A1(n10135), .A2(n10134), .A3(n11535), .ZN(n11436) );
  AND3_X1 U11569 ( .A1(n11440), .A2(n11439), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11441) );
  NAND2_X2 U11570 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n20788), .ZN(n20734) );
  NAND2_X2 U11571 ( .A1(n20788), .A2(n21751), .ZN(n20733) );
  BUF_X4 U11572 ( .A(n11529), .Z(n12783) );
  AND3_X1 U11573 ( .A1(n10705), .A2(n10704), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11389) );
  AND2_X1 U11574 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12851), .ZN(
        n12861) );
  INV_X4 U11575 ( .A(n18273), .ZN(n9723) );
  NAND2_X1 U11576 ( .A1(n13663), .A2(n13666), .ZN(n10722) );
  AND2_X2 U11577 ( .A1(n16789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11529) );
  NAND2_X2 U11578 ( .A1(n13664), .A2(n13654), .ZN(n10739) );
  CLKBUF_X1 U11579 ( .A(n11430), .Z(n12666) );
  AND2_X2 U11580 ( .A1(n10753), .A2(n10756), .ZN(n13321) );
  AND2_X2 U11581 ( .A1(n10754), .A2(n10756), .ZN(n13327) );
  AND2_X1 U11582 ( .A1(n17398), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13664) );
  AND2_X2 U11583 ( .A1(n10757), .A2(n10755), .ZN(n10773) );
  AND2_X1 U11584 ( .A1(n10744), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10754) );
  AND2_X1 U11585 ( .A1(n17414), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13666) );
  AND2_X1 U11586 ( .A1(n10449), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10753) );
  AND2_X1 U11587 ( .A1(n10745), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10554) );
  INV_X1 U11588 ( .A(n17420), .ZN(n13910) );
  NOR2_X1 U11589 ( .A1(n12852), .A2(n14264), .ZN(n12851) );
  AND2_X1 U11590 ( .A1(n11537), .A2(n11651), .ZN(n12784) );
  AND2_X1 U11591 ( .A1(n11537), .A2(n11651), .ZN(n9739) );
  NOR2_X1 U11592 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13655) );
  INV_X1 U11593 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11377) );
  INV_X1 U11594 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14264) );
  AND2_X1 U11595 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13660) );
  AND2_X2 U11596 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17415) );
  INV_X2 U11597 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20825) );
  INV_X1 U11598 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10745) );
  NOR2_X2 U11599 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10757) );
  XNOR2_X2 U11600 ( .A(n14682), .B(n12287), .ZN(n12509) );
  NOR4_X1 U11601 ( .A1(n19943), .A2(n19355), .A3(n16952), .A4(n19830), .ZN(
        n18501) );
  AOI22_X1 U11602 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10791) );
  NOR2_X1 U11603 ( .A1(n17105), .A2(n19163), .ZN(n18931) );
  NAND2_X2 U11604 ( .A1(n10529), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n17105) );
  AND2_X2 U11605 ( .A1(n10756), .A2(n14012), .ZN(n9748) );
  AND2_X2 U11610 ( .A1(n13663), .A2(n17403), .ZN(n13684) );
  AND2_X4 U11611 ( .A1(n17414), .A2(n10418), .ZN(n17403) );
  NAND2_X1 U11612 ( .A1(n10129), .A2(n16451), .ZN(n9981) );
  NAND2_X1 U11613 ( .A1(n16451), .A2(n11932), .ZN(n16416) );
  AND2_X1 U11614 ( .A1(n11537), .A2(n11651), .ZN(n9728) );
  AND2_X1 U11615 ( .A1(n11537), .A2(n11651), .ZN(n9729) );
  AND2_X2 U11616 ( .A1(n11651), .A2(n16788), .ZN(n9731) );
  AND2_X2 U11617 ( .A1(n11470), .A2(n12028), .ZN(n11892) );
  AND2_X1 U11618 ( .A1(n11651), .A2(n16788), .ZN(n9730) );
  AND2_X2 U11619 ( .A1(n11651), .A2(n16788), .ZN(n12639) );
  AND2_X1 U11620 ( .A1(n11651), .A2(n16788), .ZN(n9732) );
  AND2_X1 U11621 ( .A1(n16789), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9736) );
  NOR2_X1 U11622 ( .A1(n13683), .A2(n13682), .ZN(n9733) );
  NOR2_X2 U11623 ( .A1(n13683), .A2(n13682), .ZN(n19383) );
  AND2_X4 U11624 ( .A1(n12073), .A2(n20807), .ZN(n12386) );
  NOR4_X2 U11625 ( .A1(n19820), .A2(n19936), .A3(n19819), .A4(n19818), .ZN(
        n19831) );
  AND2_X1 U11626 ( .A1(n13663), .A2(n17403), .ZN(n9738) );
  AND2_X1 U11627 ( .A1(n10757), .A2(n10755), .ZN(n9740) );
  AOI211_X1 U11628 ( .C1(n19232), .C2(n17329), .A(n17328), .B(n17327), .ZN(
        n17335) );
  NOR2_X4 U11629 ( .A1(n15015), .A2(n14959), .ZN(n14960) );
  AOI21_X2 U11631 ( .B1(n16500), .B2(n16509), .A(n16240), .ZN(n16506) );
  AOI211_X2 U11632 ( .C1(n19288), .C2(n19074), .A(n19290), .B(n19073), .ZN(
        n19077) );
  AND2_X1 U11633 ( .A1(n11537), .A2(n11651), .ZN(n9742) );
  AND2_X1 U11634 ( .A1(n11537), .A2(n11651), .ZN(n9743) );
  INV_X1 U11635 ( .A(n10864), .ZN(n9744) );
  INV_X4 U11636 ( .A(n10864), .ZN(n11217) );
  BUF_X2 U11638 ( .A(n12826), .Z(n9746) );
  XNOR2_X1 U11639 ( .A(n10459), .B(n11036), .ZN(n12826) );
  AND2_X1 U11640 ( .A1(n10756), .A2(n14012), .ZN(n9749) );
  AND2_X1 U11641 ( .A1(n10756), .A2(n14012), .ZN(n10954) );
  NAND2_X2 U11642 ( .A1(n12804), .A2(n13634), .ZN(n11227) );
  AOI21_X1 U11643 ( .B1(n16589), .B2(n17606), .A(n16588), .ZN(n16590) );
  INV_X1 U11644 ( .A(n20822), .ZN(n13550) );
  INV_X1 U11645 ( .A(n11010), .ZN(n10158) );
  INV_X1 U11646 ( .A(n9941), .ZN(n10408) );
  NAND2_X1 U11647 ( .A1(n10040), .A2(n9833), .ZN(n10623) );
  INV_X1 U11648 ( .A(n11472), .ZN(n12023) );
  AND2_X1 U11649 ( .A1(n12520), .A2(n16887), .ZN(n13939) );
  AND2_X1 U11650 ( .A1(n11939), .A2(n11932), .ZN(n10129) );
  NAND2_X1 U11651 ( .A1(n16418), .A2(n16701), .ZN(n11935) );
  NAND2_X1 U11652 ( .A1(n10193), .A2(n16418), .ZN(n11934) );
  NAND2_X1 U11653 ( .A1(n11513), .A2(n11514), .ZN(n9985) );
  AND2_X1 U11654 ( .A1(n20135), .A2(n16873), .ZN(n9970) );
  NAND2_X1 U11655 ( .A1(n18985), .A2(n17072), .ZN(n17076) );
  OAI211_X1 U11656 ( .C1(n17503), .C2(n11208), .A(n10186), .B(n9846), .ZN(
        n10183) );
  OR2_X1 U11657 ( .A1(n15665), .A2(n15613), .ZN(n10001) );
  NAND2_X1 U11658 ( .A1(n10479), .A2(n9773), .ZN(n10635) );
  NAND2_X1 U11659 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10347) );
  NAND2_X1 U11660 ( .A1(n11035), .A2(n11036), .ZN(n11010) );
  NOR2_X1 U11661 ( .A1(n10402), .A2(n9760), .ZN(n10034) );
  NAND2_X1 U11662 ( .A1(n10406), .A2(n10405), .ZN(n10409) );
  NAND2_X1 U11663 ( .A1(n11930), .A2(n14606), .ZN(n10405) );
  NOR2_X1 U11664 ( .A1(n10288), .A2(n10285), .ZN(n10630) );
  NAND2_X1 U11665 ( .A1(n10287), .A2(n10286), .ZN(n10285) );
  NAND2_X1 U11666 ( .A1(n20148), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10286) );
  INV_X2 U11667 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11651) );
  INV_X1 U11668 ( .A(n11463), .ZN(n11454) );
  NAND2_X1 U11669 ( .A1(n13788), .A2(n17708), .ZN(n13900) );
  NAND2_X1 U11670 ( .A1(n11067), .A2(n11066), .ZN(n10379) );
  NAND2_X1 U11671 ( .A1(n10221), .A2(n10220), .ZN(n11113) );
  AND3_X1 U11672 ( .A1(n10969), .A2(n10968), .A3(n10967), .ZN(n10973) );
  OR2_X1 U11673 ( .A1(n16774), .A2(n12029), .ZN(n16802) );
  NAND2_X1 U11674 ( .A1(n10122), .A2(n11768), .ZN(n10121) );
  INV_X1 U11675 ( .A(n10653), .ZN(n10122) );
  OR2_X1 U11676 ( .A1(n10656), .A2(n11777), .ZN(n10655) );
  AND2_X1 U11677 ( .A1(n14040), .A2(n11736), .ZN(n10658) );
  NOR2_X1 U11678 ( .A1(n11674), .A2(n10117), .ZN(n10116) );
  AND2_X1 U11679 ( .A1(n12503), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10591) );
  NOR2_X1 U11680 ( .A1(n12073), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12072) );
  NOR2_X1 U11681 ( .A1(n14703), .A2(n10620), .ZN(n10619) );
  INV_X1 U11682 ( .A(n14356), .ZN(n10620) );
  INV_X1 U11683 ( .A(n16280), .ZN(n10476) );
  INV_X1 U11684 ( .A(n10437), .ZN(n10258) );
  NOR2_X1 U11685 ( .A1(n10258), .A2(n9767), .ZN(n10083) );
  INV_X1 U11686 ( .A(n10435), .ZN(n10084) );
  AOI21_X1 U11687 ( .B1(n10437), .B2(n10441), .A(n10436), .ZN(n10435) );
  INV_X1 U11688 ( .A(n16352), .ZN(n10436) );
  NOR2_X1 U11689 ( .A1(n16205), .A2(n14318), .ZN(n10733) );
  NAND2_X1 U11690 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U11691 ( .A1(n12072), .A2(n9726), .ZN(n12220) );
  INV_X1 U11692 ( .A(n11521), .ZN(n10383) );
  NAND2_X1 U11693 ( .A1(n10040), .A2(n15977), .ZN(n10022) );
  NAND2_X1 U11694 ( .A1(n11453), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U11695 ( .A1(n10273), .A2(n11535), .ZN(n10272) );
  AND2_X2 U11696 ( .A1(n13915), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13663) );
  AND2_X2 U11697 ( .A1(n10426), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13654) );
  INV_X1 U11698 ( .A(n10421), .ZN(n10420) );
  OAI21_X1 U11699 ( .B1(n13780), .B2(n19365), .A(n13795), .ZN(n10421) );
  INV_X1 U11700 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10418) );
  INV_X1 U11701 ( .A(n21572), .ZN(n14240) );
  NAND2_X1 U11702 ( .A1(n13354), .A2(n13353), .ZN(n13992) );
  INV_X1 U11703 ( .A(n13932), .ZN(n13346) );
  NOR2_X1 U11704 ( .A1(n9828), .A2(n10699), .ZN(n10698) );
  INV_X1 U11705 ( .A(n14796), .ZN(n10699) );
  NAND2_X1 U11706 ( .A1(n10461), .A2(n10462), .ZN(n12801) );
  NAND2_X1 U11707 ( .A1(n11129), .A2(n10637), .ZN(n10461) );
  NAND2_X1 U11708 ( .A1(n12802), .A2(n10735), .ZN(n10252) );
  NAND2_X1 U11709 ( .A1(n9766), .A2(n15190), .ZN(n12802) );
  AND2_X1 U11710 ( .A1(n11356), .A2(n11355), .ZN(n14464) );
  INV_X1 U11711 ( .A(n16803), .ZN(n16895) );
  OR2_X1 U11712 ( .A1(n11793), .A2(n10655), .ZN(n11780) );
  NAND2_X1 U11713 ( .A1(n12419), .A2(n16341), .ZN(n14696) );
  NAND2_X1 U11714 ( .A1(n16226), .A2(n16225), .ZN(n16216) );
  INV_X1 U11715 ( .A(n15676), .ZN(n12010) );
  INV_X1 U11716 ( .A(n15675), .ZN(n12011) );
  OR3_X1 U11717 ( .A1(n11852), .A2(n14606), .A3(n16514), .ZN(n16252) );
  NOR2_X1 U11718 ( .A1(n10474), .A2(n10403), .ZN(n10402) );
  INV_X1 U11719 ( .A(n16273), .ZN(n10403) );
  INV_X1 U11720 ( .A(n10081), .ZN(n11752) );
  OAI21_X1 U11721 ( .B1(n16388), .B2(n9865), .A(n9767), .ZN(n10081) );
  INV_X1 U11722 ( .A(n10228), .ZN(n10100) );
  AND2_X1 U11723 ( .A1(n10393), .A2(n9918), .ZN(n10139) );
  INV_X1 U11724 ( .A(n16377), .ZN(n10294) );
  NAND2_X1 U11725 ( .A1(n11753), .A2(n11752), .ZN(n12415) );
  NAND2_X1 U11726 ( .A1(n11934), .A2(n16722), .ZN(n9946) );
  NOR2_X1 U11727 ( .A1(n10516), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n9975) );
  INV_X1 U11728 ( .A(n9975), .ZN(n9973) );
  NOR2_X1 U11729 ( .A1(n12539), .A2(n10106), .ZN(n10105) );
  NAND2_X1 U11730 ( .A1(n11875), .A2(n11874), .ZN(n16894) );
  OR2_X1 U11731 ( .A1(n11902), .A2(n20033), .ZN(n11874) );
  AND3_X2 U11732 ( .A1(n13893), .A2(n15977), .A3(n11518), .ZN(n20103) );
  INV_X1 U11733 ( .A(n20494), .ZN(n20619) );
  INV_X2 U11734 ( .A(n13703), .ZN(n17027) );
  NOR2_X1 U11735 ( .A1(n18509), .A2(n19355), .ZN(n10231) );
  INV_X1 U11736 ( .A(n13791), .ZN(n10232) );
  INV_X1 U11737 ( .A(n18891), .ZN(n17100) );
  NAND2_X1 U11738 ( .A1(n17034), .A2(n17116), .ZN(n17333) );
  OAI21_X1 U11739 ( .B1(n15173), .B2(n15370), .A(n15172), .ZN(n10550) );
  INV_X1 U11740 ( .A(n15370), .ZN(n17530) );
  AND2_X1 U11741 ( .A1(n15447), .A2(n11368), .ZN(n15427) );
  OR2_X1 U11742 ( .A1(n20791), .A2(n17509), .ZN(n12262) );
  NAND2_X1 U11743 ( .A1(n14684), .A2(n15969), .ZN(n14692) );
  NAND2_X1 U11744 ( .A1(n16689), .A2(n16454), .ZN(n10207) );
  OR2_X1 U11745 ( .A1(n16494), .A2(n16763), .ZN(n10583) );
  INV_X1 U11746 ( .A(n16492), .ZN(n10584) );
  INV_X1 U11747 ( .A(n14705), .ZN(n10683) );
  INV_X1 U11748 ( .A(n17608), .ZN(n16763) );
  NAND2_X1 U11749 ( .A1(n17194), .A2(n17336), .ZN(n17332) );
  OR2_X2 U11750 ( .A1(n17091), .A2(n17355), .ZN(n17350) );
  NOR2_X1 U11751 ( .A1(n9780), .A2(n9987), .ZN(n11613) );
  NAND2_X1 U11752 ( .A1(n20174), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n9990) );
  INV_X1 U11753 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10449) );
  INV_X1 U11754 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n9957) );
  NAND2_X1 U11755 ( .A1(n20174), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U11756 ( .A1(n11466), .A2(n10037), .ZN(n11888) );
  NAND2_X1 U11757 ( .A1(n10256), .A2(n11209), .ZN(n10253) );
  NAND2_X1 U11758 ( .A1(n10866), .A2(n12819), .ZN(n10862) );
  NAND2_X1 U11759 ( .A1(n10158), .A2(n10157), .ZN(n11087) );
  INV_X1 U11760 ( .A(n10160), .ZN(n10157) );
  OR2_X1 U11761 ( .A1(n11084), .A2(n11083), .ZN(n11097) );
  OR2_X1 U11762 ( .A1(n11006), .A2(n11005), .ZN(n11013) );
  NAND2_X1 U11763 ( .A1(n10858), .A2(n11152), .ZN(n10859) );
  NAND2_X1 U11764 ( .A1(n10868), .A2(n14290), .ZN(n10798) );
  AOI21_X1 U11765 ( .B1(n11144), .B2(n11143), .A(n11136), .ZN(n11142) );
  INV_X1 U11766 ( .A(n11171), .ZN(n10200) );
  INV_X1 U11767 ( .A(n11172), .ZN(n10199) );
  AND2_X1 U11768 ( .A1(n11169), .A2(n11173), .ZN(n10201) );
  INV_X1 U11769 ( .A(n11163), .ZN(n11155) );
  OAI21_X1 U11770 ( .B1(n20178), .B2(n11722), .A(n10390), .ZN(n11723) );
  NAND2_X1 U11771 ( .A1(n9938), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11772 ( .A1(n11897), .A2(n9940), .ZN(n9939) );
  NOR2_X1 U11773 ( .A1(n11461), .A2(n10202), .ZN(n11896) );
  INV_X1 U11774 ( .A(n11473), .ZN(n10202) );
  NAND2_X1 U11775 ( .A1(n11459), .A2(n11458), .ZN(n11472) );
  AND2_X1 U11776 ( .A1(n11332), .A2(n11331), .ZN(n11345) );
  NAND2_X1 U11777 ( .A1(n14770), .A2(n10701), .ZN(n10700) );
  INV_X1 U11778 ( .A(n14784), .ZN(n10701) );
  AND2_X1 U11779 ( .A1(n10694), .A2(n10695), .ZN(n10693) );
  INV_X1 U11780 ( .A(n14834), .ZN(n10694) );
  AND2_X1 U11781 ( .A1(n9774), .A2(n13089), .ZN(n10282) );
  INV_X1 U11782 ( .A(n14876), .ZN(n13089) );
  INV_X1 U11783 ( .A(n13300), .ZN(n13342) );
  NOR2_X1 U11784 ( .A1(n15586), .A2(n20825), .ZN(n13300) );
  NAND2_X1 U11785 ( .A1(n9812), .A2(n10690), .ZN(n10689) );
  INV_X1 U11786 ( .A(n14362), .ZN(n10066) );
  NAND2_X1 U11787 ( .A1(n10877), .A2(n10867), .ZN(n11206) );
  NAND2_X1 U11788 ( .A1(n15234), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10245) );
  NAND2_X1 U11789 ( .A1(n10643), .A2(n10642), .ZN(n10641) );
  NAND2_X1 U11790 ( .A1(n11126), .A2(n15262), .ZN(n10447) );
  NOR2_X1 U11791 ( .A1(n14894), .A2(n14906), .ZN(n10571) );
  NAND2_X1 U11792 ( .A1(n11252), .A2(n10564), .ZN(n10563) );
  INV_X1 U11793 ( .A(n14364), .ZN(n10564) );
  OR2_X1 U11794 ( .A1(n10991), .A2(n10990), .ZN(n10995) );
  NAND2_X1 U11795 ( .A1(n13628), .A2(n13634), .ZN(n10559) );
  XNOR2_X1 U11796 ( .A(n10005), .B(n10973), .ZN(n12831) );
  NAND2_X1 U11797 ( .A1(n10006), .A2(n10952), .ZN(n10005) );
  NAND3_X1 U11798 ( .A1(n10455), .A2(n10314), .A3(n20825), .ZN(n10006) );
  INV_X1 U11799 ( .A(n11206), .ZN(n11199) );
  INV_X1 U11800 ( .A(n14114), .ZN(n14115) );
  INV_X1 U11801 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21166) );
  OR2_X1 U11802 ( .A1(n21291), .A2(n21290), .ZN(n21330) );
  NAND2_X1 U11803 ( .A1(n20825), .A2(n14276), .ZN(n14414) );
  NOR2_X1 U11804 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21008), .ZN(
        n11141) );
  INV_X1 U11805 ( .A(n11167), .ZN(n11180) );
  OR2_X1 U11806 ( .A1(n11544), .A2(n11543), .ZN(n10126) );
  NOR2_X1 U11807 ( .A1(n11831), .A2(n11830), .ZN(n11832) );
  AND2_X1 U11808 ( .A1(n11763), .A2(n10649), .ZN(n10648) );
  NOR2_X1 U11809 ( .A1(n10338), .A2(n16395), .ZN(n10337) );
  INV_X1 U11810 ( .A(n16404), .ZN(n10338) );
  NAND2_X1 U11811 ( .A1(n10035), .A2(n11709), .ZN(n10650) );
  INV_X1 U11812 ( .A(n10651), .ZN(n10035) );
  INV_X1 U11813 ( .A(n11679), .ZN(n11663) );
  NAND2_X1 U11814 ( .A1(n11396), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11403) );
  INV_X1 U11815 ( .A(n12735), .ZN(n10109) );
  OR2_X1 U11816 ( .A1(n10679), .A2(n10678), .ZN(n10677) );
  INV_X1 U11817 ( .A(n16047), .ZN(n10678) );
  NAND2_X1 U11818 ( .A1(n10680), .A2(n16053), .ZN(n10679) );
  INV_X1 U11819 ( .A(n16058), .ZN(n10680) );
  NAND2_X1 U11820 ( .A1(n13938), .A2(n9876), .ZN(n16061) );
  AND2_X1 U11821 ( .A1(n15646), .A2(n12020), .ZN(n10586) );
  NOR2_X1 U11822 ( .A1(n16283), .A2(n10596), .ZN(n10595) );
  NAND2_X1 U11823 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10590) );
  INV_X1 U11824 ( .A(n11653), .ZN(n12087) );
  AOI21_X1 U11825 ( .B1(n11574), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n10030), .ZN(n11561) );
  AND2_X1 U11826 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10030) );
  NOR3_X1 U11827 ( .A1(n9771), .A2(n9824), .A3(n10025), .ZN(n10024) );
  NOR3_X1 U11828 ( .A1(n11635), .A2(n10028), .A3(n10027), .ZN(n10026) );
  NAND2_X1 U11829 ( .A1(n15651), .A2(n10382), .ZN(n11850) );
  INV_X1 U11830 ( .A(n12438), .ZN(n10601) );
  NOR2_X1 U11831 ( .A1(n12441), .A2(n15708), .ZN(n10574) );
  NOR2_X1 U11832 ( .A1(n15736), .A2(n14606), .ZN(n11819) );
  INV_X1 U11833 ( .A(n12466), .ZN(n10618) );
  NOR2_X1 U11834 ( .A1(n10396), .A2(n10209), .ZN(n10394) );
  AND3_X1 U11835 ( .A1(n12126), .A2(n12125), .A3(n12124), .ZN(n14048) );
  INV_X1 U11836 ( .A(n15918), .ZN(n10051) );
  INV_X1 U11837 ( .A(n10409), .ZN(n10048) );
  NAND2_X1 U11838 ( .A1(n11929), .A2(n16767), .ZN(n10213) );
  NAND2_X1 U11839 ( .A1(n10119), .A2(n10118), .ZN(n11674) );
  NAND2_X1 U11840 ( .A1(n11669), .A2(n20127), .ZN(n10119) );
  INV_X1 U11841 ( .A(n11516), .ZN(n10624) );
  AND2_X1 U11842 ( .A1(n13939), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12539) );
  AND2_X1 U11843 ( .A1(n13939), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12521) );
  NAND2_X1 U11844 ( .A1(n9953), .A2(n9952), .ZN(n11875) );
  NAND2_X1 U11845 ( .A1(n20808), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n9952) );
  NAND2_X1 U11846 ( .A1(n9954), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U11847 ( .A1(n11872), .A2(n9955), .ZN(n9954) );
  AND2_X1 U11848 ( .A1(n10036), .A2(n11470), .ZN(n11475) );
  NOR2_X1 U11849 ( .A1(n11473), .A2(n10037), .ZN(n10036) );
  AND2_X1 U11850 ( .A1(n20246), .A2(n20749), .ZN(n20175) );
  NAND2_X2 U11851 ( .A1(n9931), .A2(n9930), .ZN(n12028) );
  NAND2_X1 U11852 ( .A1(n17076), .A2(n17075), .ZN(n17077) );
  NOR2_X1 U11853 ( .A1(n10872), .A2(n21578), .ZN(n12842) );
  NOR2_X2 U11854 ( .A1(n13345), .A2(n14749), .ZN(n14748) );
  NAND2_X1 U11855 ( .A1(n13223), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13259) );
  NAND2_X1 U11856 ( .A1(n13181), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13221) );
  NAND2_X1 U11857 ( .A1(n13092), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13126) );
  NAND2_X1 U11858 ( .A1(n12926), .A2(n12925), .ZN(n12932) );
  AND2_X1 U11859 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12925) );
  AND4_X1 U11860 ( .A1(n12898), .A2(n12897), .A3(n12896), .A4(n12895), .ZN(
        n14367) );
  NAND2_X1 U11861 ( .A1(n10009), .A2(n9912), .ZN(n11050) );
  NAND2_X1 U11862 ( .A1(n14202), .A2(n10299), .ZN(n11052) );
  NAND2_X1 U11863 ( .A1(n10247), .A2(n10246), .ZN(n10299) );
  INV_X1 U11864 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10246) );
  NAND2_X1 U11865 ( .A1(n10009), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10247) );
  NAND2_X1 U11866 ( .A1(n9816), .A2(n10466), .ZN(n10465) );
  INV_X1 U11867 ( .A(n14722), .ZN(n10565) );
  NAND2_X1 U11869 ( .A1(n11129), .A2(n10735), .ZN(n15198) );
  NAND2_X1 U11870 ( .A1(n10178), .A2(n9840), .ZN(n15314) );
  INV_X1 U11871 ( .A(n15329), .ZN(n10178) );
  INV_X1 U11872 ( .A(n10013), .ZN(n15352) );
  INV_X1 U11873 ( .A(n11103), .ZN(n10378) );
  NAND2_X1 U11874 ( .A1(n10916), .A2(n10972), .ZN(n10153) );
  XNOR2_X1 U11875 ( .A(n14013), .B(n14275), .ZN(n13994) );
  NAND2_X1 U11876 ( .A1(n14374), .A2(n14373), .ZN(n21082) );
  INV_X1 U11877 ( .A(n21110), .ZN(n21137) );
  OAI21_X1 U11878 ( .B1(n14409), .B2(n21160), .A(n21288), .ZN(n14418) );
  CLKBUF_X1 U11879 ( .A(n10994), .Z(n14729) );
  INV_X1 U11880 ( .A(n21264), .ZN(n21258) );
  AND2_X1 U11881 ( .A1(n14113), .A2(n21287), .ZN(n21257) );
  OR2_X1 U11882 ( .A1(n14373), .A2(n9746), .ZN(n21264) );
  INV_X1 U11883 ( .A(n21330), .ZN(n21407) );
  OR2_X1 U11884 ( .A1(n14113), .A2(n14375), .ZN(n21339) );
  NOR2_X1 U11885 ( .A1(n21228), .A2(n14414), .ZN(n21376) );
  AOI21_X1 U11886 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21329), .A(n14414), 
        .ZN(n21416) );
  AND2_X1 U11887 ( .A1(n9874), .A2(n21486), .ZN(n14234) );
  AND2_X1 U11888 ( .A1(n16899), .A2(n16897), .ZN(n13422) );
  AND2_X1 U11889 ( .A1(n11902), .A2(n11901), .ZN(n16897) );
  OR2_X1 U11890 ( .A1(n11900), .A2(n11907), .ZN(n11901) );
  INV_X1 U11891 ( .A(n16802), .ZN(n16896) );
  OR2_X1 U11892 ( .A1(n15627), .A2(n10319), .ZN(n10335) );
  INV_X1 U11893 ( .A(n11845), .ZN(n15651) );
  NAND2_X1 U11894 ( .A1(n10657), .A2(n11760), .ZN(n10656) );
  INV_X1 U11895 ( .A(n11759), .ZN(n10657) );
  OR2_X1 U11896 ( .A1(n12327), .A2(n16359), .ZN(n12331) );
  INV_X1 U11897 ( .A(n11791), .ZN(n11757) );
  NAND2_X1 U11898 ( .A1(n11676), .A2(n10113), .ZN(n11712) );
  NOR2_X1 U11899 ( .A1(n10114), .A2(n10652), .ZN(n10113) );
  INV_X1 U11900 ( .A(n10116), .ZN(n10114) );
  INV_X1 U11901 ( .A(n15991), .ZN(n15951) );
  AND3_X1 U11902 ( .A1(n12155), .A2(n12154), .A3(n12153), .ZN(n14061) );
  OAI211_X1 U11903 ( .C1(n12220), .C2(n12076), .A(n12088), .B(n12075), .ZN(
        n13954) );
  OR2_X1 U11904 ( .A1(n16191), .A2(n12396), .ZN(n13952) );
  NAND2_X1 U11905 ( .A1(n16894), .A2(n16887), .ZN(n20030) );
  NAND3_X1 U11906 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12308) );
  AND2_X1 U11907 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12306) );
  INV_X1 U11908 ( .A(n14627), .ZN(n10614) );
  NAND2_X1 U11909 ( .A1(n14600), .A2(n14599), .ZN(n14603) );
  NOR2_X2 U11910 ( .A1(n15678), .A2(n15665), .ZN(n15667) );
  INV_X1 U11911 ( .A(n10709), .ZN(n10707) );
  INV_X1 U11912 ( .A(n10475), .ZN(n10474) );
  NOR2_X1 U11913 ( .A1(n11822), .A2(n10476), .ZN(n10404) );
  OAI21_X1 U11914 ( .B1(n12424), .B2(n10365), .A(n16313), .ZN(n10364) );
  NAND2_X1 U11915 ( .A1(n14695), .A2(n10086), .ZN(n10087) );
  AND2_X1 U11916 ( .A1(n10612), .A2(n16312), .ZN(n10086) );
  NOR2_X1 U11917 ( .A1(n10084), .A2(n10083), .ZN(n10082) );
  NAND2_X1 U11918 ( .A1(n10525), .A2(n10523), .ZN(n10522) );
  NAND2_X1 U11919 ( .A1(n12414), .A2(n12416), .ZN(n10523) );
  NAND2_X1 U11920 ( .A1(n10524), .A2(n12416), .ZN(n10521) );
  OR2_X1 U11921 ( .A1(n16685), .A2(n16656), .ZN(n16633) );
  NAND2_X1 U11922 ( .A1(n10166), .A2(n10165), .ZN(n10164) );
  NAND2_X1 U11923 ( .A1(n10173), .A2(n16392), .ZN(n10165) );
  OAI21_X1 U11924 ( .B1(n10170), .B2(n10169), .A(n16394), .ZN(n10166) );
  AND2_X1 U11925 ( .A1(n10395), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10392) );
  INV_X1 U11926 ( .A(n11934), .ZN(n16417) );
  NAND2_X1 U11927 ( .A1(n11705), .A2(n12207), .ZN(n10605) );
  NAND2_X1 U11928 ( .A1(n9978), .A2(n9877), .ZN(n16741) );
  NAND2_X1 U11929 ( .A1(n9979), .A2(n10431), .ZN(n9978) );
  NAND2_X1 U11930 ( .A1(n9977), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9976) );
  INV_X1 U11931 ( .A(n10430), .ZN(n16458) );
  XNOR2_X1 U11932 ( .A(n11509), .B(n11510), .ZN(n9971) );
  NAND2_X1 U11933 ( .A1(n12255), .A2(n12047), .ZN(n12052) );
  NAND2_X1 U11934 ( .A1(n12527), .A2(n12526), .ZN(n12529) );
  INV_X1 U11935 ( .A(n20174), .ZN(n20178) );
  OR2_X1 U11936 ( .A1(n11603), .A2(n20489), .ZN(n10130) );
  NAND2_X1 U11937 ( .A1(n16856), .A2(n20750), .ZN(n20396) );
  INV_X1 U11938 ( .A(n20746), .ZN(n20453) );
  INV_X1 U11939 ( .A(n20517), .ZN(n10016) );
  NAND2_X1 U11940 ( .A1(n20762), .A2(n20750), .ZN(n20535) );
  AND2_X2 U11941 ( .A1(n16842), .A2(n16841), .ZN(n20494) );
  NAND2_X1 U11942 ( .A1(n16938), .A2(n20808), .ZN(n16842) );
  INV_X1 U11943 ( .A(n13902), .ZN(n19789) );
  NOR2_X1 U11944 ( .A1(n17762), .A2(n17761), .ZN(n17760) );
  NAND2_X1 U11945 ( .A1(n10496), .A2(n10495), .ZN(n17782) );
  NAND2_X1 U11946 ( .A1(n18098), .A2(n17732), .ZN(n10495) );
  INV_X1 U11947 ( .A(n17796), .ZN(n10497) );
  NOR2_X1 U11948 ( .A1(n17839), .A2(n18098), .ZN(n17829) );
  NOR2_X1 U11949 ( .A1(n17858), .A2(n18098), .ZN(n17848) );
  INV_X1 U11950 ( .A(n17869), .ZN(n17859) );
  NOR2_X1 U11951 ( .A1(n17859), .A2(n18847), .ZN(n17858) );
  AND2_X1 U11952 ( .A1(n17213), .A2(n10499), .ZN(n17166) );
  AND2_X1 U11953 ( .A1(n10500), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10499) );
  NAND2_X1 U11954 ( .A1(n18629), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n10429) );
  NOR2_X1 U11955 ( .A1(n18502), .A2(n19373), .ZN(n17397) );
  INV_X1 U11956 ( .A(n19355), .ZN(n18651) );
  NAND2_X1 U11957 ( .A1(n17213), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17734) );
  AND2_X1 U11958 ( .A1(n17100), .A2(n9778), .ZN(n18814) );
  INV_X1 U11959 ( .A(n18895), .ZN(n10506) );
  INV_X1 U11960 ( .A(n17139), .ZN(n17137) );
  INV_X1 U11961 ( .A(n17058), .ZN(n10054) );
  NAND2_X1 U11962 ( .A1(n9716), .A2(n18811), .ZN(n18809) );
  OR2_X2 U11963 ( .A1(n13765), .A2(n13764), .ZN(n18707) );
  NAND2_X1 U11964 ( .A1(n18792), .A2(n10041), .ZN(n18783) );
  AND2_X1 U11965 ( .A1(n17085), .A2(n10061), .ZN(n10041) );
  INV_X1 U11966 ( .A(n17068), .ZN(n10046) );
  INV_X1 U11967 ( .A(n18986), .ZN(n10045) );
  NAND2_X1 U11968 ( .A1(n19237), .A2(n19314), .ZN(n19121) );
  NOR2_X1 U11969 ( .A1(n17723), .A2(n13770), .ZN(n17425) );
  OR2_X1 U11970 ( .A1(n14245), .A2(n14243), .ZN(n15047) );
  OR2_X1 U11971 ( .A1(n14245), .A2(n14238), .ZN(n20894) );
  INV_X1 U11972 ( .A(n15151), .ZN(n15156) );
  INV_X1 U11973 ( .A(n10548), .ZN(n10547) );
  OR2_X1 U11974 ( .A1(n13304), .A2(n13305), .ZN(n13306) );
  NAND2_X1 U11975 ( .A1(n20829), .A2(n13313), .ZN(n17533) );
  INV_X1 U11976 ( .A(n17533), .ZN(n17517) );
  NAND2_X1 U11977 ( .A1(n13307), .A2(n21420), .ZN(n15370) );
  NAND2_X1 U11978 ( .A1(n15375), .A2(n10195), .ZN(n12816) );
  NOR2_X1 U11979 ( .A1(n10196), .A2(n12812), .ZN(n10195) );
  NOR2_X1 U11980 ( .A1(n15563), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10196) );
  NAND2_X1 U11981 ( .A1(n12801), .A2(n13308), .ZN(n11130) );
  NAND2_X1 U11982 ( .A1(n12816), .A2(n10194), .ZN(n11374) );
  NAND2_X1 U11983 ( .A1(n12813), .A2(n12812), .ZN(n10194) );
  XNOR2_X1 U11984 ( .A(n9821), .B(n13309), .ZN(n15379) );
  OAI21_X1 U11985 ( .B1(n15463), .B2(n15244), .A(n10191), .ZN(n15447) );
  OR2_X1 U11986 ( .A1(n11365), .A2(n15477), .ZN(n10191) );
  AND2_X1 U11987 ( .A1(n15480), .A2(n15479), .ZN(n15506) );
  INV_X1 U11988 ( .A(n15304), .ZN(n10375) );
  NAND2_X1 U11989 ( .A1(n15306), .A2(n15305), .ZN(n10376) );
  OR2_X1 U11990 ( .A1(n15533), .A2(n14134), .ZN(n14135) );
  CLKBUF_X1 U11991 ( .A(n11212), .Z(n11213) );
  AND2_X1 U11992 ( .A1(n11354), .A2(n11326), .ZN(n20998) );
  INV_X1 U11993 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21329) );
  INV_X1 U11994 ( .A(n21420), .ZN(n21418) );
  INV_X1 U11995 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21409) );
  INV_X1 U11996 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13446) );
  OAI21_X1 U11997 ( .B1(n11191), .B2(n11188), .A(n11187), .ZN(n11193) );
  AND2_X1 U11998 ( .A1(n11186), .A2(n11189), .ZN(n11188) );
  NAND2_X1 U11999 ( .A1(n13422), .A2(n20026), .ZN(n20805) );
  NAND2_X1 U12000 ( .A1(n10327), .A2(n10325), .ZN(n15617) );
  AND2_X1 U12001 ( .A1(n10328), .A2(n10326), .ZN(n10325) );
  OR2_X1 U12002 ( .A1(n15967), .A2(n16230), .ZN(n10328) );
  NAND2_X1 U12003 ( .A1(n10331), .A2(n10330), .ZN(n10329) );
  INV_X1 U12004 ( .A(n15622), .ZN(n10330) );
  NAND2_X1 U12005 ( .A1(n16493), .A2(n12388), .ZN(n10331) );
  NAND3_X1 U12006 ( .A1(n9923), .A2(n10480), .A3(n11500), .ZN(n9922) );
  NAND2_X1 U12007 ( .A1(n10319), .A2(n19994), .ZN(n15969) );
  XNOR2_X1 U12008 ( .A(n15616), .B(n12799), .ZN(n16473) );
  INV_X1 U12009 ( .A(n20762), .ZN(n16856) );
  NAND2_X1 U12010 ( .A1(n13532), .A2(n16799), .ZN(n12797) );
  INV_X1 U12011 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U12013 ( .A1(n10073), .A2(n14598), .ZN(n11854) );
  NAND2_X1 U12014 ( .A1(n10386), .A2(n16660), .ZN(n10385) );
  OR2_X1 U12015 ( .A1(n10173), .A2(n10169), .ZN(n10168) );
  INV_X1 U12016 ( .A(n16672), .ZN(n10352) );
  AOI21_X1 U12017 ( .B1(n16416), .B2(n11933), .A(n9973), .ZN(n16693) );
  INV_X1 U12018 ( .A(n16414), .ZN(n10206) );
  AND2_X1 U12019 ( .A1(n17599), .A2(n12268), .ZN(n16454) );
  NAND2_X1 U12020 ( .A1(n17599), .A2(n13565), .ZN(n16448) );
  NAND2_X1 U12021 ( .A1(n13424), .A2(n12267), .ZN(n17599) );
  INV_X1 U12022 ( .A(n16448), .ZN(n17586) );
  INV_X1 U12023 ( .A(n16454), .ZN(n17589) );
  OR2_X1 U12024 ( .A1(n14680), .A2(n10716), .ZN(n14681) );
  NAND2_X1 U12025 ( .A1(n10416), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U12026 ( .A1(n10415), .A2(n16217), .ZN(n10414) );
  XNOR2_X1 U12027 ( .A(n10473), .B(n9818), .ZN(n16484) );
  NAND2_X1 U12028 ( .A1(n16216), .A2(n16224), .ZN(n10473) );
  INV_X1 U12029 ( .A(n16229), .ZN(n9965) );
  AND2_X1 U12030 ( .A1(n16515), .A2(n12061), .ZN(n16491) );
  INV_X1 U12031 ( .A(n14598), .ZN(n10072) );
  INV_X1 U12032 ( .A(n10074), .ZN(n10073) );
  OAI21_X1 U12033 ( .B1(n14600), .B2(n14601), .A(n14599), .ZN(n10074) );
  NOR2_X1 U12034 ( .A1(n11854), .A2(n14630), .ZN(n12261) );
  NAND2_X1 U12035 ( .A1(n16255), .A2(n9844), .ZN(n16522) );
  NAND2_X1 U12036 ( .A1(n12433), .A2(n12434), .ZN(n10265) );
  NAND2_X1 U12037 ( .A1(n9944), .A2(n9878), .ZN(n9943) );
  OAI21_X1 U12038 ( .B1(n16363), .B2(n9789), .A(n10684), .ZN(n9983) );
  NAND2_X1 U12039 ( .A1(n16615), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10684) );
  NAND2_X1 U12040 ( .A1(n10517), .A2(n9779), .ZN(n10518) );
  INV_X1 U12041 ( .A(n16345), .ZN(n10517) );
  NAND2_X1 U12042 ( .A1(n16377), .A2(n12416), .ZN(n10132) );
  NAND2_X1 U12043 ( .A1(n12415), .A2(n12414), .ZN(n16376) );
  AND2_X1 U12044 ( .A1(n10173), .A2(n10170), .ZN(n10161) );
  AND2_X1 U12045 ( .A1(n12255), .A2(n20789), .ZN(n17606) );
  NAND2_X1 U12046 ( .A1(n12255), .A2(n12026), .ZN(n16764) );
  AND2_X1 U12047 ( .A1(n12255), .A2(n12254), .ZN(n17608) );
  INV_X1 U12048 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20766) );
  INV_X1 U12049 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20758) );
  NAND2_X1 U12050 ( .A1(n20762), .A2(n20769), .ZN(n20752) );
  NAND2_X1 U12051 ( .A1(n19958), .A2(n18651), .ZN(n19956) );
  INV_X1 U12052 ( .A(n17747), .ZN(n10512) );
  NOR2_X1 U12053 ( .A1(n10511), .A2(n10510), .ZN(n10509) );
  NOR2_X1 U12054 ( .A1(n18096), .A2(n17749), .ZN(n10510) );
  INV_X1 U12055 ( .A(n17748), .ZN(n10511) );
  NOR2_X1 U12056 ( .A1(n17760), .A2(n18098), .ZN(n17751) );
  INV_X1 U12057 ( .A(n18113), .ZN(n18091) );
  INV_X1 U12058 ( .A(n18076), .ZN(n18112) );
  OR3_X1 U12059 ( .A1(n13676), .A2(n13675), .A3(n13674), .ZN(n13683) );
  NOR2_X1 U12060 ( .A1(n16973), .A2(n10429), .ZN(n18617) );
  INV_X1 U12061 ( .A(n18618), .ZN(n18643) );
  INV_X1 U12062 ( .A(n18625), .ZN(n18645) );
  INV_X1 U12063 ( .A(n18632), .ZN(n18625) );
  NOR2_X1 U12064 ( .A1(n17379), .A2(n18966), .ZN(n10235) );
  NAND2_X1 U12065 ( .A1(n17332), .A2(n10536), .ZN(n17334) );
  INV_X1 U12066 ( .A(n10537), .ZN(n10536) );
  OAI21_X1 U12067 ( .B1(n17350), .B2(n17333), .A(n17331), .ZN(n10537) );
  AND2_X1 U12068 ( .A1(n17344), .A2(n17343), .ZN(n19106) );
  NOR2_X1 U12069 ( .A1(n19137), .A2(n10489), .ZN(n19123) );
  NOR2_X1 U12070 ( .A1(n19237), .A2(n10490), .ZN(n10489) );
  NOR2_X1 U12071 ( .A1(n19111), .A2(n19110), .ZN(n10490) );
  OAI21_X1 U12072 ( .B1(n10488), .B2(n10486), .A(n19156), .ZN(n19135) );
  NAND2_X1 U12073 ( .A1(n10487), .A2(n19122), .ZN(n10486) );
  INV_X1 U12074 ( .A(n19123), .ZN(n10488) );
  NAND2_X1 U12075 ( .A1(n19234), .A2(n19124), .ZN(n10487) );
  AND2_X1 U12076 ( .A1(n13826), .A2(n19938), .ZN(n19323) );
  INV_X1 U12077 ( .A(n19323), .ZN(n19336) );
  AOI21_X1 U12078 ( .B1(n9801), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n10020), .ZN(n11612) );
  INV_X1 U12079 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10021) );
  AOI22_X1 U12080 ( .A1(n11603), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11604), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11608) );
  NAND2_X1 U12081 ( .A1(n11154), .A2(n11153), .ZN(n11163) );
  NAND2_X1 U12082 ( .A1(n20766), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11660) );
  NAND2_X1 U12083 ( .A1(n20103), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10390) );
  NAND2_X1 U12084 ( .A1(n20249), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U12085 ( .A1(n20336), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U12086 ( .A1(n11604), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U12087 ( .A1(n20212), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10287) );
  INV_X1 U12088 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n9958) );
  NOR2_X1 U12089 ( .A1(n16887), .A2(n11890), .ZN(n9940) );
  NOR2_X1 U12090 ( .A1(n16792), .A2(n20808), .ZN(n10077) );
  AND2_X1 U12091 ( .A1(n11064), .A2(n11063), .ZN(n11066) );
  CLKBUF_X1 U12092 ( .A(n10955), .Z(n13292) );
  AND2_X1 U12093 ( .A1(n10281), .A2(n10553), .ZN(n11016) );
  INV_X1 U12094 ( .A(n15176), .ZN(n10639) );
  AND2_X1 U12095 ( .A1(n11008), .A2(n11007), .ZN(n11065) );
  INV_X1 U12096 ( .A(n17482), .ZN(n13348) );
  NOR2_X1 U12097 ( .A1(n10946), .A2(n20825), .ZN(n10949) );
  NOR2_X1 U12098 ( .A1(n10880), .A2(n20825), .ZN(n10446) );
  NAND2_X1 U12099 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10853) );
  AOI22_X1 U12100 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10741), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U12101 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10925), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U12102 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10811), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U12103 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10761) );
  AOI22_X1 U12104 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10788) );
  XNOR2_X1 U12105 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11664) );
  AOI21_X1 U12106 ( .B1(n11574), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n10031), .ZN(n11575) );
  AND2_X1 U12107 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10031) );
  INV_X1 U12108 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10277) );
  NAND2_X1 U12109 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10029) );
  INV_X1 U12110 ( .A(n11628), .ZN(n10027) );
  NAND2_X1 U12111 ( .A1(n11626), .A2(n11627), .ZN(n10025) );
  AOI22_X1 U12112 ( .A1(n11603), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11604), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11714) );
  NAND2_X1 U12113 ( .A1(n16862), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10017) );
  INV_X1 U12114 ( .A(n10022), .ZN(n10019) );
  NAND2_X1 U12115 ( .A1(n10249), .A2(n10388), .ZN(n10387) );
  INV_X1 U12116 ( .A(n11731), .ZN(n10249) );
  NAND2_X1 U12117 ( .A1(n20103), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U12118 ( .A1(n10040), .A2(n9842), .ZN(n10629) );
  NAND2_X1 U12119 ( .A1(n16862), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10627) );
  NAND2_X1 U12120 ( .A1(n10040), .A2(n9834), .ZN(n10626) );
  AOI22_X1 U12121 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20524), .B1(
        n11605), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U12122 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11603), .B1(
        n20212), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11549) );
  NAND2_X1 U12123 ( .A1(n16862), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10513) );
  NAND2_X1 U12124 ( .A1(n16884), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10471) );
  NAND2_X1 U12125 ( .A1(n10040), .A2(n9781), .ZN(n9992) );
  NAND2_X1 U12126 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20786), .ZN(
        n11858) );
  AOI21_X1 U12127 ( .B1(n12366), .B2(P2_EBX_REG_1__SCAN_IN), .A(n9883), .ZN(
        n10078) );
  INV_X1 U12128 ( .A(n9956), .ZN(n9955) );
  OAI21_X1 U12129 ( .B1(n11683), .B2(n11898), .A(n11902), .ZN(n9956) );
  NOR2_X1 U12130 ( .A1(n11513), .A2(n10204), .ZN(n11521) );
  NAND2_X1 U12131 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10705) );
  NAND2_X1 U12132 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10704) );
  NAND2_X1 U12133 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U12134 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10348) );
  AOI21_X1 U12135 ( .B1(n9739), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10349) );
  NAND2_X1 U12136 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10134) );
  NAND2_X1 U12137 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10135) );
  NAND2_X1 U12138 ( .A1(n11536), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11439) );
  NAND2_X1 U12139 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11440) );
  NOR2_X1 U12140 ( .A1(n17215), .A2(n18110), .ZN(n10502) );
  NAND2_X1 U12141 ( .A1(n16990), .A2(n17114), .ZN(n17059) );
  NOR2_X1 U12142 ( .A1(n13811), .A2(n13812), .ZN(n13810) );
  NAND2_X1 U12143 ( .A1(n13778), .A2(n13816), .ZN(n13780) );
  AND2_X1 U12144 ( .A1(n11142), .A2(n11141), .ZN(n11179) );
  AND2_X1 U12145 ( .A1(n10692), .A2(n10693), .ZN(n10691) );
  INV_X1 U12146 ( .A(n14824), .ZN(n10692) );
  AND2_X1 U12147 ( .A1(n9838), .A2(n14403), .ZN(n10283) );
  INV_X1 U12148 ( .A(n14904), .ZN(n10688) );
  NAND2_X1 U12149 ( .A1(n11088), .A2(n11107), .ZN(n12868) );
  CLKBUF_X1 U12150 ( .A(n11016), .Z(n11017) );
  AND2_X1 U12151 ( .A1(n13308), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10467) );
  AND2_X1 U12152 ( .A1(n10638), .A2(n10467), .ZN(n10466) );
  NOR2_X1 U12153 ( .A1(n10154), .A2(n11372), .ZN(n10637) );
  AND2_X1 U12154 ( .A1(n10639), .A2(n15381), .ZN(n10181) );
  INV_X1 U12155 ( .A(n14761), .ZN(n10566) );
  NOR2_X1 U12156 ( .A1(n14778), .A2(n10568), .ZN(n10567) );
  INV_X1 U12157 ( .A(n14782), .ZN(n10568) );
  NOR2_X1 U12158 ( .A1(n14878), .A2(n10570), .ZN(n10569) );
  INV_X1 U12159 ( .A(n10571), .ZN(n10570) );
  NAND2_X1 U12160 ( .A1(n15291), .A2(n15305), .ZN(n15277) );
  INV_X1 U12161 ( .A(n14455), .ZN(n10562) );
  OR2_X1 U12162 ( .A1(n11121), .A2(n11120), .ZN(n15278) );
  NAND2_X1 U12163 ( .A1(n12883), .A2(n13621), .ZN(n11101) );
  NAND2_X1 U12164 ( .A1(n11047), .A2(n11046), .ZN(n14127) );
  NAND2_X1 U12165 ( .A1(n10185), .A2(n14290), .ZN(n10184) );
  INV_X1 U12166 ( .A(n11198), .ZN(n10185) );
  NAND2_X1 U12167 ( .A1(n17503), .A2(n10187), .ZN(n10186) );
  AND2_X1 U12168 ( .A1(n11197), .A2(n10281), .ZN(n10187) );
  OR2_X1 U12169 ( .A1(n10931), .A2(n10930), .ZN(n11024) );
  INV_X1 U12170 ( .A(n10949), .ZN(n11105) );
  AND2_X1 U12171 ( .A1(n10872), .A2(n10915), .ZN(n10452) );
  INV_X1 U12172 ( .A(n10889), .ZN(n10453) );
  NOR2_X1 U12173 ( .A1(n10873), .A2(n10888), .ZN(n10218) );
  OAI211_X1 U12174 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n13446), .A(n15604), 
        .B(n21475), .ZN(n14276) );
  NAND2_X1 U12175 ( .A1(n13994), .A2(n20825), .ZN(n10180) );
  OR2_X1 U12176 ( .A1(n11218), .A2(n20825), .ZN(n10980) );
  NOR2_X1 U12177 ( .A1(n9776), .A2(n9831), .ZN(n10198) );
  NAND2_X1 U12178 ( .A1(n11683), .A2(n11899), .ZN(n9961) );
  NAND2_X1 U12179 ( .A1(n11848), .A2(n11843), .ZN(n11845) );
  NAND2_X1 U12180 ( .A1(n15695), .A2(n15967), .ZN(n10318) );
  NAND2_X1 U12181 ( .A1(n10654), .A2(n9869), .ZN(n10653) );
  INV_X1 U12182 ( .A(n10655), .ZN(n10654) );
  NAND2_X1 U12183 ( .A1(n11713), .A2(n11732), .ZN(n10651) );
  AND2_X1 U12184 ( .A1(n10343), .A2(n10342), .ZN(n10341) );
  INV_X1 U12185 ( .A(n17585), .ZN(n10342) );
  AND2_X1 U12186 ( .A1(n15816), .A2(n14699), .ZN(n10578) );
  CLKBUF_X1 U12187 ( .A(n12644), .Z(n12781) );
  CLKBUF_X1 U12188 ( .A(n12639), .Z(n12785) );
  CLKBUF_X1 U12189 ( .A(n12640), .Z(n12782) );
  NOR2_X1 U12190 ( .A1(n15730), .A2(n15751), .ZN(n10602) );
  NOR2_X1 U12191 ( .A1(n10112), .A2(n10670), .ZN(n10111) );
  NAND2_X1 U12192 ( .A1(n10671), .A2(n16074), .ZN(n10670) );
  INV_X1 U12193 ( .A(n12551), .ZN(n10112) );
  INV_X1 U12194 ( .A(n10673), .ZN(n10671) );
  OR2_X1 U12195 ( .A1(n12353), .A2(n16242), .ZN(n12356) );
  INV_X1 U12196 ( .A(n13397), .ZN(n11975) );
  INV_X1 U12197 ( .A(n13396), .ZN(n11976) );
  INV_X1 U12198 ( .A(n13942), .ZN(n10580) );
  NOR2_X1 U12199 ( .A1(n10710), .A2(n16556), .ZN(n10708) );
  INV_X1 U12200 ( .A(n14610), .ZN(n10585) );
  NAND2_X1 U12201 ( .A1(n10150), .A2(n10034), .ZN(n10479) );
  AND2_X1 U12202 ( .A1(n10616), .A2(n9866), .ZN(n10615) );
  INV_X1 U12203 ( .A(n12249), .ZN(n10616) );
  INV_X1 U12204 ( .A(n16238), .ZN(n11844) );
  NOR2_X1 U12205 ( .A1(n10381), .A2(n9909), .ZN(n10380) );
  NAND2_X1 U12206 ( .A1(n9927), .A2(n16260), .ZN(n9926) );
  INV_X1 U12207 ( .A(n10034), .ZN(n9927) );
  OR2_X1 U12208 ( .A1(n15679), .A2(n14606), .ZN(n11836) );
  NOR2_X1 U12209 ( .A1(n16525), .A2(n16539), .ZN(n10709) );
  INV_X1 U12210 ( .A(n9909), .ZN(n10229) );
  NOR2_X1 U12211 ( .A1(n10706), .A2(n16305), .ZN(n10482) );
  NOR2_X1 U12212 ( .A1(n11991), .A2(n10577), .ZN(n10576) );
  OR2_X1 U12213 ( .A1(n15770), .A2(n12465), .ZN(n11991) );
  INV_X1 U12214 ( .A(n10578), .ZN(n10577) );
  AND2_X1 U12215 ( .A1(n9873), .A2(n15767), .ZN(n10617) );
  AND2_X1 U12216 ( .A1(n11965), .A2(n9997), .ZN(n9996) );
  INV_X1 U12217 ( .A(n14148), .ZN(n9997) );
  NOR2_X1 U12218 ( .A1(n9764), .A2(n10600), .ZN(n10599) );
  INV_X1 U12219 ( .A(n14053), .ZN(n10600) );
  NAND2_X1 U12220 ( .A1(n10515), .A2(n11939), .ZN(n10395) );
  NAND2_X1 U12221 ( .A1(n10075), .A2(n10409), .ZN(n10049) );
  INV_X1 U12222 ( .A(n19982), .ZN(n9977) );
  NOR2_X1 U12223 ( .A1(n11690), .A2(n10432), .ZN(n10431) );
  NOR2_X1 U12224 ( .A1(n10433), .A2(n14606), .ZN(n10432) );
  NOR2_X1 U12225 ( .A1(n11624), .A2(n11623), .ZN(n12105) );
  AND2_X1 U12226 ( .A1(n12104), .A2(n12103), .ZN(n14318) );
  AND2_X1 U12227 ( .A1(n12539), .A2(n10104), .ZN(n10103) );
  NAND2_X1 U12228 ( .A1(n12538), .A2(n16839), .ZN(n10104) );
  AND2_X1 U12229 ( .A1(n10014), .A2(n11487), .ZN(n11488) );
  NAND2_X1 U12230 ( .A1(n12541), .A2(n20800), .ZN(n12537) );
  AND2_X1 U12231 ( .A1(n13939), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U12232 ( .A1(n9762), .A2(n16887), .ZN(n16775) );
  AND4_X1 U12233 ( .A1(n11905), .A2(n11904), .A3(n12033), .A4(n11903), .ZN(
        n13533) );
  INV_X1 U12234 ( .A(n11384), .ZN(n9950) );
  NAND2_X1 U12235 ( .A1(n11420), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9933) );
  NAND2_X1 U12236 ( .A1(n11425), .A2(n11535), .ZN(n9932) );
  NAND2_X1 U12237 ( .A1(n20619), .A2(n20767), .ZN(n16848) );
  INV_X1 U12238 ( .A(n11464), .ZN(n11897) );
  INV_X1 U12239 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18272) );
  INV_X1 U12240 ( .A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18401) );
  NAND2_X1 U12241 ( .A1(n13666), .A2(n13660), .ZN(n13703) );
  NAND2_X1 U12242 ( .A1(n13666), .A2(n13654), .ZN(n18273) );
  NAND2_X1 U12243 ( .A1(n13782), .A2(n13780), .ZN(n13791) );
  NOR2_X1 U12244 ( .A1(n10501), .A2(n17182), .ZN(n10500) );
  INV_X1 U12245 ( .A(n10502), .ZN(n10501) );
  AND2_X1 U12246 ( .A1(n17244), .A2(n10505), .ZN(n10504) );
  AND2_X1 U12247 ( .A1(n17122), .A2(n17114), .ZN(n17121) );
  NOR2_X1 U12248 ( .A1(n10533), .A2(n18799), .ZN(n10532) );
  NAND2_X1 U12249 ( .A1(n18873), .A2(n17284), .ZN(n10533) );
  NOR2_X1 U12250 ( .A1(n19383), .A2(n19365), .ZN(n13782) );
  INV_X1 U12251 ( .A(n17077), .ZN(n10528) );
  XNOR2_X1 U12252 ( .A(n17124), .B(n10535), .ZN(n17051) );
  NOR2_X1 U12253 ( .A1(n13821), .A2(n19377), .ZN(n13851) );
  NOR2_X1 U12254 ( .A1(n13818), .A2(n13820), .ZN(n13902) );
  NAND2_X1 U12255 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13740) );
  AOI211_X1 U12256 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n13691), .B(n13690), .ZN(n13693) );
  NOR2_X1 U12257 ( .A1(n13898), .A2(n13791), .ZN(n14484) );
  INV_X1 U12258 ( .A(n13901), .ZN(n18650) );
  INV_X1 U12259 ( .A(n10888), .ZN(n13545) );
  INV_X1 U12260 ( .A(n15047), .ZN(n20857) );
  OR3_X1 U12261 ( .A1(n21572), .A2(n17539), .A3(n14236), .ZN(n15008) );
  AND2_X1 U12262 ( .A1(n11280), .A2(n11279), .ZN(n14931) );
  INV_X1 U12263 ( .A(n15096), .ZN(n14274) );
  NAND2_X1 U12264 ( .A1(n13318), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14227) );
  AOI22_X1 U12265 ( .A1(n14727), .A2(n14232), .B1(n13303), .B2(n13302), .ZN(
        n13305) );
  INV_X1 U12266 ( .A(n13221), .ZN(n13222) );
  OAI21_X1 U12267 ( .B1(n15202), .B2(n9867), .A(n13242), .ZN(n14784) );
  INV_X1 U12268 ( .A(n13179), .ZN(n13180) );
  NAND2_X1 U12269 ( .A1(n13203), .A2(n13202), .ZN(n14810) );
  OR2_X1 U12270 ( .A1(n15222), .A2(n9867), .ZN(n13203) );
  INV_X1 U12271 ( .A(n13126), .ZN(n13127) );
  OR2_X1 U12272 ( .A1(n15237), .A2(n9867), .ZN(n13150) );
  NOR2_X1 U12273 ( .A1(n13112), .A2(n10696), .ZN(n10695) );
  INV_X1 U12274 ( .A(n14854), .ZN(n10696) );
  INV_X1 U12275 ( .A(n13090), .ZN(n13091) );
  AND2_X1 U12276 ( .A1(n13111), .A2(n13110), .ZN(n14865) );
  OR2_X1 U12277 ( .A1(n15254), .A2(n9867), .ZN(n13111) );
  NOR2_X2 U12278 ( .A1(n13052), .A2(n14907), .ZN(n13053) );
  OR2_X1 U12279 ( .A1(n15271), .A2(n9867), .ZN(n13072) );
  INV_X1 U12280 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U12281 ( .A1(n13018), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13019) );
  OAI21_X1 U12282 ( .B1(n14960), .B2(n10067), .A(n9898), .ZN(n14963) );
  NOR2_X1 U12283 ( .A1(n15015), .A2(n14996), .ZN(n10067) );
  NAND2_X1 U12284 ( .A1(n12933), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12977) );
  AND4_X1 U12285 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n15016) );
  INV_X1 U12286 ( .A(n12909), .ZN(n12926) );
  AND2_X1 U12287 ( .A1(n14335), .A2(n10065), .ZN(n10064) );
  INV_X1 U12288 ( .A(n14367), .ZN(n10065) );
  NAND2_X1 U12289 ( .A1(n12877), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12909) );
  CLKBUF_X1 U12290 ( .A(n14105), .Z(n14106) );
  NAND2_X1 U12291 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12852) );
  OR2_X1 U12292 ( .A1(n14724), .A2(n12804), .ZN(n12807) );
  NAND2_X1 U12293 ( .A1(n14724), .A2(n12805), .ZN(n12806) );
  NAND2_X1 U12294 ( .A1(n14781), .A2(n10567), .ZN(n14776) );
  OR3_X1 U12295 ( .A1(n15428), .A2(n15399), .A3(n15199), .ZN(n15390) );
  AND2_X1 U12296 ( .A1(n11304), .A2(n11303), .ZN(n14819) );
  AND2_X1 U12297 ( .A1(n11301), .A2(n11300), .ZN(n14837) );
  NAND2_X1 U12298 ( .A1(n10174), .A2(n10156), .ZN(n15234) );
  AND2_X1 U12299 ( .A1(n11125), .A2(n9917), .ZN(n10356) );
  AND2_X1 U12300 ( .A1(n11286), .A2(n10569), .ZN(n14877) );
  NAND2_X1 U12301 ( .A1(n10735), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15262) );
  INV_X1 U12302 ( .A(n10447), .ZN(n15273) );
  AND2_X1 U12303 ( .A1(n11290), .A2(n11289), .ZN(n14894) );
  NAND2_X1 U12304 ( .A1(n11286), .A2(n10571), .ZN(n14892) );
  NAND2_X1 U12305 ( .A1(n14933), .A2(n14919), .ZN(n14918) );
  AND2_X1 U12306 ( .A1(n11278), .A2(n11277), .ZN(n14949) );
  NOR2_X2 U12307 ( .A1(n14968), .A2(n14949), .ZN(n14948) );
  INV_X1 U12308 ( .A(n15279), .ZN(n10012) );
  AND2_X1 U12309 ( .A1(n21003), .A2(n11357), .ZN(n15525) );
  NAND2_X1 U12310 ( .A1(n15313), .A2(n10179), .ZN(n15329) );
  AND2_X1 U12311 ( .A1(n11269), .A2(n11268), .ZN(n14999) );
  INV_X1 U12312 ( .A(n15278), .ZN(n15363) );
  NAND2_X1 U12313 ( .A1(n10154), .A2(n11112), .ZN(n14458) );
  XNOR2_X1 U12314 ( .A(n11102), .B(n17537), .ZN(n17512) );
  NAND2_X1 U12315 ( .A1(n17513), .A2(n17512), .ZN(n17511) );
  INV_X1 U12316 ( .A(n14211), .ZN(n10557) );
  CLKBUF_X1 U12317 ( .A(n14127), .Z(n14200) );
  INV_X1 U12318 ( .A(n14102), .ZN(n10555) );
  NAND2_X1 U12319 ( .A1(n10470), .A2(n12850), .ZN(n10248) );
  AND2_X1 U12320 ( .A1(n12848), .A2(n13621), .ZN(n10470) );
  CLKBUF_X1 U12321 ( .A(n11323), .Z(n11324) );
  CLKBUF_X1 U12322 ( .A(n11209), .Z(n11210) );
  NOR2_X1 U12323 ( .A1(n10918), .A2(n10354), .ZN(n10353) );
  INV_X1 U12324 ( .A(n10886), .ZN(n10354) );
  NAND2_X2 U12325 ( .A1(n10368), .A2(n10369), .ZN(n10314) );
  NAND2_X1 U12326 ( .A1(n10176), .A2(n10886), .ZN(n10369) );
  NAND2_X1 U12327 ( .A1(n10886), .A2(n10884), .ZN(n10454) );
  INV_X1 U12328 ( .A(n10904), .ZN(n10687) );
  INV_X1 U12329 ( .A(n12832), .ZN(n12833) );
  INV_X1 U12330 ( .A(n12831), .ZN(n12834) );
  NAND2_X1 U12331 ( .A1(n12850), .A2(n12848), .ZN(n14373) );
  OR2_X1 U12332 ( .A1(n14113), .A2(n21287), .ZN(n21109) );
  AND3_X1 U12333 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20825), .A3(n14276), 
        .ZN(n14307) );
  INV_X1 U12334 ( .A(n21225), .ZN(n21368) );
  INV_X1 U12335 ( .A(n14414), .ZN(n14305) );
  NOR2_X2 U12336 ( .A1(n15370), .A2(n14274), .ZN(n14304) );
  AND2_X1 U12337 ( .A1(n11140), .A2(n11139), .ZN(n11189) );
  NAND2_X1 U12338 ( .A1(n10125), .A2(n10124), .ZN(n11883) );
  NAND2_X1 U12339 ( .A1(n11683), .A2(n11855), .ZN(n10124) );
  MUX2_X1 U12340 ( .A(n11856), .B(n11918), .S(n12386), .Z(n11885) );
  NAND2_X1 U12341 ( .A1(n10319), .A2(n9785), .ZN(n10326) );
  AOI21_X1 U12342 ( .B1(n15681), .B2(n15967), .A(n16249), .ZN(n15662) );
  NAND2_X1 U12343 ( .A1(n10318), .A2(n10315), .ZN(n15681) );
  NOR2_X1 U12344 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  NOR2_X1 U12345 ( .A1(n10319), .A2(n15694), .ZN(n10317) );
  OAI21_X1 U12346 ( .B1(n15718), .B2(n15719), .A(n12347), .ZN(n15710) );
  AOI21_X1 U12347 ( .B1(n11843), .B2(n10646), .A(n9872), .ZN(n10645) );
  NAND2_X1 U12348 ( .A1(n10120), .A2(n11843), .ZN(n10123) );
  INV_X1 U12349 ( .A(n10648), .ZN(n10646) );
  NAND2_X1 U12350 ( .A1(n11824), .A2(n11843), .ZN(n11823) );
  NAND2_X1 U12351 ( .A1(n15737), .A2(n16297), .ZN(n15718) );
  NOR2_X1 U12352 ( .A1(n15755), .A2(n16308), .ZN(n15737) );
  OR2_X1 U12353 ( .A1(n11765), .A2(n11763), .ZN(n11764) );
  NOR2_X1 U12354 ( .A1(n11793), .A2(n11759), .ZN(n11773) );
  AND2_X1 U12355 ( .A1(n11800), .A2(n11799), .ZN(n15831) );
  NAND2_X1 U12356 ( .A1(n11755), .A2(n11754), .ZN(n11782) );
  INV_X1 U12357 ( .A(n16382), .ZN(n10336) );
  NAND2_X1 U12358 ( .A1(n15863), .A2(n10337), .ZN(n15846) );
  NAND2_X1 U12359 ( .A1(n10592), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12323) );
  NAND2_X1 U12360 ( .A1(n15863), .A2(n16404), .ZN(n15852) );
  NOR2_X1 U12361 ( .A1(n11674), .A2(n11680), .ZN(n10115) );
  NOR2_X1 U12362 ( .A1(n19991), .A2(n10344), .ZN(n10343) );
  INV_X1 U12363 ( .A(n15940), .ZN(n10344) );
  NAND2_X1 U12364 ( .A1(n11509), .A2(n11510), .ZN(n10002) );
  XNOR2_X1 U12365 ( .A(n11943), .B(n11506), .ZN(n11507) );
  OAI21_X1 U12366 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_0__SCAN_IN), .A(n10321), .ZN(n15963) );
  NAND2_X1 U12367 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10321) );
  AND2_X1 U12368 ( .A1(n15815), .A2(n15816), .ZN(n14698) );
  OR2_X1 U12369 ( .A1(n10674), .A2(n12552), .ZN(n10673) );
  NAND2_X1 U12370 ( .A1(n16087), .A2(n10675), .ZN(n10674) );
  OR2_X1 U12371 ( .A1(n12123), .A2(n12122), .ZN(n14216) );
  NAND2_X1 U12372 ( .A1(n12796), .A2(n16895), .ZN(n13532) );
  NOR2_X1 U12373 ( .A1(n10663), .A2(n10668), .ZN(n10661) );
  NAND2_X1 U12374 ( .A1(n16000), .A2(n10662), .ZN(n10664) );
  NOR2_X1 U12375 ( .A1(n10663), .A2(n16001), .ZN(n10662) );
  NAND2_X1 U12376 ( .A1(n10665), .A2(n10666), .ZN(n10102) );
  NAND2_X1 U12377 ( .A1(n16000), .A2(n12767), .ZN(n10666) );
  OR2_X1 U12378 ( .A1(n10677), .A2(n16043), .ZN(n10676) );
  AND2_X1 U12379 ( .A1(n12236), .A2(n12235), .ZN(n12438) );
  CLKBUF_X1 U12380 ( .A(n12435), .Z(n12436) );
  NOR2_X1 U12381 ( .A1(n16056), .A2(n10679), .ZN(n16051) );
  NOR2_X1 U12382 ( .A1(n16056), .A2(n16058), .ZN(n16057) );
  AND2_X1 U12383 ( .A1(n12226), .A2(n12225), .ZN(n12466) );
  AND2_X1 U12384 ( .A1(n12224), .A2(n12223), .ZN(n14703) );
  NAND2_X1 U12385 ( .A1(n14270), .A2(n10619), .ZN(n14701) );
  NAND2_X1 U12386 ( .A1(n12393), .A2(n12392), .ZN(n13526) );
  AND3_X1 U12387 ( .A1(n11465), .A2(n11892), .A3(n20135), .ZN(n12040) );
  XNOR2_X1 U12388 ( .A(n12302), .B(n12301), .ZN(n14621) );
  NOR2_X1 U12389 ( .A1(n12356), .A2(n21876), .ZN(n12358) );
  NAND2_X1 U12390 ( .A1(n12341), .A2(n9787), .ZN(n12350) );
  AND2_X1 U12391 ( .A1(n12341), .A2(n9889), .ZN(n12352) );
  NAND2_X1 U12392 ( .A1(n12341), .A2(n10595), .ZN(n12348) );
  NAND2_X1 U12393 ( .A1(n12341), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12345) );
  AND2_X1 U12394 ( .A1(n12334), .A2(n9890), .ZN(n12342) );
  NAND2_X1 U12395 ( .A1(n12334), .A2(n9788), .ZN(n12339) );
  NOR2_X1 U12396 ( .A1(n9758), .A2(n10594), .ZN(n10593) );
  INV_X1 U12397 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10594) );
  NOR2_X1 U12398 ( .A1(n12319), .A2(n9758), .ZN(n12328) );
  NAND2_X1 U12399 ( .A1(n10592), .A2(n9755), .ZN(n12325) );
  INV_X1 U12400 ( .A(n16392), .ZN(n10169) );
  NAND2_X1 U12401 ( .A1(n10588), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10587) );
  INV_X1 U12402 ( .A(n10590), .ZN(n10588) );
  NAND2_X1 U12403 ( .A1(n10589), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12315) );
  INV_X1 U12404 ( .A(n12312), .ZN(n10589) );
  OR2_X2 U12405 ( .A1(n11566), .A2(n11565), .ZN(n13563) );
  NAND2_X1 U12406 ( .A1(n15657), .A2(n10615), .ZN(n14628) );
  NAND2_X1 U12407 ( .A1(n14598), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14605) );
  OR2_X1 U12408 ( .A1(n15640), .A2(n14606), .ZN(n14601) );
  AND2_X1 U12409 ( .A1(n11853), .A2(n16252), .ZN(n14599) );
  NOR2_X1 U12410 ( .A1(n12433), .A2(n10023), .ZN(n16240) );
  INV_X1 U12411 ( .A(n10380), .ZN(n10023) );
  INV_X1 U12412 ( .A(n11840), .ZN(n16253) );
  NOR2_X1 U12413 ( .A1(n10573), .A2(n10575), .ZN(n10572) );
  INV_X1 U12414 ( .A(n15700), .ZN(n10575) );
  INV_X1 U12415 ( .A(n10574), .ZN(n10573) );
  NAND2_X1 U12416 ( .A1(n16270), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16262) );
  NAND2_X1 U12417 ( .A1(n12440), .A2(n12001), .ZN(n15709) );
  INV_X1 U12418 ( .A(n11822), .ZN(n10478) );
  AND2_X1 U12419 ( .A1(n16292), .A2(n16290), .ZN(n12427) );
  NAND2_X1 U12420 ( .A1(n10607), .A2(n10609), .ZN(n16291) );
  INV_X1 U12421 ( .A(n10610), .ZN(n10609) );
  OAI21_X1 U12422 ( .B1(n10612), .B2(n10611), .A(n12425), .ZN(n10610) );
  CLKBUF_X1 U12423 ( .A(n15748), .Z(n15749) );
  AND2_X1 U12424 ( .A1(n14270), .A2(n9873), .ZN(n15768) );
  AND2_X1 U12425 ( .A1(n10483), .A2(n16567), .ZN(n10481) );
  NOR2_X1 U12426 ( .A1(n10613), .A2(n12459), .ZN(n10612) );
  INV_X1 U12427 ( .A(n12422), .ZN(n10613) );
  NOR2_X1 U12428 ( .A1(n16364), .A2(n16356), .ZN(n16355) );
  INV_X1 U12429 ( .A(n16366), .ZN(n10438) );
  INV_X1 U12430 ( .A(n10522), .ZN(n10439) );
  AND3_X1 U12431 ( .A1(n12195), .A2(n12194), .A3(n12193), .ZN(n13393) );
  AND3_X1 U12432 ( .A1(n12180), .A2(n12179), .A3(n12178), .ZN(n14084) );
  CLKBUF_X1 U12433 ( .A(n14051), .Z(n14085) );
  NOR2_X1 U12434 ( .A1(n16393), .A2(n10171), .ZN(n10170) );
  OR2_X1 U12435 ( .A1(n16423), .A2(n10095), .ZN(n10094) );
  INV_X1 U12436 ( .A(n16391), .ZN(n10095) );
  NAND2_X1 U12437 ( .A1(n10579), .A2(n9999), .ZN(n9998) );
  INV_X1 U12438 ( .A(n14067), .ZN(n9999) );
  OR2_X1 U12439 ( .A1(n16728), .A2(n12055), .ZN(n16716) );
  CLKBUF_X1 U12440 ( .A(n14046), .Z(n14047) );
  NAND2_X1 U12441 ( .A1(n16766), .A2(n16751), .ZN(n16728) );
  INV_X1 U12442 ( .A(n17615), .ZN(n16568) );
  AND3_X1 U12443 ( .A1(n12101), .A2(n12100), .A3(n12099), .ZN(n16205) );
  AND3_X1 U12444 ( .A1(n10480), .A2(n11500), .A3(n11943), .ZN(n13944) );
  INV_X1 U12445 ( .A(n11929), .ZN(n10203) );
  NAND2_X1 U12446 ( .A1(n10703), .A2(n11591), .ZN(n10136) );
  OR2_X1 U12447 ( .A1(n12252), .A2(n16774), .ZN(n16803) );
  NAND2_X1 U12448 ( .A1(n13585), .A2(n13584), .ZN(n13587) );
  NAND2_X1 U12449 ( .A1(n11478), .A2(n9830), .ZN(n12022) );
  XNOR2_X1 U12450 ( .A(n12530), .B(n12531), .ZN(n13606) );
  AND2_X1 U12451 ( .A1(n16787), .A2(n11518), .ZN(n9991) );
  NOR2_X1 U12452 ( .A1(n20453), .A2(n20244), .ZN(n20179) );
  NOR2_X1 U12453 ( .A1(n11604), .A2(n20458), .ZN(n20462) );
  NOR2_X1 U12454 ( .A1(n20494), .A2(n20800), .ZN(n20136) );
  NOR2_X1 U12455 ( .A1(n17724), .A2(n17723), .ZN(n19788) );
  NOR2_X1 U12456 ( .A1(n17782), .A2(n18098), .ZN(n17774) );
  NOR2_X1 U12457 ( .A1(n17775), .A2(n17774), .ZN(n17773) );
  OR2_X1 U12458 ( .A1(n17848), .A2(n18837), .ZN(n10498) );
  NAND2_X1 U12459 ( .A1(n17742), .A2(n10720), .ZN(n17869) );
  INV_X1 U12460 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17983) );
  INV_X1 U12461 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17998) );
  NOR2_X1 U12462 ( .A1(n21671), .A2(n18973), .ZN(n10505) );
  NAND2_X1 U12463 ( .A1(n18191), .A2(n9795), .ZN(n18177) );
  NOR2_X1 U12464 ( .A1(n17834), .A2(n10149), .ZN(n10148) );
  INV_X1 U12465 ( .A(n17455), .ZN(n10144) );
  NOR2_X1 U12466 ( .A1(n18657), .A2(n10423), .ZN(n10422) );
  AND2_X1 U12467 ( .A1(n18592), .A2(n9792), .ZN(n18550) );
  NOR2_X1 U12468 ( .A1(n21685), .A2(n10425), .ZN(n10424) );
  OR2_X1 U12469 ( .A1(n17033), .A2(n17032), .ZN(n17116) );
  OR2_X1 U12470 ( .A1(n17004), .A2(n17003), .ZN(n17115) );
  AOI21_X1 U12471 ( .B1(n17419), .B2(n10715), .A(n13908), .ZN(n16954) );
  NOR2_X1 U12472 ( .A1(n18705), .A2(n18650), .ZN(n18676) );
  NAND2_X1 U12473 ( .A1(n17213), .A2(n10500), .ZN(n17187) );
  NOR3_X1 U12474 ( .A1(n17998), .A2(n17983), .A3(n17971), .ZN(n17244) );
  INV_X1 U12475 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17227) );
  NOR2_X1 U12476 ( .A1(n17227), .A2(n17952), .ZN(n18925) );
  NAND2_X1 U12477 ( .A1(n10504), .A2(n17261), .ZN(n18894) );
  NAND2_X1 U12478 ( .A1(n17261), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18006) );
  XNOR2_X1 U12479 ( .A(n10059), .B(n17056), .ZN(n19026) );
  NAND2_X1 U12480 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19007) );
  NAND2_X1 U12481 ( .A1(n17163), .A2(n10308), .ZN(n10307) );
  AND2_X1 U12482 ( .A1(n18771), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17363) );
  AND2_X1 U12483 ( .A1(n18910), .A2(n19070), .ZN(n10042) );
  INV_X1 U12484 ( .A(n10533), .ZN(n18795) );
  NAND2_X1 U12485 ( .A1(n18889), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10543) );
  AND2_X1 U12486 ( .A1(n18910), .A2(n10542), .ZN(n10541) );
  NAND2_X1 U12487 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U12488 ( .A1(n10313), .A2(n10309), .ZN(n18906) );
  AND2_X1 U12489 ( .A1(n17222), .A2(n19213), .ZN(n10309) );
  NAND2_X1 U12490 ( .A1(n18976), .A2(n17077), .ZN(n10529) );
  NAND2_X1 U12491 ( .A1(n17105), .A2(n17222), .ZN(n17268) );
  NAND2_X1 U12492 ( .A1(n17049), .A2(n17050), .ZN(n19036) );
  XNOR2_X1 U12493 ( .A(n17051), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19037) );
  NAND2_X1 U12494 ( .A1(n19037), .A2(n19036), .ZN(n19035) );
  NAND2_X1 U12495 ( .A1(n19951), .A2(n14484), .ZN(n19314) );
  NAND2_X1 U12496 ( .A1(n9808), .A2(n13849), .ZN(n17050) );
  NAND2_X1 U12497 ( .A1(n13786), .A2(n10419), .ZN(n13904) );
  INV_X1 U12498 ( .A(n13781), .ZN(n10419) );
  INV_X1 U12499 ( .A(n19314), .ZN(n19787) );
  NAND2_X1 U12500 ( .A1(n17425), .A2(n13905), .ZN(n17419) );
  INV_X1 U12501 ( .A(n13904), .ZN(n13905) );
  NOR2_X2 U12502 ( .A1(n13671), .A2(n13670), .ZN(n19373) );
  INV_X1 U12503 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21661) );
  NAND2_X1 U12504 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  NAND2_X1 U12505 ( .A1(n19786), .A2(n9870), .ZN(n10240) );
  NAND2_X1 U12506 ( .A1(n14226), .A2(n14225), .ZN(n21572) );
  INV_X1 U12507 ( .A(n20894), .ZN(n20909) );
  OR2_X1 U12508 ( .A1(n14245), .A2(n14244), .ZN(n20883) );
  AND2_X1 U12509 ( .A1(n20936), .A2(n14730), .ZN(n20931) );
  NAND2_X1 U12510 ( .A1(n13632), .A2(n13631), .ZN(n20936) );
  OR3_X1 U12511 ( .A1(n17503), .A2(n20822), .A3(n13990), .ZN(n13632) );
  INV_X1 U12512 ( .A(n20931), .ZN(n20925) );
  NOR2_X1 U12513 ( .A1(n15156), .A2(n13858), .ZN(n15158) );
  OR2_X1 U12514 ( .A1(n13630), .A2(n10888), .ZN(n13357) );
  NAND2_X1 U12515 ( .A1(n13992), .A2(n13550), .ZN(n13358) );
  INV_X1 U12516 ( .A(n15158), .ZN(n15153) );
  NAND2_X1 U12517 ( .A1(n13592), .A2(n13591), .ZN(n20940) );
  OR3_X1 U12518 ( .A1(n17497), .A2(n20822), .A3(n14003), .ZN(n13591) );
  INV_X2 U12519 ( .A(n14256), .ZN(n20993) );
  AOI22_X1 U12520 ( .A1(n12842), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13346), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13347) );
  XNOR2_X1 U12521 ( .A(n10223), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15168) );
  NAND2_X1 U12522 ( .A1(n10458), .A2(n10456), .ZN(n15193) );
  NAND2_X1 U12523 ( .A1(n15191), .A2(n11121), .ZN(n10458) );
  NAND2_X1 U12524 ( .A1(n15427), .A2(n10188), .ZN(n15412) );
  NOR2_X1 U12525 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  NOR2_X1 U12526 ( .A1(n11370), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10190) );
  INV_X1 U12527 ( .A(n11369), .ZN(n10189) );
  NAND2_X1 U12528 ( .A1(n11363), .A2(n11364), .ZN(n15463) );
  INV_X1 U12529 ( .A(n15509), .ZN(n10373) );
  NAND2_X1 U12530 ( .A1(n15352), .A2(n10155), .ZN(n15344) );
  OR2_X1 U12531 ( .A1(n14336), .A2(n14337), .ZN(n14365) );
  AND2_X1 U12532 ( .A1(n13884), .A2(n13883), .ZN(n15535) );
  NAND2_X1 U12533 ( .A1(n13635), .A2(n13634), .ZN(n13637) );
  XNOR2_X1 U12534 ( .A(n10560), .B(n13628), .ZN(n13635) );
  NAND2_X1 U12535 ( .A1(n10242), .A2(n14013), .ZN(n21291) );
  INV_X1 U12536 ( .A(n11035), .ZN(n10459) );
  INV_X1 U12537 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21008) );
  CLKBUF_X1 U12538 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n15602) );
  INV_X1 U12539 ( .A(n10871), .ZN(n13997) );
  NAND2_X1 U12540 ( .A1(n17503), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15604) );
  OAI22_X1 U12541 ( .A1(n21014), .A2(n21013), .B1(n21171), .B2(n21112), .ZN(
        n21033) );
  OAI211_X1 U12542 ( .C1(n21014), .C2(n21012), .A(n21236), .B(n21011), .ZN(
        n21034) );
  INV_X1 U12543 ( .A(n21058), .ZN(n21061) );
  OAI22_X1 U12544 ( .A1(n14385), .A2(n14379), .B1(n14410), .B2(n21171), .ZN(
        n21070) );
  INV_X1 U12545 ( .A(n21070), .ZN(n14401) );
  AND2_X1 U12546 ( .A1(n21076), .A2(n21225), .ZN(n21104) );
  OAI211_X1 U12547 ( .C1(n21088), .C2(n21087), .A(n21416), .B(n21086), .ZN(
        n21105) );
  OAI21_X1 U12548 ( .B1(n9906), .B2(n21116), .A(n21376), .ZN(n21133) );
  OAI211_X1 U12549 ( .C1(n14420), .C2(n21706), .A(n21376), .B(n14419), .ZN(
        n14447) );
  INV_X1 U12550 ( .A(n14449), .ZN(n14311) );
  OAI211_X1 U12551 ( .C1(n21177), .C2(n21176), .A(n21236), .B(n21175), .ZN(
        n21196) );
  INV_X1 U12552 ( .A(n21178), .ZN(n21195) );
  OAI211_X1 U12553 ( .C1(n9907), .C2(n21706), .A(n21376), .B(n21299), .ZN(
        n21324) );
  INV_X1 U12554 ( .A(n21366), .ZN(n21322) );
  AOI22_X1 U12555 ( .A1(n21298), .A2(n21295), .B1(n21293), .B2(n21292), .ZN(
        n21328) );
  OAI211_X1 U12556 ( .C1(n21401), .C2(n21377), .A(n21376), .B(n21375), .ZN(
        n21402) );
  INV_X1 U12557 ( .A(n14443), .ZN(n21412) );
  AND2_X1 U12558 ( .A1(n14305), .A2(n15141), .ZN(n21411) );
  INV_X1 U12559 ( .A(n14439), .ZN(n21426) );
  AND2_X1 U12560 ( .A1(n14305), .A2(n15129), .ZN(n21431) );
  INV_X1 U12561 ( .A(n21019), .ZN(n21432) );
  AND2_X1 U12562 ( .A1(n14305), .A2(n15124), .ZN(n21437) );
  INV_X1 U12563 ( .A(n21022), .ZN(n21438) );
  INV_X1 U12564 ( .A(n14428), .ZN(n21444) );
  AND2_X1 U12565 ( .A1(n14305), .A2(n15121), .ZN(n21443) );
  INV_X1 U12566 ( .A(n14432), .ZN(n21452) );
  AND2_X1 U12567 ( .A1(n14305), .A2(n15116), .ZN(n21451) );
  AND2_X1 U12568 ( .A1(n14305), .A2(n15112), .ZN(n21457) );
  INV_X1 U12569 ( .A(n21029), .ZN(n21458) );
  INV_X1 U12570 ( .A(n21449), .ZN(n21468) );
  INV_X1 U12571 ( .A(n14421), .ZN(n21466) );
  AND2_X1 U12572 ( .A1(n14305), .A2(n15108), .ZN(n21464) );
  INV_X2 U12573 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21578) );
  NAND2_X1 U12574 ( .A1(n13446), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21475) );
  AOI221_X1 U12575 ( .B1(n20825), .B2(n13446), .C1(n17498), .C2(n13446), .A(
        n17578), .ZN(n17580) );
  OR2_X1 U12576 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21483), .ZN(n21570) );
  AND2_X1 U12577 ( .A1(n11838), .A2(n11843), .ZN(n15670) );
  OR2_X1 U12578 ( .A1(n11793), .A2(n10656), .ZN(n11778) );
  NAND2_X1 U12579 ( .A1(n20805), .A2(n12296), .ZN(n15970) );
  NAND2_X1 U12580 ( .A1(n11748), .A2(n14040), .ZN(n11737) );
  NAND2_X1 U12581 ( .A1(n15938), .A2(n15940), .ZN(n19990) );
  INV_X1 U12582 ( .A(n16947), .ZN(n19994) );
  NAND2_X1 U12583 ( .A1(n15938), .A2(n10343), .ZN(n19993) );
  INV_X1 U12584 ( .A(n15970), .ZN(n19985) );
  NAND2_X1 U12585 ( .A1(n15967), .A2(n19994), .ZN(n15991) );
  AND2_X1 U12586 ( .A1(n15970), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19981) );
  NAND2_X1 U12587 ( .A1(n10323), .A2(n10322), .ZN(n16778) );
  NAND2_X1 U12588 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10322) );
  NAND2_X1 U12589 ( .A1(n20808), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10323) );
  OR2_X1 U12590 ( .A1(n12152), .A2(n12151), .ZN(n14032) );
  INV_X1 U12591 ( .A(n16080), .ZN(n16070) );
  INV_X1 U12592 ( .A(n20769), .ZN(n20750) );
  NAND2_X1 U12593 ( .A1(n16006), .A2(n16008), .ZN(n16007) );
  INV_X1 U12594 ( .A(n16184), .ZN(n16193) );
  OR2_X1 U12595 ( .A1(n16191), .A2(n9969), .ZN(n16184) );
  NAND2_X1 U12596 ( .A1(n12408), .A2(n16847), .ZN(n16197) );
  NOR2_X1 U12597 ( .A1(n12530), .A2(n13612), .ZN(n16855) );
  AND4_X1 U12598 ( .A1(n10271), .A2(n13611), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20800), .ZN(n13612) );
  INV_X1 U12599 ( .A(n16202), .ZN(n20020) );
  INV_X1 U12600 ( .A(n20002), .ZN(n20016) );
  AND2_X1 U12601 ( .A1(n20032), .A2(n20031), .ZN(n20082) );
  NOR2_X1 U12602 ( .A1(n20778), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20086) );
  BUF_X1 U12603 ( .A(n20086), .Z(n20799) );
  INV_X1 U12604 ( .A(n20028), .ZN(n13520) );
  OAI21_X1 U12605 ( .B1(n16029), .B2(n20812), .A(n13428), .ZN(n13452) );
  NAND2_X1 U12606 ( .A1(n10634), .A2(n12484), .ZN(n10633) );
  INV_X1 U12607 ( .A(n12501), .ZN(n10634) );
  NAND2_X1 U12608 ( .A1(n16473), .A2(n16454), .ZN(n16220) );
  NAND2_X1 U12609 ( .A1(n10686), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10685) );
  INV_X1 U12610 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16359) );
  INV_X1 U12611 ( .A(n17599), .ZN(n16445) );
  NAND2_X1 U12612 ( .A1(n12509), .A2(n17608), .ZN(n10632) );
  XNOR2_X1 U12613 ( .A(n12508), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14618) );
  AND2_X1 U12614 ( .A1(n12494), .A2(n16215), .ZN(n12495) );
  AND2_X1 U12615 ( .A1(n10633), .A2(n17602), .ZN(n10631) );
  AND2_X1 U12616 ( .A1(n16524), .A2(n16526), .ZN(n16515) );
  INV_X1 U12617 ( .A(n10402), .ZN(n10400) );
  NAND2_X1 U12618 ( .A1(n10401), .A2(n10474), .ZN(n16274) );
  AND2_X1 U12619 ( .A1(n12432), .A2(n17606), .ZN(n10097) );
  AND2_X1 U12620 ( .A1(n10039), .A2(n12433), .ZN(n16589) );
  NAND2_X1 U12621 ( .A1(n16304), .A2(n16305), .ZN(n10039) );
  XNOR2_X1 U12622 ( .A(n10366), .B(n16303), .ZN(n16591) );
  NAND2_X1 U12623 ( .A1(n10087), .A2(n10363), .ZN(n10366) );
  INV_X1 U12624 ( .A(n10364), .ZN(n10363) );
  XNOR2_X1 U12625 ( .A(n10260), .B(n10259), .ZN(n16606) );
  NAND2_X1 U12626 ( .A1(n16313), .A2(n16312), .ZN(n10259) );
  NAND2_X1 U12627 ( .A1(n10608), .A2(n12424), .ZN(n10260) );
  NAND2_X1 U12628 ( .A1(n14695), .A2(n10612), .ZN(n10608) );
  NAND2_X1 U12629 ( .A1(n9943), .A2(n9942), .ZN(n9945) );
  AND2_X1 U12630 ( .A1(n12458), .A2(n10712), .ZN(n9942) );
  XNOR2_X1 U12631 ( .A(n9980), .B(n10527), .ZN(n16332) );
  INV_X1 U12632 ( .A(n12459), .ZN(n10527) );
  NAND2_X1 U12633 ( .A1(n14695), .A2(n12422), .ZN(n9980) );
  NAND2_X1 U12634 ( .A1(n9986), .A2(n10521), .ZN(n16367) );
  NAND2_X1 U12635 ( .A1(n12415), .A2(n10522), .ZN(n9986) );
  INV_X1 U12636 ( .A(n16363), .ZN(n16378) );
  INV_X1 U12637 ( .A(n10386), .ZN(n16671) );
  OAI21_X1 U12638 ( .B1(n16416), .B2(n9973), .A(n9972), .ZN(n9974) );
  AOI21_X1 U12639 ( .B1(n9975), .B2(n10515), .A(n16748), .ZN(n9972) );
  XNOR2_X1 U12640 ( .A(n10088), .B(n16419), .ZN(n16712) );
  NOR2_X1 U12641 ( .A1(n16435), .A2(n9843), .ZN(n10088) );
  INV_X1 U12642 ( .A(n16423), .ZN(n16434) );
  CLKBUF_X1 U12643 ( .A(n16449), .Z(n16450) );
  NAND2_X1 U12644 ( .A1(n10434), .A2(n16456), .ZN(n16457) );
  OR2_X1 U12645 ( .A1(n9959), .A2(n17603), .ZN(n14670) );
  NOR2_X1 U12646 ( .A1(n12052), .A2(n13579), .ZN(n9959) );
  NOR2_X1 U12647 ( .A1(n12255), .A2(n16754), .ZN(n17603) );
  INV_X1 U12648 ( .A(n16855), .ZN(n20781) );
  CLKBUF_X1 U12649 ( .A(n12022), .Z(n16904) );
  NAND2_X1 U12650 ( .A1(n12523), .A2(n12534), .ZN(n13867) );
  AND2_X1 U12651 ( .A1(n16894), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16938) );
  INV_X1 U12652 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16924) );
  AND2_X1 U12653 ( .A1(n10389), .A2(n20800), .ZN(n20101) );
  OR2_X1 U12654 ( .A1(n20103), .A2(n20489), .ZN(n10389) );
  AND2_X1 U12655 ( .A1(n20152), .A2(n20149), .ZN(n20169) );
  OAI21_X1 U12656 ( .B1(n20215), .B2(n20210), .A(n20209), .ZN(n20240) );
  INV_X1 U12657 ( .A(n20253), .ZN(n20271) );
  NAND2_X1 U12658 ( .A1(n10131), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20281) );
  OR2_X1 U12659 ( .A1(n11603), .A2(n20280), .ZN(n10131) );
  OAI21_X1 U12660 ( .B1(n20283), .B2(n20279), .A(n20278), .ZN(n20309) );
  NAND2_X1 U12661 ( .A1(n10130), .A2(n20800), .ZN(n20277) );
  NAND2_X1 U12662 ( .A1(n16846), .A2(n16845), .ZN(n20329) );
  AOI211_X2 U12663 ( .C1(n16865), .C2(n16864), .A(n20494), .B(n16863), .ZN(
        n20393) );
  OAI21_X1 U12664 ( .B1(n20404), .B2(n20403), .A(n20402), .ZN(n20428) );
  NAND2_X1 U12665 ( .A1(n16882), .A2(n10472), .ZN(n16883) );
  OAI21_X1 U12666 ( .B1(n20455), .B2(n16886), .A(n16885), .ZN(n20448) );
  NOR2_X1 U12667 ( .A1(n20556), .A2(n20453), .ZN(n20475) );
  INV_X1 U12668 ( .A(n20475), .ZN(n20485) );
  OAI21_X1 U12669 ( .B1(n20517), .B2(n20800), .A(n20496), .ZN(n20521) );
  AOI21_X1 U12670 ( .B1(n20528), .B2(n20489), .A(n20527), .ZN(n20551) );
  AOI22_X1 U12671 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20133), .ZN(n20578) );
  NAND2_X1 U12672 ( .A1(n20136), .A2(n10037), .ZN(n20587) );
  NAND2_X1 U12673 ( .A1(n9994), .A2(n9993), .ZN(n20563) );
  NOR2_X1 U12674 ( .A1(n20565), .A2(n20749), .ZN(n9993) );
  OAI21_X1 U12675 ( .B1(n20568), .B2(n20567), .A(n20566), .ZN(n20606) );
  INV_X1 U12676 ( .A(n20559), .ZN(n20604) );
  NOR2_X1 U12677 ( .A1(n20556), .A2(n20752), .ZN(n20622) );
  INV_X1 U12678 ( .A(n20572), .ZN(n20627) );
  INV_X1 U12679 ( .A(n20577), .ZN(n20633) );
  INV_X1 U12680 ( .A(n20587), .ZN(n20645) );
  INV_X1 U12681 ( .A(n20592), .ZN(n20651) );
  INV_X1 U12682 ( .A(n20597), .ZN(n20657) );
  AND2_X1 U12683 ( .A1(n20099), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20663) );
  INV_X1 U12684 ( .A(n20602), .ZN(n20664) );
  INV_X1 U12685 ( .A(n19958), .ZN(n19954) );
  INV_X1 U12686 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n17725) );
  INV_X1 U12687 ( .A(n18706), .ZN(n18704) );
  NOR2_X1 U12688 ( .A1(n18117), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19955) );
  NAND2_X1 U12689 ( .A1(n17805), .A2(n10497), .ZN(n10494) );
  NOR2_X1 U12690 ( .A1(n17795), .A2(n17796), .ZN(n17794) );
  NOR2_X1 U12691 ( .A1(n17805), .A2(n18098), .ZN(n17795) );
  NOR2_X1 U12692 ( .A1(n17807), .A2(n17806), .ZN(n17805) );
  NOR2_X1 U12693 ( .A1(n17818), .A2(n18098), .ZN(n17806) );
  NOR2_X1 U12694 ( .A1(n18778), .A2(n17819), .ZN(n17818) );
  OAI22_X1 U12695 ( .A1(n17848), .A2(n9871), .B1(n17742), .B2(n18825), .ZN(
        n17839) );
  INV_X1 U12696 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17952) );
  INV_X1 U12697 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17971) );
  AND2_X1 U12698 ( .A1(n17261), .A2(n10505), .ZN(n17993) );
  INV_X1 U12699 ( .A(n18096), .ZN(n18099) );
  OR2_X1 U12700 ( .A1(n17728), .A2(n17727), .ZN(n18113) );
  OAI21_X1 U12701 ( .B1(n10143), .B2(n18498), .A(n9881), .ZN(n18168) );
  NOR2_X1 U12702 ( .A1(n18177), .A2(n17803), .ZN(n18181) );
  NOR2_X1 U12703 ( .A1(n18123), .A2(n18224), .ZN(n18191) );
  NOR2_X1 U12704 ( .A1(n18261), .A2(n18595), .ZN(n18244) );
  NOR2_X1 U12705 ( .A1(n21753), .A2(n18298), .ZN(n10147) );
  NAND2_X1 U12706 ( .A1(n18299), .A2(n10145), .ZN(n18261) );
  NOR2_X1 U12707 ( .A1(n10146), .A2(n17875), .ZN(n10145) );
  INV_X1 U12708 ( .A(n10147), .ZN(n10146) );
  NAND2_X1 U12709 ( .A1(n18299), .A2(P3_EBX_REG_17__SCAN_IN), .ZN(n18280) );
  NOR2_X1 U12710 ( .A1(n17906), .A2(n18337), .ZN(n18299) );
  NOR2_X1 U12711 ( .A1(n18355), .A2(n21674), .ZN(n18338) );
  NAND2_X1 U12712 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n18338), .ZN(n18337) );
  NAND2_X1 U12713 ( .A1(n9761), .A2(P3_EBX_REG_13__SCAN_IN), .ZN(n18355) );
  NAND2_X1 U12714 ( .A1(n9725), .A2(n17457), .ZN(n18477) );
  INV_X1 U12715 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n18478) );
  INV_X1 U12716 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n18486) );
  INV_X1 U12717 ( .A(n19383), .ZN(n18595) );
  INV_X1 U12718 ( .A(n18520), .ZN(n18515) );
  NAND2_X1 U12719 ( .A1(n18532), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n18528) );
  NOR2_X1 U12720 ( .A1(n18721), .A2(n18539), .ZN(n18532) );
  OR2_X1 U12721 ( .A1(n18719), .A2(n18538), .ZN(n18539) );
  NOR2_X1 U12722 ( .A1(n18545), .A2(n18717), .ZN(n18544) );
  NAND2_X1 U12723 ( .A1(n18592), .A2(n9791), .ZN(n18582) );
  INV_X1 U12724 ( .A(n18551), .ZN(n18580) );
  AND2_X1 U12725 ( .A1(n18592), .A2(n10424), .ZN(n18586) );
  NAND2_X1 U12726 ( .A1(n18592), .A2(P3_EAX_REG_14__SCAN_IN), .ZN(n18591) );
  NOR2_X1 U12727 ( .A1(n10429), .A2(n9900), .ZN(n10428) );
  INV_X1 U12728 ( .A(n18626), .ZN(n18648) );
  NOR2_X2 U12730 ( .A1(n18755), .A2(n19943), .ZN(n18756) );
  NAND2_X1 U12731 ( .A1(n10538), .A2(n17337), .ZN(n17194) );
  NAND2_X1 U12732 ( .A1(n17350), .A2(n18910), .ZN(n10538) );
  INV_X1 U12733 ( .A(n19049), .ZN(n17104) );
  NAND2_X1 U12734 ( .A1(n17100), .A2(n9756), .ZN(n18844) );
  NAND2_X1 U12735 ( .A1(n17100), .A2(n17099), .ZN(n18882) );
  AND2_X1 U12736 ( .A1(n19051), .A2(n18624), .ZN(n18946) );
  INV_X1 U12737 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21671) );
  NOR2_X1 U12738 ( .A1(n19007), .A2(n19022), .ZN(n19000) );
  INV_X1 U12739 ( .A(n19690), .ZN(n19730) );
  NAND2_X1 U12740 ( .A1(n19591), .A2(n19407), .ZN(n19690) );
  NAND2_X1 U12741 ( .A1(n18792), .A2(n17085), .ZN(n18785) );
  OR2_X1 U12742 ( .A1(n13903), .A2(n13897), .ZN(n10230) );
  AND2_X1 U12743 ( .A1(n19308), .A2(n17382), .ZN(n19263) );
  NAND2_X1 U12744 ( .A1(n10043), .A2(n17068), .ZN(n18987) );
  NAND2_X1 U12745 ( .A1(n18999), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10043) );
  INV_X1 U12746 ( .A(n19329), .ZN(n19290) );
  INV_X1 U12747 ( .A(n19786), .ZN(n19321) );
  INV_X1 U12748 ( .A(n19335), .ZN(n19285) );
  AND2_X1 U12749 ( .A1(n19786), .A2(n19323), .ZN(n19335) );
  INV_X1 U12750 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19587) );
  NOR3_X1 U12751 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19942), .ZN(n19407) );
  INV_X1 U12752 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19806) );
  INV_X1 U12753 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19814) );
  INV_X2 U12754 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17398) );
  INV_X1 U12755 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18649) );
  NOR2_X1 U12756 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19923), .ZN(
        n19821) );
  NOR2_X1 U12757 ( .A1(n17725), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19835) );
  OAI211_X1 U12758 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19853), .B(n21587), .ZN(n19941) );
  INV_X1 U12759 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19853) );
  CLKBUF_X1 U12760 ( .A(n19909), .Z(n21587) );
  NAND2_X1 U12761 ( .A1(n19853), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19933) );
  INV_X2 U12762 ( .A(n19933), .ZN(n21589) );
  INV_X1 U12764 ( .A(U212), .ZN(n17658) );
  CLKBUF_X1 U12765 ( .A(n17698), .Z(n17699) );
  AOI211_X1 U12766 ( .C1(n20919), .C2(n14727), .A(n14726), .B(n14725), .ZN(
        n14728) );
  INV_X1 U12767 ( .A(n10550), .ZN(n10549) );
  AND2_X1 U12768 ( .A1(n11131), .A2(n17531), .ZN(n10546) );
  OAI21_X1 U12769 ( .B1(n15379), .B2(n20829), .A(n9845), .ZN(P1_U2970) );
  NAND2_X1 U12770 ( .A1(n10010), .A2(n15311), .ZN(P1_U2984) );
  NAND2_X1 U12771 ( .A1(n10011), .A2(n17531), .ZN(n10010) );
  OAI21_X1 U12772 ( .B1(n10548), .B2(n10468), .A(n11376), .ZN(P1_U3001) );
  NAND2_X1 U12773 ( .A1(n11131), .A2(n20999), .ZN(n10468) );
  NAND2_X1 U12774 ( .A1(n10374), .A2(n10371), .ZN(P1_U3016) );
  AND2_X1 U12775 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  NAND2_X1 U12776 ( .A1(n10011), .A2(n20999), .ZN(n10374) );
  NAND2_X1 U12777 ( .A1(n15510), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10372) );
  AOI21_X1 U12778 ( .B1(n14683), .B2(n14692), .A(n14691), .ZN(n14694) );
  NAND2_X1 U12779 ( .A1(n14690), .A2(n14689), .ZN(n14691) );
  AOI21_X1 U12780 ( .B1(n10333), .B2(n10332), .A(n10329), .ZN(n15623) );
  NAND2_X1 U12781 ( .A1(n15618), .A2(n15969), .ZN(n10332) );
  NOR2_X1 U12782 ( .A1(n15948), .A2(n10226), .ZN(n15949) );
  NOR2_X1 U12783 ( .A1(n10717), .A2(n10723), .ZN(n12800) );
  OAI21_X1 U12784 ( .B1(n16480), .B2(n20002), .A(n14716), .ZN(n14717) );
  NAND2_X1 U12785 ( .A1(n12265), .A2(n17587), .ZN(n12278) );
  NAND2_X1 U12786 ( .A1(n11854), .A2(n14630), .ZN(n12265) );
  OAI211_X1 U12787 ( .C1(n16522), .C2(n16472), .A(n16259), .B(n10410), .ZN(
        P2_U2989) );
  AOI21_X1 U12788 ( .B1(n16519), .B2(n16454), .A(n16257), .ZN(n10410) );
  INV_X1 U12789 ( .A(n10278), .ZN(n16300) );
  AOI21_X1 U12790 ( .B1(n16566), .B2(n16454), .A(n16299), .ZN(n10279) );
  OAI21_X1 U12791 ( .B1(n10518), .B2(n17594), .A(n10397), .ZN(P2_U2999) );
  INV_X1 U12792 ( .A(n10398), .ZN(n10397) );
  INV_X1 U12793 ( .A(n16350), .ZN(n10399) );
  AOI21_X1 U12794 ( .B1(n16664), .B2(n16454), .A(n16398), .ZN(n10384) );
  AND2_X1 U12795 ( .A1(n10351), .A2(n10350), .ZN(n16407) );
  AOI21_X1 U12796 ( .B1(n16676), .B2(n16454), .A(n16406), .ZN(n10350) );
  AOI21_X1 U12797 ( .B1(n10208), .B2(n16405), .A(n10205), .ZN(n16415) );
  NAND2_X1 U12798 ( .A1(n10207), .A2(n10206), .ZN(n10205) );
  NOR2_X1 U12799 ( .A1(n16693), .A2(n17594), .ZN(n10208) );
  OAI21_X1 U12800 ( .B1(n10442), .B2(n16484), .A(n16483), .ZN(P2_U3016) );
  OAI211_X1 U12801 ( .C1(n16496), .C2(n10442), .A(n10581), .B(n10133), .ZN(
        P2_U3017) );
  AOI21_X1 U12802 ( .B1(n16493), .B2(n17604), .A(n10582), .ZN(n10581) );
  NAND2_X1 U12803 ( .A1(n10584), .A2(n10583), .ZN(n10582) );
  OAI211_X1 U12804 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n10073), .A(
        n10071), .B(n17602), .ZN(n10070) );
  NAND2_X1 U12805 ( .A1(n10072), .A2(n14630), .ZN(n10071) );
  INV_X1 U12806 ( .A(n10263), .ZN(n16578) );
  NOR2_X1 U12807 ( .A1(n16576), .A2(n9826), .ZN(n10264) );
  AND2_X1 U12808 ( .A1(n9943), .A2(n12458), .ZN(n14707) );
  OAI21_X1 U12809 ( .B1(n10518), .B2(n16748), .A(n10519), .ZN(P2_U3031) );
  INV_X1 U12810 ( .A(n10520), .ZN(n10519) );
  OAI21_X1 U12811 ( .B1(n16617), .B2(n10442), .A(n16616), .ZN(n10520) );
  NAND2_X1 U12812 ( .A1(n16644), .A2(n17606), .ZN(n16653) );
  NAND2_X1 U12813 ( .A1(n10167), .A2(n10162), .ZN(n16670) );
  OAI21_X1 U12814 ( .B1(n17751), .B2(n9897), .A(n10507), .ZN(P3_U2640) );
  AOI21_X1 U12815 ( .B1(n17757), .B2(n18129), .A(n10508), .ZN(n10507) );
  NAND2_X1 U12816 ( .A1(n10512), .A2(n10509), .ZN(n10508) );
  OAI21_X1 U12817 ( .B1(n10142), .B2(n21832), .A(n10140), .ZN(P3_U2674) );
  AOI21_X1 U12818 ( .B1(n18167), .B2(n21832), .A(n10141), .ZN(n10140) );
  INV_X1 U12819 ( .A(n18168), .ZN(n10142) );
  NOR2_X1 U12820 ( .A1(n18484), .A2(n18518), .ZN(n10141) );
  NAND2_X1 U12821 ( .A1(n10427), .A2(n18629), .ZN(n18619) );
  NAND2_X1 U12822 ( .A1(n17221), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10233) );
  NOR2_X1 U12823 ( .A1(n10235), .A2(n17220), .ZN(n10234) );
  OR4_X2 U12824 ( .A1(n18798), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n18773), .A4(n18799), .ZN(n10236) );
  OR2_X1 U12825 ( .A1(n17353), .A2(n10539), .ZN(P3_U2834) );
  OR2_X1 U12826 ( .A1(n17351), .A2(n17352), .ZN(n10539) );
  NAND2_X1 U12827 ( .A1(n19135), .A2(n10485), .ZN(n19127) );
  OR2_X1 U12828 ( .A1(n19125), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10485) );
  INV_X2 U12829 ( .A(n10932), .ZN(n13186) );
  AND2_X1 U12830 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n9755) );
  NAND2_X1 U12831 ( .A1(n11520), .A2(n10225), .ZN(n10266) );
  AND2_X1 U12832 ( .A1(n9769), .A2(n10730), .ZN(n9756) );
  INV_X1 U12833 ( .A(n14524), .ZN(n13831) );
  NAND2_X1 U12834 ( .A1(n10756), .A2(n13977), .ZN(n10762) );
  INV_X1 U12835 ( .A(n18193), .ZN(n13748) );
  NAND2_X1 U12836 ( .A1(n14270), .A2(n14356), .ZN(n14355) );
  NAND2_X1 U12837 ( .A1(n14781), .A2(n14782), .ZN(n14775) );
  NOR2_X1 U12838 ( .A1(n14402), .A2(n9807), .ZN(n14903) );
  NAND2_X1 U12839 ( .A1(n13345), .A2(n13306), .ZN(n14742) );
  NAND2_X1 U12840 ( .A1(n15657), .A2(n9866), .ZN(n12248) );
  AND4_X1 U12841 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n9757) );
  NAND2_X1 U12842 ( .A1(n9755), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9758) );
  OR3_X1 U12843 ( .A1(n12482), .A2(n14606), .A3(n16217), .ZN(n9759) );
  NAND2_X1 U12844 ( .A1(n10644), .A2(n11125), .ZN(n15241) );
  INV_X1 U12845 ( .A(n11522), .ZN(n10215) );
  OR2_X1 U12846 ( .A1(n9775), .A2(n16261), .ZN(n9760) );
  AND2_X1 U12847 ( .A1(n9725), .A2(n9895), .ZN(n9761) );
  BUF_X2 U12848 ( .A(n11517), .Z(n13893) );
  NAND2_X1 U12849 ( .A1(n11895), .A2(n11462), .ZN(n9762) );
  AND3_X1 U12850 ( .A1(n11552), .A2(n11551), .A3(n9992), .ZN(n9763) );
  OR2_X1 U12851 ( .A1(n14043), .A2(n14061), .ZN(n9764) );
  AND2_X1 U12852 ( .A1(n11844), .A2(n11839), .ZN(n9765) );
  INV_X1 U12853 ( .A(n16322), .ZN(n9944) );
  AND2_X1 U12854 ( .A1(n10640), .A2(n10181), .ZN(n9766) );
  AND4_X1 U12855 ( .A1(n16386), .A2(n16390), .A3(n16400), .A4(n16409), .ZN(
        n9767) );
  AND4_X1 U12856 ( .A1(n10806), .A2(n10805), .A3(n10804), .A4(n10803), .ZN(
        n9768) );
  AND2_X1 U12857 ( .A1(n17099), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9769) );
  AND4_X1 U12858 ( .A1(n10810), .A2(n10809), .A3(n10808), .A4(n10807), .ZN(
        n9770) );
  INV_X1 U12859 ( .A(n10669), .ZN(n16073) );
  INV_X1 U12860 ( .A(n18172), .ZN(n10143) );
  AND2_X1 U12861 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n9771) );
  OR2_X1 U12862 ( .A1(n14783), .A2(n10700), .ZN(n9772) );
  AND3_X1 U12863 ( .A1(n9765), .A2(n9860), .A3(n16260), .ZN(n9773) );
  AND2_X1 U12864 ( .A1(n10283), .A2(n9899), .ZN(n9774) );
  NOR2_X1 U12865 ( .A1(n11828), .A2(n16539), .ZN(n9775) );
  AND3_X1 U12866 ( .A1(n10200), .A2(n11173), .A3(n10199), .ZN(n9776) );
  NOR2_X1 U12867 ( .A1(n12433), .A2(n9911), .ZN(n16228) );
  OR2_X1 U12868 ( .A1(n14683), .A2(n15991), .ZN(n9777) );
  AND2_X1 U12869 ( .A1(n9756), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9778) );
  OR2_X1 U12870 ( .A1(n16355), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9779) );
  AND2_X1 U12871 ( .A1(n20103), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9780) );
  AND2_X1 U12872 ( .A1(n10597), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9781) );
  INV_X1 U12873 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16397) );
  AND4_X1 U12874 ( .A1(n13750), .A2(n13746), .A3(n13749), .A4(n13745), .ZN(
        n9782) );
  OR2_X1 U12875 ( .A1(n10914), .A2(n10913), .ZN(n10916) );
  AND2_X1 U12876 ( .A1(n12420), .A2(n12424), .ZN(n9783) );
  AND2_X1 U12877 ( .A1(n10714), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n9784) );
  INV_X1 U12878 ( .A(n12041), .ZN(n12039) );
  NAND2_X1 U12879 ( .A1(n10580), .A2(n11949), .ZN(n13959) );
  AND2_X1 U12880 ( .A1(n10334), .A2(n15628), .ZN(n9785) );
  AND2_X1 U12881 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9786) );
  AND2_X1 U12882 ( .A1(n10595), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9787) );
  AND2_X1 U12883 ( .A1(n9786), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9788) );
  INV_X1 U12884 ( .A(n10865), .ZN(n10281) );
  INV_X1 U12885 ( .A(n11671), .ZN(n10117) );
  NAND2_X1 U12886 ( .A1(n13852), .A2(n13851), .ZN(n19791) );
  INV_X1 U12887 ( .A(n19791), .ZN(n10239) );
  AND2_X1 U12888 ( .A1(n12234), .A2(n12233), .ZN(n15730) );
  NAND2_X1 U12889 ( .A1(n17606), .A2(n10686), .ZN(n9789) );
  AND2_X1 U12890 ( .A1(n12486), .A2(n11846), .ZN(n9790) );
  INV_X1 U12891 ( .A(n15994), .ZN(n10663) );
  NAND2_X1 U12892 ( .A1(n11234), .A2(n11233), .ZN(n13875) );
  AND2_X1 U12893 ( .A1(n10424), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n9791) );
  AND2_X1 U12894 ( .A1(n9791), .A2(n9910), .ZN(n9792) );
  INV_X1 U12895 ( .A(n20804), .ZN(n20749) );
  NAND2_X1 U12896 ( .A1(n10229), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9793) );
  INV_X1 U12897 ( .A(n10416), .ZN(n10415) );
  NAND2_X1 U12898 ( .A1(n9794), .A2(n10417), .ZN(n10416) );
  AND2_X1 U12899 ( .A1(n10708), .A2(n10709), .ZN(n9794) );
  INV_X1 U12900 ( .A(n16370), .ZN(n10339) );
  AND2_X1 U12901 ( .A1(n10148), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n9795) );
  AND2_X1 U12902 ( .A1(n10422), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n9796) );
  AND2_X1 U12903 ( .A1(n10636), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9797) );
  NAND2_X2 U12904 ( .A1(n13951), .A2(n12072), .ZN(n12090) );
  NAND2_X2 U12905 ( .A1(n10280), .A2(n11218), .ZN(n11235) );
  NAND2_X2 U12906 ( .A1(n17403), .A2(n13660), .ZN(n18285) );
  NOR2_X1 U12907 ( .A1(n14402), .A2(n10689), .ZN(n9798) );
  AND2_X2 U12908 ( .A1(n16789), .A2(n12642), .ZN(n11559) );
  NAND2_X1 U12909 ( .A1(n15815), .A2(n10578), .ZN(n12463) );
  NAND2_X2 U12910 ( .A1(n13912), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9799) );
  NAND2_X1 U12911 ( .A1(n15241), .A2(n15273), .ZN(n15243) );
  NAND2_X1 U12912 ( .A1(n13890), .A2(n12545), .ZN(n13938) );
  NOR2_X1 U12913 ( .A1(n14862), .A2(n13112), .ZN(n14853) );
  NAND2_X1 U12914 ( .A1(n10123), .A2(n10645), .ZN(n11831) );
  NAND2_X1 U12915 ( .A1(n11536), .A2(n11535), .ZN(n9800) );
  NOR2_X2 U12916 ( .A1(n13395), .A2(n15829), .ZN(n15815) );
  NOR2_X1 U12917 ( .A1(n12312), .A2(n10590), .ZN(n12314) );
  NAND2_X1 U12918 ( .A1(n14368), .A2(n10283), .ZN(n14889) );
  NOR2_X1 U12919 ( .A1(n16056), .A2(n10676), .ZN(n16026) );
  AND2_X1 U12920 ( .A1(n14105), .A2(n14122), .ZN(n14121) );
  NAND2_X1 U12921 ( .A1(n10863), .A2(n11152), .ZN(n11195) );
  NOR2_X1 U12922 ( .A1(n14783), .A2(n14784), .ZN(n14769) );
  NAND2_X1 U12923 ( .A1(n15667), .A2(n10586), .ZN(n12371) );
  AND2_X1 U12924 ( .A1(n18191), .A2(n10148), .ZN(n9802) );
  AND2_X1 U12925 ( .A1(n18191), .A2(P3_EBX_REG_22__SCAN_IN), .ZN(n9803) );
  AND2_X1 U12926 ( .A1(n10335), .A2(n15628), .ZN(n9804) );
  AND2_X1 U12927 ( .A1(n18532), .A2(n10422), .ZN(n9805) );
  NAND2_X1 U12928 ( .A1(n11845), .A2(n11846), .ZN(n9806) );
  OR2_X1 U12929 ( .A1(n10689), .A2(n13035), .ZN(n9807) );
  INV_X1 U12930 ( .A(n20237), .ZN(n20270) );
  INV_X1 U12931 ( .A(n12678), .ZN(n12712) );
  AND2_X1 U12932 ( .A1(n17127), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n9808) );
  NOR2_X1 U12933 ( .A1(n12308), .A2(n16466), .ZN(n12307) );
  AND2_X1 U12934 ( .A1(n10337), .A2(n10336), .ZN(n9809) );
  NAND2_X1 U12935 ( .A1(n15365), .A2(n11118), .ZN(n10644) );
  AND4_X1 U12936 ( .A1(n10815), .A2(n10814), .A3(n10813), .A4(n10812), .ZN(
        n9810) );
  OR2_X1 U12937 ( .A1(n14742), .A2(n15370), .ZN(n9811) );
  NOR3_X1 U12938 ( .A1(n14947), .A2(n14936), .A3(n13016), .ZN(n9812) );
  INV_X1 U12939 ( .A(n10262), .ZN(n11478) );
  AND2_X1 U12940 ( .A1(n10110), .A2(n10109), .ZN(n16000) );
  AND2_X1 U12941 ( .A1(n11930), .A2(n10382), .ZN(n9813) );
  AND2_X1 U12942 ( .A1(n11549), .A2(n10513), .ZN(n9814) );
  INV_X1 U12943 ( .A(n15977), .ZN(n10597) );
  AND2_X1 U12944 ( .A1(n12527), .A2(n11513), .ZN(n9815) );
  INV_X1 U12945 ( .A(n10441), .ZN(n10440) );
  NAND2_X1 U12946 ( .A1(n10521), .A2(n16365), .ZN(n10441) );
  NAND2_X1 U12947 ( .A1(n10477), .A2(n11821), .ZN(n16279) );
  AND2_X1 U12948 ( .A1(n10003), .A2(n10450), .ZN(n17518) );
  NAND2_X1 U12949 ( .A1(n17511), .A2(n11103), .ZN(n14457) );
  AND2_X1 U12950 ( .A1(n15216), .A2(n9797), .ZN(n9816) );
  OR2_X1 U12951 ( .A1(n11793), .A2(n10653), .ZN(n9817) );
  AND2_X1 U12952 ( .A1(n16215), .A2(n9759), .ZN(n9818) );
  OR2_X1 U12953 ( .A1(n16261), .A2(n10033), .ZN(n9819) );
  AND2_X1 U12954 ( .A1(n10251), .A2(n10252), .ZN(n9821) );
  NAND2_X1 U12955 ( .A1(n14121), .A2(n14335), .ZN(n14359) );
  NAND2_X1 U12956 ( .A1(n11663), .A2(n11678), .ZN(n11675) );
  NAND2_X1 U12957 ( .A1(n14863), .A2(n10695), .ZN(n14833) );
  NAND2_X1 U12958 ( .A1(n14682), .A2(n14681), .ZN(n16480) );
  NAND2_X1 U12959 ( .A1(n14368), .A2(n9774), .ZN(n9822) );
  AND4_X1 U12960 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n9823) );
  NAND2_X1 U12961 ( .A1(n9810), .A2(n9770), .ZN(n10553) );
  INV_X1 U12962 ( .A(n10553), .ZN(n10280) );
  AND2_X1 U12963 ( .A1(n11568), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n9824) );
  AND2_X2 U12964 ( .A1(n11430), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11637) );
  AND2_X1 U12965 ( .A1(n11932), .A2(n11939), .ZN(n9825) );
  NAND2_X2 U12966 ( .A1(n9935), .A2(n9934), .ZN(n12035) );
  AND2_X1 U12967 ( .A1(n16577), .A2(n17608), .ZN(n9826) );
  AND2_X1 U12968 ( .A1(n10404), .A2(n16273), .ZN(n9827) );
  OR2_X1 U12969 ( .A1(n14758), .A2(n10700), .ZN(n9828) );
  NAND2_X1 U12970 ( .A1(n14863), .A2(n10693), .ZN(n10697) );
  AND2_X1 U12971 ( .A1(n10576), .A2(n15753), .ZN(n9829) );
  INV_X1 U12972 ( .A(n11930), .ZN(n10388) );
  AND2_X1 U12973 ( .A1(n9995), .A2(n13529), .ZN(n9830) );
  AND2_X1 U12974 ( .A1(n11175), .A2(n11174), .ZN(n9831) );
  AND2_X1 U12975 ( .A1(n9996), .A2(n14141), .ZN(n9832) );
  INV_X2 U12976 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11535) );
  NOR2_X1 U12977 ( .A1(n10597), .A2(n9958), .ZN(n9833) );
  NOR2_X1 U12978 ( .A1(n10597), .A2(n9957), .ZN(n9834) );
  AND2_X1 U12979 ( .A1(n10465), .A2(n10463), .ZN(n9835) );
  NAND2_X1 U12980 ( .A1(n10530), .A2(n10531), .ZN(n9836) );
  INV_X1 U12981 ( .A(n10515), .ZN(n11933) );
  AND2_X1 U12982 ( .A1(n11892), .A2(n12386), .ZN(n9837) );
  INV_X1 U12983 ( .A(n16260), .ZN(n10033) );
  NOR2_X1 U12984 ( .A1(n9807), .A2(n10688), .ZN(n9838) );
  AND2_X1 U12985 ( .A1(n12440), .A2(n10574), .ZN(n9839) );
  AND2_X1 U12986 ( .A1(n15325), .A2(n15327), .ZN(n9840) );
  NOR2_X1 U12987 ( .A1(n11065), .A2(n11066), .ZN(n9841) );
  AND2_X1 U12988 ( .A1(n11514), .A2(n11512), .ZN(n12527) );
  INV_X1 U12989 ( .A(n12527), .ZN(n10204) );
  AND2_X1 U12990 ( .A1(n10597), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n9842) );
  AND2_X1 U12991 ( .A1(n16416), .A2(n16417), .ZN(n9843) );
  OR2_X1 U12992 ( .A1(n16236), .A2(n16256), .ZN(n9844) );
  INV_X1 U12993 ( .A(n14043), .ZN(n12142) );
  AND3_X1 U12994 ( .A1(n12141), .A2(n12140), .A3(n12139), .ZN(n14043) );
  AND2_X1 U12995 ( .A1(n9811), .A2(n13317), .ZN(n9845) );
  AND2_X1 U12996 ( .A1(n15672), .A2(n12243), .ZN(n15657) );
  AND2_X1 U12997 ( .A1(n13988), .A2(n10184), .ZN(n9846) );
  AND2_X1 U12998 ( .A1(n11074), .A2(n11050), .ZN(n9847) );
  NAND2_X1 U12999 ( .A1(n12440), .A2(n10572), .ZN(n15675) );
  INV_X1 U13000 ( .A(n16745), .ZN(n16743) );
  AND2_X1 U13001 ( .A1(n10128), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16745) );
  AND2_X1 U13002 ( .A1(n14458), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9848) );
  OR2_X1 U13003 ( .A1(n11694), .A2(n10651), .ZN(n9849) );
  INV_X1 U13004 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12321) );
  INV_X1 U13005 ( .A(n10525), .ZN(n10524) );
  OAI21_X1 U13006 ( .B1(n12414), .B2(n12416), .A(n16374), .ZN(n10525) );
  OR2_X1 U13007 ( .A1(n14724), .A2(n14723), .ZN(n14741) );
  NAND2_X1 U13008 ( .A1(n12232), .A2(n12231), .ZN(n15729) );
  AND2_X1 U13009 ( .A1(n13827), .A2(n10492), .ZN(n9850) );
  INV_X1 U13010 ( .A(n10876), .ZN(n10895) );
  INV_X1 U13011 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16437) );
  NAND2_X1 U13012 ( .A1(n12232), .A2(n10602), .ZN(n12437) );
  AND2_X1 U13013 ( .A1(n13752), .A2(n13744), .ZN(n9851) );
  NOR2_X1 U13014 ( .A1(n11517), .A2(n16787), .ZN(n9852) );
  OR2_X1 U13015 ( .A1(n17325), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9853) );
  AND3_X1 U13016 ( .A1(n12507), .A2(n12506), .A3(n10632), .ZN(n9854) );
  NOR2_X1 U13017 ( .A1(n10563), .A2(n10562), .ZN(n9855) );
  AND2_X1 U13018 ( .A1(n12432), .A2(n16470), .ZN(n9856) );
  INV_X1 U13019 ( .A(n10120), .ZN(n11765) );
  OR2_X1 U13020 ( .A1(n11793), .A2(n10121), .ZN(n10120) );
  AND2_X1 U13021 ( .A1(n20113), .A2(n16873), .ZN(n9857) );
  INV_X1 U13022 ( .A(n11939), .ZN(n10516) );
  NAND2_X1 U13023 ( .A1(n11023), .A2(n10974), .ZN(n9858) );
  INV_X1 U13024 ( .A(n10000), .ZN(n15612) );
  NOR3_X1 U13025 ( .A1(n15678), .A2(n15665), .A3(n9864), .ZN(n10000) );
  AND2_X1 U13026 ( .A1(n16745), .A2(n10388), .ZN(n9859) );
  NAND2_X1 U13027 ( .A1(n14601), .A2(n12485), .ZN(n9860) );
  AND2_X1 U13028 ( .A1(n9809), .A2(n16370), .ZN(n9861) );
  INV_X1 U13029 ( .A(n10551), .ZN(n10448) );
  NOR2_X1 U13030 ( .A1(n10447), .A2(n9913), .ZN(n10551) );
  INV_X1 U13031 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13659) );
  NAND2_X1 U13032 ( .A1(n10972), .A2(n11015), .ZN(n9862) );
  AOI21_X1 U13033 ( .B1(n14621), .B2(n20808), .A(n10591), .ZN(n12347) );
  INV_X1 U13034 ( .A(n12077), .ZN(n12196) );
  INV_X1 U13035 ( .A(n17559), .ZN(n20999) );
  NAND2_X1 U13036 ( .A1(n18814), .A2(n10726), .ZN(n17733) );
  INV_X1 U13037 ( .A(n11530), .ZN(n12641) );
  INV_X1 U13038 ( .A(n11707), .ZN(n14606) );
  INV_X1 U13039 ( .A(n12538), .ZN(n10106) );
  OAI21_X1 U13040 ( .B1(n16954), .B2(n16953), .A(n19938), .ZN(n16973) );
  NOR2_X1 U13041 ( .A1(n13392), .A2(n13393), .ZN(n13391) );
  AND2_X1 U13042 ( .A1(n13938), .A2(n10111), .ZN(n16066) );
  NAND2_X1 U13043 ( .A1(n13938), .A2(n12551), .ZN(n14143) );
  OR2_X1 U13044 ( .A1(n16061), .A2(n16062), .ZN(n16056) );
  OR2_X1 U13045 ( .A1(n16056), .A2(n10677), .ZN(n9863) );
  INV_X1 U13046 ( .A(n17602), .ZN(n10442) );
  NAND2_X1 U13047 ( .A1(n11676), .A2(n10116), .ZN(n11694) );
  NAND2_X1 U13048 ( .A1(n14068), .A2(n14339), .ZN(n14219) );
  NAND2_X1 U13049 ( .A1(n14035), .A2(n9832), .ZN(n13396) );
  NAND2_X1 U13050 ( .A1(n12334), .A2(n9786), .ZN(n12336) );
  NAND2_X1 U13051 ( .A1(n10586), .A2(n10585), .ZN(n9864) );
  NAND3_X1 U13052 ( .A1(n16421), .A2(n11734), .A3(n16432), .ZN(n9865) );
  NOR2_X1 U13053 ( .A1(n14042), .A2(n9764), .ZN(n14052) );
  AND2_X1 U13054 ( .A1(n14035), .A2(n9996), .ZN(n14140) );
  NOR2_X1 U13055 ( .A1(n15019), .A2(n15020), .ZN(n14998) );
  NAND2_X1 U13056 ( .A1(n10580), .A2(n10579), .ZN(n14066) );
  AND2_X1 U13057 ( .A1(n15815), .A2(n10576), .ZN(n15752) );
  NAND2_X1 U13058 ( .A1(n14075), .A2(n12097), .ZN(n14317) );
  NAND2_X1 U13059 ( .A1(n10598), .A2(n12142), .ZN(n14041) );
  INV_X1 U13060 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20786) );
  NOR2_X1 U13061 ( .A1(n14219), .A2(n14220), .ZN(n14035) );
  AND2_X1 U13062 ( .A1(n15645), .A2(n15659), .ZN(n9866) );
  OR2_X1 U13063 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n9867) );
  AND2_X1 U13064 ( .A1(n12342), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12341) );
  NOR2_X1 U13065 ( .A1(n12312), .A2(n10587), .ZN(n12317) );
  AND2_X1 U13066 ( .A1(n12358), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12357) );
  AND2_X1 U13067 ( .A1(n12334), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12333) );
  MUX2_X1 U13068 ( .A(n11880), .B(n15955), .S(n12290), .Z(n11682) );
  NOR2_X1 U13069 ( .A1(n13942), .A2(n9998), .ZN(n14068) );
  AND2_X1 U13070 ( .A1(n14998), .A2(n14999), .ZN(n14982) );
  NAND2_X1 U13071 ( .A1(n14035), .A2(n11965), .ZN(n14034) );
  AND2_X1 U13072 ( .A1(n11591), .A2(n11546), .ZN(n9868) );
  OR2_X1 U13073 ( .A1(n20127), .A2(n11762), .ZN(n9869) );
  INV_X1 U13074 ( .A(n13372), .ZN(n10254) );
  AND2_X1 U13075 ( .A1(n14729), .A2(n11217), .ZN(n13621) );
  AND2_X1 U13076 ( .A1(n13809), .A2(n13818), .ZN(n9870) );
  INV_X1 U13077 ( .A(n10735), .ZN(n11121) );
  OR2_X1 U13078 ( .A1(n18825), .A2(n18837), .ZN(n9871) );
  OR2_X1 U13079 ( .A1(n11712), .A2(n12290), .ZN(n11843) );
  INV_X1 U13080 ( .A(n11843), .ZN(n10647) );
  AND2_X1 U13081 ( .A1(n12290), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U13082 ( .A1(n11286), .A2(n11285), .ZN(n14891) );
  OAI21_X1 U13083 ( .B1(n12867), .B2(n13014), .A(n12866), .ZN(n14122) );
  NAND2_X1 U13084 ( .A1(n10318), .A2(n15694), .ZN(n15680) );
  OR2_X1 U13085 ( .A1(n14143), .A2(n14350), .ZN(n14351) );
  NAND2_X1 U13086 ( .A1(n12819), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13014) );
  INV_X1 U13087 ( .A(n13014), .ZN(n12993) );
  AND2_X1 U13088 ( .A1(n10619), .A2(n10618), .ZN(n9873) );
  AND3_X1 U13089 ( .A1(n16929), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n20026) );
  NOR2_X1 U13090 ( .A1(n11841), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15650) );
  INV_X1 U13091 ( .A(n12441), .ZN(n12001) );
  OR2_X1 U13092 ( .A1(n14306), .A2(n20825), .ZN(n10981) );
  XOR2_X1 U13093 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .Z(n9874) );
  INV_X1 U13094 ( .A(n12424), .ZN(n10611) );
  INV_X1 U13095 ( .A(n19237), .ZN(n19226) );
  AND2_X1 U13096 ( .A1(n13896), .A2(n10230), .ZN(n19237) );
  NAND2_X1 U13097 ( .A1(n17213), .A2(n10502), .ZN(n10503) );
  INV_X1 U13098 ( .A(n14906), .ZN(n11285) );
  AND2_X1 U13099 ( .A1(n10494), .A2(n17742), .ZN(n9875) );
  AND2_X1 U13100 ( .A1(n10111), .A2(n16067), .ZN(n9876) );
  AND2_X1 U13101 ( .A1(n11692), .A2(n9976), .ZN(n9877) );
  OR2_X1 U13102 ( .A1(n17606), .A2(n14664), .ZN(n9878) );
  AND2_X1 U13103 ( .A1(n11757), .A2(n11754), .ZN(n9879) );
  OR2_X1 U13104 ( .A1(n14143), .A2(n10673), .ZN(n10669) );
  AND2_X1 U13105 ( .A1(n18299), .A2(n10147), .ZN(n9880) );
  INV_X1 U13106 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18843) );
  INV_X1 U13107 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16379) );
  OR2_X1 U13108 ( .A1(n18495), .A2(n18122), .ZN(n9881) );
  AND2_X1 U13109 ( .A1(n12230), .A2(n12229), .ZN(n15751) );
  INV_X1 U13110 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20808) );
  INV_X1 U13111 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18110) );
  INV_X1 U13112 ( .A(n10672), .ZN(n16085) );
  OR2_X1 U13113 ( .A1(n14143), .A2(n10674), .ZN(n10672) );
  NAND2_X1 U13114 ( .A1(n10115), .A2(n11663), .ZN(n9882) );
  INV_X1 U13115 ( .A(n16394), .ZN(n10173) );
  NOR2_X1 U13116 ( .A1(n11704), .A2(n11703), .ZN(n12109) );
  AND2_X1 U13117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9883) );
  AND2_X1 U13118 ( .A1(n10540), .A2(n10543), .ZN(n9884) );
  NOR2_X1 U13119 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9885) );
  AND2_X1 U13120 ( .A1(n10602), .A2(n10601), .ZN(n9886) );
  AND2_X1 U13121 ( .A1(n10569), .A2(n14866), .ZN(n9887) );
  INV_X1 U13122 ( .A(n16312), .ZN(n10365) );
  AND2_X1 U13124 ( .A1(n10615), .A2(n10614), .ZN(n9888) );
  AND2_X1 U13125 ( .A1(n9787), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9889) );
  AND2_X1 U13126 ( .A1(n9788), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9890) );
  AND2_X1 U13127 ( .A1(n17732), .A2(n10497), .ZN(n9891) );
  AND2_X1 U13128 ( .A1(n9868), .A2(n11918), .ZN(n9892) );
  AND2_X1 U13129 ( .A1(n10164), .A2(n17587), .ZN(n9893) );
  INV_X1 U13130 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14004) );
  AND2_X1 U13131 ( .A1(n12406), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16847)
         );
  NAND2_X1 U13132 ( .A1(n17503), .A2(n13311), .ZN(n20829) );
  INV_X1 U13133 ( .A(n20829), .ZN(n17531) );
  INV_X1 U13134 ( .A(n19785), .ZN(n10238) );
  AND3_X1 U13135 ( .A1(n11234), .A2(n11233), .A3(n10555), .ZN(n14101) );
  OR2_X1 U13136 ( .A1(n17333), .A2(n17330), .ZN(n18830) );
  INV_X1 U13137 ( .A(n18830), .ZN(n18910) );
  AND2_X1 U13138 ( .A1(n10567), .A2(n10566), .ZN(n9894) );
  OR2_X1 U13139 ( .A1(n11602), .A2(n11601), .ZN(n11918) );
  AND2_X1 U13140 ( .A1(n12266), .A2(n16029), .ZN(n16470) );
  AND2_X1 U13141 ( .A1(n10144), .A2(n17457), .ZN(n9895) );
  INV_X1 U13142 ( .A(n16266), .ZN(n10316) );
  XNOR2_X1 U13143 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n16456), .ZN(
        n9896) );
  OR2_X1 U13144 ( .A1(n18055), .A2(n17752), .ZN(n9897) );
  AND2_X1 U13145 ( .A1(n14964), .A2(n14962), .ZN(n9898) );
  NAND2_X1 U13146 ( .A1(n20808), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16839) );
  AND2_X1 U13147 ( .A1(n13072), .A2(n13071), .ZN(n9899) );
  INV_X1 U13148 ( .A(n9969), .ZN(n13951) );
  NAND2_X1 U13149 ( .A1(n9720), .A2(n16873), .ZN(n9969) );
  INV_X1 U13150 ( .A(n16230), .ZN(n10334) );
  NAND3_X1 U13151 ( .A1(n18600), .A2(P3_EAX_REG_11__SCAN_IN), .A3(
        P3_EAX_REG_12__SCAN_IN), .ZN(n9900) );
  INV_X1 U13152 ( .A(n10668), .ZN(n10667) );
  NAND2_X1 U13153 ( .A1(n16008), .A2(n12767), .ZN(n10668) );
  INV_X1 U13154 ( .A(n14606), .ZN(n10382) );
  OR2_X1 U13155 ( .A1(n17082), .A2(n18907), .ZN(n9901) );
  NAND3_X1 U13156 ( .A1(n15491), .A2(n21704), .A3(n11281), .ZN(n9902) );
  AND2_X1 U13157 ( .A1(n10498), .A2(n17742), .ZN(n9903) );
  AND2_X1 U13158 ( .A1(n9894), .A2(n10565), .ZN(n9904) );
  AND2_X1 U13159 ( .A1(n9790), .A2(n12478), .ZN(n9905) );
  INV_X1 U13160 ( .A(n14337), .ZN(n11252) );
  AND2_X1 U13161 ( .A1(n11251), .A2(n11250), .ZN(n14337) );
  NOR2_X1 U13162 ( .A1(n21294), .A2(n21136), .ZN(n9906) );
  NOR2_X1 U13163 ( .A1(n21294), .A2(n21408), .ZN(n9907) );
  AND2_X1 U13164 ( .A1(n13664), .A2(n13665), .ZN(n18193) );
  INV_X1 U13165 ( .A(n18193), .ZN(n13705) );
  INV_X1 U13166 ( .A(n19213), .ZN(n10312) );
  INV_X1 U13167 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10209) );
  INV_X1 U13168 ( .A(n14350), .ZN(n10675) );
  AND2_X1 U13169 ( .A1(n17100), .A2(n9769), .ZN(n9908) );
  OR2_X1 U13170 ( .A1(n21805), .A2(n12434), .ZN(n9909) );
  NOR2_X1 U13171 ( .A1(n18989), .A2(n18990), .ZN(n17261) );
  INV_X1 U13172 ( .A(n16485), .ZN(n10417) );
  INV_X1 U13173 ( .A(n12062), .ZN(n10710) );
  AND2_X1 U13174 ( .A1(n10725), .A2(P3_EAX_REG_19__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U13175 ( .A1(n15863), .A2(n9809), .ZN(n10340) );
  NAND2_X1 U13176 ( .A1(n10380), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9911) );
  NAND2_X1 U13177 ( .A1(n10341), .A2(n15938), .ZN(n10345) );
  AND2_X1 U13178 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U13179 ( .A1(n11127), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9913) );
  OR2_X1 U13180 ( .A1(n10685), .A2(n12416), .ZN(n9914) );
  NOR2_X1 U13181 ( .A1(n16614), .A2(n16356), .ZN(n9915) );
  INV_X1 U13182 ( .A(n16567), .ZN(n10706) );
  AND2_X1 U13183 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9916) );
  NOR2_X1 U13184 ( .A1(n15242), .A2(n10641), .ZN(n9917) );
  AND2_X1 U13185 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9918) );
  INV_X1 U13186 ( .A(n10686), .ZN(n10293) );
  AND2_X1 U13187 ( .A1(n9915), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10686) );
  NOR2_X1 U13188 ( .A1(n10707), .A2(n16556), .ZN(n9919) );
  INV_X1 U13189 ( .A(n11372), .ZN(n10636) );
  INV_X1 U13190 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10643) );
  INV_X1 U13191 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10061) );
  INV_X1 U13192 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10542) );
  INV_X1 U13193 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n10425) );
  INV_X1 U13194 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10642) );
  INV_X1 U13195 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10596) );
  INV_X1 U13196 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20800) );
  INV_X1 U13197 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13570) );
  INV_X1 U13198 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n10423) );
  INV_X1 U13199 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n10149) );
  INV_X1 U13200 ( .A(n10320), .ZN(n15965) );
  OR2_X1 U13201 ( .A1(n16778), .A2(n15963), .ZN(n10320) );
  INV_X1 U13202 ( .A(n12452), .ZN(n10396) );
  INV_X1 U13203 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10649) );
  INV_X1 U13204 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10220) );
  AND2_X1 U13205 ( .A1(n20800), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n9920) );
  AOI22_X1 U13206 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20133), .ZN(n9921) );
  NOR2_X2 U13207 ( .A1(n16849), .A2(n16848), .ZN(n20134) );
  NOR2_X2 U13208 ( .A1(n16847), .A2(n16848), .ZN(n20133) );
  INV_X1 U13209 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19923) );
  NOR4_X2 U13210 ( .A1(n17719), .A2(n17718), .A3(n17717), .A4(n17716), .ZN(
        n19928) );
  NOR3_X2 U13211 ( .A1(n19688), .A2(n19806), .A3(n19475), .ZN(n19446) );
  NAND3_X2 U13212 ( .A1(n9924), .A2(n10361), .A3(n9922), .ZN(n11517) );
  INV_X1 U13213 ( .A(n11507), .ZN(n9923) );
  NAND2_X1 U13214 ( .A1(n9925), .A2(n11507), .ZN(n9924) );
  INV_X1 U13215 ( .A(n10480), .ZN(n9925) );
  NAND4_X1 U13216 ( .A1(n11614), .A2(n11613), .A3(n11611), .A4(n11612), .ZN(
        n9928) );
  NAND4_X1 U13217 ( .A1(n11390), .A2(n11389), .A3(n11391), .A4(n11388), .ZN(
        n9930) );
  NAND2_X1 U13218 ( .A1(n9823), .A2(n9951), .ZN(n9931) );
  NAND2_X2 U13219 ( .A1(n9933), .A2(n9932), .ZN(n11455) );
  NAND4_X1 U13220 ( .A1(n11438), .A2(n11436), .A3(n11437), .A4(n11435), .ZN(
        n9934) );
  NAND4_X1 U13221 ( .A1(n11443), .A2(n11441), .A3(n11442), .A4(n11444), .ZN(
        n9935) );
  NAND2_X2 U13222 ( .A1(n9937), .A2(n9936), .ZN(n20118) );
  OAI21_X1 U13223 ( .B1(n9947), .B2(n9948), .A(n11535), .ZN(n9936) );
  NAND3_X1 U13224 ( .A1(n9939), .A2(n13529), .A3(n9995), .ZN(n9938) );
  NAND2_X2 U13225 ( .A1(n11475), .A2(n10038), .ZN(n13529) );
  XNOR2_X2 U13226 ( .A(n10407), .B(n9941), .ZN(n10128) );
  AND3_X2 U13227 ( .A1(n10703), .A2(n9892), .A3(n9968), .ZN(n10407) );
  NAND2_X1 U13228 ( .A1(n9945), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12473) );
  NAND3_X1 U13229 ( .A1(n11379), .A2(n11381), .A3(n11378), .ZN(n9947) );
  INV_X1 U13230 ( .A(n11380), .ZN(n9948) );
  NAND3_X1 U13231 ( .A1(n11383), .A2(n11382), .A3(n11385), .ZN(n9949) );
  NAND2_X1 U13232 ( .A1(n10262), .A2(n10714), .ZN(n11502) );
  NAND2_X1 U13233 ( .A1(n11916), .A2(n11915), .ZN(n9960) );
  INV_X1 U13234 ( .A(n9961), .ZN(n11868) );
  NAND2_X1 U13235 ( .A1(n11654), .A2(n9961), .ZN(n11880) );
  NAND2_X1 U13236 ( .A1(n10262), .A2(n9784), .ZN(n9962) );
  AND3_X2 U13237 ( .A1(n9963), .A2(n10078), .A3(n9962), .ZN(n10359) );
  NAND2_X1 U13238 ( .A1(n11492), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9963) );
  NOR2_X2 U13239 ( .A1(n16716), .A2(n12056), .ZN(n16687) );
  NOR2_X2 U13240 ( .A1(n14321), .A2(n14325), .ZN(n16766) );
  NAND2_X1 U13241 ( .A1(n16495), .A2(n17606), .ZN(n10133) );
  AND2_X2 U13242 ( .A1(n9966), .A2(n9965), .ZN(n16495) );
  NAND2_X1 U13243 ( .A1(n9967), .A2(n16490), .ZN(n9966) );
  NAND2_X1 U13244 ( .A1(n16228), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9967) );
  NAND2_X1 U13245 ( .A1(n9968), .A2(n11546), .ZN(n10137) );
  NAND3_X1 U13246 ( .A1(n10703), .A2(n9968), .A3(n9868), .ZN(n10214) );
  NAND4_X1 U13247 ( .A1(n11465), .A2(n11892), .A3(n11655), .A4(n9970), .ZN(
        n9995) );
  XNOR2_X2 U13248 ( .A(n11508), .B(n9971), .ZN(n11522) );
  NOR2_X1 U13249 ( .A1(n16692), .A2(n9974), .ZN(n16694) );
  NAND2_X1 U13250 ( .A1(n10275), .A2(n15943), .ZN(n9979) );
  XNOR2_X2 U13251 ( .A(n10136), .B(n10137), .ZN(n10275) );
  NAND3_X1 U13252 ( .A1(n12419), .A2(n16341), .A3(n12420), .ZN(n14695) );
  NAND2_X1 U13253 ( .A1(n10139), .A2(n9981), .ZN(n16364) );
  NAND2_X1 U13254 ( .A1(n9983), .A2(n14706), .ZN(n9982) );
  INV_X1 U13255 ( .A(n10682), .ZN(n9984) );
  NAND3_X1 U13256 ( .A1(n11484), .A2(n11483), .A3(n11490), .ZN(n11511) );
  NAND2_X1 U13257 ( .A1(n11489), .A2(n11488), .ZN(n10212) );
  XNOR2_X2 U13258 ( .A(n10359), .B(n10360), .ZN(n11513) );
  AND3_X2 U13259 ( .A1(n13893), .A2(n15977), .A3(n11520), .ZN(n20249) );
  AND3_X2 U13260 ( .A1(n13893), .A2(n16787), .A3(n11520), .ZN(n16837) );
  INV_X1 U13261 ( .A(n16837), .ZN(n11719) );
  INV_X1 U13262 ( .A(n20249), .ZN(n11720) );
  NAND3_X1 U13263 ( .A1(n9990), .A2(n9989), .A3(n9988), .ZN(n9987) );
  NAND2_X1 U13264 ( .A1(n16837), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n9988) );
  NAND2_X1 U13265 ( .A1(n20249), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n9989) );
  NAND2_X1 U13266 ( .A1(n9801), .A2(n20800), .ZN(n9994) );
  NOR2_X2 U13267 ( .A1(n12433), .A2(n9793), .ZN(n16270) );
  NAND2_X2 U13268 ( .A1(n10099), .A2(n10411), .ZN(n12433) );
  NAND3_X1 U13269 ( .A1(n10003), .A2(n17520), .A3(n10450), .ZN(n10298) );
  NAND3_X1 U13270 ( .A1(n9847), .A2(n11052), .A3(n11051), .ZN(n10003) );
  NAND2_X1 U13271 ( .A1(n12832), .A2(n12831), .ZN(n10004) );
  NAND3_X1 U13272 ( .A1(n21037), .A2(n20825), .A3(n10971), .ZN(n10007) );
  NAND2_X2 U13273 ( .A1(n10244), .A2(n10243), .ZN(n10971) );
  NAND2_X1 U13274 ( .A1(n10970), .A2(n10314), .ZN(n21037) );
  INV_X1 U13275 ( .A(n10009), .ZN(n11049) );
  AOI21_X1 U13276 ( .B1(n14201), .B2(n10009), .A(n10008), .ZN(n14204) );
  AND2_X1 U13277 ( .A1(n14200), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10008) );
  XNOR2_X1 U13278 ( .A(n14201), .B(n10009), .ZN(n14269) );
  NAND2_X2 U13279 ( .A1(n10250), .A2(n10377), .ZN(n15365) );
  NOR2_X1 U13280 ( .A1(n10266), .A2(n10021), .ZN(n10015) );
  AND2_X1 U13281 ( .A1(n10022), .A2(n10016), .ZN(n20495) );
  NAND2_X1 U13282 ( .A1(n10019), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10018) );
  NAND3_X1 U13283 ( .A1(n10026), .A2(n11647), .A3(n10024), .ZN(n11707) );
  NAND3_X1 U13284 ( .A1(n11629), .A2(n11636), .A3(n10029), .ZN(n10028) );
  AND2_X2 U13285 ( .A1(n12642), .A2(n16788), .ZN(n12632) );
  NAND3_X1 U13286 ( .A1(n9827), .A2(n11753), .A3(n11752), .ZN(n10150) );
  NAND4_X1 U13287 ( .A1(n9827), .A2(n11753), .A3(n11752), .A4(n16260), .ZN(
        n10032) );
  NAND2_X2 U13288 ( .A1(n16387), .A2(n10367), .ZN(n11753) );
  NAND2_X2 U13289 ( .A1(n11755), .A2(n9879), .ZN(n11793) );
  INV_X4 U13290 ( .A(n11456), .ZN(n16887) );
  INV_X1 U13291 ( .A(n16228), .ZN(n10151) );
  XNOR2_X1 U13292 ( .A(n10535), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13849) );
  NAND2_X4 U13293 ( .A1(n10053), .A2(n10052), .ZN(n10535) );
  NAND2_X2 U13294 ( .A1(n13665), .A2(n13666), .ZN(n18301) );
  INV_X2 U13295 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n17414) );
  NAND3_X1 U13296 ( .A1(n10540), .A2(n19143), .A3(n10543), .ZN(n10060) );
  INV_X2 U13297 ( .A(n11517), .ZN(n10225) );
  NOR2_X1 U13298 ( .A1(n12041), .A2(n20808), .ZN(n10047) );
  NAND2_X1 U13299 ( .A1(n9837), .A2(n12039), .ZN(n16799) );
  NAND2_X1 U13300 ( .A1(n10048), .A2(n15918), .ZN(n10050) );
  AND4_X2 U13301 ( .A1(n13841), .A2(n13846), .A3(n13848), .A4(n13842), .ZN(
        n10052) );
  AND4_X2 U13302 ( .A1(n13845), .A2(n13844), .A3(n13847), .A4(n13843), .ZN(
        n10053) );
  OR2_X2 U13303 ( .A1(n13836), .A2(n13837), .ZN(n17127) );
  NAND2_X1 U13304 ( .A1(n19018), .A2(n17062), .ZN(n17067) );
  OAI21_X1 U13305 ( .B1(n19035), .B2(n17056), .A(n10055), .ZN(n10058) );
  INV_X1 U13306 ( .A(n17053), .ZN(n10056) );
  NAND2_X1 U13307 ( .A1(n10059), .A2(n17057), .ZN(n17058) );
  NAND2_X1 U13308 ( .A1(n19035), .A2(n17053), .ZN(n10059) );
  NAND2_X2 U13309 ( .A1(n10060), .A2(n18830), .ZN(n18792) );
  NAND3_X1 U13310 ( .A1(n10066), .A2(n14121), .A3(n14335), .ZN(n14360) );
  NAND2_X2 U13311 ( .A1(n10068), .A2(n11683), .ZN(n20810) );
  INV_X1 U13312 ( .A(n11465), .ZN(n10068) );
  AND2_X2 U13313 ( .A1(n10407), .A2(n10408), .ZN(n11731) );
  NAND3_X1 U13314 ( .A1(n10069), .A2(n11503), .A3(n11504), .ZN(n11943) );
  OAI21_X1 U13315 ( .B1(n12261), .B2(n10070), .A(n12260), .ZN(P2_U3019) );
  AND2_X1 U13316 ( .A1(n20801), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10079) );
  INV_X1 U13317 ( .A(n10085), .ZN(n10257) );
  INV_X1 U13318 ( .A(n14696), .ZN(n12421) );
  NAND2_X1 U13319 ( .A1(n10091), .A2(n10089), .ZN(n16449) );
  NAND2_X1 U13320 ( .A1(n10702), .A2(n10090), .ZN(n10089) );
  INV_X1 U13321 ( .A(n10138), .ZN(n10090) );
  AOI21_X1 U13322 ( .B1(n10138), .B2(n10092), .A(n9859), .ZN(n10091) );
  INV_X1 U13323 ( .A(n11931), .ZN(n10092) );
  NOR2_X2 U13324 ( .A1(n16744), .A2(n10261), .ZN(n10138) );
  NAND2_X2 U13325 ( .A1(n16449), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16451) );
  OAI21_X2 U13326 ( .B1(n10275), .B2(n14315), .A(n11927), .ZN(n11928) );
  NOR2_X1 U13327 ( .A1(n10128), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10261) );
  OAI21_X2 U13328 ( .B1(n11928), .B2(n10096), .A(n10213), .ZN(n16744) );
  NAND2_X1 U13329 ( .A1(n16298), .A2(n21805), .ZN(n10098) );
  NAND2_X1 U13330 ( .A1(n10098), .A2(n10097), .ZN(n12451) );
  NAND2_X1 U13331 ( .A1(n10098), .A2(n9856), .ZN(n12515) );
  NAND2_X1 U13332 ( .A1(n10099), .A2(n10481), .ZN(n16304) );
  NAND2_X1 U13333 ( .A1(n10099), .A2(n9919), .ZN(n10227) );
  NAND2_X2 U13334 ( .A1(n16451), .A2(n9825), .ZN(n10099) );
  AND3_X2 U13335 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11530) );
  INV_X1 U13336 ( .A(n10102), .ZN(n10101) );
  NAND2_X1 U13337 ( .A1(n10102), .A2(n15994), .ZN(n15995) );
  OR2_X1 U13338 ( .A1(n13893), .A2(n16839), .ZN(n10107) );
  NOR2_X2 U13339 ( .A1(n16000), .A2(n10108), .ZN(n16006) );
  NAND2_X1 U13340 ( .A1(n12290), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10118) );
  INV_X1 U13341 ( .A(n10126), .ZN(n11545) );
  NAND2_X1 U13342 ( .A1(n10126), .A2(n12386), .ZN(n10125) );
  AOI22_X1 U13343 ( .A1(n12207), .A2(n10126), .B1(n12283), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n12104) );
  NAND3_X1 U13344 ( .A1(n12510), .A2(n9854), .A3(n10127), .ZN(P2_U3015) );
  NAND3_X1 U13345 ( .A1(n12500), .A2(n10631), .A3(n12499), .ZN(n10127) );
  AND2_X2 U13346 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11910) );
  NAND2_X1 U13347 ( .A1(n10128), .A2(n14606), .ZN(n11673) );
  AND2_X4 U13348 ( .A1(n11910), .A2(n16905), .ZN(n11536) );
  NAND2_X1 U13349 ( .A1(n10138), .A2(n16743), .ZN(n16747) );
  NAND2_X1 U13350 ( .A1(n10152), .A2(n10153), .ZN(n10460) );
  NAND3_X1 U13351 ( .A1(n14013), .A2(n10242), .A3(n20825), .ZN(n10152) );
  NAND2_X1 U13352 ( .A1(n10154), .A2(n15536), .ZN(n15327) );
  NAND2_X1 U13353 ( .A1(n10154), .A2(n11114), .ZN(n15325) );
  NAND2_X1 U13354 ( .A1(n10154), .A2(n15524), .ZN(n10179) );
  NAND2_X1 U13355 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U13356 ( .A1(n10154), .A2(n11349), .ZN(n11126) );
  NAND2_X1 U13357 ( .A1(n10154), .A2(n21704), .ZN(n15305) );
  NOR2_X1 U13358 ( .A1(n10735), .A2(n9916), .ZN(n10728) );
  NAND2_X1 U13359 ( .A1(n10154), .A2(n15399), .ZN(n15197) );
  INV_X4 U13360 ( .A(n10735), .ZN(n10154) );
  NOR2_X1 U13361 ( .A1(n10735), .A2(n15556), .ZN(n10155) );
  NAND3_X1 U13362 ( .A1(n11118), .A2(n10551), .A3(n15365), .ZN(n10156) );
  NAND2_X2 U13363 ( .A1(n10159), .A2(n10158), .ZN(n11107) );
  NOR2_X2 U13364 ( .A1(n10160), .A2(n10742), .ZN(n10159) );
  NAND3_X1 U13365 ( .A1(n10167), .A2(n9893), .A3(n10163), .ZN(n10172) );
  NAND2_X1 U13366 ( .A1(n16410), .A2(n10161), .ZN(n10167) );
  AND2_X1 U13367 ( .A1(n10163), .A2(n10164), .ZN(n10162) );
  INV_X1 U13368 ( .A(n16409), .ZN(n10171) );
  OAI211_X1 U13369 ( .C1(n16655), .C2(n17594), .A(n10172), .B(n10384), .ZN(
        P2_U3003) );
  INV_X1 U13370 ( .A(n10175), .ZN(n10174) );
  OAI21_X1 U13371 ( .B1(n11125), .B2(n10448), .A(n10154), .ZN(n10175) );
  NAND2_X1 U13372 ( .A1(n10296), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U13373 ( .A1(n10177), .A2(n15602), .ZN(n10903) );
  NAND2_X1 U13374 ( .A1(n10177), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10355) );
  NAND2_X1 U13375 ( .A1(n10177), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10979) );
  NAND2_X2 U13376 ( .A1(n10180), .A2(n10992), .ZN(n14114) );
  NAND3_X1 U13377 ( .A1(n9766), .A2(n15190), .A3(n9885), .ZN(n10729) );
  NAND2_X1 U13378 ( .A1(n15174), .A2(n15399), .ZN(n10638) );
  NAND2_X2 U13379 ( .A1(n10182), .A2(n10638), .ZN(n15190) );
  NAND3_X1 U13380 ( .A1(n10193), .A2(n11935), .A3(n10192), .ZN(n11938) );
  NAND2_X1 U13381 ( .A1(n11170), .A2(n10201), .ZN(n10197) );
  NAND2_X1 U13382 ( .A1(n10197), .A2(n10198), .ZN(n11177) );
  NOR2_X2 U13383 ( .A1(n12432), .A2(n10416), .ZN(n16229) );
  NAND2_X1 U13384 ( .A1(n11928), .A2(n10203), .ZN(n16461) );
  NAND2_X1 U13385 ( .A1(n10211), .A2(n10210), .ZN(n11512) );
  INV_X1 U13386 ( .A(n11511), .ZN(n10210) );
  INV_X1 U13387 ( .A(n10212), .ZN(n10211) );
  NAND4_X1 U13388 ( .A1(n12069), .A2(n9720), .A3(n12035), .A4(n11457), .ZN(
        n12041) );
  INV_X1 U13389 ( .A(n10224), .ZN(n11524) );
  NAND2_X2 U13390 ( .A1(n10245), .A2(n10154), .ZN(n15216) );
  NAND2_X1 U13391 ( .A1(n13351), .A2(n10216), .ZN(n11212) );
  NAND2_X1 U13392 ( .A1(n11323), .A2(n11217), .ZN(n10216) );
  NAND2_X1 U13394 ( .A1(n10861), .A2(n11218), .ZN(n10217) );
  NAND3_X1 U13395 ( .A1(n10876), .A2(n10219), .A3(n10218), .ZN(n13351) );
  NAND3_X1 U13396 ( .A1(n10862), .A2(n10872), .A3(n10280), .ZN(n10873) );
  INV_X1 U13397 ( .A(n10295), .ZN(n10219) );
  NAND2_X1 U13398 ( .A1(n10859), .A2(n10872), .ZN(n11203) );
  NAND3_X1 U13399 ( .A1(n17513), .A2(n17512), .A3(n11113), .ZN(n10250) );
  INV_X1 U13400 ( .A(n14458), .ZN(n10221) );
  NAND2_X1 U13401 ( .A1(n10222), .A2(n9835), .ZN(n10223) );
  NAND3_X1 U13402 ( .A1(n10251), .A2(n10252), .A3(n12803), .ZN(n10222) );
  NOR2_X1 U13403 ( .A1(n10224), .A2(n11517), .ZN(n11605) );
  NAND2_X1 U13404 ( .A1(n11518), .A2(n10225), .ZN(n11519) );
  NAND2_X1 U13405 ( .A1(n16454), .A2(n10225), .ZN(n14330) );
  AND2_X1 U13406 ( .A1(n11525), .A2(n10225), .ZN(n20401) );
  NOR2_X1 U13407 ( .A1(n11517), .A2(n19987), .ZN(n10226) );
  INV_X1 U13408 ( .A(n12801), .ZN(n10251) );
  NAND2_X1 U13409 ( .A1(n10301), .A2(n10530), .ZN(n17211) );
  NOR2_X2 U13410 ( .A1(n17337), .A2(n17087), .ZN(n17162) );
  NAND2_X1 U13411 ( .A1(n11012), .A2(n11067), .ZN(n10544) );
  INV_X1 U13412 ( .A(n14934), .ZN(n15015) );
  AOI21_X2 U13413 ( .B1(n16525), .B2(n16262), .A(n16239), .ZN(n16534) );
  NAND2_X2 U13414 ( .A1(n10232), .A2(n10231), .ZN(n18706) );
  NAND3_X1 U13415 ( .A1(n10236), .A2(n10234), .A3(n10233), .ZN(P3_U2804) );
  NAND2_X2 U13416 ( .A1(n19820), .A2(n19938), .ZN(n17710) );
  NAND2_X2 U13417 ( .A1(n10240), .A2(n10237), .ZN(n19820) );
  AND2_X2 U13418 ( .A1(n19183), .A2(n19943), .ZN(n19786) );
  OAI21_X1 U13419 ( .B1(n10970), .B2(n10314), .A(n10901), .ZN(n10241) );
  NAND3_X1 U13420 ( .A1(n10971), .A2(n10901), .A3(n10687), .ZN(n10242) );
  INV_X1 U13421 ( .A(n10314), .ZN(n10243) );
  INV_X1 U13422 ( .A(n10970), .ZN(n10244) );
  NOR2_X2 U13423 ( .A1(n11212), .A2(n10253), .ZN(n10882) );
  INV_X1 U13424 ( .A(n13972), .ZN(n10255) );
  NAND2_X1 U13425 ( .A1(n11323), .A2(n9874), .ZN(n10256) );
  OAI21_X1 U13426 ( .B1(n11753), .B2(n10258), .A(n10257), .ZN(n16342) );
  NAND2_X1 U13427 ( .A1(n16342), .A2(n12418), .ZN(n12419) );
  OAI21_X1 U13428 ( .B1(n16745), .B2(n10261), .A(n16744), .ZN(n16746) );
  NAND2_X1 U13429 ( .A1(n16884), .A2(n9920), .ZN(n10472) );
  NAND2_X1 U13430 ( .A1(n10267), .A2(n11535), .ZN(n10268) );
  NAND4_X1 U13431 ( .A1(n11433), .A2(n11432), .A3(n11434), .A4(n11431), .ZN(
        n10267) );
  NAND2_X1 U13432 ( .A1(n10270), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10269) );
  NAND4_X1 U13433 ( .A1(n11428), .A2(n11429), .A3(n11427), .A4(n11426), .ZN(
        n10270) );
  NAND4_X1 U13434 ( .A1(n11447), .A2(n11448), .A3(n11446), .A4(n11445), .ZN(
        n10273) );
  OAI21_X1 U13435 ( .B1(n10275), .B2(n10382), .A(n15943), .ZN(n10430) );
  XNOR2_X1 U13436 ( .A(n10275), .B(n10274), .ZN(n14332) );
  INV_X1 U13437 ( .A(n14315), .ZN(n10274) );
  INV_X1 U13438 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10276) );
  NAND4_X1 U13439 ( .A1(n10893), .A2(n10894), .A3(n10887), .A4(n10896), .ZN(
        n10918) );
  NAND2_X1 U13440 ( .A1(n12819), .A2(n10871), .ZN(n11338) );
  NAND2_X1 U13441 ( .A1(n14368), .A2(n10282), .ZN(n14862) );
  NAND4_X1 U13442 ( .A1(n12251), .A2(n11895), .A3(n11462), .A4(n10734), .ZN(
        n11469) );
  NAND4_X1 U13443 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10288) );
  AND2_X2 U13444 ( .A1(n13893), .A2(n11524), .ZN(n20336) );
  NAND2_X1 U13445 ( .A1(n10295), .A2(n10867), .ZN(n10874) );
  NAND2_X1 U13446 ( .A1(n10296), .A2(n10446), .ZN(n10445) );
  NAND3_X1 U13447 ( .A1(n10882), .A2(n10879), .A3(n11200), .ZN(n10296) );
  OR2_X1 U13448 ( .A1(n14202), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10297) );
  NAND3_X1 U13449 ( .A1(n14127), .A2(n11048), .A3(n10297), .ZN(n11051) );
  NAND2_X1 U13450 ( .A1(n17211), .A2(n10300), .ZN(n17091) );
  NAND2_X1 U13451 ( .A1(n18759), .A2(n18910), .ZN(n18764) );
  NAND2_X1 U13452 ( .A1(n18759), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10530) );
  AND2_X1 U13453 ( .A1(n10531), .A2(n17374), .ZN(n10301) );
  INV_X1 U13454 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13915) );
  NAND2_X1 U13455 ( .A1(n10302), .A2(n17058), .ZN(n19016) );
  NAND2_X1 U13456 ( .A1(n19026), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10302) );
  NAND2_X1 U13457 ( .A1(n10304), .A2(n10303), .ZN(P3_U2833) );
  NAND2_X1 U13458 ( .A1(n17316), .A2(n19255), .ZN(n10304) );
  NAND2_X1 U13459 ( .A1(n10307), .A2(n10306), .ZN(n10305) );
  NAND2_X1 U13460 ( .A1(n17162), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10306) );
  INV_X1 U13461 ( .A(n17162), .ZN(n10308) );
  NOR2_X1 U13462 ( .A1(n19147), .A2(n10312), .ZN(n10311) );
  NAND2_X1 U13463 ( .A1(n10314), .A2(n10455), .ZN(n14590) );
  NAND3_X1 U13464 ( .A1(n10314), .A2(n10455), .A3(n20825), .ZN(n11023) );
  NAND2_X1 U13465 ( .A1(n15278), .A2(n10324), .ZN(n11122) );
  NAND2_X1 U13466 ( .A1(n10735), .A2(n9902), .ZN(n10324) );
  AND2_X4 U13467 ( .A1(n11107), .A2(n11106), .ZN(n10735) );
  NAND2_X1 U13468 ( .A1(n15627), .A2(n9785), .ZN(n10327) );
  INV_X1 U13469 ( .A(n15617), .ZN(n10333) );
  NAND2_X1 U13470 ( .A1(n15863), .A2(n9861), .ZN(n15825) );
  NAND3_X1 U13471 ( .A1(n10341), .A2(n15938), .A3(n16447), .ZN(n15901) );
  INV_X1 U13472 ( .A(n10345), .ZN(n15912) );
  NAND3_X1 U13473 ( .A1(n10352), .A2(n10386), .A3(n16470), .ZN(n10351) );
  NAND2_X1 U13474 ( .A1(n10644), .A2(n10356), .ZN(n11128) );
  NAND2_X1 U13475 ( .A1(n10358), .A2(n10359), .ZN(n10357) );
  INV_X1 U13476 ( .A(n10360), .ZN(n10358) );
  NAND2_X1 U13477 ( .A1(n11507), .A2(n10362), .ZN(n10361) );
  INV_X1 U13478 ( .A(n11500), .ZN(n10362) );
  XNOR2_X2 U13479 ( .A(n10370), .B(n10900), .ZN(n10970) );
  NAND2_X1 U13480 ( .A1(n10445), .A2(n10881), .ZN(n10370) );
  AOI21_X2 U13481 ( .B1(n11113), .B2(n10378), .A(n9848), .ZN(n10377) );
  NAND4_X1 U13482 ( .A1(n11035), .A2(n11036), .A3(n11011), .A4(n14114), .ZN(
        n11067) );
  NAND2_X1 U13483 ( .A1(n11087), .A2(n10379), .ZN(n12867) );
  INV_X1 U13484 ( .A(n9794), .ZN(n10381) );
  NAND3_X1 U13485 ( .A1(n11753), .A2(n11752), .A3(n10404), .ZN(n10401) );
  NAND3_X1 U13486 ( .A1(n11753), .A2(n11752), .A3(n10478), .ZN(n10477) );
  NAND3_X1 U13487 ( .A1(n10408), .A2(n10407), .A3(n14606), .ZN(n10406) );
  NAND2_X1 U13488 ( .A1(n10515), .A2(n11939), .ZN(n10483) );
  AND2_X2 U13489 ( .A1(n10483), .A2(n10482), .ZN(n10411) );
  OAI211_X1 U13490 ( .C1(n12432), .C2(n10414), .A(n10413), .B(n10412), .ZN(
        n16482) );
  NAND2_X1 U13491 ( .A1(n12432), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10412) );
  AND2_X2 U13492 ( .A1(n13654), .A2(n17403), .ZN(n18254) );
  AND4_X2 U13493 ( .A1(n9782), .A2(n9851), .A3(n13747), .A4(n13751), .ZN(
        n19355) );
  NAND2_X1 U13494 ( .A1(n18532), .A2(n9796), .ZN(n18520) );
  INV_X2 U13495 ( .A(n13729), .ZN(n17446) );
  NAND2_X2 U13496 ( .A1(n13665), .A2(n17415), .ZN(n13729) );
  AND2_X2 U13497 ( .A1(n10426), .A2(n13659), .ZN(n13665) );
  INV_X2 U13498 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10426) );
  INV_X1 U13499 ( .A(n16973), .ZN(n10427) );
  NAND2_X1 U13500 ( .A1(n10427), .A2(n10428), .ZN(n18596) );
  INV_X1 U13501 ( .A(n15943), .ZN(n10433) );
  NAND2_X1 U13502 ( .A1(n16458), .A2(n12032), .ZN(n10434) );
  XNOR2_X1 U13503 ( .A(n16458), .B(n9896), .ZN(n14334) );
  OAI21_X1 U13504 ( .B1(n12415), .B2(n10441), .A(n10437), .ZN(n16353) );
  AOI21_X2 U13505 ( .B1(n10440), .B2(n10439), .A(n10438), .ZN(n10437) );
  OAI21_X1 U13506 ( .B1(n10443), .B2(n10442), .A(n10683), .ZN(n10682) );
  NAND2_X1 U13507 ( .A1(n14695), .A2(n10444), .ZN(n10443) );
  NAND2_X1 U13508 ( .A1(n14696), .A2(n14697), .ZN(n10444) );
  NAND4_X1 U13509 ( .A1(n10745), .A2(n10880), .A3(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10469) );
  NAND3_X1 U13510 ( .A1(n11051), .A2(n11052), .A3(n11050), .ZN(n17525) );
  INV_X1 U13511 ( .A(n11074), .ZN(n10451) );
  NAND2_X2 U13512 ( .A1(n10772), .A2(n10771), .ZN(n10994) );
  AND2_X2 U13513 ( .A1(n10795), .A2(n10794), .ZN(n12819) );
  NAND3_X1 U13514 ( .A1(n15198), .A2(n15190), .A3(n10735), .ZN(n10456) );
  XNOR2_X2 U13515 ( .A(n10460), .B(n10917), .ZN(n11035) );
  NAND2_X1 U13516 ( .A1(n9816), .A2(n10638), .ZN(n10462) );
  NAND2_X1 U13517 ( .A1(n11129), .A2(n10464), .ZN(n10463) );
  AND2_X1 U13518 ( .A1(n10467), .A2(n10637), .ZN(n10464) );
  NAND2_X1 U13519 ( .A1(n11204), .A2(n10866), .ZN(n10860) );
  NAND3_X1 U13520 ( .A1(n12819), .A2(n10994), .A3(n10866), .ZN(n11204) );
  INV_X2 U13521 ( .A(n10469), .ZN(n10919) );
  AOI22_X1 U13522 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10919), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10790) );
  NOR2_X2 U13523 ( .A1(n19204), .A2(n10484), .ZN(n18933) );
  NAND2_X2 U13524 ( .A1(n17266), .A2(n17141), .ZN(n17339) );
  OAI21_X1 U13525 ( .B1(n18455), .B2(n14535), .A(n10493), .ZN(n10491) );
  INV_X1 U13526 ( .A(n10491), .ZN(n10492) );
  NAND3_X1 U13527 ( .A1(n13654), .A2(n17403), .A3(
        P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10493) );
  XNOR2_X2 U13528 ( .A(n17103), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17742) );
  NAND2_X1 U13529 ( .A1(n17805), .A2(n9891), .ZN(n10496) );
  INV_X1 U13530 ( .A(n10498), .ZN(n17847) );
  INV_X1 U13531 ( .A(n10503), .ZN(n17214) );
  NAND3_X1 U13532 ( .A1(n10504), .A2(n10506), .A3(n17261), .ZN(n18891) );
  NAND2_X1 U13533 ( .A1(n10514), .A2(n11929), .ZN(n16462) );
  INV_X1 U13534 ( .A(n11928), .ZN(n10514) );
  NAND3_X1 U13535 ( .A1(n10526), .A2(n12473), .A3(n12472), .ZN(P2_U3029) );
  NAND2_X1 U13536 ( .A1(n18783), .A2(n10532), .ZN(n18759) );
  INV_X1 U13537 ( .A(n10535), .ZN(n17048) );
  NOR2_X1 U13538 ( .A1(n10535), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17128) );
  NAND2_X1 U13539 ( .A1(n17124), .A2(n10535), .ZN(n17054) );
  NAND2_X1 U13540 ( .A1(n17127), .A2(n10535), .ZN(n17125) );
  MUX2_X1 U13541 ( .A(n10534), .B(n10535), .S(n17127), .Z(n17129) );
  AOI21_X1 U13542 ( .B1(n10535), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10534) );
  AND2_X4 U13543 ( .A1(n10753), .A2(n10757), .ZN(n13211) );
  OAI22_X2 U13544 ( .A1(n10544), .A2(n11104), .B1(n11014), .B2(n17492), .ZN(
        n14202) );
  NAND2_X1 U13545 ( .A1(n10545), .A2(n10549), .ZN(P1_U2969) );
  NAND2_X1 U13546 ( .A1(n10546), .A2(n10547), .ZN(n10545) );
  CLKBUF_X1 U13547 ( .A(n10553), .Z(n10552) );
  NAND2_X1 U13548 ( .A1(n10867), .A2(n10552), .ZN(n11040) );
  NAND2_X1 U13549 ( .A1(n10889), .A2(n10552), .ZN(n10890) );
  NAND2_X1 U13550 ( .A1(n14307), .A2(n10552), .ZN(n21022) );
  AND2_X2 U13551 ( .A1(n10554), .A2(n10755), .ZN(n10811) );
  NAND3_X1 U13552 ( .A1(n11234), .A2(n10556), .A3(n11233), .ZN(n14210) );
  INV_X1 U13553 ( .A(n14210), .ZN(n11246) );
  NAND2_X1 U13554 ( .A1(n10559), .A2(n10560), .ZN(n13877) );
  INV_X1 U13555 ( .A(n14336), .ZN(n10561) );
  NAND2_X1 U13556 ( .A1(n10561), .A2(n9855), .ZN(n14454) );
  NOR2_X1 U13557 ( .A1(n14336), .A2(n10563), .ZN(n14363) );
  NAND2_X1 U13558 ( .A1(n14781), .A2(n9894), .ZN(n14759) );
  AND2_X2 U13559 ( .A1(n14781), .A2(n9904), .ZN(n14724) );
  NAND2_X1 U13560 ( .A1(n11286), .A2(n9887), .ZN(n14849) );
  AND2_X1 U13561 ( .A1(n15667), .A2(n15646), .ZN(n12019) );
  INV_X1 U13562 ( .A(n12319), .ZN(n10592) );
  NAND2_X1 U13563 ( .A1(n10592), .A2(n10593), .ZN(n12327) );
  INV_X1 U13564 ( .A(n14042), .ZN(n10598) );
  NAND2_X1 U13565 ( .A1(n10598), .A2(n10599), .ZN(n14051) );
  NAND2_X1 U13566 ( .A1(n10603), .A2(n10605), .ZN(n14059) );
  NAND3_X1 U13567 ( .A1(n14075), .A2(n10733), .A3(n10604), .ZN(n10603) );
  INV_X1 U13568 ( .A(n12097), .ZN(n10606) );
  NAND3_X1 U13569 ( .A1(n10733), .A2(n14075), .A3(n12097), .ZN(n15932) );
  NAND2_X1 U13570 ( .A1(n12421), .A2(n9783), .ZN(n10607) );
  AND2_X1 U13571 ( .A1(n15657), .A2(n15659), .ZN(n15644) );
  AND2_X2 U13572 ( .A1(n15657), .A2(n9888), .ZN(n15611) );
  NAND2_X1 U13573 ( .A1(n14270), .A2(n10617), .ZN(n15748) );
  NAND3_X1 U13574 ( .A1(n11527), .A2(n10627), .A3(n10626), .ZN(n10625) );
  NAND3_X1 U13575 ( .A1(n12500), .A2(n12499), .A3(n10633), .ZN(n14625) );
  NAND2_X1 U13576 ( .A1(n11840), .A2(n11839), .ZN(n16236) );
  NAND2_X1 U13577 ( .A1(n11765), .A2(n10648), .ZN(n11824) );
  NAND2_X1 U13578 ( .A1(n11765), .A2(n11763), .ZN(n11770) );
  NAND2_X1 U13579 ( .A1(n11845), .A2(n9790), .ZN(n12477) );
  NAND2_X1 U13580 ( .A1(n11845), .A2(n9905), .ZN(n12476) );
  INV_X1 U13581 ( .A(n11732), .ZN(n10652) );
  NAND2_X1 U13582 ( .A1(n11748), .A2(n10658), .ZN(n11784) );
  NAND2_X1 U13583 ( .A1(n13609), .A2(n12533), .ZN(n13866) );
  INV_X1 U13584 ( .A(n13866), .ZN(n10659) );
  NAND2_X1 U13585 ( .A1(n13865), .A2(n12534), .ZN(n13889) );
  NAND3_X1 U13586 ( .A1(n12523), .A2(n10659), .A3(n12534), .ZN(n13865) );
  AOI21_X1 U13587 ( .B1(n16006), .B2(n10661), .A(n12771), .ZN(n10660) );
  NAND2_X1 U13588 ( .A1(n16006), .A2(n10667), .ZN(n10665) );
  NAND2_X1 U13589 ( .A1(n10664), .A2(n10660), .ZN(n12795) );
  OAI21_X1 U13590 ( .B1(n14707), .B2(n14706), .A(n10681), .ZN(P2_U3030) );
  NOR2_X1 U13591 ( .A1(n14402), .A2(n15016), .ZN(n14934) );
  INV_X1 U13592 ( .A(n15016), .ZN(n10690) );
  INV_X1 U13593 ( .A(n10697), .ZN(n14822) );
  NAND2_X1 U13594 ( .A1(n14795), .A2(n14796), .ZN(n14783) );
  CLKBUF_X1 U13595 ( .A(n14336), .Z(n17552) );
  CLKBUF_X1 U13596 ( .A(n14454), .Z(n15574) );
  INV_X1 U13597 ( .A(n14454), .ZN(n11263) );
  INV_X1 U13598 ( .A(n14046), .ZN(n12128) );
  INV_X1 U13599 ( .A(n14051), .ZN(n12182) );
  INV_X1 U13600 ( .A(n14835), .ZN(n14851) );
  INV_X1 U13601 ( .A(n12471), .ZN(n12472) );
  NAND2_X1 U13602 ( .A1(n12307), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12312) );
  OAI21_X1 U13603 ( .B1(n12275), .B2(n17594), .A(n12274), .ZN(n12276) );
  OAI21_X1 U13604 ( .B1(n12275), .B2(n16748), .A(n12258), .ZN(n12259) );
  NAND2_X1 U13605 ( .A1(n13889), .A2(n13892), .ZN(n13890) );
  AOI21_X1 U13606 ( .B1(n15056), .B2(n20909), .A(n14646), .ZN(n14647) );
  INV_X1 U13607 ( .A(n9746), .ZN(n14374) );
  NAND2_X1 U13608 ( .A1(n14114), .A2(n9746), .ZN(n21415) );
  AND2_X2 U13609 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13977) );
  OAI211_X1 U13610 ( .C1(n12364), .C2(n12363), .A(n12362), .B(n9777), .ZN(
        n12365) );
  OAI211_X1 U13611 ( .C1(n12090), .C2(n19973), .A(n12071), .B(n12070), .ZN(
        n13953) );
  CLKBUF_X1 U13612 ( .A(n11910), .Z(n16821) );
  NAND2_X1 U13613 ( .A1(n10993), .A2(n14114), .ZN(n11009) );
  AND2_X2 U13614 ( .A1(n9729), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11568) );
  AOI22_X1 U13615 ( .A1(n12644), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12784), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11394) );
  AND2_X1 U13616 ( .A1(n9746), .A2(n14115), .ZN(n21139) );
  NAND2_X1 U13617 ( .A1(n11010), .A2(n14115), .ZN(n12848) );
  AND2_X1 U13618 ( .A1(n20936), .A2(n10872), .ZN(n20932) );
  AND2_X1 U13619 ( .A1(n12450), .A2(n12449), .ZN(n10711) );
  OR2_X1 U13620 ( .A1(n17615), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10712) );
  AND2_X1 U13621 ( .A1(n12451), .A2(n10711), .ZN(n10713) );
  AND2_X1 U13622 ( .A1(n12255), .A2(n11917), .ZN(n17602) );
  AND2_X1 U13623 ( .A1(n16887), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10714) );
  OR2_X1 U13624 ( .A1(n18706), .A2(n19943), .ZN(n10715) );
  NAND2_X1 U13625 ( .A1(n12285), .A2(n12284), .ZN(n10716) );
  AND2_X1 U13626 ( .A1(n16473), .A2(n16080), .ZN(n10717) );
  AND2_X1 U13627 ( .A1(n12829), .A2(n12828), .ZN(n10718) );
  AND2_X1 U13628 ( .A1(n12515), .A2(n12514), .ZN(n10719) );
  OR2_X1 U13629 ( .A1(n18810), .A2(n17911), .ZN(n10720) );
  OR2_X1 U13630 ( .A1(n17397), .A2(n19226), .ZN(n10721) );
  INV_X1 U13631 ( .A(n17425), .ZN(n13903) );
  INV_X1 U13632 ( .A(n11333), .ZN(n12804) );
  AND2_X1 U13633 ( .A1(n16078), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10723) );
  INV_X1 U13634 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11842) );
  AND2_X1 U13635 ( .A1(n11693), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10724) );
  INV_X1 U13636 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n21483) );
  OR2_X1 U13637 ( .A1(n20244), .A2(n20535), .ZN(n20306) );
  INV_X1 U13638 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12311) );
  AND4_X1 U13639 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(P3_EAX_REG_20__SCAN_IN), .ZN(n10725)
         );
  AND3_X1 U13640 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10726) );
  AND3_X1 U13641 ( .A1(n12998), .A2(n12997), .A3(n12996), .ZN(n10727) );
  INV_X1 U13642 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15295) );
  OR2_X1 U13643 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20684), .ZN(n20818) );
  AND2_X1 U13644 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10730) );
  NAND2_X1 U13645 ( .A1(n12028), .A2(n12073), .ZN(n10731) );
  OR2_X1 U13646 ( .A1(n16022), .A2(n16014), .ZN(n10732) );
  AND2_X1 U13647 ( .A1(n20807), .A2(n20118), .ZN(n10734) );
  INV_X1 U13648 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20395) );
  INV_X1 U13649 ( .A(n20904), .ZN(n17539) );
  AND3_X1 U13650 ( .A1(n16030), .A2(n16028), .A3(n16031), .ZN(n10736) );
  NAND2_X2 U13651 ( .A1(n9725), .A2(n18595), .ZN(n18484) );
  AND2_X1 U13652 ( .A1(n16032), .A2(n16030), .ZN(n10737) );
  AND2_X1 U13653 ( .A1(n15709), .A2(n15708), .ZN(n10738) );
  INV_X1 U13654 ( .A(n12440), .ZN(n15733) );
  INV_X1 U13655 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10884) );
  NAND2_X1 U13656 ( .A1(n10752), .A2(n13977), .ZN(n10820) );
  AND2_X1 U13657 ( .A1(n11086), .A2(n11085), .ZN(n10742) );
  NOR2_X2 U13658 ( .A1(n21415), .A2(n21339), .ZN(n10743) );
  INV_X1 U13659 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10746) );
  AND2_X1 U13660 ( .A1(n11105), .A2(n10973), .ZN(n10974) );
  INV_X1 U13661 ( .A(n11157), .ZN(n11145) );
  NAND2_X1 U13662 ( .A1(n11135), .A2(n11134), .ZN(n11144) );
  OR2_X1 U13663 ( .A1(n10951), .A2(n10950), .ZN(n10952) );
  INV_X1 U13664 ( .A(n11858), .ZN(n11649) );
  AND4_X1 U13665 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11614) );
  NOR2_X1 U13666 ( .A1(n20113), .A2(n20808), .ZN(n11460) );
  NAND2_X1 U13667 ( .A1(n11661), .A2(n11660), .ZN(n11665) );
  INV_X1 U13668 ( .A(n10862), .ZN(n10863) );
  INV_X1 U13669 ( .A(n12855), .ZN(n12827) );
  NOR2_X1 U13670 ( .A1(n15277), .A2(n10728), .ZN(n11117) );
  NOR2_X2 U13671 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U13672 ( .A1(n11430), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11399) );
  INV_X1 U13673 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11736) );
  AND4_X1 U13674 ( .A1(n11717), .A2(n11716), .A3(n11715), .A4(n11714), .ZN(
        n11728) );
  OR3_X1 U13675 ( .A1(n11871), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n11668), .ZN(n11856) );
  NAND2_X1 U13676 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10829) );
  INV_X1 U13677 ( .A(n14865), .ZN(n13112) );
  INV_X1 U13678 ( .A(n12932), .ZN(n12933) );
  OR2_X1 U13679 ( .A1(n11062), .A2(n11061), .ZN(n11070) );
  OR2_X1 U13680 ( .A1(n11138), .A2(n11137), .ZN(n11140) );
  OR2_X1 U13681 ( .A1(n10965), .A2(n10964), .ZN(n11015) );
  INV_X1 U13682 ( .A(n11010), .ZN(n10993) );
  INV_X1 U13683 ( .A(n14048), .ZN(n12127) );
  INV_X1 U13684 ( .A(n14094), .ZN(n11953) );
  INV_X1 U13685 ( .A(n15751), .ZN(n12231) );
  NAND2_X1 U13686 ( .A1(n11667), .A2(n11666), .ZN(n11871) );
  AOI22_X1 U13687 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11383) );
  OR2_X1 U13688 ( .A1(n17071), .A2(n19270), .ZN(n17072) );
  AOI21_X1 U13689 ( .B1(n19806), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n13810), .ZN(n13802) );
  INV_X1 U13690 ( .A(n15573), .ZN(n11262) );
  INV_X1 U13691 ( .A(n14917), .ZN(n13035) );
  INV_X1 U13692 ( .A(n13017), .ZN(n13018) );
  INV_X1 U13693 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12981) );
  AND2_X1 U13694 ( .A1(n11267), .A2(n11266), .ZN(n15020) );
  INV_X1 U13695 ( .A(n17550), .ZN(n11245) );
  INV_X1 U13696 ( .A(n10916), .ZN(n11039) );
  INV_X1 U13697 ( .A(n10948), .ZN(n11022) );
  AND2_X1 U13698 ( .A1(n12544), .A2(n12543), .ZN(n12545) );
  INV_X1 U13699 ( .A(n12713), .ZN(n12696) );
  INV_X1 U13700 ( .A(n14036), .ZN(n11965) );
  INV_X1 U13701 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16466) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12416) );
  INV_X1 U13703 ( .A(n14084), .ZN(n12181) );
  AOI21_X1 U13704 ( .B1(n11871), .B2(n11870), .A(n11869), .ZN(n11902) );
  OAI22_X1 U13705 ( .A1(n13806), .A2(n13805), .B1(n21661), .B2(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n13814) );
  AND2_X1 U13706 ( .A1(n13127), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13128) );
  INV_X1 U13707 ( .A(n14227), .ZN(n14228) );
  NAND2_X1 U13708 ( .A1(n13053), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13090) );
  NAND2_X1 U13709 ( .A1(n12950), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13017) );
  INV_X1 U13710 ( .A(n12842), .ZN(n13047) );
  NAND2_X1 U13711 ( .A1(n11167), .A2(n13621), .ZN(n11187) );
  OR2_X1 U13712 ( .A1(n15520), .A2(n15525), .ZN(n15480) );
  INV_X1 U13713 ( .A(n13621), .ZN(n11104) );
  OR3_X1 U13714 ( .A1(n13993), .A2(n13992), .A3(n13991), .ZN(n14595) );
  NAND2_X1 U13715 ( .A1(n10979), .A2(n10978), .ZN(n14275) );
  INV_X1 U13716 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16346) );
  INV_X1 U13717 ( .A(n11755), .ZN(n11739) );
  OR2_X1 U13718 ( .A1(n12732), .A2(n12736), .ZN(n12766) );
  OR2_X1 U13719 ( .A1(n12638), .A2(n12637), .ZN(n12676) );
  AND3_X1 U13720 ( .A1(n12108), .A2(n12107), .A3(n12106), .ZN(n15933) );
  INV_X1 U13721 ( .A(n16254), .ZN(n11839) );
  AND2_X1 U13722 ( .A1(n12240), .A2(n12239), .ZN(n15691) );
  AND2_X1 U13723 ( .A1(n12046), .A2(n12045), .ZN(n16816) );
  NAND2_X1 U13724 ( .A1(n19377), .A2(n14481), .ZN(n13898) );
  INV_X1 U13725 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18328) );
  AND2_X1 U13726 ( .A1(n14483), .A2(n13769), .ZN(n13770) );
  AOI21_X1 U13727 ( .B1(n13808), .B2(n13807), .A(n13814), .ZN(n13818) );
  INV_X1 U13728 ( .A(n13280), .ZN(n13318) );
  NAND2_X1 U13729 ( .A1(n13128), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13179) );
  NAND2_X1 U13730 ( .A1(n14228), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14230) );
  INV_X1 U13731 ( .A(n20912), .ZN(n20882) );
  INV_X1 U13732 ( .A(n14274), .ZN(n15086) );
  OR2_X1 U13733 ( .A1(n13019), .A2(n15295), .ZN(n13052) );
  AND2_X1 U13734 ( .A1(n12870), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12877) );
  INV_X1 U13735 ( .A(n12808), .ZN(n12809) );
  INV_X1 U13736 ( .A(n15277), .ZN(n15293) );
  OR2_X1 U13737 ( .A1(n21082), .A2(n21081), .ZN(n21113) );
  NAND2_X1 U13738 ( .A1(n21139), .A2(n21225), .ZN(n14449) );
  NOR2_X1 U13739 ( .A1(n21293), .A2(n14414), .ZN(n21236) );
  XNOR2_X1 U13740 ( .A(n12840), .B(n12839), .ZN(n14375) );
  AND2_X1 U13741 ( .A1(n14113), .A2(n14375), .ZN(n21225) );
  INV_X1 U13742 ( .A(n12798), .ZN(n12799) );
  AND2_X1 U13743 ( .A1(n12280), .A2(n12279), .ZN(n14627) );
  INV_X1 U13744 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16306) );
  INV_X1 U13745 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16316) );
  AND2_X1 U13746 ( .A1(n13520), .A2(n12297), .ZN(n13388) );
  INV_X1 U13747 ( .A(n14715), .ZN(n14716) );
  NOR2_X1 U13748 ( .A1(n10000), .A2(n15614), .ZN(n15615) );
  OR2_X1 U13749 ( .A1(n16633), .A2(n12461), .ZN(n16620) );
  NAND2_X1 U13750 ( .A1(n16723), .A2(n16700), .ZN(n16685) );
  AND4_X1 U13752 ( .A1(n12263), .A2(n13533), .A3(n11914), .A4(n11913), .ZN(
        n11915) );
  OR2_X1 U13753 ( .A1(n20148), .A2(n20147), .ZN(n20152) );
  OR2_X1 U13754 ( .A1(n20453), .A2(n20205), .ZN(n20237) );
  OR2_X1 U13755 ( .A1(n20205), .A2(n20535), .ZN(n20298) );
  NOR2_X1 U13756 ( .A1(n20762), .A2(n20750), .ZN(n20746) );
  OR2_X1 U13757 ( .A1(n11605), .A2(n20611), .ZN(n20618) );
  NOR2_X1 U13758 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20801) );
  NOR2_X1 U13759 ( .A1(n18791), .A2(n17829), .ZN(n17828) );
  INV_X1 U13760 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17907) );
  NOR2_X1 U13761 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17977), .ZN(n17976) );
  INV_X1 U13762 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n18020) );
  NOR2_X1 U13763 ( .A1(n14481), .A2(n18595), .ZN(n14482) );
  INV_X1 U13764 ( .A(n19373), .ZN(n18509) );
  INV_X1 U13765 ( .A(n18855), .ZN(n18896) );
  INV_X1 U13766 ( .A(n18624), .ZN(n17330) );
  AOI21_X1 U13767 ( .B1(n19341), .B2(n19842), .A(n19821), .ZN(n19352) );
  INV_X1 U13768 ( .A(n19200), .ZN(n19232) );
  INV_X1 U13769 ( .A(n19591), .ZN(n19635) );
  OR2_X1 U13770 ( .A1(n21475), .A2(n20825), .ZN(n20822) );
  OR2_X1 U13771 ( .A1(n14240), .A2(n10867), .ZN(n14245) );
  XNOR2_X1 U13772 ( .A(n14230), .B(n14229), .ZN(n15164) );
  INV_X1 U13773 ( .A(n20851), .ZN(n20879) );
  INV_X1 U13774 ( .A(n20883), .ZN(n20907) );
  INV_X1 U13775 ( .A(n20936), .ZN(n15075) );
  INV_X1 U13776 ( .A(n15138), .ZN(n15128) );
  NOR2_X2 U13777 ( .A1(n20988), .A2(n14157), .ZN(n20980) );
  INV_X1 U13778 ( .A(n17527), .ZN(n20933) );
  INV_X1 U13779 ( .A(n17524), .ZN(n17528) );
  OR2_X1 U13780 ( .A1(n15560), .A2(n17546), .ZN(n17540) );
  NAND2_X1 U13781 ( .A1(n14136), .A2(n14135), .ZN(n17555) );
  INV_X1 U13782 ( .A(n14378), .ZN(n21369) );
  NOR2_X1 U13783 ( .A1(n13556), .A2(n14157), .ZN(n17468) );
  NOR2_X1 U13784 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n17567) );
  INV_X1 U13785 ( .A(n21074), .ZN(n21055) );
  OAI211_X1 U13786 ( .C1(n14385), .C2(n14384), .A(n21236), .B(n14383), .ZN(
        n21071) );
  INV_X1 U13787 ( .A(n21113), .ZN(n21132) );
  AND2_X1 U13788 ( .A1(n21139), .A2(n14408), .ZN(n21160) );
  OAI211_X1 U13789 ( .C1(n21420), .C2(n14412), .A(n21416), .B(n14281), .ZN(
        n14312) );
  INV_X1 U13790 ( .A(n21109), .ZN(n21165) );
  NOR2_X2 U13791 ( .A1(n21264), .A2(n21339), .ZN(n21252) );
  NOR2_X2 U13792 ( .A1(n21264), .A2(n21368), .ZN(n21283) );
  INV_X1 U13793 ( .A(n21300), .ZN(n21323) );
  OAI21_X1 U13794 ( .B1(n21338), .B2(n21337), .A(n21416), .ZN(n21363) );
  AND2_X1 U13795 ( .A1(n14305), .A2(n15134), .ZN(n21425) );
  INV_X1 U13796 ( .A(n21472), .ZN(n21446) );
  INV_X1 U13797 ( .A(n21367), .ZN(n21467) );
  INV_X1 U13798 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21486) );
  AND2_X1 U13799 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21583), .ZN(n21533) );
  NAND2_X1 U13800 ( .A1(n20800), .A2(n20489), .ZN(n20804) );
  INV_X1 U13801 ( .A(n19987), .ZN(n12388) );
  AND2_X1 U13802 ( .A1(n13415), .A2(n12292), .ZN(n15984) );
  OR2_X1 U13803 ( .A1(n13413), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16464) );
  AND2_X1 U13804 ( .A1(n13415), .A2(n16932), .ZN(n15982) );
  INV_X1 U13805 ( .A(n19981), .ZN(n15968) );
  OR2_X1 U13806 ( .A1(n12206), .A2(n12205), .ZN(n16087) );
  OR2_X1 U13807 ( .A1(n12165), .A2(n12164), .ZN(n14151) );
  INV_X1 U13808 ( .A(n16072), .ZN(n16086) );
  OR2_X1 U13809 ( .A1(n13411), .A2(n11478), .ZN(n13427) );
  BUF_X1 U13810 ( .A(n16387), .Z(n16444) );
  INV_X1 U13811 ( .A(n16764), .ZN(n17604) );
  AOI21_X1 U13812 ( .B1(n16614), .B2(n12457), .A(n16608), .ZN(n12458) );
  NOR2_X1 U13813 ( .A1(n16768), .A2(n12049), .ZN(n16723) );
  OAI21_X1 U13814 ( .B1(n20215), .B2(n20214), .A(n20213), .ZN(n20239) );
  INV_X1 U13815 ( .A(n20306), .ZN(n20275) );
  OAI21_X1 U13816 ( .B1(n20283), .B2(n20282), .A(n20281), .ZN(n20308) );
  INV_X1 U13817 ( .A(n20298), .ZN(n20312) );
  NOR2_X1 U13818 ( .A1(n20556), .A2(n20396), .ZN(n20394) );
  AOI21_X1 U13819 ( .B1(n20489), .B2(n20459), .A(n20462), .ZN(n20481) );
  OAI211_X1 U13820 ( .C1(n20534), .C2(n20562), .A(n20619), .B(n20533), .ZN(
        n20552) );
  INV_X1 U13821 ( .A(n20571), .ZN(n20621) );
  INV_X1 U13822 ( .A(n20582), .ZN(n20639) );
  AND2_X1 U13823 ( .A1(n20808), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16838) );
  INV_X1 U13824 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21751) );
  NAND2_X1 U13825 ( .A1(n19938), .A2(n19789), .ZN(n18705) );
  NOR2_X1 U13826 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17814), .ZN(n17793) );
  NOR2_X1 U13827 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17852), .ZN(n17840) );
  NOR2_X1 U13828 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17874), .ZN(n17856) );
  NOR2_X1 U13829 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17900), .ZN(n17880) );
  NOR2_X1 U13830 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17968), .ZN(n17953) );
  NOR2_X1 U13831 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18075), .ZN(n18053) );
  NOR2_X2 U13832 ( .A1(n19956), .A2(n19823), .ZN(n18093) );
  NAND4_X1 U13833 ( .A1(n19156), .A2(n19954), .A3(n19839), .A4(n19828), .ZN(
        n18116) );
  AOI22_X1 U13834 ( .A1(n9870), .A2(n14484), .B1(n14483), .B2(n14482), .ZN(
        n16952) );
  OR2_X1 U13835 ( .A1(n17047), .A2(n17046), .ZN(n18624) );
  OAI211_X1 U13836 ( .C1(n19944), .C2(n19943), .A(n18704), .B(n18703), .ZN(
        n18734) );
  NOR2_X1 U13837 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19352), .ZN(n19591) );
  AND2_X1 U13838 ( .A1(n19213), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n19210) );
  INV_X1 U13839 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17241) );
  AND2_X1 U13840 ( .A1(n19331), .A2(n18624), .ZN(n19255) );
  AND2_X1 U13841 ( .A1(n19323), .A2(n10239), .ZN(n19331) );
  NAND2_X1 U13842 ( .A1(n17425), .A2(n13904), .ZN(n19337) );
  CLKBUF_X1 U13843 ( .A(n19481), .Z(n19493) );
  INV_X1 U13844 ( .A(n19537), .ZN(n19539) );
  INV_X1 U13845 ( .A(n19557), .ZN(n19561) );
  INV_X1 U13846 ( .A(n19633), .ZN(n19626) );
  NOR2_X1 U13847 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19923), .ZN(n19688) );
  INV_X1 U13848 ( .A(n19830), .ZN(n19938) );
  NAND2_X1 U13849 ( .A1(n17503), .A2(n13444), .ZN(n14226) );
  INV_X1 U13850 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21173) );
  INV_X1 U13851 ( .A(n20889), .ZN(n20917) );
  INV_X1 U13852 ( .A(n15349), .ZN(n15155) );
  NAND2_X1 U13853 ( .A1(n13358), .A2(n13357), .ZN(n15151) );
  INV_X1 U13854 ( .A(n20940), .ZN(n20969) );
  NOR2_X1 U13855 ( .A1(n14226), .A2(n14156), .ZN(n14169) );
  NAND2_X1 U13856 ( .A1(n17533), .A2(n13624), .ZN(n17524) );
  INV_X1 U13857 ( .A(n20998), .ZN(n15576) );
  OR2_X1 U13858 ( .A1(n17544), .A2(n15558), .ZN(n17538) );
  OR2_X1 U13859 ( .A1(n11216), .A2(n11215), .ZN(n17559) );
  OR2_X1 U13860 ( .A1(n14020), .A2(n14305), .ZN(n21007) );
  INV_X1 U13861 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17569) );
  OR2_X1 U13862 ( .A1(n21082), .A2(n21109), .ZN(n21058) );
  OR2_X1 U13863 ( .A1(n21082), .A2(n21339), .ZN(n21074) );
  AOI22_X1 U13864 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21080), .B1(n21084), 
        .B2(n21087), .ZN(n21108) );
  NAND2_X1 U13865 ( .A1(n21139), .A2(n21165), .ZN(n21164) );
  AOI22_X1 U13866 ( .A1(n14418), .A2(n14415), .B1(n21293), .B2(n14411), .ZN(
        n14453) );
  NAND2_X1 U13867 ( .A1(n21139), .A2(n21257), .ZN(n21178) );
  NAND2_X1 U13868 ( .A1(n21258), .A2(n21165), .ZN(n21223) );
  AOI22_X1 U13869 ( .A1(n21232), .A2(n21229), .B1(n21228), .B2(n21370), .ZN(
        n21256) );
  NAND2_X1 U13870 ( .A1(n21258), .A2(n21257), .ZN(n21300) );
  INV_X1 U13871 ( .A(n21437), .ZN(n21312) );
  OR2_X1 U13872 ( .A1(n21335), .A2(n21287), .ZN(n21366) );
  OR2_X1 U13873 ( .A1(n21415), .A2(n21368), .ZN(n21449) );
  OR2_X1 U13874 ( .A1(n21415), .A2(n21081), .ZN(n21472) );
  INV_X1 U13875 ( .A(n21560), .ZN(n21477) );
  INV_X1 U13876 ( .A(n21530), .ZN(n21547) );
  INV_X1 U13877 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20675) );
  NAND2_X1 U13878 ( .A1(n12264), .A2(n20026), .ZN(n13424) );
  NAND2_X1 U13879 ( .A1(n15993), .A2(n12388), .ZN(n12389) );
  OR2_X1 U13880 ( .A1(n20805), .A2(n12387), .ZN(n19987) );
  INV_X1 U13881 ( .A(n15982), .ZN(n19983) );
  NAND2_X1 U13882 ( .A1(n12797), .A2(n20026), .ZN(n16078) );
  INV_X1 U13883 ( .A(n16078), .ZN(n16080) );
  NAND2_X1 U13884 ( .A1(n16080), .A2(n16873), .ZN(n16072) );
  OR2_X1 U13885 ( .A1(n16191), .A2(n11466), .ZN(n16202) );
  INV_X1 U13886 ( .A(n16191), .ZN(n20001) );
  AND2_X1 U13887 ( .A1(n16202), .A2(n20002), .ZN(n16213) );
  AND2_X1 U13888 ( .A1(n16184), .A2(n13952), .ZN(n20024) );
  NAND2_X1 U13889 ( .A1(n20082), .A2(n20034), .ZN(n20061) );
  OR2_X1 U13890 ( .A1(n20082), .A2(n20799), .ZN(n20084) );
  OR2_X1 U13891 ( .A1(n13427), .A2(n16887), .ZN(n20028) );
  INV_X1 U13892 ( .A(n12276), .ZN(n12277) );
  INV_X1 U13893 ( .A(n16470), .ZN(n17594) );
  INV_X1 U13894 ( .A(n12259), .ZN(n12260) );
  INV_X1 U13895 ( .A(n17606), .ZN(n16748) );
  AOI21_X1 U13896 ( .B1(n16925), .B2(n20026), .A(n13537), .ZN(n16833) );
  OR2_X1 U13897 ( .A1(n20396), .A2(n20244), .ZN(n20173) );
  INV_X1 U13898 ( .A(n20179), .ZN(n20243) );
  AOI211_X2 U13899 ( .C1(n20335), .C2(n20338), .A(n20494), .B(n20334), .ZN(
        n20365) );
  INV_X1 U13900 ( .A(n20394), .ZN(n20426) );
  INV_X1 U13901 ( .A(n20668), .ZN(n20625) );
  INV_X1 U13902 ( .A(n20622), .ZN(n20672) );
  INV_X1 U13903 ( .A(n20745), .ZN(n20674) );
  NOR2_X1 U13904 ( .A1(n19788), .A2(n18705), .ZN(n19958) );
  AOI211_X1 U13905 ( .C1(n17756), .C2(n18101), .A(n17755), .B(n17754), .ZN(
        n17759) );
  INV_X1 U13906 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18881) );
  INV_X1 U13907 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n18375) );
  INV_X1 U13908 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18990) );
  NAND2_X1 U13909 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n18116), .ZN(n18096) );
  NOR2_X2 U13910 ( .A1(n9734), .A2(n16973), .ZN(n18618) );
  NOR2_X1 U13911 ( .A1(n17019), .A2(n17018), .ZN(n18635) );
  NOR3_X1 U13912 ( .A1(n18504), .A2(n18697), .A3(n18505), .ZN(n18642) );
  INV_X1 U13913 ( .A(n18676), .ZN(n18701) );
  INV_X1 U13914 ( .A(n18756), .ZN(n18750) );
  INV_X1 U13915 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19022) );
  INV_X1 U13916 ( .A(n19048), .ZN(n19040) );
  INV_X1 U13917 ( .A(n19255), .ZN(n19249) );
  OR2_X1 U13918 ( .A1(n19323), .A2(n19268), .ZN(n19329) );
  NOR2_X1 U13919 ( .A1(n19354), .A2(n13909), .ZN(n17439) );
  INV_X1 U13920 ( .A(n19667), .ZN(n19741) );
  NAND2_X1 U13921 ( .A1(n19835), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19830) );
  INV_X1 U13922 ( .A(n18101), .ZN(n19839) );
  INV_X1 U13923 ( .A(n19920), .ZN(n19917) );
  INV_X1 U13924 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n21816) );
  NAND2_X1 U13925 ( .A1(n21589), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19909) );
  AND2_X1 U13926 ( .A1(n13369), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15096)
         );
  NOR2_X1 U13927 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13383), .ZN(n17694)
         );
  INV_X1 U13928 ( .A(n17656), .ZN(n17660) );
  INV_X1 U13929 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10744) );
  NOR2_X4 U13930 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13931 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10750) );
  AND2_X2 U13932 ( .A1(n10746), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10756) );
  AND2_X4 U13933 ( .A1(n10755), .A2(n10752), .ZN(n10955) );
  AOI22_X1 U13934 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10748) );
  INV_X2 U13935 ( .A(n10820), .ZN(n13040) );
  AOI22_X1 U13936 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10747) );
  AND2_X4 U13937 ( .A1(n10753), .A2(n10752), .ZN(n13326) );
  AOI22_X1 U13938 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10760) );
  AND2_X2 U13939 ( .A1(n10754), .A2(n10757), .ZN(n10924) );
  AOI22_X1 U13940 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10759) );
  AND2_X2 U13941 ( .A1(n10757), .A2(n13977), .ZN(n10937) );
  AOI22_X1 U13942 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13943 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U13944 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10765) );
  INV_X2 U13945 ( .A(n10762), .ZN(n13165) );
  AOI22_X1 U13946 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U13947 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10763) );
  AOI22_X1 U13948 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13949 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13950 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13951 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10767) );
  AOI22_X1 U13952 ( .A1(n13326), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10776) );
  AOI22_X1 U13953 ( .A1(n13165), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10775) );
  AOI22_X1 U13954 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10825), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10783) );
  AOI22_X1 U13955 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10782) );
  NAND2_X1 U13956 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10779) );
  NAND2_X1 U13957 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10778) );
  AOI22_X1 U13958 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U13959 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13960 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9740), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13961 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10786) );
  AOI22_X1 U13962 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13963 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10792) );
  NOR2_X1 U13964 ( .A1(n11152), .A2(n14290), .ZN(n10796) );
  NAND2_X1 U13965 ( .A1(n10858), .A2(n10796), .ZN(n10797) );
  AOI22_X1 U13966 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n13291), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13967 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13968 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10800) );
  AOI22_X1 U13969 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10799) );
  AOI22_X1 U13970 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13971 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13972 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10773), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10804) );
  AOI22_X1 U13973 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13974 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10810) );
  AOI22_X1 U13975 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10809) );
  AOI22_X1 U13976 ( .A1(n9740), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10937), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10808) );
  AOI22_X1 U13977 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13978 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10815) );
  AOI22_X1 U13979 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10814) );
  AOI22_X1 U13980 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10813) );
  AOI22_X1 U13981 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10812) );
  NAND2_X1 U13982 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10819) );
  NAND2_X1 U13983 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10818) );
  NAND2_X1 U13984 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10817) );
  NAND2_X1 U13985 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10816) );
  NAND2_X1 U13986 ( .A1(n10925), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10824) );
  NAND2_X1 U13987 ( .A1(n13326), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10823) );
  NAND2_X1 U13988 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10822) );
  NAND2_X1 U13989 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10821) );
  NAND2_X1 U13990 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10828) );
  NAND2_X1 U13991 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10827) );
  NAND2_X1 U13992 ( .A1(n10924), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10826) );
  NAND2_X1 U13993 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10833) );
  NAND2_X1 U13994 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10832) );
  NAND2_X1 U13995 ( .A1(n13165), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10831) );
  NAND2_X1 U13996 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10830) );
  NAND2_X1 U13997 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10841) );
  NAND2_X1 U13998 ( .A1(n10825), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10840) );
  NAND2_X1 U13999 ( .A1(n10811), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10839) );
  NAND2_X1 U14000 ( .A1(n10924), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10838) );
  NAND2_X1 U14001 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10845) );
  NAND2_X1 U14002 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10844) );
  NAND2_X1 U14003 ( .A1(n13165), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10843) );
  NAND2_X1 U14004 ( .A1(n10955), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14005 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10849) );
  NAND2_X1 U14006 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10848) );
  NAND2_X1 U14007 ( .A1(n10937), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10847) );
  NAND2_X1 U14008 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U14009 ( .A1(n13326), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10852) );
  NAND2_X1 U14010 ( .A1(n10741), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10851) );
  NAND2_X1 U14011 ( .A1(n13040), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10850) );
  NAND2_X1 U14013 ( .A1(n11016), .A2(n10872), .ZN(n11194) );
  INV_X1 U14014 ( .A(n11194), .ZN(n10861) );
  INV_X4 U14015 ( .A(n10867), .ZN(n11218) );
  NAND2_X1 U14017 ( .A1(n13356), .A2(n13545), .ZN(n13972) );
  NAND2_X1 U14018 ( .A1(n10858), .A2(n10872), .ZN(n13372) );
  NAND2_X1 U14019 ( .A1(n10864), .A2(n11218), .ZN(n17492) );
  NAND2_X1 U14020 ( .A1(n10867), .A2(n11217), .ZN(n14239) );
  NAND2_X1 U14021 ( .A1(n14290), .A2(n11218), .ZN(n11328) );
  OR2_X1 U14022 ( .A1(n10868), .A2(n11224), .ZN(n10869) );
  NOR2_X1 U14023 ( .A1(n10892), .A2(n10871), .ZN(n10879) );
  NAND2_X1 U14024 ( .A1(n11199), .A2(n10873), .ZN(n10875) );
  NAND2_X1 U14025 ( .A1(n10895), .A2(n15586), .ZN(n10878) );
  NAND2_X1 U14026 ( .A1(n21409), .A2(n21329), .ZN(n21294) );
  NAND2_X1 U14027 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21405) );
  NAND2_X1 U14028 ( .A1(n21294), .A2(n21405), .ZN(n21233) );
  INV_X1 U14029 ( .A(n21233), .ZN(n21169) );
  NAND2_X1 U14030 ( .A1(n17567), .A2(n20825), .ZN(n13312) );
  INV_X1 U14031 ( .A(n13312), .ZN(n10977) );
  AND2_X1 U14032 ( .A1(n21475), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10897) );
  AOI21_X1 U14033 ( .B1(n21169), .B2(n10977), .A(n10897), .ZN(n10881) );
  INV_X1 U14034 ( .A(n10882), .ZN(n10883) );
  INV_X1 U14035 ( .A(n21475), .ZN(n10885) );
  MUX2_X1 U14036 ( .A(n10885), .B(n13312), .S(n21329), .Z(n10886) );
  INV_X1 U14037 ( .A(n17492), .ZN(n11110) );
  AND2_X1 U14038 ( .A1(n10888), .A2(n11224), .ZN(n14745) );
  AOI22_X1 U14039 ( .A1(n11203), .A2(n11110), .B1(n14745), .B2(n10890), .ZN(
        n10894) );
  NAND3_X1 U14040 ( .A1(n11338), .A2(n17567), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10891) );
  NOR2_X1 U14041 ( .A1(n10892), .A2(n10891), .ZN(n10893) );
  NAND3_X1 U14042 ( .A1(n10895), .A2(n11217), .A3(n15586), .ZN(n10896) );
  INV_X1 U14043 ( .A(n10897), .ZN(n10898) );
  NAND2_X1 U14044 ( .A1(n10898), .A2(n10880), .ZN(n10899) );
  NAND2_X1 U14045 ( .A1(n10900), .A2(n10899), .ZN(n10901) );
  XNOR2_X1 U14046 ( .A(n21405), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14380) );
  AOI22_X1 U14047 ( .A1(n10977), .A2(n14380), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n21475), .ZN(n10902) );
  INV_X1 U14048 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n21720) );
  AOI22_X1 U14049 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U14050 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10907) );
  AOI22_X1 U14051 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10906) );
  AOI22_X1 U14052 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10905) );
  NAND4_X1 U14053 ( .A1(n10908), .A2(n10907), .A3(n10906), .A4(n10905), .ZN(
        n10914) );
  AOI22_X1 U14054 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U14055 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U14056 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U14057 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10909) );
  NAND4_X1 U14058 ( .A1(n10912), .A2(n10911), .A3(n10910), .A4(n10909), .ZN(
        n10913) );
  INV_X1 U14059 ( .A(n10980), .ZN(n10966) );
  AOI22_X1 U14060 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10966), .B2(n10916), .ZN(n10917) );
  NAND2_X1 U14061 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10945) );
  AOI22_X1 U14062 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13320), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U14063 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U14064 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U14065 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10920) );
  NAND4_X1 U14066 ( .A1(n10923), .A2(n10922), .A3(n10921), .A4(n10920), .ZN(
        n10931) );
  AOI22_X1 U14067 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n10924), .B1(
        n13995), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10929) );
  INV_X1 U14068 ( .A(n13165), .ZN(n10932) );
  AOI22_X1 U14069 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13293), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10928) );
  AOI22_X1 U14070 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9754), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10927) );
  AOI22_X1 U14071 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10926) );
  NAND4_X1 U14072 ( .A1(n10929), .A2(n10928), .A3(n10927), .A4(n10926), .ZN(
        n10930) );
  AOI21_X1 U14073 ( .B1(n10867), .B2(n11024), .A(n20825), .ZN(n10944) );
  AOI22_X1 U14074 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U14075 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10924), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10935) );
  AOI22_X1 U14076 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U14077 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10933) );
  NAND4_X1 U14078 ( .A1(n10936), .A2(n10935), .A3(n10934), .A4(n10933), .ZN(
        n10943) );
  AOI22_X1 U14079 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U14080 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14081 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14082 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10938) );
  NAND4_X1 U14083 ( .A1(n10941), .A2(n10940), .A3(n10939), .A4(n10938), .ZN(
        n10942) );
  NAND2_X1 U14084 ( .A1(n10866), .A2(n11109), .ZN(n10946) );
  NAND3_X1 U14085 ( .A1(n10945), .A2(n10944), .A3(n10946), .ZN(n12839) );
  INV_X1 U14086 ( .A(n12839), .ZN(n10951) );
  NOR2_X1 U14087 ( .A1(n10981), .A2(n11109), .ZN(n10953) );
  INV_X1 U14088 ( .A(n11024), .ZN(n10947) );
  MUX2_X1 U14089 ( .A(n10953), .B(n10949), .S(n10947), .Z(n10948) );
  AND2_X1 U14090 ( .A1(n11022), .A2(n11105), .ZN(n10950) );
  INV_X1 U14091 ( .A(n10953), .ZN(n10969) );
  NAND2_X1 U14092 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10968) );
  AOI22_X1 U14093 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14094 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U14095 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14096 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14097 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10965) );
  AOI22_X1 U14098 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U14099 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U14100 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U14101 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10960) );
  NAND4_X1 U14102 ( .A1(n10963), .A2(n10962), .A3(n10961), .A4(n10960), .ZN(
        n10964) );
  NAND2_X1 U14103 ( .A1(n10966), .A2(n11015), .ZN(n10967) );
  INV_X1 U14104 ( .A(n10981), .ZN(n10972) );
  INV_X1 U14105 ( .A(n21405), .ZN(n21078) );
  INV_X1 U14106 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21234) );
  NAND2_X1 U14107 ( .A1(n21234), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n21136) );
  INV_X1 U14108 ( .A(n21136), .ZN(n10975) );
  NAND2_X1 U14109 ( .A1(n21078), .A2(n10975), .ZN(n14308) );
  OAI21_X1 U14110 ( .B1(n21405), .B2(n21166), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U14111 ( .A1(n14308), .A2(n10976), .ZN(n21168) );
  AOI22_X1 U14112 ( .A1(n21168), .A2(n10977), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n21475), .ZN(n10978) );
  AOI22_X1 U14113 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14114 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14115 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10983) );
  AOI22_X1 U14116 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10982) );
  NAND4_X1 U14117 ( .A1(n10985), .A2(n10984), .A3(n10983), .A4(n10982), .ZN(
        n10991) );
  AOI22_X1 U14118 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10954), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10989) );
  AOI22_X1 U14119 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10988) );
  AOI22_X1 U14120 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10987) );
  INV_X2 U14121 ( .A(n10820), .ZN(n13284) );
  AOI22_X1 U14122 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10986) );
  NAND4_X1 U14123 ( .A1(n10989), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n10990) );
  AOI22_X1 U14124 ( .A1(n11186), .A2(n10995), .B1(n11167), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10992) );
  NAND2_X1 U14125 ( .A1(n11015), .A2(n11024), .ZN(n11038) );
  NAND2_X1 U14126 ( .A1(n11038), .A2(n11039), .ZN(n11037) );
  NAND2_X1 U14127 ( .A1(n11037), .A2(n10995), .ZN(n11069) );
  OAI211_X1 U14128 ( .C1(n10995), .C2(n11037), .A(n11069), .B(n11110), .ZN(
        n10996) );
  AOI22_X1 U14129 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14130 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14131 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14132 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10997) );
  NAND4_X1 U14133 ( .A1(n11000), .A2(n10999), .A3(n10998), .A4(n10997), .ZN(
        n11006) );
  AOI22_X1 U14134 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14135 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11003) );
  INV_X1 U14136 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21813) );
  AOI22_X1 U14137 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14138 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11001) );
  NAND4_X1 U14139 ( .A1(n11004), .A2(n11003), .A3(n11002), .A4(n11001), .ZN(
        n11005) );
  NAND2_X1 U14140 ( .A1(n11186), .A2(n11013), .ZN(n11008) );
  NAND2_X1 U14141 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U14142 ( .A1(n11009), .A2(n11065), .ZN(n11012) );
  INV_X1 U14143 ( .A(n11065), .ZN(n11011) );
  INV_X1 U14144 ( .A(n11013), .ZN(n11068) );
  XNOR2_X1 U14145 ( .A(n11069), .B(n11068), .ZN(n11014) );
  NAND2_X1 U14146 ( .A1(n12832), .A2(n11217), .ZN(n11021) );
  XNOR2_X1 U14147 ( .A(n11015), .B(n11024), .ZN(n11018) );
  OAI211_X1 U14148 ( .C1(n11018), .C2(n17492), .A(n11017), .B(n14729), .ZN(
        n11019) );
  INV_X1 U14149 ( .A(n11019), .ZN(n11020) );
  NAND2_X1 U14150 ( .A1(n11021), .A2(n11020), .ZN(n11032) );
  NAND2_X1 U14151 ( .A1(n12840), .A2(n12839), .ZN(n11030) );
  OR2_X1 U14152 ( .A1(n17492), .A2(n11024), .ZN(n11025) );
  NAND2_X1 U14153 ( .A1(n11025), .A2(n11040), .ZN(n13620) );
  INV_X1 U14154 ( .A(n12840), .ZN(n11028) );
  NOR2_X1 U14155 ( .A1(n12839), .A2(n13620), .ZN(n11027) );
  OAI21_X1 U14156 ( .B1(n13620), .B2(n13621), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11026) );
  AOI21_X1 U14157 ( .B1(n11028), .B2(n11027), .A(n11026), .ZN(n11029) );
  OAI21_X1 U14158 ( .B1(n11030), .B2(n13620), .A(n11029), .ZN(n11031) );
  XNOR2_X1 U14159 ( .A(n11032), .B(n11031), .ZN(n13633) );
  NAND2_X1 U14160 ( .A1(n13633), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11034) );
  INV_X1 U14161 ( .A(n11031), .ZN(n13622) );
  NAND2_X1 U14162 ( .A1(n11032), .A2(n13622), .ZN(n11033) );
  NAND2_X1 U14163 ( .A1(n11034), .A2(n11033), .ZN(n11045) );
  XNOR2_X1 U14164 ( .A(n11045), .B(n13885), .ZN(n13872) );
  NAND2_X1 U14165 ( .A1(n9746), .A2(n13621), .ZN(n11044) );
  OAI21_X1 U14166 ( .B1(n11039), .B2(n11038), .A(n11037), .ZN(n11042) );
  INV_X1 U14167 ( .A(n11040), .ZN(n11041) );
  AOI21_X1 U14168 ( .B1(n11042), .B2(n11110), .A(n11041), .ZN(n11043) );
  NAND2_X1 U14169 ( .A1(n11044), .A2(n11043), .ZN(n13871) );
  NAND2_X1 U14170 ( .A1(n13872), .A2(n13871), .ZN(n11047) );
  NAND2_X1 U14171 ( .A1(n11045), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11046) );
  INV_X1 U14172 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U14173 ( .A1(n11049), .A2(n14128), .ZN(n11048) );
  AOI22_X1 U14174 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U14175 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13293), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U14176 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U14177 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11053) );
  NAND4_X1 U14178 ( .A1(n11056), .A2(n11055), .A3(n11054), .A4(n11053), .ZN(
        n11062) );
  AOI22_X1 U14179 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14180 ( .A1(n10954), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11059) );
  AOI22_X1 U14181 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U14182 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11057) );
  NAND4_X1 U14183 ( .A1(n11060), .A2(n11059), .A3(n11058), .A4(n11057), .ZN(
        n11061) );
  NAND2_X1 U14184 ( .A1(n11186), .A2(n11070), .ZN(n11064) );
  NAND2_X1 U14185 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11063) );
  NOR2_X1 U14186 ( .A1(n11069), .A2(n11068), .ZN(n11071) );
  NAND2_X1 U14187 ( .A1(n11071), .A2(n11070), .ZN(n11096) );
  OAI211_X1 U14188 ( .C1(n11071), .C2(n11070), .A(n11096), .B(n11110), .ZN(
        n11072) );
  OAI21_X1 U14189 ( .B1(n12867), .B2(n11104), .A(n11072), .ZN(n11073) );
  INV_X1 U14190 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21873) );
  XNOR2_X1 U14191 ( .A(n11073), .B(n21873), .ZN(n17526) );
  NAND2_X1 U14192 ( .A1(n11073), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11074) );
  AOI22_X1 U14193 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14194 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14195 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14196 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11075) );
  NAND4_X1 U14197 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11084) );
  AOI22_X1 U14198 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14199 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14200 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14201 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11079) );
  NAND4_X1 U14202 ( .A1(n11082), .A2(n11081), .A3(n11080), .A4(n11079), .ZN(
        n11083) );
  NAND2_X1 U14203 ( .A1(n11186), .A2(n11097), .ZN(n11086) );
  NAND2_X1 U14204 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14205 ( .A1(n11087), .A2(n10742), .ZN(n11088) );
  OR2_X1 U14206 ( .A1(n12868), .A2(n11104), .ZN(n11091) );
  XNOR2_X1 U14207 ( .A(n11096), .B(n11097), .ZN(n11089) );
  NAND2_X1 U14208 ( .A1(n11089), .A2(n11110), .ZN(n11090) );
  NAND2_X1 U14209 ( .A1(n11091), .A2(n11090), .ZN(n11092) );
  NAND2_X1 U14210 ( .A1(n11092), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17519) );
  NAND2_X1 U14211 ( .A1(n11186), .A2(n11109), .ZN(n11094) );
  NAND2_X1 U14212 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11093) );
  NAND2_X1 U14213 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  INV_X1 U14214 ( .A(n11096), .ZN(n11098) );
  NAND2_X1 U14215 ( .A1(n11098), .A2(n11097), .ZN(n11108) );
  XNOR2_X1 U14216 ( .A(n11108), .B(n11109), .ZN(n11099) );
  NAND2_X1 U14217 ( .A1(n11099), .A2(n11110), .ZN(n11100) );
  NAND2_X1 U14218 ( .A1(n11101), .A2(n11100), .ZN(n11102) );
  INV_X1 U14219 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17537) );
  NAND2_X1 U14220 ( .A1(n11102), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11103) );
  NOR2_X1 U14221 ( .A1(n11105), .A2(n11104), .ZN(n11106) );
  INV_X1 U14222 ( .A(n11108), .ZN(n11111) );
  NAND3_X1 U14223 ( .A1(n11111), .A2(n11110), .A3(n11109), .ZN(n11112) );
  INV_X1 U14224 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15524) );
  INV_X1 U14225 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15536) );
  NAND2_X1 U14226 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11114) );
  INV_X1 U14227 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15515) );
  AND2_X1 U14228 ( .A1(n10154), .A2(n15515), .ZN(n11115) );
  NOR2_X2 U14229 ( .A1(n15314), .A2(n11115), .ZN(n15281) );
  OR2_X1 U14230 ( .A1(n11121), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15283) );
  NAND2_X1 U14231 ( .A1(n15283), .A2(n11116), .ZN(n15291) );
  INV_X1 U14232 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21704) );
  OR2_X1 U14233 ( .A1(n11121), .A2(n15536), .ZN(n15326) );
  NOR2_X1 U14234 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11119) );
  OR2_X1 U14235 ( .A1(n11121), .A2(n11119), .ZN(n15323) );
  NAND2_X1 U14236 ( .A1(n15326), .A2(n15323), .ZN(n15279) );
  INV_X1 U14237 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15491) );
  INV_X1 U14238 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11281) );
  INV_X1 U14239 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11120) );
  OR2_X1 U14240 ( .A1(n10154), .A2(n15515), .ZN(n11123) );
  NAND2_X1 U14241 ( .A1(n15313), .A2(n11123), .ZN(n15280) );
  NOR2_X2 U14242 ( .A1(n11124), .A2(n15280), .ZN(n11125) );
  INV_X1 U14243 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11349) );
  NAND2_X1 U14244 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15244) );
  INV_X1 U14245 ( .A(n15244), .ZN(n11127) );
  INV_X1 U14246 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15456) );
  NAND2_X1 U14247 ( .A1(n15456), .A2(n11349), .ZN(n15242) );
  NAND2_X1 U14248 ( .A1(n11128), .A2(n10735), .ZN(n15233) );
  NAND3_X1 U14249 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15399) );
  INV_X1 U14250 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15209) );
  INV_X1 U14251 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15398) );
  INV_X1 U14252 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11305) );
  NAND3_X1 U14253 ( .A1(n15209), .A2(n15398), .A3(n11305), .ZN(n15176) );
  NOR2_X1 U14254 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15381) );
  NAND2_X1 U14255 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11372) );
  AND2_X1 U14256 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13308) );
  INV_X1 U14257 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12812) );
  NAND3_X1 U14258 ( .A1(n11130), .A2(n12812), .A3(n10729), .ZN(n11131) );
  XNOR2_X1 U14259 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14260 ( .A1(n21329), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11157) );
  NAND2_X1 U14261 ( .A1(n11146), .A2(n11145), .ZN(n11133) );
  NAND2_X1 U14262 ( .A1(n21409), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14263 ( .A1(n11133), .A2(n11132), .ZN(n11148) );
  XNOR2_X1 U14264 ( .A(n15602), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14265 ( .A1(n11148), .A2(n11147), .ZN(n11135) );
  NAND2_X1 U14266 ( .A1(n21166), .A2(n15602), .ZN(n11134) );
  XNOR2_X1 U14267 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11143) );
  NOR2_X1 U14268 ( .A1(n14004), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11136) );
  INV_X1 U14269 ( .A(n11142), .ZN(n11138) );
  NOR2_X1 U14270 ( .A1(n17569), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11137) );
  INV_X1 U14271 ( .A(n11141), .ZN(n11139) );
  XNOR2_X1 U14272 ( .A(n11144), .B(n11143), .ZN(n11174) );
  XNOR2_X1 U14273 ( .A(n11146), .B(n11145), .ZN(n11156) );
  XNOR2_X1 U14274 ( .A(n11148), .B(n11147), .ZN(n11151) );
  NOR4_X1 U14275 ( .A1(n11179), .A2(n11174), .A3(n11156), .A4(n11151), .ZN(
        n11149) );
  NOR2_X1 U14276 ( .A1(n11189), .A2(n11149), .ZN(n13555) );
  NAND2_X1 U14277 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21574) );
  AND2_X1 U14278 ( .A1(n13555), .A2(n21574), .ZN(n13352) );
  OAI21_X1 U14279 ( .B1(n14157), .B2(n14234), .A(n13352), .ZN(n11198) );
  NAND2_X1 U14280 ( .A1(n11152), .A2(n11218), .ZN(n11150) );
  NAND2_X1 U14281 ( .A1(n11150), .A2(n10864), .ZN(n11172) );
  INV_X1 U14282 ( .A(n11151), .ZN(n11168) );
  NAND2_X1 U14283 ( .A1(n11186), .A2(n11168), .ZN(n11171) );
  NAND2_X1 U14284 ( .A1(n11186), .A2(n11217), .ZN(n11154) );
  NAND2_X1 U14285 ( .A1(n11152), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U14286 ( .A1(n11155), .A2(n11217), .ZN(n11178) );
  INV_X1 U14287 ( .A(n11156), .ZN(n11166) );
  OAI21_X1 U14288 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21329), .A(
        n11157), .ZN(n11158) );
  INV_X1 U14289 ( .A(n11158), .ZN(n11159) );
  OAI211_X1 U14290 ( .C1(n10868), .C2(n10867), .A(n11172), .B(n11159), .ZN(
        n11162) );
  NAND2_X1 U14291 ( .A1(n11186), .A2(n11159), .ZN(n11160) );
  NAND2_X1 U14292 ( .A1(n11187), .A2(n11160), .ZN(n11161) );
  OAI211_X1 U14293 ( .C1(n11163), .C2(n11166), .A(n11162), .B(n11161), .ZN(
        n11165) );
  NAND2_X1 U14294 ( .A1(n11163), .A2(n11166), .ZN(n11164) );
  OAI211_X1 U14295 ( .C1(n11178), .C2(n11166), .A(n11165), .B(n11164), .ZN(
        n11170) );
  OAI211_X1 U14296 ( .C1(n11168), .C2(n11180), .A(n11171), .B(n11172), .ZN(
        n11169) );
  NAND2_X1 U14297 ( .A1(n11180), .A2(n11174), .ZN(n11173) );
  INV_X1 U14298 ( .A(n11187), .ZN(n11175) );
  NAND2_X1 U14299 ( .A1(n11180), .A2(n11179), .ZN(n11176) );
  NAND2_X1 U14300 ( .A1(n11177), .A2(n11176), .ZN(n11185) );
  INV_X1 U14301 ( .A(n11178), .ZN(n11183) );
  INV_X1 U14302 ( .A(n11179), .ZN(n11181) );
  NOR2_X1 U14303 ( .A1(n11181), .A2(n11180), .ZN(n11182) );
  AOI22_X1 U14304 ( .A1(n11183), .A2(n11182), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20825), .ZN(n11184) );
  NAND2_X1 U14305 ( .A1(n11185), .A2(n11184), .ZN(n11191) );
  INV_X1 U14306 ( .A(n11189), .ZN(n11190) );
  NAND2_X1 U14307 ( .A1(n11191), .A2(n11190), .ZN(n11192) );
  NOR2_X1 U14308 ( .A1(n11194), .A2(n11195), .ZN(n13986) );
  INV_X1 U14309 ( .A(n13986), .ZN(n13973) );
  INV_X1 U14310 ( .A(n21574), .ZN(n21478) );
  NOR2_X1 U14311 ( .A1(n13973), .A2(n21478), .ZN(n17493) );
  OAI22_X1 U14312 ( .A1(n17493), .A2(n10867), .B1(n14234), .B2(n17492), .ZN(
        n11196) );
  NAND2_X1 U14313 ( .A1(n11196), .A2(n13372), .ZN(n11197) );
  NAND2_X1 U14314 ( .A1(n11200), .A2(n11199), .ZN(n13556) );
  NAND2_X1 U14315 ( .A1(n10889), .A2(n11218), .ZN(n11201) );
  NAND2_X1 U14316 ( .A1(n11201), .A2(n17492), .ZN(n11202) );
  NAND2_X1 U14317 ( .A1(n10895), .A2(n11202), .ZN(n11337) );
  INV_X1 U14318 ( .A(n11203), .ZN(n11205) );
  AND2_X1 U14319 ( .A1(n11205), .A2(n11204), .ZN(n11334) );
  NAND3_X1 U14320 ( .A1(n11334), .A2(n11017), .A3(n11206), .ZN(n17482) );
  NAND2_X1 U14321 ( .A1(n11337), .A2(n13348), .ZN(n11207) );
  NAND2_X1 U14322 ( .A1(n13556), .A2(n11207), .ZN(n13988) );
  NOR2_X1 U14323 ( .A1(n15586), .A2(n14157), .ZN(n11344) );
  INV_X1 U14324 ( .A(n11344), .ZN(n11208) );
  INV_X1 U14325 ( .A(n11354), .ZN(n11216) );
  NAND2_X1 U14326 ( .A1(n10868), .A2(n10888), .ZN(n11211) );
  NAND2_X1 U14327 ( .A1(n13348), .A2(n11211), .ZN(n13551) );
  OAI21_X1 U14328 ( .B1(n10866), .B2(n11210), .A(n13551), .ZN(n11214) );
  NOR2_X1 U14329 ( .A1(n11214), .A2(n11213), .ZN(n11215) );
  AND2_X4 U14330 ( .A1(n11218), .A2(n11217), .ZN(n13634) );
  INV_X1 U14331 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11219) );
  NAND2_X1 U14332 ( .A1(n11235), .A2(n11219), .ZN(n11222) );
  INV_X1 U14333 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n11220) );
  NAND2_X1 U14334 ( .A1(n13634), .A2(n11220), .ZN(n11221) );
  NAND3_X1 U14335 ( .A1(n11222), .A2(n11333), .A3(n11221), .ZN(n11223) );
  NAND2_X1 U14336 ( .A1(n11235), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n11226) );
  BUF_X4 U14337 ( .A(n11224), .Z(n11333) );
  INV_X1 U14338 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14246) );
  NAND2_X1 U14339 ( .A1(n9747), .A2(n14246), .ZN(n11225) );
  NAND2_X1 U14340 ( .A1(n11226), .A2(n11225), .ZN(n13628) );
  INV_X1 U14341 ( .A(n13877), .ZN(n11234) );
  INV_X2 U14342 ( .A(n11227), .ZN(n11314) );
  INV_X1 U14343 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n11228) );
  NAND2_X1 U14344 ( .A1(n11314), .A2(n11228), .ZN(n11232) );
  NAND2_X1 U14345 ( .A1(n11235), .A2(n13885), .ZN(n11230) );
  NAND2_X1 U14346 ( .A1(n13634), .A2(n11228), .ZN(n11229) );
  NAND3_X1 U14347 ( .A1(n11230), .A2(n11333), .A3(n11229), .ZN(n11231) );
  MUX2_X1 U14348 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n11236) );
  OAI21_X1 U14349 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13629), .A(
        n11236), .ZN(n14102) );
  NAND2_X1 U14350 ( .A1(n9747), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11237) );
  NAND2_X1 U14351 ( .A1(n11235), .A2(n11237), .ZN(n11240) );
  INV_X1 U14352 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U14353 ( .A1(n13634), .A2(n11238), .ZN(n11239) );
  NAND2_X1 U14354 ( .A1(n11240), .A2(n11239), .ZN(n11241) );
  OAI21_X1 U14355 ( .B1(n11227), .B2(P1_EBX_REG_4__SCAN_IN), .A(n11241), .ZN(
        n14211) );
  NAND2_X1 U14356 ( .A1(n9747), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11243) );
  OAI211_X1 U14357 ( .C1(n11242), .C2(P1_EBX_REG_5__SCAN_IN), .A(n11235), .B(
        n11243), .ZN(n11244) );
  OAI21_X1 U14358 ( .B1(n11311), .B2(P1_EBX_REG_5__SCAN_IN), .A(n11244), .ZN(
        n17550) );
  NAND2_X1 U14359 ( .A1(n11246), .A2(n11245), .ZN(n14336) );
  INV_X1 U14360 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n11247) );
  NAND2_X1 U14361 ( .A1(n11314), .A2(n11247), .ZN(n11251) );
  NAND2_X1 U14362 ( .A1(n11333), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14363 ( .A1(n11235), .A2(n11248), .ZN(n11249) );
  OAI21_X1 U14364 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(n11242), .A(n11249), .ZN(
        n11250) );
  NAND2_X1 U14365 ( .A1(n9747), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11253) );
  OAI211_X1 U14366 ( .C1(n11242), .C2(P1_EBX_REG_7__SCAN_IN), .A(n11235), .B(
        n11253), .ZN(n11254) );
  OAI21_X1 U14367 ( .B1(n11311), .B2(P1_EBX_REG_7__SCAN_IN), .A(n11254), .ZN(
        n14364) );
  NAND2_X1 U14368 ( .A1(n11333), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11255) );
  NAND2_X1 U14369 ( .A1(n11235), .A2(n11255), .ZN(n11258) );
  INV_X1 U14370 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U14371 ( .A1(n13634), .A2(n11256), .ZN(n11257) );
  NAND2_X1 U14372 ( .A1(n11258), .A2(n11257), .ZN(n11259) );
  OAI21_X1 U14373 ( .B1(n11227), .B2(P1_EBX_REG_8__SCAN_IN), .A(n11259), .ZN(
        n14455) );
  NAND2_X1 U14374 ( .A1(n11333), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11260) );
  OAI211_X1 U14375 ( .C1(n11242), .C2(P1_EBX_REG_9__SCAN_IN), .A(n11235), .B(
        n11260), .ZN(n11261) );
  OAI21_X1 U14376 ( .B1(n11311), .B2(P1_EBX_REG_9__SCAN_IN), .A(n11261), .ZN(
        n15573) );
  NAND2_X1 U14377 ( .A1(n11263), .A2(n11262), .ZN(n15019) );
  INV_X1 U14378 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15081) );
  NAND2_X1 U14379 ( .A1(n11314), .A2(n15081), .ZN(n11267) );
  INV_X1 U14380 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15556) );
  NAND2_X1 U14381 ( .A1(n11235), .A2(n15556), .ZN(n11265) );
  NAND2_X1 U14382 ( .A1(n13634), .A2(n15081), .ZN(n11264) );
  NAND3_X1 U14383 ( .A1(n11265), .A2(n11333), .A3(n11264), .ZN(n11266) );
  MUX2_X1 U14384 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11269) );
  OR2_X1 U14385 ( .A1(n13629), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14386 ( .A1(n9747), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11270) );
  NAND2_X1 U14387 ( .A1(n11235), .A2(n11270), .ZN(n11272) );
  INV_X1 U14388 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15078) );
  NAND2_X1 U14389 ( .A1(n13634), .A2(n15078), .ZN(n11271) );
  NAND2_X1 U14390 ( .A1(n11272), .A2(n11271), .ZN(n11273) );
  OAI21_X1 U14391 ( .B1(n11227), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11273), .ZN(
        n14983) );
  NAND2_X1 U14392 ( .A1(n14982), .A2(n14983), .ZN(n14965) );
  MUX2_X1 U14393 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n11274) );
  OAI21_X1 U14394 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n13629), .A(
        n11274), .ZN(n14966) );
  OR2_X2 U14395 ( .A1(n14965), .A2(n14966), .ZN(n14968) );
  INV_X1 U14396 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U14397 ( .A1(n11314), .A2(n11275), .ZN(n11278) );
  NAND2_X1 U14398 ( .A1(n11235), .A2(n15515), .ZN(n11276) );
  OAI211_X1 U14399 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n11242), .A(n11276), .B(
        n9747), .ZN(n11277) );
  MUX2_X1 U14400 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11280) );
  OR2_X1 U14401 ( .A1(n13629), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11279) );
  AND2_X2 U14402 ( .A1(n14948), .A2(n14931), .ZN(n14933) );
  NAND2_X1 U14403 ( .A1(n11235), .A2(n11281), .ZN(n11282) );
  OAI211_X1 U14404 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n11242), .A(n11282), .B(
        n9747), .ZN(n11283) );
  OAI21_X1 U14405 ( .B1(P1_EBX_REG_16__SCAN_IN), .B2(n11227), .A(n11283), .ZN(
        n14919) );
  INV_X1 U14406 ( .A(n14918), .ZN(n11286) );
  MUX2_X1 U14407 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n11284) );
  OAI21_X1 U14408 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n13629), .A(
        n11284), .ZN(n14906) );
  INV_X1 U14409 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n11287) );
  NAND2_X1 U14410 ( .A1(n11314), .A2(n11287), .ZN(n11290) );
  NAND2_X1 U14411 ( .A1(n11235), .A2(n11349), .ZN(n11288) );
  OAI211_X1 U14412 ( .C1(P1_EBX_REG_18__SCAN_IN), .C2(n11242), .A(n11288), .B(
        n9747), .ZN(n11289) );
  MUX2_X1 U14413 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11291) );
  OAI21_X1 U14414 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n13629), .A(
        n11291), .ZN(n14878) );
  NAND2_X1 U14415 ( .A1(n9747), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11292) );
  NAND2_X1 U14416 ( .A1(n11235), .A2(n11292), .ZN(n11295) );
  INV_X1 U14417 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n11293) );
  NAND2_X1 U14418 ( .A1(n13634), .A2(n11293), .ZN(n11294) );
  NAND2_X1 U14419 ( .A1(n11295), .A2(n11294), .ZN(n11296) );
  OAI21_X1 U14420 ( .B1(n11227), .B2(P1_EBX_REG_20__SCAN_IN), .A(n11296), .ZN(
        n14866) );
  MUX2_X1 U14421 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n11297) );
  OAI21_X1 U14422 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n13629), .A(
        n11297), .ZN(n14850) );
  NOR2_X2 U14423 ( .A1(n14849), .A2(n14850), .ZN(n14835) );
  INV_X1 U14424 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n11298) );
  NAND2_X1 U14425 ( .A1(n11314), .A2(n11298), .ZN(n11301) );
  INV_X1 U14426 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U14427 ( .A1(n11235), .A2(n15435), .ZN(n11299) );
  OAI211_X1 U14428 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n11242), .A(n11299), .B(
        n9747), .ZN(n11300) );
  INV_X1 U14429 ( .A(n14837), .ZN(n11302) );
  AND2_X2 U14430 ( .A1(n14835), .A2(n11302), .ZN(n14836) );
  MUX2_X1 U14431 ( .A(n11311), .B(n9747), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11304) );
  OR2_X1 U14432 ( .A1(n13629), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11303) );
  AND2_X2 U14433 ( .A1(n14836), .A2(n14819), .ZN(n14821) );
  NAND2_X1 U14434 ( .A1(n11235), .A2(n11305), .ZN(n11306) );
  OAI211_X1 U14435 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n11242), .A(n11306), .B(
        n11333), .ZN(n11307) );
  OAI21_X1 U14436 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n11227), .A(n11307), .ZN(
        n14808) );
  NAND2_X1 U14437 ( .A1(n14821), .A2(n14808), .ZN(n14807) );
  MUX2_X1 U14438 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11308) );
  OAI21_X1 U14439 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n13629), .A(
        n11308), .ZN(n14802) );
  NOR2_X2 U14440 ( .A1(n14807), .A2(n14802), .ZN(n14781) );
  INV_X1 U14441 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15199) );
  NAND2_X1 U14442 ( .A1(n11235), .A2(n15199), .ZN(n11309) );
  OAI211_X1 U14443 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n11242), .A(n11309), .B(
        n9747), .ZN(n11310) );
  OAI21_X1 U14444 ( .B1(P1_EBX_REG_26__SCAN_IN), .B2(n11227), .A(n11310), .ZN(
        n14782) );
  MUX2_X1 U14445 ( .A(n11311), .B(n11333), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n11312) );
  OAI21_X1 U14446 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n13629), .A(
        n11312), .ZN(n14778) );
  INV_X1 U14447 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U14448 ( .A1(n11314), .A2(n11313), .ZN(n11317) );
  INV_X1 U14449 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15180) );
  NAND2_X1 U14450 ( .A1(n11235), .A2(n15180), .ZN(n11315) );
  OAI211_X1 U14451 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n11242), .A(n11315), .B(
        n9747), .ZN(n11316) );
  AND2_X1 U14452 ( .A1(n11317), .A2(n11316), .ZN(n14761) );
  INV_X1 U14453 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14743) );
  NAND2_X1 U14454 ( .A1(n13634), .A2(n14743), .ZN(n11319) );
  OR2_X1 U14455 ( .A1(n13629), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U14456 ( .A1(n11318), .A2(n11319), .ZN(n11320) );
  MUX2_X1 U14457 ( .A(n11319), .B(n11320), .S(n11333), .Z(n14722) );
  OAI22_X1 U14458 ( .A1(n14724), .A2(n9747), .B1(n14759), .B2(n11320), .ZN(
        n11322) );
  AND2_X1 U14459 ( .A1(n11242), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11321) );
  AOI21_X1 U14460 ( .B1(n13629), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11321), .ZN(
        n12805) );
  XNOR2_X1 U14461 ( .A(n11322), .B(n12805), .ZN(n15059) );
  NAND2_X1 U14462 ( .A1(n11324), .A2(n14157), .ZN(n11325) );
  OAI21_X1 U14463 ( .B1(n11210), .B2(n14306), .A(n11325), .ZN(n11326) );
  INV_X1 U14464 ( .A(n11017), .ZN(n11327) );
  NAND2_X1 U14465 ( .A1(n11327), .A2(n13629), .ZN(n11332) );
  INV_X1 U14466 ( .A(n14239), .ZN(n11330) );
  INV_X1 U14467 ( .A(n11328), .ZN(n11329) );
  AOI21_X1 U14468 ( .B1(n11330), .B2(n10868), .A(n11329), .ZN(n11331) );
  OAI21_X1 U14469 ( .B1(n11334), .B2(n11333), .A(n11345), .ZN(n11335) );
  INV_X1 U14470 ( .A(n11335), .ZN(n11336) );
  AND3_X1 U14471 ( .A1(n11337), .A2(n10887), .A3(n11336), .ZN(n13975) );
  NAND2_X1 U14472 ( .A1(n13975), .A2(n11338), .ZN(n11339) );
  NAND3_X1 U14473 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11341) );
  NAND2_X1 U14474 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11340) );
  NOR2_X1 U14475 ( .A1(n11341), .A2(n11340), .ZN(n15551) );
  AND2_X1 U14476 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14477 ( .A1(n15551), .A2(n11342), .ZN(n15514) );
  NAND2_X1 U14478 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17556) );
  NOR2_X1 U14479 ( .A1(n21873), .A2(n17556), .ZN(n14460) );
  INV_X1 U14480 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13885) );
  NOR2_X1 U14481 ( .A1(n13885), .A2(n11219), .ZN(n14131) );
  NAND2_X1 U14482 ( .A1(n14460), .A2(n14131), .ZN(n14462) );
  NOR2_X1 U14483 ( .A1(n15514), .A2(n14462), .ZN(n11357) );
  AND2_X1 U14484 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11357), .ZN(
        n11343) );
  NAND2_X1 U14485 ( .A1(n13882), .A2(n11343), .ZN(n11348) );
  NAND2_X1 U14486 ( .A1(n11345), .A2(n11344), .ZN(n13990) );
  INV_X1 U14487 ( .A(n13990), .ZN(n13553) );
  INV_X1 U14488 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21835) );
  OAI21_X1 U14489 ( .B1(n21835), .B2(n11219), .A(n13885), .ZN(n14133) );
  NAND2_X1 U14490 ( .A1(n14133), .A2(n14460), .ZN(n15557) );
  NOR2_X1 U14491 ( .A1(n15514), .A2(n15557), .ZN(n11360) );
  INV_X1 U14492 ( .A(n11360), .ZN(n11346) );
  OR2_X1 U14493 ( .A1(n15533), .A2(n11346), .ZN(n11347) );
  NAND2_X1 U14494 ( .A1(n11348), .A2(n11347), .ZN(n15520) );
  NAND2_X1 U14495 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15478) );
  NOR2_X1 U14496 ( .A1(n15478), .A2(n11349), .ZN(n11350) );
  AND3_X1 U14497 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15473) );
  NAND2_X1 U14498 ( .A1(n11350), .A2(n15473), .ZN(n11362) );
  INV_X1 U14499 ( .A(n11362), .ZN(n11351) );
  NAND2_X1 U14500 ( .A1(n15480), .A2(n11351), .ZN(n15466) );
  NOR2_X1 U14501 ( .A1(n15466), .A2(n15244), .ZN(n15439) );
  NAND2_X1 U14502 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11367) );
  INV_X1 U14503 ( .A(n11367), .ZN(n11352) );
  NAND2_X1 U14504 ( .A1(n15439), .A2(n11352), .ZN(n15428) );
  INV_X1 U14505 ( .A(n15390), .ZN(n15371) );
  NAND3_X1 U14506 ( .A1(n15371), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10636), .ZN(n12813) );
  INV_X1 U14507 ( .A(n15533), .ZN(n13873) );
  OR2_X2 U14508 ( .A1(n17547), .A2(n13873), .ZN(n15477) );
  INV_X1 U14509 ( .A(n15477), .ZN(n15563) );
  INV_X1 U14510 ( .A(n13882), .ZN(n11353) );
  NAND2_X1 U14511 ( .A1(n11353), .A2(n15533), .ZN(n21001) );
  INV_X1 U14512 ( .A(n21001), .ZN(n11370) );
  NAND2_X1 U14513 ( .A1(n13882), .A2(n21835), .ZN(n11356) );
  OR2_X2 U14514 ( .A1(n13312), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20904) );
  OR2_X1 U14515 ( .A1(n11354), .A2(n17539), .ZN(n11355) );
  INV_X1 U14516 ( .A(n11357), .ZN(n11358) );
  NAND2_X1 U14517 ( .A1(n17547), .A2(n11358), .ZN(n11359) );
  OAI211_X1 U14518 ( .C1(n11360), .C2(n15533), .A(n14464), .B(n11359), .ZN(
        n11361) );
  INV_X1 U14519 ( .A(n11361), .ZN(n11364) );
  NAND2_X1 U14520 ( .A1(n15477), .A2(n11362), .ZN(n11363) );
  INV_X1 U14521 ( .A(n14464), .ZN(n11365) );
  NOR2_X1 U14522 ( .A1(n15533), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11366) );
  AOI21_X1 U14523 ( .B1(n15477), .B2(n11367), .A(n11366), .ZN(n11368) );
  AOI22_X1 U14524 ( .A1(n21003), .A2(n15399), .B1(n13882), .B2(n15209), .ZN(
        n11369) );
  NOR2_X1 U14525 ( .A1(n15412), .A2(n15477), .ZN(n12811) );
  INV_X1 U14526 ( .A(n12811), .ZN(n11371) );
  NOR2_X1 U14527 ( .A1(n15412), .A2(n15199), .ZN(n15402) );
  AOI21_X1 U14528 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15402), .A(
        n12811), .ZN(n15393) );
  AOI21_X1 U14529 ( .B1(n11372), .B2(n11371), .A(n15393), .ZN(n15375) );
  INV_X1 U14530 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21550) );
  NOR2_X1 U14531 ( .A1(n20904), .A2(n21550), .ZN(n15171) );
  INV_X1 U14532 ( .A(n15171), .ZN(n11373) );
  NAND2_X1 U14533 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  AOI21_X1 U14534 ( .B1(n15059), .B2(n20998), .A(n11375), .ZN(n11376) );
  INV_X2 U14535 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16905) );
  AND2_X4 U14536 ( .A1(n16805), .A2(n16905), .ZN(n12640) );
  AOI22_X1 U14537 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11381) );
  INV_X2 U14538 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16792) );
  NOR2_X2 U14539 ( .A1(n16792), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16788) );
  AND2_X4 U14540 ( .A1(n11538), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12644) );
  AOI22_X1 U14541 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11380) );
  NOR2_X2 U14542 ( .A1(n11377), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16789) );
  AND2_X2 U14543 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14544 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9739), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14545 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14546 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14547 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14548 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14549 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14550 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14551 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14552 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14553 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14554 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11395) );
  AOI22_X1 U14555 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14556 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12640), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11392) );
  NAND4_X1 U14557 ( .A1(n11395), .A2(n11394), .A3(n11393), .A4(n11392), .ZN(
        n11396) );
  AOI22_X1 U14558 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14559 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12640), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14560 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11397) );
  NAND4_X1 U14561 ( .A1(n11400), .A2(n11399), .A3(n11398), .A4(n11397), .ZN(
        n11401) );
  NAND2_X1 U14562 ( .A1(n11401), .A2(n11535), .ZN(n11402) );
  AOI22_X1 U14563 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12640), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14564 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14565 ( .A1(n11430), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14566 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U14567 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11408) );
  NAND2_X1 U14568 ( .A1(n11408), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11415) );
  AOI22_X1 U14569 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14570 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14571 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14572 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14573 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11413) );
  NAND2_X1 U14574 ( .A1(n11413), .A2(n11535), .ZN(n11414) );
  AOI22_X1 U14575 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12640), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14576 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14577 ( .A1(n11430), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9728), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14578 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11416) );
  NAND4_X1 U14579 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n11420) );
  AOI22_X1 U14580 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9737), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14581 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14582 ( .A1(n11430), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14583 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14584 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11425) );
  AOI22_X1 U14585 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14586 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14587 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12784), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14588 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14589 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14590 ( .A1(n9730), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14591 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11432) );
  AOI22_X1 U14592 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14593 ( .A1(n9731), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11438) );
  AOI22_X1 U14594 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12784), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11437) );
  AOI22_X1 U14595 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11435) );
  AOI22_X1 U14596 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14597 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14598 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12784), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14599 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14600 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14601 ( .A1(n11529), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9742), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14602 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14603 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12644), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14604 ( .A1(n12640), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11430), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14605 ( .A1(n9736), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9729), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14606 ( .A1(n11530), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11536), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11449) );
  NAND4_X1 U14607 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n11453) );
  INV_X1 U14608 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20692) );
  NAND2_X1 U14609 ( .A1(n11466), .A2(n20118), .ZN(n11459) );
  NAND2_X1 U14610 ( .A1(n11896), .A2(n12035), .ZN(n11895) );
  AND2_X1 U14611 ( .A1(n11888), .A2(n16873), .ZN(n11462) );
  NOR2_X2 U14612 ( .A1(n11463), .A2(n11473), .ZN(n11887) );
  NAND4_X1 U14613 ( .A1(n12251), .A2(n11470), .A3(n12039), .A4(n20807), .ZN(
        n11468) );
  NAND3_X1 U14614 ( .A1(n12041), .A2(n11465), .A3(n11466), .ZN(n11467) );
  NAND3_X1 U14615 ( .A1(n11469), .A2(n11468), .A3(n11467), .ZN(n11477) );
  NAND3_X1 U14616 ( .A1(n11470), .A2(n12035), .A3(n20135), .ZN(n11471) );
  NAND2_X1 U14617 ( .A1(n11472), .A2(n11471), .ZN(n11474) );
  NAND3_X1 U14618 ( .A1(n11474), .A2(n12028), .A3(n11473), .ZN(n11476) );
  NAND2_X1 U14619 ( .A1(n11475), .A2(n9857), .ZN(n13538) );
  NAND3_X1 U14620 ( .A1(n11476), .A2(n11890), .A3(n13538), .ZN(n12044) );
  INV_X1 U14621 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19973) );
  NAND2_X1 U14622 ( .A1(n12366), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n11481) );
  INV_X1 U14623 ( .A(n20801), .ZN(n11501) );
  NAND2_X1 U14624 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11479) );
  AND2_X1 U14625 ( .A1(n11501), .A2(n11479), .ZN(n11480) );
  OAI211_X1 U14626 ( .C1(n11502), .C2(n19973), .A(n11481), .B(n11480), .ZN(
        n11482) );
  INV_X1 U14627 ( .A(n11482), .ZN(n11484) );
  NAND2_X1 U14628 ( .A1(n11492), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11483) );
  AND2_X1 U14629 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11485) );
  OAI22_X1 U14630 ( .A1(n11486), .A2(n9837), .B1(n11485), .B2(n12366), .ZN(
        n11489) );
  NAND2_X1 U14631 ( .A1(n20801), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11487) );
  AOI21_X1 U14632 ( .B1(n20808), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11491) );
  INV_X1 U14633 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20694) );
  NAND2_X1 U14634 ( .A1(n12366), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U14635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11493) );
  OAI211_X1 U14636 ( .C1(n11502), .C2(n20694), .A(n11494), .B(n11493), .ZN(
        n11495) );
  INV_X1 U14637 ( .A(n11495), .ZN(n11496) );
  INV_X1 U14638 ( .A(n11510), .ZN(n11499) );
  INV_X1 U14639 ( .A(n11509), .ZN(n11498) );
  NAND2_X1 U14640 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  OAI22_X1 U14641 ( .A1(n11490), .A2(n11535), .B1(n11501), .B2(n20758), .ZN(
        n11506) );
  BUF_X2 U14642 ( .A(n11502), .Z(n12382) );
  INV_X1 U14643 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U14644 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11504) );
  AOI22_X1 U14645 ( .A1(n12366), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11503) );
  INV_X1 U14646 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11515) );
  AND2_X2 U14647 ( .A1(n13893), .A2(n11523), .ZN(n11603) );
  AOI22_X1 U14648 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n11603), .B1(
        n20401), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14650 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11534) );
  AND2_X4 U14651 ( .A1(n12783), .A2(n11535), .ZN(n12625) );
  AOI22_X1 U14652 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11533) );
  AND2_X2 U14653 ( .A1(n12640), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12583) );
  AOI22_X1 U14654 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11532) );
  INV_X1 U14655 ( .A(n11536), .ZN(n12645) );
  AND2_X2 U14656 ( .A1(n11530), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11630) );
  AOI22_X1 U14657 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11531) );
  NAND4_X1 U14658 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11544) );
  AND2_X2 U14659 ( .A1(n12644), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11596) );
  AND2_X2 U14660 ( .A1(n12644), .A2(n11535), .ZN(n11573) );
  AOI22_X1 U14661 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U14662 ( .A1(n11530), .A2(n11535), .ZN(n11634) );
  INV_X2 U14663 ( .A(n9800), .ZN(n12626) );
  AOI22_X1 U14664 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11541) );
  NOR2_X2 U14665 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12642) );
  AOI22_X1 U14666 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11540) );
  AOI22_X1 U14667 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11539) );
  NAND4_X1 U14668 ( .A1(n11542), .A2(n11541), .A3(n11540), .A4(n11539), .ZN(
        n11543) );
  NAND2_X1 U14669 ( .A1(n11545), .A2(n16029), .ZN(n11546) );
  AOI22_X1 U14670 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20148), .B1(
        n11605), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14671 ( .A1(n16837), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20336), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14672 ( .A1(n20249), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11552) );
  NAND2_X1 U14673 ( .A1(n20174), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11551) );
  INV_X1 U14674 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16892) );
  AOI21_X1 U14675 ( .B1(n20401), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n16029), .ZN(n11554) );
  NAND2_X1 U14676 ( .A1(n20103), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11553) );
  AOI22_X1 U14677 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11558) );
  AOI22_X1 U14678 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n11909), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11557) );
  AOI22_X1 U14679 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14680 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12626), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11555) );
  NAND4_X1 U14681 ( .A1(n11558), .A2(n11557), .A3(n11556), .A4(n11555), .ZN(
        n11566) );
  AOI22_X1 U14682 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11596), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11564) );
  INV_X2 U14683 ( .A(n11634), .ZN(n12588) );
  AOI22_X1 U14684 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12588), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14685 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n11559), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U14686 ( .A1(n11564), .A2(n11563), .A3(n11562), .A4(n11561), .ZN(
        n11565) );
  AOI22_X1 U14687 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14688 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12625), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14689 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14690 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11630), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11569) );
  NAND4_X1 U14691 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11580) );
  AOI22_X1 U14692 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11573), .B1(
        n11596), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14693 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12626), .B1(
        n12588), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14694 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11559), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14695 ( .A1(n11578), .A2(n11577), .A3(n11576), .A4(n11575), .ZN(
        n11579) );
  NAND3_X1 U14696 ( .A1(n16029), .A2(n13563), .A3(n12080), .ZN(n11922) );
  AOI22_X1 U14697 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14698 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14699 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14700 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14701 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AOI22_X1 U14702 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14703 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14704 ( .A1(n11560), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14705 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11559), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14706 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  NAND2_X1 U14707 ( .A1(n11922), .A2(n12087), .ZN(n11591) );
  AOI22_X1 U14708 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14709 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14710 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14711 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14712 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11602) );
  AOI22_X1 U14713 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14714 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14715 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14716 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11597) );
  NAND4_X1 U14717 ( .A1(n11600), .A2(n11599), .A3(n11598), .A4(n11597), .ZN(
        n11601) );
  INV_X1 U14718 ( .A(n11918), .ZN(n12098) );
  AOI22_X1 U14719 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20212), .B1(
        n20401), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14720 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20148), .B1(
        n20524), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14721 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20336), .B1(
        n11605), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11606) );
  INV_X1 U14722 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11610) );
  INV_X1 U14723 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14089) );
  AOI22_X1 U14724 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n16884), .B1(
        n16862), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14725 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14726 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14727 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14728 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11615) );
  NAND4_X1 U14729 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11624) );
  AOI22_X1 U14730 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14731 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14732 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14733 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11619) );
  NAND4_X1 U14734 ( .A1(n11622), .A2(n11621), .A3(n11620), .A4(n11619), .ZN(
        n11623) );
  NAND2_X1 U14735 ( .A1(n12105), .A2(n16029), .ZN(n11625) );
  AOI22_X1 U14736 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14737 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14738 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11627) );
  NAND2_X1 U14739 ( .A1(n11573), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11626) );
  INV_X1 U14740 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11633) );
  INV_X1 U14741 ( .A(n11630), .ZN(n11632) );
  INV_X1 U14742 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11631) );
  OAI22_X1 U14743 ( .A1(n11634), .A2(n11633), .B1(n11632), .B2(n11631), .ZN(
        n11635) );
  NAND2_X1 U14744 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11636) );
  INV_X1 U14745 ( .A(n12625), .ZN(n11640) );
  INV_X1 U14746 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11639) );
  INV_X1 U14747 ( .A(n11637), .ZN(n11638) );
  INV_X1 U14748 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12778) );
  OAI22_X1 U14749 ( .A1(n11640), .A2(n11639), .B1(n11638), .B2(n12778), .ZN(
        n11646) );
  INV_X1 U14750 ( .A(n11641), .ZN(n11644) );
  INV_X1 U14751 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11643) );
  INV_X1 U14752 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11642) );
  OAI22_X1 U14753 ( .A1(n11644), .A2(n11643), .B1(n9800), .B2(n11642), .ZN(
        n11645) );
  NOR2_X1 U14754 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  INV_X4 U14755 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20776) );
  NAND2_X1 U14756 ( .A1(n20776), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11650) );
  NAND2_X1 U14757 ( .A1(n16792), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11648) );
  AND2_X1 U14758 ( .A1(n11650), .A2(n11648), .ZN(n11857) );
  NAND2_X1 U14759 ( .A1(n11649), .A2(n11857), .ZN(n11859) );
  NAND2_X1 U14760 ( .A1(n11859), .A2(n11650), .ZN(n11659) );
  NAND2_X1 U14761 ( .A1(n11651), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11652) );
  NAND2_X1 U14762 ( .A1(n11660), .A2(n11652), .ZN(n11657) );
  XNOR2_X1 U14763 ( .A(n11659), .B(n11657), .ZN(n11899) );
  NAND2_X1 U14764 ( .A1(n11653), .A2(n12386), .ZN(n11654) );
  INV_X1 U14765 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n15955) );
  NOR2_X1 U14766 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n11656) );
  MUX2_X1 U14767 ( .A(n11656), .B(n12080), .S(n20127), .Z(n11684) );
  NAND2_X1 U14768 ( .A1(n11682), .A2(n11684), .ZN(n11679) );
  INV_X1 U14769 ( .A(n11657), .ZN(n11658) );
  NAND2_X1 U14770 ( .A1(n11659), .A2(n11658), .ZN(n11661) );
  INV_X1 U14771 ( .A(n11664), .ZN(n11662) );
  XNOR2_X1 U14772 ( .A(n11665), .B(n11662), .ZN(n11855) );
  INV_X1 U14773 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n15944) );
  MUX2_X1 U14774 ( .A(n11883), .B(n15944), .S(n12290), .Z(n11678) );
  NAND2_X1 U14775 ( .A1(n11665), .A2(n11664), .ZN(n11667) );
  NAND2_X1 U14776 ( .A1(n20758), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11666) );
  INV_X1 U14777 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n11668) );
  INV_X1 U14778 ( .A(n11885), .ZN(n11669) );
  INV_X1 U14779 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13962) );
  INV_X1 U14780 ( .A(n12105), .ZN(n11670) );
  MUX2_X1 U14781 ( .A(n13962), .B(n11670), .S(n20127), .Z(n11671) );
  NAND2_X1 U14782 ( .A1(n9882), .A2(n10117), .ZN(n11672) );
  NAND2_X1 U14783 ( .A1(n11694), .A2(n11672), .ZN(n15929) );
  NAND2_X1 U14784 ( .A1(n11673), .A2(n15929), .ZN(n11693) );
  INV_X1 U14785 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16752) );
  XNOR2_X1 U14786 ( .A(n11693), .B(n16752), .ZN(n16740) );
  INV_X1 U14787 ( .A(n11674), .ZN(n11677) );
  INV_X1 U14788 ( .A(n11675), .ZN(n11676) );
  XNOR2_X1 U14789 ( .A(n11677), .B(n11676), .ZN(n19982) );
  INV_X1 U14790 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16767) );
  INV_X1 U14791 ( .A(n11678), .ZN(n11680) );
  NAND2_X1 U14792 ( .A1(n11680), .A2(n11679), .ZN(n11681) );
  NAND2_X1 U14793 ( .A1(n11675), .A2(n11681), .ZN(n15943) );
  XNOR2_X1 U14794 ( .A(n11682), .B(n11684), .ZN(n15959) );
  XNOR2_X1 U14795 ( .A(n15959), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14656) );
  OAI21_X1 U14796 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20786), .A(
        n11858), .ZN(n11908) );
  INV_X1 U14797 ( .A(n11908), .ZN(n11861) );
  MUX2_X1 U14798 ( .A(n13563), .B(n11861), .S(n11683), .Z(n11879) );
  MUX2_X1 U14799 ( .A(P2_EBX_REG_0__SCAN_IN), .B(n11879), .S(n20127), .Z(
        n15983) );
  NAND2_X1 U14800 ( .A1(n15983), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13573) );
  INV_X1 U14801 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13580) );
  AND2_X1 U14802 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U14803 ( .A1(n15983), .A2(n13579), .ZN(n11687) );
  INV_X1 U14804 ( .A(n11684), .ZN(n11686) );
  NAND3_X1 U14805 ( .A1(n12290), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n11685) );
  NAND2_X1 U14806 ( .A1(n11686), .A2(n11685), .ZN(n15971) );
  AOI22_X1 U14807 ( .A1(n13573), .A2(n13580), .B1(n11687), .B2(n15971), .ZN(
        n14657) );
  NAND2_X1 U14808 ( .A1(n14656), .A2(n14657), .ZN(n14677) );
  INV_X1 U14809 ( .A(n15959), .ZN(n11688) );
  NAND2_X1 U14810 ( .A1(n11688), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11689) );
  NAND2_X1 U14811 ( .A1(n14677), .A2(n11689), .ZN(n16456) );
  NAND2_X1 U14812 ( .A1(n19982), .A2(n16767), .ZN(n11691) );
  OAI21_X1 U14813 ( .B1(n16456), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n11691), .ZN(n11690) );
  NAND3_X1 U14814 ( .A1(n11691), .A2(n16456), .A3(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n11692) );
  AOI21_X2 U14815 ( .B1(n16740), .B2(n16741), .A(n10724), .ZN(n16387) );
  INV_X1 U14816 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n11706) );
  AOI22_X1 U14817 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14818 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11697) );
  AOI22_X1 U14819 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11696) );
  AOI22_X1 U14820 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11695) );
  NAND4_X1 U14821 ( .A1(n11698), .A2(n11697), .A3(n11696), .A4(n11695), .ZN(
        n11704) );
  AOI22_X1 U14822 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11702) );
  AOI22_X1 U14823 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14824 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14825 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11699) );
  NAND4_X1 U14826 ( .A1(n11702), .A2(n11701), .A3(n11700), .A4(n11699), .ZN(
        n11703) );
  INV_X1 U14827 ( .A(n12109), .ZN(n11705) );
  MUX2_X1 U14828 ( .A(n11706), .B(n11705), .S(n20127), .Z(n11732) );
  INV_X1 U14829 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n11708) );
  MUX2_X1 U14830 ( .A(n11708), .B(n11707), .S(n20127), .Z(n11713) );
  NAND2_X1 U14831 ( .A1(n12290), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n11709) );
  INV_X1 U14832 ( .A(n11709), .ZN(n11710) );
  NAND2_X1 U14833 ( .A1(n9849), .A2(n11710), .ZN(n11711) );
  NAND2_X1 U14834 ( .A1(n11746), .A2(n11711), .ZN(n15895) );
  NOR2_X1 U14835 ( .A1(n15895), .A2(n14606), .ZN(n11740) );
  NAND2_X1 U14836 ( .A1(n11740), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16421) );
  XNOR2_X1 U14837 ( .A(n11712), .B(n11713), .ZN(n15905) );
  NAND2_X1 U14838 ( .A1(n15905), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16432) );
  AND2_X1 U14839 ( .A1(n16421), .A2(n16432), .ZN(n16391) );
  AOI22_X1 U14840 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20524), .B1(
        n20401), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14841 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20336), .B1(
        n11605), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14842 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20212), .B1(
        n20148), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11715) );
  INV_X1 U14843 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11721) );
  INV_X1 U14844 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11718) );
  OAI22_X1 U14845 ( .A1(n11721), .A2(n11720), .B1(n11719), .B2(n11718), .ZN(
        n11724) );
  INV_X1 U14846 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11722) );
  NOR2_X1 U14847 ( .A1(n11724), .A2(n11723), .ZN(n11727) );
  AOI22_X1 U14848 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n16884), .B1(
        n9801), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11725) );
  NAND4_X1 U14849 ( .A1(n11728), .A2(n11727), .A3(n11726), .A4(n11725), .ZN(
        n11730) );
  NAND2_X1 U14850 ( .A1(n12109), .A2(n16029), .ZN(n11729) );
  NAND2_X1 U14851 ( .A1(n11694), .A2(n10652), .ZN(n11733) );
  NAND2_X1 U14852 ( .A1(n11712), .A2(n11733), .ZN(n15918) );
  INV_X1 U14853 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11734) );
  INV_X1 U14854 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11735) );
  NOR2_X4 U14855 ( .A1(n11746), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11748) );
  INV_X1 U14856 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n14040) );
  NAND3_X1 U14857 ( .A1(n11737), .A2(n12290), .A3(P2_EBX_REG_11__SCAN_IN), 
        .ZN(n11738) );
  NAND2_X1 U14858 ( .A1(n11739), .A2(n11738), .ZN(n15859) );
  INV_X1 U14859 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16660) );
  OAI21_X1 U14860 ( .B1(n15859), .B2(n14606), .A(n16660), .ZN(n16386) );
  INV_X1 U14861 ( .A(n11740), .ZN(n11741) );
  INV_X1 U14862 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16701) );
  NAND2_X1 U14863 ( .A1(n11741), .A2(n16701), .ZN(n16420) );
  INV_X1 U14864 ( .A(n15905), .ZN(n11742) );
  INV_X1 U14865 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16722) );
  NAND2_X1 U14866 ( .A1(n11742), .A2(n16722), .ZN(n16431) );
  AND2_X1 U14867 ( .A1(n16420), .A2(n16431), .ZN(n16390) );
  NAND2_X1 U14868 ( .A1(n12290), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11743) );
  MUX2_X1 U14869 ( .A(n11743), .B(P2_EBX_REG_10__SCAN_IN), .S(n11748), .Z(
        n11744) );
  AND2_X1 U14870 ( .A1(n11744), .A2(n11843), .ZN(n15867) );
  NAND2_X1 U14871 ( .A1(n15867), .A2(n10382), .ZN(n11745) );
  INV_X1 U14872 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16674) );
  NAND2_X1 U14873 ( .A1(n11745), .A2(n16674), .ZN(n16400) );
  NAND2_X1 U14874 ( .A1(n12290), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11747) );
  MUX2_X1 U14875 ( .A(n12290), .B(n11747), .S(n11746), .Z(n11750) );
  INV_X1 U14876 ( .A(n11748), .ZN(n11749) );
  NAND2_X1 U14877 ( .A1(n15877), .A2(n10382), .ZN(n11751) );
  NAND2_X1 U14878 ( .A1(n11751), .A2(n10209), .ZN(n16409) );
  INV_X1 U14879 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n21785) );
  NOR2_X1 U14880 ( .A1(n20127), .A2(n21785), .ZN(n11783) );
  INV_X1 U14881 ( .A(n11783), .ZN(n11754) );
  INV_X1 U14882 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n11756) );
  NOR2_X1 U14883 ( .A1(n20127), .A2(n11756), .ZN(n11791) );
  NOR2_X1 U14884 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n11758) );
  NOR2_X1 U14885 ( .A1(n20127), .A2(n11758), .ZN(n11759) );
  NAND2_X1 U14886 ( .A1(n12290), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n11760) );
  INV_X1 U14887 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11761) );
  NOR2_X1 U14888 ( .A1(n20127), .A2(n11761), .ZN(n11777) );
  INV_X1 U14889 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n11762) );
  NAND2_X1 U14890 ( .A1(n12290), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n11768) );
  INV_X1 U14891 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n11763) );
  MUX2_X1 U14892 ( .A(n11764), .B(n10120), .S(n20127), .Z(n11766) );
  NAND2_X1 U14893 ( .A1(n11766), .A2(n11770), .ZN(n15736) );
  INV_X1 U14894 ( .A(n11819), .ZN(n11767) );
  INV_X1 U14895 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12434) );
  NAND2_X1 U14896 ( .A1(n11767), .A2(n12434), .ZN(n16292) );
  XNOR2_X1 U14897 ( .A(n9817), .B(n11768), .ZN(n15758) );
  NAND2_X1 U14898 ( .A1(n15758), .A2(n10382), .ZN(n11805) );
  INV_X1 U14899 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16305) );
  NAND2_X1 U14900 ( .A1(n11805), .A2(n16305), .ZN(n16301) );
  XNOR2_X1 U14901 ( .A(n11780), .B(n9869), .ZN(n15773) );
  NAND2_X1 U14902 ( .A1(n15773), .A2(n10382), .ZN(n11769) );
  INV_X1 U14903 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U14904 ( .A1(n11769), .A2(n11941), .ZN(n16313) );
  AND2_X1 U14905 ( .A1(n16301), .A2(n16313), .ZN(n16290) );
  AND3_X1 U14906 ( .A1(n11770), .A2(n12290), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n11771) );
  NOR2_X1 U14907 ( .A1(n11823), .A2(n11771), .ZN(n15722) );
  NAND2_X1 U14908 ( .A1(n15722), .A2(n10382), .ZN(n11804) );
  INV_X1 U14909 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n21805) );
  NAND2_X1 U14910 ( .A1(n11804), .A2(n21805), .ZN(n12428) );
  INV_X1 U14911 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11772) );
  NAND2_X1 U14912 ( .A1(n11773), .A2(n11772), .ZN(n11775) );
  INV_X1 U14913 ( .A(n11773), .ZN(n11788) );
  NAND3_X1 U14914 ( .A1(n11788), .A2(n12290), .A3(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n11774) );
  NAND3_X1 U14915 ( .A1(n11775), .A2(n11774), .A3(n11843), .ZN(n15801) );
  NOR2_X1 U14916 ( .A1(n15801), .A2(n14606), .ZN(n11807) );
  INV_X1 U14917 ( .A(n11807), .ZN(n11776) );
  XNOR2_X1 U14918 ( .A(n11776), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12420) );
  NAND2_X1 U14919 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  AND2_X1 U14920 ( .A1(n11780), .A2(n11779), .ZN(n15794) );
  NAND2_X1 U14921 ( .A1(n15794), .A2(n10382), .ZN(n11781) );
  INV_X1 U14922 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16323) );
  NAND2_X1 U14923 ( .A1(n11781), .A2(n16323), .ZN(n12424) );
  NAND2_X1 U14924 ( .A1(n11784), .A2(n11783), .ZN(n11785) );
  NAND2_X1 U14925 ( .A1(n11782), .A2(n11785), .ZN(n15840) );
  OR2_X1 U14926 ( .A1(n15840), .A2(n14606), .ZN(n16374) );
  INV_X1 U14927 ( .A(n16374), .ZN(n11795) );
  INV_X1 U14928 ( .A(n11793), .ZN(n11797) );
  INV_X1 U14929 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n16091) );
  NAND2_X1 U14930 ( .A1(n11797), .A2(n16091), .ZN(n11799) );
  INV_X1 U14931 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11786) );
  NOR2_X1 U14932 ( .A1(n20127), .A2(n11786), .ZN(n11787) );
  NAND2_X1 U14933 ( .A1(n11799), .A2(n11787), .ZN(n11789) );
  NAND2_X1 U14934 ( .A1(n11789), .A2(n11788), .ZN(n15821) );
  OR2_X1 U14935 ( .A1(n15821), .A2(n14606), .ZN(n11790) );
  INV_X1 U14936 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16614) );
  NAND2_X1 U14937 ( .A1(n11790), .A2(n16614), .ZN(n16341) );
  NAND2_X1 U14938 ( .A1(n11782), .A2(n11791), .ZN(n11792) );
  NAND2_X1 U14939 ( .A1(n11793), .A2(n11792), .ZN(n13390) );
  NOR2_X1 U14940 ( .A1(n13390), .A2(n14606), .ZN(n11813) );
  INV_X1 U14941 ( .A(n11813), .ZN(n11794) );
  INV_X1 U14942 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U14943 ( .A1(n11794), .A2(n16638), .ZN(n16365) );
  OAI211_X1 U14944 ( .C1(n11795), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16341), .B(n16365), .ZN(n11796) );
  INV_X1 U14945 ( .A(n11796), .ZN(n11802) );
  NAND2_X1 U14946 ( .A1(n12290), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11798) );
  MUX2_X1 U14947 ( .A(n11798), .B(n12290), .S(n11797), .Z(n11800) );
  NAND2_X1 U14948 ( .A1(n15831), .A2(n10382), .ZN(n11801) );
  INV_X1 U14949 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16356) );
  NAND2_X1 U14950 ( .A1(n11801), .A2(n16356), .ZN(n16352) );
  AND4_X1 U14951 ( .A1(n12420), .A2(n12424), .A3(n11802), .A4(n16352), .ZN(
        n11803) );
  NAND3_X1 U14952 ( .A1(n12427), .A2(n12428), .A3(n11803), .ZN(n11822) );
  OR2_X1 U14953 ( .A1(n11804), .A2(n21805), .ZN(n12429) );
  OR2_X1 U14954 ( .A1(n11805), .A2(n16305), .ZN(n16302) );
  AND2_X1 U14955 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14956 ( .A1(n15773), .A2(n11806), .ZN(n16312) );
  AND2_X1 U14957 ( .A1(n16302), .A2(n16312), .ZN(n12425) );
  NAND2_X1 U14958 ( .A1(n11807), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12422) );
  NOR2_X1 U14959 ( .A1(n16374), .A2(n12416), .ZN(n11812) );
  AND2_X1 U14960 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U14961 ( .A1(n15867), .A2(n11808), .ZN(n16399) );
  AND2_X1 U14962 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14963 ( .A1(n15877), .A2(n11809), .ZN(n16408) );
  AND2_X1 U14964 ( .A1(n16399), .A2(n16408), .ZN(n16392) );
  INV_X1 U14965 ( .A(n15859), .ZN(n11811) );
  AND2_X1 U14966 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14967 ( .A1(n11811), .A2(n11810), .ZN(n16385) );
  NAND2_X1 U14968 ( .A1(n16392), .A2(n16385), .ZN(n12413) );
  NOR2_X1 U14969 ( .A1(n11812), .A2(n12413), .ZN(n11815) );
  NAND2_X1 U14970 ( .A1(n11813), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16366) );
  AND2_X1 U14971 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U14972 ( .A1(n15794), .A2(n11814), .ZN(n12423) );
  NAND4_X1 U14973 ( .A1(n12422), .A2(n11815), .A3(n16366), .A4(n12423), .ZN(
        n11818) );
  AND2_X1 U14974 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14975 ( .A1(n15831), .A2(n11816), .ZN(n16351) );
  NAND2_X1 U14976 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11817) );
  OR2_X1 U14977 ( .A1(n15821), .A2(n11817), .ZN(n16340) );
  NAND2_X1 U14978 ( .A1(n16351), .A2(n16340), .ZN(n12417) );
  NOR2_X1 U14979 ( .A1(n11818), .A2(n12417), .ZN(n11820) );
  NAND2_X1 U14980 ( .A1(n11819), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16293) );
  AND4_X1 U14981 ( .A1(n12429), .A2(n12425), .A3(n11820), .A4(n16293), .ZN(
        n11821) );
  NAND2_X1 U14982 ( .A1(n11824), .A2(n9872), .ZN(n11825) );
  NAND2_X1 U14983 ( .A1(n11831), .A2(n11825), .ZN(n15715) );
  OR2_X1 U14984 ( .A1(n15715), .A2(n14606), .ZN(n11826) );
  INV_X1 U14985 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16556) );
  NAND2_X1 U14986 ( .A1(n11826), .A2(n16556), .ZN(n16280) );
  INV_X1 U14987 ( .A(n11826), .ZN(n11827) );
  NAND2_X1 U14988 ( .A1(n11827), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16281) );
  NAND2_X1 U14989 ( .A1(n12290), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n11829) );
  XNOR2_X1 U14990 ( .A(n11831), .B(n11829), .ZN(n15704) );
  NAND2_X1 U14991 ( .A1(n15704), .A2(n10382), .ZN(n11828) );
  XNOR2_X1 U14992 ( .A(n11828), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16273) );
  INV_X1 U14993 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16539) );
  INV_X1 U14994 ( .A(n11829), .ZN(n11830) );
  INV_X1 U14995 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n16035) );
  NAND2_X1 U14996 ( .A1(n11832), .A2(n16035), .ZN(n11841) );
  INV_X1 U14997 ( .A(n11832), .ZN(n11834) );
  NOR2_X1 U14998 ( .A1(n20127), .A2(n16035), .ZN(n11833) );
  AOI21_X1 U14999 ( .B1(n11834), .B2(n11833), .A(n10647), .ZN(n11835) );
  NAND2_X1 U15000 ( .A1(n11841), .A2(n11835), .ZN(n15679) );
  INV_X1 U15001 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16525) );
  NOR2_X1 U15002 ( .A1(n11836), .A2(n16525), .ZN(n16261) );
  NAND2_X1 U15003 ( .A1(n11836), .A2(n16525), .ZN(n16260) );
  NAND2_X1 U15004 ( .A1(n12290), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11837) );
  MUX2_X1 U15005 ( .A(P2_EBX_REG_25__SCAN_IN), .B(n11837), .S(n11841), .Z(
        n11838) );
  AOI21_X1 U15006 ( .B1(n15670), .B2(n10382), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16254) );
  NAND2_X1 U15007 ( .A1(n15650), .A2(n11842), .ZN(n11848) );
  INV_X1 U15008 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16500) );
  XNOR2_X1 U15009 ( .A(n11850), .B(n16500), .ZN(n16238) );
  NAND2_X1 U15010 ( .A1(n12290), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n11846) );
  INV_X1 U15011 ( .A(n11846), .ZN(n11847) );
  NAND2_X1 U15012 ( .A1(n11848), .A2(n11847), .ZN(n11849) );
  NAND2_X1 U15013 ( .A1(n9806), .A2(n11849), .ZN(n15640) );
  INV_X1 U15014 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U15015 ( .A1(n11851), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11853) );
  INV_X1 U15016 ( .A(n15670), .ZN(n11852) );
  INV_X1 U15017 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16514) );
  INV_X1 U15018 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14630) );
  INV_X1 U15019 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n20684) );
  NAND2_X1 U15020 ( .A1(n21751), .A2(n20684), .ZN(n19961) );
  OAI211_X1 U15021 ( .C1(n21751), .C2(n20684), .A(n20675), .B(n19961), .ZN(
        n20806) );
  NAND2_X1 U15022 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20812) );
  INV_X1 U15023 ( .A(n20812), .ZN(n20686) );
  NOR2_X1 U15024 ( .A1(n20806), .A2(n20686), .ZN(n13527) );
  NAND2_X1 U15025 ( .A1(n20113), .A2(n13527), .ZN(n11877) );
  AND2_X1 U15026 ( .A1(n11856), .A2(n11855), .ZN(n11898) );
  NAND2_X1 U15027 ( .A1(n20807), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20033) );
  AOI21_X1 U15028 ( .B1(n20033), .B2(n16887), .A(n11899), .ZN(n11867) );
  NAND2_X1 U15029 ( .A1(n11465), .A2(n11899), .ZN(n11865) );
  INV_X1 U15030 ( .A(n11857), .ZN(n11862) );
  NAND2_X1 U15031 ( .A1(n11858), .A2(n11862), .ZN(n11878) );
  NAND2_X1 U15032 ( .A1(n11859), .A2(n11878), .ZN(n11900) );
  INV_X1 U15033 ( .A(n11900), .ZN(n11860) );
  OAI211_X1 U15034 ( .C1(n16887), .C2(n11861), .A(n11890), .B(n11860), .ZN(
        n11864) );
  OAI21_X1 U15035 ( .B1(n11908), .B2(n11862), .A(n12386), .ZN(n11863) );
  NAND3_X1 U15036 ( .A1(n11865), .A2(n11864), .A3(n11863), .ZN(n11866) );
  OAI211_X1 U15037 ( .C1(n11868), .C2(n11867), .A(n11866), .B(n11898), .ZN(
        n11872) );
  NAND2_X1 U15038 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16924), .ZN(
        n11870) );
  NOR2_X1 U15039 ( .A1(n16924), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n11869) );
  AOI21_X1 U15040 ( .B1(n11875), .B2(n11890), .A(n12035), .ZN(n11873) );
  INV_X1 U15041 ( .A(n11873), .ZN(n11876) );
  MUX2_X1 U15042 ( .A(n11877), .B(n11876), .S(n20030), .Z(n11916) );
  NAND2_X1 U15043 ( .A1(n11879), .A2(n11878), .ZN(n11882) );
  INV_X1 U15044 ( .A(n11880), .ZN(n11881) );
  NAND2_X1 U15045 ( .A1(n11882), .A2(n11881), .ZN(n11884) );
  NAND3_X1 U15046 ( .A1(n11885), .A2(n11884), .A3(n11883), .ZN(n11886) );
  AND2_X1 U15047 ( .A1(n11886), .A2(n11902), .ZN(n20793) );
  AND2_X1 U15048 ( .A1(n16029), .A2(n20807), .ZN(n12289) );
  AND2_X1 U15049 ( .A1(n11887), .A2(n12289), .ZN(n20789) );
  NAND2_X1 U15050 ( .A1(n20793), .A2(n20789), .ZN(n12263) );
  NAND2_X1 U15051 ( .A1(n11888), .A2(n12028), .ZN(n11889) );
  NAND2_X1 U15052 ( .A1(n13529), .A2(n11889), .ZN(n11905) );
  OAI21_X1 U15053 ( .B1(n12035), .B2(n16887), .A(n11890), .ZN(n11891) );
  NAND2_X1 U15054 ( .A1(n11891), .A2(n16873), .ZN(n11893) );
  AOI21_X1 U15055 ( .B1(n11893), .B2(n12028), .A(n11892), .ZN(n11894) );
  AND2_X1 U15056 ( .A1(n11895), .A2(n11894), .ZN(n11904) );
  OAI21_X1 U15057 ( .B1(n11896), .B2(n12069), .A(n12289), .ZN(n12033) );
  NAND2_X1 U15058 ( .A1(n11899), .A2(n11898), .ZN(n11907) );
  NAND3_X1 U15059 ( .A1(n11897), .A2(n13527), .A3(n16897), .ZN(n11903) );
  MUX2_X1 U15060 ( .A(n11897), .B(n20113), .S(n16029), .Z(n11906) );
  NAND3_X1 U15061 ( .A1(n11906), .A2(n20812), .A3(n16897), .ZN(n11914) );
  OAI21_X1 U15062 ( .B1(n11908), .B2(n11907), .A(n16897), .ZN(n11912) );
  INV_X1 U15063 ( .A(n11909), .ZN(n11911) );
  AOI21_X1 U15064 ( .B1(n16821), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13539) );
  AOI21_X1 U15065 ( .B1(n11911), .B2(n13539), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n20779) );
  MUX2_X1 U15066 ( .A(n11912), .B(n20779), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n17509) );
  INV_X1 U15067 ( .A(n17509), .ZN(n20790) );
  NAND3_X1 U15068 ( .A1(n11887), .A2(n16887), .A3(n20790), .ZN(n11913) );
  INV_X1 U15069 ( .A(n20026), .ZN(n13423) );
  NAND2_X1 U15070 ( .A1(n11887), .A2(n12386), .ZN(n20791) );
  INV_X1 U15071 ( .A(n20791), .ZN(n11917) );
  INV_X1 U15072 ( .A(n13563), .ZN(n12076) );
  NAND3_X1 U15073 ( .A1(n12076), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n12080), .ZN(n11921) );
  NOR2_X1 U15074 ( .A1(n13563), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11919) );
  XNOR2_X1 U15075 ( .A(n11919), .B(n12080), .ZN(n13568) );
  NAND2_X1 U15076 ( .A1(n13568), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U15077 ( .A1(n11921), .A2(n11920), .ZN(n11923) );
  XOR2_X1 U15078 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11923), .Z(
        n14655) );
  XNOR2_X1 U15079 ( .A(n11922), .B(n12087), .ZN(n14653) );
  NAND2_X1 U15080 ( .A1(n14655), .A2(n14653), .ZN(n11925) );
  NAND2_X1 U15081 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11923), .ZN(
        n11924) );
  NAND2_X1 U15082 ( .A1(n11925), .A2(n11924), .ZN(n11926) );
  XNOR2_X1 U15083 ( .A(n11926), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14315) );
  NAND2_X1 U15084 ( .A1(n11926), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11927) );
  INV_X1 U15085 ( .A(n16418), .ZN(n11936) );
  NAND2_X1 U15086 ( .A1(n11936), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11937) );
  AND2_X2 U15087 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  AND2_X1 U15088 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12452) );
  NAND2_X1 U15089 ( .A1(n12452), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16656) );
  AND2_X1 U15090 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U15091 ( .A1(n12460), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11940) );
  NOR2_X1 U15092 ( .A1(n16656), .A2(n11940), .ZN(n12454) );
  AND2_X1 U15093 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12462) );
  NAND2_X1 U15094 ( .A1(n12462), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16592) );
  NOR2_X1 U15095 ( .A1(n16592), .A2(n11941), .ZN(n11942) );
  AND2_X1 U15096 ( .A1(n12454), .A2(n11942), .ZN(n16567) );
  AND2_X1 U15097 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12062) );
  OAI21_X1 U15098 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16240), .A(
        n10151), .ZN(n12275) );
  INV_X1 U15099 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n16465) );
  NAND2_X1 U15100 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11945) );
  AOI22_X1 U15101 ( .A1(n12378), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11944) );
  OAI211_X1 U15102 ( .C1(n12382), .C2(n16465), .A(n11945), .B(n11944), .ZN(
        n13943) );
  NAND2_X1 U15103 ( .A1(n13944), .A2(n13943), .ZN(n13942) );
  INV_X1 U15104 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15925) );
  NAND2_X1 U15105 ( .A1(n12378), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n11947) );
  NAND2_X1 U15106 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11946) );
  OAI211_X1 U15107 ( .C1(n12382), .C2(n15925), .A(n11947), .B(n11946), .ZN(
        n11948) );
  AOI21_X1 U15108 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n12377), .A(
        n11948), .ZN(n13960) );
  INV_X1 U15109 ( .A(n13960), .ZN(n11949) );
  INV_X1 U15110 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20698) );
  NAND2_X1 U15111 ( .A1(n12378), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U15112 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11950) );
  OAI211_X1 U15113 ( .C1(n12382), .C2(n20698), .A(n11951), .B(n11950), .ZN(
        n11952) );
  AOI21_X1 U15114 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n12377), .A(
        n11952), .ZN(n14094) );
  INV_X1 U15115 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20700) );
  NAND2_X1 U15116 ( .A1(n12378), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n11955) );
  NAND2_X1 U15117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11954) );
  OAI211_X1 U15118 ( .C1(n12382), .C2(n20700), .A(n11955), .B(n11954), .ZN(
        n11956) );
  AOI21_X1 U15119 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n12377), .A(
        n11956), .ZN(n14067) );
  INV_X1 U15120 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20702) );
  NAND2_X1 U15121 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11958) );
  AOI22_X1 U15122 ( .A1(n12378), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11957) );
  OAI211_X1 U15123 ( .C1(n12382), .C2(n20702), .A(n11958), .B(n11957), .ZN(
        n14339) );
  INV_X1 U15124 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n15879) );
  NAND2_X1 U15125 ( .A1(n12378), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n11960) );
  NAND2_X1 U15126 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11959) );
  OAI211_X1 U15127 ( .C1(n12382), .C2(n15879), .A(n11960), .B(n11959), .ZN(
        n11961) );
  AOI21_X1 U15128 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n12377), .A(
        n11961), .ZN(n14220) );
  INV_X1 U15129 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20705) );
  NAND2_X1 U15130 ( .A1(n12378), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11963) );
  NAND2_X1 U15131 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11962) );
  OAI211_X1 U15132 ( .C1(n12382), .C2(n20705), .A(n11963), .B(n11962), .ZN(
        n11964) );
  AOI21_X1 U15133 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n12377), .A(
        n11964), .ZN(n14036) );
  INV_X1 U15134 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n21738) );
  NAND2_X1 U15135 ( .A1(n12378), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n11967) );
  NAND2_X1 U15136 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11966) );
  OAI211_X1 U15137 ( .C1(n12382), .C2(n21738), .A(n11967), .B(n11966), .ZN(
        n11968) );
  AOI21_X1 U15138 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n12377), .A(
        n11968), .ZN(n14148) );
  INV_X1 U15139 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20708) );
  NAND2_X1 U15140 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11970) );
  AOI22_X1 U15141 ( .A1(n12378), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n11969) );
  OAI211_X1 U15142 ( .C1(n12382), .C2(n20708), .A(n11970), .B(n11969), .ZN(
        n14141) );
  INV_X1 U15143 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U15144 ( .A1(n12378), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11972) );
  NAND2_X1 U15145 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11971) );
  OAI211_X1 U15146 ( .C1(n12382), .C2(n11973), .A(n11972), .B(n11971), .ZN(
        n11974) );
  AOI21_X1 U15147 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n12377), .A(
        n11974), .ZN(n13397) );
  NAND2_X1 U15148 ( .A1(n11976), .A2(n11975), .ZN(n13395) );
  INV_X1 U15149 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n15833) );
  NAND2_X1 U15150 ( .A1(n12378), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11978) );
  NAND2_X1 U15151 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11977) );
  OAI211_X1 U15152 ( .C1(n12382), .C2(n15833), .A(n11978), .B(n11977), .ZN(
        n11979) );
  AOI21_X1 U15153 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n12377), .A(
        n11979), .ZN(n15829) );
  INV_X1 U15154 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20712) );
  NAND2_X1 U15155 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11981) );
  AOI22_X1 U15156 ( .A1(n12378), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n11980) );
  OAI211_X1 U15157 ( .C1(n12382), .C2(n20712), .A(n11981), .B(n11980), .ZN(
        n15816) );
  INV_X1 U15158 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15798) );
  NAND2_X1 U15159 ( .A1(n11982), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11984) );
  AOI22_X1 U15160 ( .A1(n12378), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n11983) );
  OAI211_X1 U15161 ( .C1(n12382), .C2(n15798), .A(n11984), .B(n11983), .ZN(
        n14699) );
  INV_X1 U15162 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U15163 ( .A1(n12378), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11986) );
  NAND2_X1 U15164 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11985) );
  OAI211_X1 U15165 ( .C1(n12382), .C2(n12228), .A(n11986), .B(n11985), .ZN(
        n11987) );
  AOI21_X1 U15166 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n12377), .A(
        n11987), .ZN(n15770) );
  INV_X1 U15167 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20715) );
  NAND2_X1 U15168 ( .A1(n12378), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U15169 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11988) );
  OAI211_X1 U15170 ( .C1(n12382), .C2(n20715), .A(n11989), .B(n11988), .ZN(
        n11990) );
  AOI21_X1 U15171 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n12377), .A(
        n11990), .ZN(n12465) );
  INV_X1 U15172 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U15173 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11993) );
  AOI22_X1 U15174 ( .A1(n12378), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n11992) );
  OAI211_X1 U15175 ( .C1(n12382), .C2(n20718), .A(n11993), .B(n11992), .ZN(
        n15753) );
  INV_X1 U15176 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11996) );
  NAND2_X1 U15177 ( .A1(n12378), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n11995) );
  NAND2_X1 U15178 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11994) );
  OAI211_X1 U15179 ( .C1(n12376), .C2(n11996), .A(n11995), .B(n11994), .ZN(
        n11997) );
  AOI21_X1 U15180 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n12377), .A(
        n11997), .ZN(n15734) );
  INV_X1 U15181 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n21847) );
  NAND2_X1 U15182 ( .A1(n12378), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U15183 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n11998) );
  OAI211_X1 U15184 ( .C1(n12376), .C2(n21847), .A(n11999), .B(n11998), .ZN(
        n12000) );
  AOI21_X1 U15185 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n12377), .A(
        n12000), .ZN(n12441) );
  INV_X1 U15186 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12238) );
  NAND2_X1 U15187 ( .A1(n12378), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12003) );
  NAND2_X1 U15188 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12002) );
  OAI211_X1 U15189 ( .C1(n12376), .C2(n12238), .A(n12003), .B(n12002), .ZN(
        n12004) );
  AOI21_X1 U15190 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n12377), .A(
        n12004), .ZN(n15708) );
  INV_X1 U15191 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n21725) );
  NAND2_X1 U15192 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12006) );
  AOI22_X1 U15193 ( .A1(n12378), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12005) );
  OAI211_X1 U15194 ( .C1(n12376), .C2(n21725), .A(n12006), .B(n12005), .ZN(
        n15700) );
  INV_X1 U15195 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n21822) );
  NAND2_X1 U15196 ( .A1(n12366), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12008) );
  NAND2_X1 U15197 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12007) );
  OAI211_X1 U15198 ( .C1(n12376), .C2(n21822), .A(n12008), .B(n12007), .ZN(
        n12009) );
  AOI21_X1 U15199 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n12377), .A(
        n12009), .ZN(n15676) );
  INV_X1 U15200 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20725) );
  NAND2_X1 U15201 ( .A1(n12366), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12013) );
  NAND2_X1 U15202 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12012) );
  OAI211_X1 U15203 ( .C1(n12376), .C2(n20725), .A(n12013), .B(n12012), .ZN(
        n12014) );
  AOI21_X1 U15204 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n12377), .A(
        n12014), .ZN(n15665) );
  INV_X1 U15205 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20726) );
  NAND2_X1 U15206 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12016) );
  AOI22_X1 U15207 ( .A1(n12378), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12015) );
  OAI211_X1 U15208 ( .C1(n12376), .C2(n20726), .A(n12016), .B(n12015), .ZN(
        n15646) );
  INV_X1 U15209 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20729) );
  NAND2_X1 U15210 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12018) );
  AOI22_X1 U15211 ( .A1(n12378), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12017) );
  OAI211_X1 U15212 ( .C1(n12376), .C2(n20729), .A(n12018), .B(n12017), .ZN(
        n12020) );
  OR2_X1 U15213 ( .A1(n12019), .A2(n12020), .ZN(n12021) );
  NAND2_X1 U15214 ( .A1(n16904), .A2(n16029), .ZN(n12025) );
  OAI211_X1 U15215 ( .C1(n12024), .C2(n20118), .A(n12023), .B(n20810), .ZN(
        n16774) );
  INV_X1 U15216 ( .A(n11892), .ZN(n12036) );
  OR2_X1 U15217 ( .A1(n16774), .A2(n12036), .ZN(n16800) );
  NAND2_X1 U15218 ( .A1(n12025), .A2(n16800), .ZN(n12026) );
  NAND2_X1 U15219 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16565) );
  INV_X1 U15220 ( .A(n16565), .ZN(n12027) );
  AND2_X1 U15221 ( .A1(n16567), .A2(n12027), .ZN(n12443) );
  NAND2_X1 U15222 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n12443), .ZN(
        n12057) );
  INV_X1 U15223 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12032) );
  NAND3_X1 U15224 ( .A1(n16029), .A2(n12028), .A3(n20127), .ZN(n12029) );
  NAND2_X1 U15225 ( .A1(n12255), .A2(n16896), .ZN(n12453) );
  NAND2_X1 U15226 ( .A1(n13579), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12030) );
  NAND2_X1 U15227 ( .A1(n12453), .A2(n12030), .ZN(n12031) );
  INV_X1 U15228 ( .A(n13579), .ZN(n14665) );
  INV_X1 U15229 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12053) );
  NAND2_X1 U15230 ( .A1(n14665), .A2(n12053), .ZN(n12050) );
  NAND2_X1 U15231 ( .A1(n12031), .A2(n12050), .ZN(n14316) );
  NOR2_X1 U15232 ( .A1(n12032), .A2(n14316), .ZN(n16749) );
  NAND2_X1 U15233 ( .A1(n16775), .A2(n12033), .ZN(n12034) );
  NAND2_X1 U15234 ( .A1(n12034), .A2(n20118), .ZN(n12046) );
  INV_X1 U15235 ( .A(n20810), .ZN(n12038) );
  NAND2_X1 U15236 ( .A1(n12036), .A2(n12035), .ZN(n12037) );
  AOI22_X1 U15237 ( .A1(n12038), .A2(n12037), .B1(n20807), .B2(n20113), .ZN(
        n12043) );
  NAND2_X1 U15238 ( .A1(n12040), .A2(n12039), .ZN(n12394) );
  INV_X1 U15239 ( .A(n11466), .ZN(n12074) );
  OAI211_X1 U15240 ( .C1(n12074), .C2(n16887), .A(n12041), .B(n11892), .ZN(
        n12042) );
  AND4_X1 U15241 ( .A1(n12044), .A2(n12043), .A3(n12394), .A4(n12042), .ZN(
        n12045) );
  NAND2_X1 U15242 ( .A1(n16816), .A2(n16799), .ZN(n12047) );
  NAND2_X1 U15243 ( .A1(n16749), .A2(n16568), .ZN(n16768) );
  NAND2_X1 U15244 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16732) );
  INV_X1 U15245 ( .A(n16732), .ZN(n12048) );
  NAND2_X1 U15246 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12048), .ZN(
        n12049) );
  NOR2_X1 U15247 ( .A1(n16701), .A2(n16722), .ZN(n16700) );
  NOR2_X1 U15248 ( .A1(n12057), .A2(n16685), .ZN(n16540) );
  NAND3_X1 U15249 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n16540), .ZN(n12064) );
  INV_X1 U15250 ( .A(n12064), .ZN(n16511) );
  NAND2_X1 U15251 ( .A1(n16511), .A2(n16525), .ZN(n16524) );
  NAND2_X1 U15252 ( .A1(n16568), .A2(n16732), .ZN(n16751) );
  NOR2_X1 U15253 ( .A1(n17615), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14325) );
  OR2_X1 U15254 ( .A1(n20804), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13413) );
  INV_X2 U15255 ( .A(n16464), .ZN(n16754) );
  INV_X1 U15256 ( .A(n14670), .ZN(n12054) );
  INV_X1 U15257 ( .A(n12453), .ZN(n14664) );
  INV_X1 U15258 ( .A(n12050), .ZN(n12051) );
  NAND2_X1 U15259 ( .A1(n14664), .A2(n12051), .ZN(n14663) );
  INV_X1 U15260 ( .A(n12052), .ZN(n12457) );
  NAND2_X1 U15261 ( .A1(n12457), .A2(n12053), .ZN(n14667) );
  NAND3_X1 U15262 ( .A1(n12054), .A2(n14663), .A3(n14667), .ZN(n14321) );
  NOR2_X1 U15263 ( .A1(n17615), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12055) );
  NOR2_X1 U15264 ( .A1(n17615), .A2(n16700), .ZN(n12056) );
  NAND2_X1 U15265 ( .A1(n16568), .A2(n12057), .ZN(n12058) );
  NAND2_X1 U15266 ( .A1(n16687), .A2(n12058), .ZN(n16538) );
  NOR2_X1 U15267 ( .A1(n16539), .A2(n16556), .ZN(n12059) );
  NOR2_X1 U15268 ( .A1(n17615), .A2(n12059), .ZN(n12060) );
  NOR2_X1 U15269 ( .A1(n16538), .A2(n12060), .ZN(n16526) );
  NAND2_X1 U15270 ( .A1(n16568), .A2(n10710), .ZN(n12061) );
  NAND2_X1 U15271 ( .A1(n12062), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12063) );
  NOR2_X1 U15272 ( .A1(n12064), .A2(n12063), .ZN(n16486) );
  NAND2_X1 U15273 ( .A1(n16754), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12271) );
  INV_X1 U15274 ( .A(n12271), .ZN(n12065) );
  AOI21_X1 U15275 ( .B1(n16486), .B2(n14630), .A(n12065), .ZN(n12066) );
  OAI21_X1 U15276 ( .B1(n16491), .B2(n14630), .A(n12066), .ZN(n12257) );
  INV_X1 U15277 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12067) );
  OAI21_X1 U15278 ( .B1(n16029), .B2(n12067), .A(n20800), .ZN(n12068) );
  INV_X1 U15279 ( .A(n12068), .ZN(n12071) );
  NAND2_X1 U15280 ( .A1(n12069), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12070) );
  NAND2_X1 U15281 ( .A1(n12074), .A2(n12077), .ZN(n12088) );
  MUX2_X1 U15282 ( .A(n16873), .B(n20786), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12075) );
  NAND2_X1 U15283 ( .A1(n13953), .A2(n13954), .ZN(n13955) );
  NOR2_X1 U15284 ( .A1(n16873), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15285 ( .A1(n12091), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12078) );
  OAI21_X1 U15286 ( .B1(n12090), .B2(n20692), .A(n12078), .ZN(n12084) );
  XNOR2_X1 U15287 ( .A(n13955), .B(n12084), .ZN(n13585) );
  NAND2_X1 U15288 ( .A1(n11466), .A2(n16873), .ZN(n12079) );
  MUX2_X1 U15289 ( .A(n12079), .B(n20776), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12083) );
  INV_X1 U15290 ( .A(n12080), .ZN(n12081) );
  OR2_X1 U15291 ( .A1(n12220), .A2(n12081), .ZN(n12082) );
  AND2_X1 U15292 ( .A1(n12083), .A2(n12082), .ZN(n13584) );
  INV_X1 U15293 ( .A(n12084), .ZN(n12085) );
  NAND2_X1 U15294 ( .A1(n13955), .A2(n12085), .ZN(n12086) );
  NAND2_X1 U15295 ( .A1(n13587), .A2(n12086), .ZN(n12096) );
  OR2_X1 U15296 ( .A1(n12220), .A2(n12087), .ZN(n12089) );
  OAI211_X1 U15297 ( .C1(n20800), .C2(n20766), .A(n12089), .B(n12088), .ZN(
        n12094) );
  XNOR2_X1 U15298 ( .A(n12096), .B(n12094), .ZN(n14073) );
  NAND2_X1 U15299 ( .A1(n12282), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15300 ( .A1(n12283), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12092) );
  AND2_X1 U15301 ( .A1(n12093), .A2(n12092), .ZN(n14072) );
  NAND2_X2 U15302 ( .A1(n14073), .A2(n14072), .ZN(n14075) );
  INV_X1 U15303 ( .A(n12094), .ZN(n12095) );
  NAND2_X1 U15304 ( .A1(n12096), .A2(n12095), .ZN(n12097) );
  NAND2_X1 U15305 ( .A1(n12282), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15306 ( .A1(n12283), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12100) );
  OR2_X1 U15307 ( .A1(n12220), .A2(n12098), .ZN(n12099) );
  INV_X1 U15308 ( .A(n12220), .ZN(n12207) );
  OAI22_X1 U15309 ( .A1(n12196), .A2(n12032), .B1(n20758), .B2(n20800), .ZN(
        n12102) );
  AOI21_X1 U15310 ( .B1(n12282), .B2(P2_REIP_REG_3__SCAN_IN), .A(n12102), .ZN(
        n12103) );
  NAND2_X1 U15311 ( .A1(n12282), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15312 ( .A1(n12283), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12107) );
  OR2_X1 U15313 ( .A1(n12220), .A2(n12105), .ZN(n12106) );
  AOI22_X1 U15314 ( .A1(n12283), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12110) );
  OAI21_X1 U15315 ( .B1(n12090), .B2(n20698), .A(n12110), .ZN(n14060) );
  NAND2_X1 U15316 ( .A1(n14059), .A2(n14060), .ZN(n12112) );
  OR2_X1 U15317 ( .A1(n12220), .A2(n14606), .ZN(n12111) );
  NAND2_X1 U15318 ( .A1(n12112), .A2(n12111), .ZN(n14057) );
  AOI22_X1 U15319 ( .A1(n12283), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12113) );
  OAI21_X1 U15320 ( .B1(n12090), .B2(n20700), .A(n12113), .ZN(n14056) );
  NAND2_X1 U15321 ( .A1(n14057), .A2(n14056), .ZN(n14046) );
  NAND2_X1 U15322 ( .A1(n12282), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12126) );
  AOI22_X1 U15323 ( .A1(n12283), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15324 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11909), .B1(
        n12625), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15325 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15326 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15327 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12626), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12114) );
  NAND4_X1 U15328 ( .A1(n12117), .A2(n12116), .A3(n12115), .A4(n12114), .ZN(
        n12123) );
  AOI22_X1 U15329 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12121) );
  AOI22_X1 U15330 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15331 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15332 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12632), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12118) );
  NAND4_X1 U15333 ( .A1(n12121), .A2(n12120), .A3(n12119), .A4(n12118), .ZN(
        n12122) );
  NAND2_X1 U15334 ( .A1(n12207), .A2(n14216), .ZN(n12124) );
  NAND2_X1 U15335 ( .A1(n12128), .A2(n12127), .ZN(n14042) );
  NAND2_X1 U15336 ( .A1(n12282), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15337 ( .A1(n12283), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12077), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15338 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11567), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15339 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15340 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12625), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12130) );
  AOI22_X1 U15341 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11641), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12129) );
  NAND4_X1 U15342 ( .A1(n12132), .A2(n12131), .A3(n12130), .A4(n12129), .ZN(
        n12138) );
  AOI22_X1 U15343 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11573), .B1(
        n11596), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12136) );
  AOI22_X1 U15344 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11630), .B1(
        n12588), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12135) );
  AOI22_X1 U15345 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11559), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12134) );
  AOI22_X1 U15346 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12632), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12133) );
  NAND4_X1 U15347 ( .A1(n12136), .A2(n12135), .A3(n12134), .A4(n12133), .ZN(
        n12137) );
  NOR2_X1 U15348 ( .A1(n12138), .A2(n12137), .ZN(n12547) );
  OR2_X1 U15349 ( .A1(n12220), .A2(n12547), .ZN(n12139) );
  NAND2_X1 U15350 ( .A1(n12282), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15351 ( .A1(n12283), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12154) );
  AOI22_X1 U15352 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15353 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15354 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15355 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12143) );
  NAND4_X1 U15356 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12152) );
  AOI22_X1 U15357 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15358 ( .A1(n12626), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15359 ( .A1(n11560), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15360 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11559), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15361 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12151) );
  NAND2_X1 U15362 ( .A1(n12207), .A2(n14032), .ZN(n12153) );
  AOI22_X1 U15363 ( .A1(n12283), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15364 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15365 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15366 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15367 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12156) );
  NAND4_X1 U15368 ( .A1(n12159), .A2(n12158), .A3(n12157), .A4(n12156), .ZN(
        n12165) );
  AOI22_X1 U15369 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15370 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15371 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15372 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12160) );
  NAND4_X1 U15373 ( .A1(n12163), .A2(n12162), .A3(n12161), .A4(n12160), .ZN(
        n12164) );
  NAND2_X1 U15374 ( .A1(n12207), .A2(n14151), .ZN(n12166) );
  OAI211_X1 U15375 ( .C1(n12090), .C2(n21738), .A(n12167), .B(n12166), .ZN(
        n14053) );
  NAND2_X1 U15376 ( .A1(n12282), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15377 ( .A1(n12283), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15378 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12625), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15379 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15380 ( .A1(n11637), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15381 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12168) );
  NAND4_X1 U15382 ( .A1(n12171), .A2(n12170), .A3(n12169), .A4(n12168), .ZN(
        n12177) );
  AOI22_X1 U15383 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15384 ( .A1(n12626), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15385 ( .A1(n11560), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15386 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11559), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12172) );
  NAND4_X1 U15387 ( .A1(n12175), .A2(n12174), .A3(n12173), .A4(n12172), .ZN(
        n12176) );
  NOR2_X1 U15388 ( .A1(n12177), .A2(n12176), .ZN(n12549) );
  OR2_X1 U15389 ( .A1(n12220), .A2(n12549), .ZN(n12178) );
  NAND2_X1 U15390 ( .A1(n12182), .A2(n12181), .ZN(n13392) );
  NAND2_X1 U15391 ( .A1(n12282), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15392 ( .A1(n12283), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15393 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15394 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15395 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15396 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12183) );
  NAND4_X1 U15397 ( .A1(n12186), .A2(n12185), .A3(n12184), .A4(n12183), .ZN(
        n12192) );
  AOI22_X1 U15398 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15399 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15400 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15401 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12187) );
  NAND4_X1 U15402 ( .A1(n12190), .A2(n12189), .A3(n12188), .A4(n12187), .ZN(
        n12191) );
  NOR2_X1 U15403 ( .A1(n12192), .A2(n12191), .ZN(n14350) );
  OR2_X1 U15404 ( .A1(n12220), .A2(n14350), .ZN(n12193) );
  AOI22_X1 U15405 ( .A1(n12283), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15406 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15407 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15408 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15409 ( .A1(n12626), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15410 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12206) );
  AOI22_X1 U15411 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15412 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11641), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15413 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15414 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12201) );
  NAND4_X1 U15415 ( .A1(n12204), .A2(n12203), .A3(n12202), .A4(n12201), .ZN(
        n12205) );
  NAND2_X1 U15416 ( .A1(n12207), .A2(n16087), .ZN(n12208) );
  OAI211_X1 U15417 ( .C1(n12090), .C2(n15833), .A(n12209), .B(n12208), .ZN(
        n14271) );
  AOI22_X1 U15418 ( .A1(n12283), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15419 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15420 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15421 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15422 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12210) );
  NAND4_X1 U15423 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12219) );
  AOI22_X1 U15424 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12217) );
  AOI22_X1 U15425 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15426 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15427 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12214) );
  NAND4_X1 U15428 ( .A1(n12217), .A2(n12216), .A3(n12215), .A4(n12214), .ZN(
        n12218) );
  NOR2_X1 U15429 ( .A1(n12219), .A2(n12218), .ZN(n12552) );
  OR2_X1 U15430 ( .A1(n12220), .A2(n12552), .ZN(n12221) );
  OAI211_X1 U15431 ( .C1(n12090), .C2(n20712), .A(n12222), .B(n12221), .ZN(
        n14356) );
  NAND2_X1 U15432 ( .A1(n12282), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15433 ( .A1(n12283), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12223) );
  NAND2_X1 U15434 ( .A1(n12282), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15435 ( .A1(n12283), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15436 ( .A1(n12283), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12227) );
  OAI21_X1 U15437 ( .B1(n12090), .B2(n12228), .A(n12227), .ZN(n15767) );
  NAND2_X1 U15438 ( .A1(n12282), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15439 ( .A1(n12283), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12229) );
  NAND2_X1 U15440 ( .A1(n12282), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12234) );
  AOI22_X1 U15441 ( .A1(n12283), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12233) );
  NAND2_X1 U15442 ( .A1(n12282), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15443 ( .A1(n12283), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15444 ( .A1(n12283), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12237) );
  OAI21_X1 U15445 ( .B1(n12090), .B2(n12238), .A(n12237), .ZN(n15707) );
  NAND2_X1 U15446 ( .A1(n12435), .A2(n15707), .ZN(n15690) );
  NAND2_X1 U15447 ( .A1(n12282), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15448 ( .A1(n12283), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12239) );
  NOR2_X2 U15449 ( .A1(n15690), .A2(n15691), .ZN(n15672) );
  NAND2_X1 U15450 ( .A1(n12282), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15451 ( .A1(n12283), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12241) );
  AND2_X1 U15452 ( .A1(n12242), .A2(n12241), .ZN(n15673) );
  INV_X1 U15453 ( .A(n15673), .ZN(n12243) );
  AOI22_X1 U15454 ( .A1(n12283), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12244) );
  OAI21_X1 U15455 ( .B1(n12090), .B2(n20725), .A(n12244), .ZN(n15659) );
  AOI22_X1 U15456 ( .A1(n12283), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12245) );
  OAI21_X1 U15457 ( .B1(n12090), .B2(n20726), .A(n12245), .ZN(n15645) );
  NAND2_X1 U15458 ( .A1(n12282), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12247) );
  AOI22_X1 U15459 ( .A1(n12283), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12246) );
  AND2_X1 U15460 ( .A1(n12247), .A2(n12246), .ZN(n12249) );
  NAND2_X1 U15461 ( .A1(n12248), .A2(n12249), .ZN(n12250) );
  NAND2_X1 U15462 ( .A1(n14628), .A2(n12250), .ZN(n16111) );
  INV_X1 U15463 ( .A(n12251), .ZN(n12252) );
  NAND2_X1 U15464 ( .A1(n13529), .A2(n11478), .ZN(n16899) );
  NAND2_X1 U15465 ( .A1(n16899), .A2(n16887), .ZN(n12253) );
  NAND2_X1 U15466 ( .A1(n16803), .A2(n12253), .ZN(n12254) );
  NOR2_X1 U15467 ( .A1(n16111), .A2(n16763), .ZN(n12256) );
  AOI211_X1 U15468 ( .C1(n16009), .C2(n17604), .A(n12257), .B(n12256), .ZN(
        n12258) );
  NAND2_X1 U15469 ( .A1(n12263), .A2(n12262), .ZN(n12264) );
  OR2_X2 U15470 ( .A1(n13424), .A2(n16029), .ZN(n16472) );
  INV_X1 U15471 ( .A(n16472), .ZN(n17587) );
  INV_X1 U15472 ( .A(n13424), .ZN(n12266) );
  NOR2_X1 U15473 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16943) );
  INV_X1 U15474 ( .A(n16943), .ZN(n20747) );
  NAND2_X1 U15475 ( .A1(n20804), .A2(n20747), .ZN(n20777) );
  NAND2_X1 U15476 ( .A1(n20777), .A2(n20808), .ZN(n12267) );
  AND2_X1 U15477 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12268) );
  INV_X1 U15478 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21876) );
  NAND2_X1 U15479 ( .A1(n12317), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12319) );
  INV_X1 U15480 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16283) );
  INV_X1 U15481 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n21644) );
  INV_X1 U15482 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16263) );
  NAND2_X1 U15483 ( .A1(n12352), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12353) );
  INV_X1 U15484 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16242) );
  AND2_X1 U15485 ( .A1(n12356), .A2(n21876), .ZN(n12269) );
  NOR2_X1 U15486 ( .A1(n12358), .A2(n12269), .ZN(n15635) );
  NAND2_X1 U15487 ( .A1(n20395), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12270) );
  NAND2_X1 U15488 ( .A1(n16839), .A2(n12270), .ZN(n13565) );
  NAND2_X1 U15489 ( .A1(n15635), .A2(n17586), .ZN(n12272) );
  OAI211_X1 U15490 ( .C1(n21876), .C2(n17599), .A(n12272), .B(n12271), .ZN(
        n12273) );
  AOI21_X1 U15491 ( .B1(n16009), .B2(n16454), .A(n12273), .ZN(n12274) );
  OAI21_X1 U15492 ( .B1(n12261), .B2(n12278), .A(n12277), .ZN(P2_U2987) );
  NAND2_X1 U15493 ( .A1(n12282), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15494 ( .A1(n12283), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12279) );
  INV_X1 U15495 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20731) );
  AOI22_X1 U15496 ( .A1(n12283), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12281) );
  OAI21_X1 U15497 ( .B1(n12090), .B2(n20731), .A(n12281), .ZN(n15610) );
  NAND2_X1 U15498 ( .A1(n15611), .A2(n15610), .ZN(n15609) );
  NAND2_X1 U15499 ( .A1(n12282), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n12285) );
  AOI22_X1 U15500 ( .A1(n12283), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12284) );
  NAND2_X1 U15501 ( .A1(n14680), .A2(n10716), .ZN(n14682) );
  INV_X1 U15502 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15503 ( .A1(n12283), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n12077), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12286) );
  OAI21_X1 U15504 ( .B1(n12090), .B2(n12381), .A(n12286), .ZN(n12287) );
  INV_X1 U15505 ( .A(n20805), .ZN(n13415) );
  NAND2_X1 U15506 ( .A1(n13527), .A2(n20395), .ZN(n12297) );
  INV_X1 U15507 ( .A(n12297), .ZN(n12288) );
  AND2_X1 U15508 ( .A1(n12289), .A2(n12288), .ZN(n16932) );
  NAND2_X1 U15509 ( .A1(n12509), .A2(n15982), .ZN(n12391) );
  NAND2_X1 U15510 ( .A1(n12290), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12486) );
  NAND2_X1 U15511 ( .A1(n12290), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12478) );
  NOR2_X1 U15512 ( .A1(n12476), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12291) );
  MUX2_X1 U15513 ( .A(n15651), .B(n12291), .S(n12290), .Z(n12480) );
  INV_X1 U15514 ( .A(n12480), .ZN(n12364) );
  NAND2_X1 U15515 ( .A1(n20812), .A2(n20395), .ZN(n13385) );
  AND3_X1 U15516 ( .A1(n12386), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n13385), .ZN(
        n12292) );
  INV_X1 U15517 ( .A(n15984), .ZN(n12363) );
  NOR2_X1 U15518 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12293) );
  NAND2_X1 U15519 ( .A1(n16838), .A2(n12293), .ZN(n16947) );
  NOR2_X1 U15520 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13406) );
  AND2_X1 U15521 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12294) );
  NAND2_X1 U15522 ( .A1(n13406), .A2(n12294), .ZN(n16934) );
  NAND2_X1 U15523 ( .A1(n16947), .A2(n16934), .ZN(n12295) );
  NOR2_X1 U15524 ( .A1(n16754), .A2(n12295), .ZN(n12296) );
  INV_X1 U15525 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12301) );
  NAND2_X1 U15526 ( .A1(n16897), .A2(n20026), .ZN(n13411) );
  AOI22_X1 U15527 ( .A1(n19985), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13388), 
        .B2(P2_EBX_REG_31__SCAN_IN), .ZN(n12298) );
  OAI21_X1 U15528 ( .B1(n15968), .B2(n12301), .A(n12298), .ZN(n12299) );
  INV_X1 U15529 ( .A(n12299), .ZN(n12362) );
  NAND2_X1 U15530 ( .A1(n12357), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12360) );
  INV_X1 U15531 ( .A(n12360), .ZN(n12300) );
  NAND2_X1 U15532 ( .A1(n12300), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12302) );
  INV_X1 U15533 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12503) );
  INV_X1 U15534 ( .A(n12306), .ZN(n12305) );
  INV_X1 U15535 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12303) );
  NAND2_X1 U15536 ( .A1(n13570), .A2(n12303), .ZN(n12304) );
  NAND2_X1 U15537 ( .A1(n12305), .A2(n12304), .ZN(n15952) );
  AND2_X1 U15538 ( .A1(n15965), .A2(n15952), .ZN(n15938) );
  OAI21_X1 U15539 ( .B1(n12306), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n12308), .ZN(n15940) );
  AND2_X1 U15540 ( .A1(n12308), .A2(n16466), .ZN(n12309) );
  NOR2_X1 U15541 ( .A1(n12307), .A2(n12309), .ZN(n19991) );
  OR2_X1 U15542 ( .A1(n12307), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12310) );
  AND2_X1 U15543 ( .A1(n12312), .A2(n12310), .ZN(n17585) );
  NAND2_X1 U15544 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  NAND2_X1 U15545 ( .A1(n12315), .A2(n12313), .ZN(n16447) );
  AND2_X1 U15546 ( .A1(n12315), .A2(n16437), .ZN(n12316) );
  NOR2_X1 U15547 ( .A1(n12314), .A2(n12316), .ZN(n16440) );
  OR2_X1 U15548 ( .A1(n15901), .A2(n16440), .ZN(n15886) );
  NOR2_X1 U15549 ( .A1(n12314), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12318) );
  OR2_X1 U15550 ( .A1(n12317), .A2(n12318), .ZN(n16427) );
  INV_X1 U15551 ( .A(n16427), .ZN(n15888) );
  NOR2_X1 U15552 ( .A1(n15886), .A2(n15888), .ZN(n15874) );
  OR2_X1 U15553 ( .A1(n12317), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12320) );
  NAND2_X1 U15554 ( .A1(n12319), .A2(n12320), .ZN(n16413) );
  AND2_X1 U15555 ( .A1(n15874), .A2(n16413), .ZN(n15863) );
  NAND2_X1 U15556 ( .A1(n12319), .A2(n12321), .ZN(n12322) );
  NAND2_X1 U15557 ( .A1(n12323), .A2(n12322), .ZN(n16404) );
  NAND2_X1 U15558 ( .A1(n12323), .A2(n16397), .ZN(n12324) );
  AND2_X1 U15559 ( .A1(n12325), .A2(n12324), .ZN(n16395) );
  AND2_X1 U15560 ( .A1(n12325), .A2(n16379), .ZN(n12326) );
  NOR2_X1 U15561 ( .A1(n12328), .A2(n12326), .ZN(n16382) );
  OR2_X1 U15562 ( .A1(n12328), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12329) );
  NAND2_X1 U15563 ( .A1(n12327), .A2(n12329), .ZN(n16370) );
  NAND2_X1 U15564 ( .A1(n12327), .A2(n16359), .ZN(n12330) );
  AND2_X1 U15565 ( .A1(n12331), .A2(n12330), .ZN(n16357) );
  OR2_X1 U15566 ( .A1(n15825), .A2(n16357), .ZN(n15811) );
  AND2_X1 U15567 ( .A1(n12331), .A2(n16346), .ZN(n12332) );
  NOR2_X1 U15568 ( .A1(n12334), .A2(n12332), .ZN(n16348) );
  OR2_X1 U15569 ( .A1(n15811), .A2(n16348), .ZN(n15803) );
  NOR2_X1 U15570 ( .A1(n12334), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12335) );
  OR2_X1 U15571 ( .A1(n12333), .A2(n12335), .ZN(n16335) );
  INV_X1 U15572 ( .A(n16335), .ZN(n15804) );
  NOR2_X1 U15573 ( .A1(n15803), .A2(n15804), .ZN(n15789) );
  OR2_X1 U15574 ( .A1(n12333), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12337) );
  NAND2_X1 U15575 ( .A1(n12336), .A2(n12337), .ZN(n16328) );
  NAND2_X1 U15576 ( .A1(n15789), .A2(n16328), .ZN(n15779) );
  NAND2_X1 U15577 ( .A1(n12336), .A2(n16316), .ZN(n12338) );
  AND2_X1 U15578 ( .A1(n12339), .A2(n12338), .ZN(n16318) );
  OR2_X1 U15579 ( .A1(n15779), .A2(n16318), .ZN(n15755) );
  AND2_X1 U15580 ( .A1(n12339), .A2(n16306), .ZN(n12340) );
  NOR2_X1 U15581 ( .A1(n12342), .A2(n12340), .ZN(n16308) );
  NOR2_X1 U15582 ( .A1(n12342), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12343) );
  OR2_X1 U15583 ( .A1(n12341), .A2(n12343), .ZN(n16297) );
  OR2_X1 U15584 ( .A1(n12341), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12344) );
  AND2_X1 U15585 ( .A1(n12345), .A2(n12344), .ZN(n15719) );
  NAND2_X1 U15586 ( .A1(n12345), .A2(n16283), .ZN(n12346) );
  NAND2_X1 U15587 ( .A1(n12348), .A2(n12346), .ZN(n16286) );
  NAND2_X1 U15588 ( .A1(n15710), .A2(n16286), .ZN(n15695) );
  NAND2_X1 U15589 ( .A1(n12348), .A2(n21644), .ZN(n12349) );
  NAND2_X1 U15590 ( .A1(n12350), .A2(n12349), .ZN(n15694) );
  AND2_X1 U15591 ( .A1(n12350), .A2(n16263), .ZN(n12351) );
  OR2_X1 U15592 ( .A1(n12351), .A2(n12352), .ZN(n16266) );
  OR2_X1 U15593 ( .A1(n12352), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12354) );
  AND2_X1 U15594 ( .A1(n12354), .A2(n12353), .ZN(n16249) );
  NAND2_X1 U15595 ( .A1(n12353), .A2(n16242), .ZN(n12355) );
  NAND2_X1 U15596 ( .A1(n12356), .A2(n12355), .ZN(n16241) );
  OAI21_X1 U15597 ( .B1(n15662), .B2(n10319), .A(n16241), .ZN(n15634) );
  AOI21_X1 U15598 ( .B1(n15634), .B2(n15967), .A(n15635), .ZN(n15627) );
  NOR2_X1 U15599 ( .A1(n12358), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12359) );
  OR2_X1 U15600 ( .A1(n12357), .A2(n12359), .ZN(n15628) );
  OR2_X1 U15601 ( .A1(n12357), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12361) );
  AND2_X1 U15602 ( .A1(n12360), .A2(n12361), .ZN(n16230) );
  XOR2_X1 U15603 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12360), .Z(
        n16221) );
  OAI21_X1 U15604 ( .B1(n15617), .B2(n10319), .A(n16221), .ZN(n14683) );
  INV_X1 U15605 ( .A(n12365), .ZN(n12390) );
  INV_X1 U15606 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12369) );
  NAND2_X1 U15607 ( .A1(n12366), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12368) );
  NAND2_X1 U15608 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12367) );
  OAI211_X1 U15609 ( .C1(n12376), .C2(n12369), .A(n12368), .B(n12367), .ZN(
        n12370) );
  AOI21_X1 U15610 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12377), .A(
        n12370), .ZN(n14610) );
  AOI22_X1 U15611 ( .A1(n12378), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12372) );
  OAI21_X1 U15612 ( .B1(n12376), .B2(n20731), .A(n12372), .ZN(n12373) );
  AOI21_X1 U15613 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n12377), .A(
        n12373), .ZN(n15613) );
  INV_X1 U15614 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n16218) );
  NAND2_X1 U15615 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12375) );
  AOI22_X1 U15616 ( .A1(n12378), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12374) );
  OAI211_X1 U15617 ( .C1(n12376), .C2(n16218), .A(n12375), .B(n12374), .ZN(
        n12798) );
  NAND2_X1 U15618 ( .A1(n15616), .A2(n12798), .ZN(n12384) );
  NAND2_X1 U15619 ( .A1(n12377), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12380) );
  AOI22_X1 U15620 ( .A1(n12378), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12379) );
  OAI211_X1 U15621 ( .C1(n12382), .C2(n12381), .A(n12380), .B(n12379), .ZN(
        n12383) );
  INV_X1 U15622 ( .A(n13385), .ZN(n12385) );
  NAND2_X1 U15623 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  NAND3_X1 U15624 ( .A1(n12391), .A2(n12390), .A3(n12389), .ZN(P2_U2824) );
  NAND2_X1 U15625 ( .A1(n16894), .A2(n16896), .ZN(n12393) );
  AND2_X1 U15626 ( .A1(n20810), .A2(n20812), .ZN(n13420) );
  NAND2_X1 U15627 ( .A1(n13422), .A2(n13420), .ZN(n12392) );
  OAI21_X4 U15628 ( .B1(n13526), .B2(n12395), .A(n20026), .ZN(n16191) );
  OR2_X1 U15629 ( .A1(n16191), .A2(n16873), .ZN(n20002) );
  NAND2_X1 U15630 ( .A1(n12509), .A2(n20016), .ZN(n12412) );
  NAND2_X1 U15631 ( .A1(n16873), .A2(n20135), .ZN(n12396) );
  NOR4_X1 U15632 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12400) );
  NOR4_X1 U15633 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n12399) );
  NOR4_X1 U15634 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12398) );
  NOR4_X1 U15635 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12397) );
  AND4_X1 U15636 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12405) );
  NOR4_X1 U15637 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12403) );
  NOR4_X1 U15638 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12402) );
  NOR4_X1 U15639 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12401) );
  INV_X1 U15640 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20696) );
  AND4_X1 U15641 ( .A1(n12403), .A2(n12402), .A3(n12401), .A4(n20696), .ZN(
        n12404) );
  NAND2_X1 U15642 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  NOR2_X2 U15643 ( .A1(n13952), .A2(n16847), .ZN(n16194) );
  AOI22_X1 U15644 ( .A1(n16194), .A2(BUF2_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n16191), .ZN(n12407) );
  INV_X1 U15645 ( .A(n12407), .ZN(n12410) );
  INV_X1 U15646 ( .A(n13952), .ZN(n12408) );
  INV_X1 U15647 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n13371) );
  NOR2_X1 U15648 ( .A1(n16197), .A2(n13371), .ZN(n12409) );
  NOR2_X1 U15649 ( .A1(n12410), .A2(n12409), .ZN(n12411) );
  NAND2_X1 U15650 ( .A1(n12412), .A2(n12411), .ZN(P2_U2888) );
  INV_X1 U15651 ( .A(n12413), .ZN(n12414) );
  INV_X1 U15652 ( .A(n12417), .ZN(n12418) );
  INV_X1 U15653 ( .A(n12420), .ZN(n14697) );
  NAND2_X1 U15654 ( .A1(n12424), .A2(n12423), .ZN(n12459) );
  INV_X1 U15655 ( .A(n16293), .ZN(n12426) );
  AOI21_X2 U15656 ( .B1(n16291), .B2(n12427), .A(n12426), .ZN(n12431) );
  NAND2_X1 U15657 ( .A1(n12429), .A2(n12428), .ZN(n12430) );
  XNOR2_X1 U15658 ( .A(n12431), .B(n12430), .ZN(n12516) );
  AND2_X1 U15659 ( .A1(n12437), .A2(n12438), .ZN(n12439) );
  NOR2_X1 U15660 ( .A1(n12436), .A2(n12439), .ZN(n16157) );
  NAND2_X1 U15661 ( .A1(n16157), .A2(n17608), .ZN(n12450) );
  NAND2_X1 U15662 ( .A1(n15733), .A2(n12441), .ZN(n12442) );
  NAND2_X1 U15663 ( .A1(n15709), .A2(n12442), .ZN(n16048) );
  INV_X1 U15664 ( .A(n16048), .ZN(n15726) );
  NAND2_X1 U15665 ( .A1(n12443), .A2(n21805), .ZN(n12447) );
  OAI21_X1 U15666 ( .B1(n17615), .B2(n12443), .A(n16687), .ZN(n12445) );
  NAND2_X1 U15667 ( .A1(n16754), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12511) );
  INV_X1 U15668 ( .A(n12511), .ZN(n12444) );
  AOI21_X1 U15669 ( .B1(n12445), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n12444), .ZN(n12446) );
  OAI21_X1 U15670 ( .B1(n16685), .B2(n12447), .A(n12446), .ZN(n12448) );
  AOI21_X1 U15671 ( .B1(n15726), .B2(n17604), .A(n12448), .ZN(n12449) );
  OAI21_X1 U15672 ( .B1(n12516), .B2(n10442), .A(n10713), .ZN(P2_U3025) );
  INV_X1 U15673 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14706) );
  INV_X1 U15674 ( .A(n12454), .ZN(n12455) );
  NAND2_X1 U15675 ( .A1(n16568), .A2(n12455), .ZN(n12456) );
  NAND2_X1 U15676 ( .A1(n16687), .A2(n12456), .ZN(n16608) );
  INV_X1 U15677 ( .A(n12460), .ZN(n12461) );
  NOR2_X1 U15678 ( .A1(n16620), .A2(n16356), .ZN(n16615) );
  AOI22_X1 U15679 ( .A1(n16322), .A2(n17606), .B1(n12462), .B2(n16615), .ZN(
        n12470) );
  OR2_X1 U15680 ( .A1(n12463), .A2(n12465), .ZN(n15771) );
  INV_X1 U15681 ( .A(n15771), .ZN(n12464) );
  AOI21_X1 U15682 ( .B1(n12465), .B2(n12463), .A(n12464), .ZN(n16324) );
  NOR2_X1 U15683 ( .A1(n16464), .A2(n20715), .ZN(n16325) );
  AOI21_X1 U15684 ( .B1(n16324), .B2(n17604), .A(n16325), .ZN(n12469) );
  AND2_X1 U15685 ( .A1(n14701), .A2(n12466), .ZN(n12467) );
  NOR2_X1 U15686 ( .A1(n15768), .A2(n12467), .ZN(n16187) );
  NAND2_X1 U15687 ( .A1(n16187), .A2(n17608), .ZN(n12468) );
  OAI211_X1 U15688 ( .C1(n12470), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n12469), .B(n12468), .ZN(n12471) );
  INV_X1 U15689 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n12474) );
  NOR2_X1 U15690 ( .A1(n20127), .A2(n12474), .ZN(n12475) );
  XNOR2_X1 U15691 ( .A(n12476), .B(n12475), .ZN(n12482) );
  INV_X1 U15692 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16217) );
  XNOR2_X1 U15693 ( .A(n12477), .B(n12478), .ZN(n15619) );
  AND2_X1 U15694 ( .A1(n10382), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12479) );
  NAND2_X1 U15695 ( .A1(n15619), .A2(n12479), .ZN(n16224) );
  AND2_X1 U15696 ( .A1(n9759), .A2(n16224), .ZN(n12498) );
  INV_X1 U15697 ( .A(n12498), .ZN(n12481) );
  NAND2_X1 U15698 ( .A1(n12480), .A2(n10382), .ZN(n12493) );
  AOI21_X1 U15699 ( .B1(n12503), .B2(n12481), .A(n12493), .ZN(n12501) );
  INV_X1 U15700 ( .A(n12482), .ZN(n14685) );
  NAND2_X1 U15701 ( .A1(n14685), .A2(n10382), .ZN(n12483) );
  NAND2_X1 U15702 ( .A1(n12483), .A2(n16217), .ZN(n16215) );
  OAI21_X1 U15703 ( .B1(n16215), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12493), .ZN(n12484) );
  AND2_X1 U15704 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16487) );
  INV_X1 U15705 ( .A(n16487), .ZN(n12485) );
  INV_X1 U15706 ( .A(n12486), .ZN(n12487) );
  NAND2_X1 U15707 ( .A1(n9806), .A2(n12487), .ZN(n12488) );
  NAND2_X1 U15708 ( .A1(n12477), .A2(n12488), .ZN(n15626) );
  OAI21_X1 U15709 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n10382), .ZN(n12489) );
  OAI21_X1 U15710 ( .B1(n15626), .B2(n12489), .A(n14599), .ZN(n12490) );
  INV_X1 U15711 ( .A(n12490), .ZN(n12491) );
  NAND2_X1 U15712 ( .A1(n15619), .A2(n10382), .ZN(n12492) );
  INV_X1 U15713 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16490) );
  NAND2_X1 U15714 ( .A1(n12492), .A2(n16490), .ZN(n16225) );
  INV_X1 U15715 ( .A(n16216), .ZN(n12496) );
  XNOR2_X1 U15716 ( .A(n12493), .B(n12503), .ZN(n12497) );
  INV_X1 U15717 ( .A(n12497), .ZN(n12494) );
  NAND2_X1 U15718 ( .A1(n12496), .A2(n12495), .ZN(n12500) );
  NAND3_X1 U15719 ( .A1(n16216), .A2(n12498), .A3(n12497), .ZN(n12499) );
  NAND2_X1 U15720 ( .A1(n15993), .A2(n17604), .ZN(n12507) );
  NAND2_X1 U15721 ( .A1(n16487), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16485) );
  OAI21_X1 U15722 ( .B1(n17615), .B2(n10417), .A(n16491), .ZN(n16477) );
  AOI21_X1 U15723 ( .B1(n16568), .B2(n16217), .A(n16477), .ZN(n12504) );
  NAND2_X1 U15724 ( .A1(n16754), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14620) );
  NAND4_X1 U15725 ( .A1(n16486), .A2(n10417), .A3(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n12503), .ZN(n12502) );
  OAI211_X1 U15726 ( .C1(n12504), .C2(n12503), .A(n14620), .B(n12502), .ZN(
        n12505) );
  INV_X1 U15727 ( .A(n12505), .ZN(n12506) );
  NAND2_X1 U15728 ( .A1(n16229), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12508) );
  NAND2_X1 U15729 ( .A1(n14618), .A2(n17606), .ZN(n12510) );
  OAI21_X1 U15730 ( .B1(n17599), .B2(n10596), .A(n12511), .ZN(n12513) );
  NOR2_X1 U15731 ( .A1(n16048), .A2(n17589), .ZN(n12512) );
  AOI211_X1 U15732 ( .C1(n17586), .C2(n15719), .A(n12513), .B(n12512), .ZN(
        n12514) );
  OAI21_X1 U15733 ( .B1(n12516), .B2(n16472), .A(n10719), .ZN(P2_U2993) );
  NAND2_X1 U15734 ( .A1(n20135), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12541) );
  NAND2_X1 U15735 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12535) );
  NAND2_X1 U15736 ( .A1(n12535), .A2(n20766), .ZN(n12517) );
  NOR2_X1 U15737 ( .A1(n20766), .A2(n20776), .ZN(n20557) );
  NAND2_X1 U15738 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20557), .ZN(
        n20098) );
  NAND2_X1 U15739 ( .A1(n12517), .A2(n20098), .ZN(n20245) );
  NOR2_X1 U15740 ( .A1(n20245), .A2(n20804), .ZN(n12518) );
  AOI21_X1 U15741 ( .B1(n12537), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12518), .ZN(n12519) );
  NOR2_X1 U15742 ( .A1(n20135), .A2(n20808), .ZN(n12520) );
  INV_X1 U15743 ( .A(n16839), .ZN(n12526) );
  NAND2_X1 U15744 ( .A1(n16787), .A2(n12526), .ZN(n12525) );
  NAND2_X1 U15745 ( .A1(n20776), .A2(n20786), .ZN(n20247) );
  AND2_X1 U15746 ( .A1(n20247), .A2(n12535), .ZN(n20246) );
  AOI21_X1 U15747 ( .B1(n12537), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n20175), .ZN(n12524) );
  NAND2_X1 U15748 ( .A1(n12525), .A2(n12524), .ZN(n13607) );
  AOI22_X1 U15749 ( .A1(n12537), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20749), .B2(n20786), .ZN(n12528) );
  INV_X1 U15750 ( .A(n12530), .ZN(n16780) );
  INV_X1 U15751 ( .A(n12531), .ZN(n12532) );
  NAND2_X1 U15752 ( .A1(n16780), .A2(n12532), .ZN(n12533) );
  INV_X1 U15753 ( .A(n12535), .ZN(n20457) );
  NAND2_X1 U15754 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20758), .ZN(
        n20274) );
  INV_X1 U15755 ( .A(n20274), .ZN(n20276) );
  NAND2_X1 U15756 ( .A1(n20457), .A2(n20276), .ZN(n16859) );
  NAND2_X1 U15757 ( .A1(n20098), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12536) );
  AOI21_X1 U15758 ( .B1(n16859), .B2(n12536), .A(n20804), .ZN(n20486) );
  AOI21_X1 U15759 ( .B1(n12537), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n20486), .ZN(n12538) );
  INV_X1 U15760 ( .A(n12541), .ZN(n12542) );
  NAND2_X1 U15761 ( .A1(n12542), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12543) );
  NAND2_X1 U15762 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14065) );
  NAND2_X1 U15763 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12546) );
  NOR2_X1 U15764 ( .A1(n14065), .A2(n12546), .ZN(n12548) );
  INV_X1 U15765 ( .A(n12547), .ZN(n14218) );
  NAND4_X1 U15766 ( .A1(n13939), .A2(n12548), .A3(n14218), .A4(n14216), .ZN(
        n14028) );
  INV_X1 U15767 ( .A(n12549), .ZN(n14144) );
  NAND3_X1 U15768 ( .A1(n14144), .A2(n14151), .A3(n14032), .ZN(n12550) );
  NOR2_X1 U15769 ( .A1(n14028), .A2(n12550), .ZN(n12551) );
  INV_X1 U15770 ( .A(n12552), .ZN(n16082) );
  AOI22_X1 U15771 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11567), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15772 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15773 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n12625), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12554) );
  AOI22_X1 U15774 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12553) );
  NAND4_X1 U15775 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12562) );
  AOI22_X1 U15776 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n11596), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U15777 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15778 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15779 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n12632), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12557) );
  NAND4_X1 U15780 ( .A1(n12560), .A2(n12559), .A3(n12558), .A4(n12557), .ZN(
        n12561) );
  OR2_X1 U15781 ( .A1(n12562), .A2(n12561), .ZN(n16074) );
  AOI22_X1 U15782 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n11567), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U15783 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15784 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12625), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15785 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11641), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12563) );
  NAND4_X1 U15786 ( .A1(n12566), .A2(n12565), .A3(n12564), .A4(n12563), .ZN(
        n12572) );
  AOI22_X1 U15787 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11573), .B1(
        n11596), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15788 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11630), .B1(
        n12588), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15789 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n11559), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12568) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12632), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12567) );
  NAND4_X1 U15791 ( .A1(n12570), .A2(n12569), .A3(n12568), .A4(n12567), .ZN(
        n12571) );
  OR2_X1 U15792 ( .A1(n12572), .A2(n12571), .ZN(n16067) );
  AOI22_X1 U15793 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12576) );
  AOI22_X1 U15794 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12575) );
  AOI22_X1 U15795 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12574) );
  AOI22_X1 U15796 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12573) );
  NAND4_X1 U15797 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12582) );
  AOI22_X1 U15798 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12580) );
  AOI22_X1 U15799 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12579) );
  AOI22_X1 U15800 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15801 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12577) );
  NAND4_X1 U15802 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12581) );
  NOR2_X1 U15803 ( .A1(n12582), .A2(n12581), .ZN(n16062) );
  AOI22_X1 U15804 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12587) );
  AOI22_X1 U15805 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12586) );
  AOI22_X1 U15806 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12585) );
  AOI22_X1 U15807 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12584) );
  NAND4_X1 U15808 ( .A1(n12587), .A2(n12586), .A3(n12585), .A4(n12584), .ZN(
        n12594) );
  AOI22_X1 U15809 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12592) );
  AOI22_X1 U15810 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15811 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12590) );
  AOI22_X1 U15812 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12589) );
  NAND4_X1 U15813 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n12593) );
  NOR2_X1 U15814 ( .A1(n12594), .A2(n12593), .ZN(n16058) );
  AOI22_X1 U15815 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12598) );
  AOI22_X1 U15816 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15817 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15818 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U15819 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12604) );
  AOI22_X1 U15820 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12602) );
  AOI22_X1 U15821 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12601) );
  AOI22_X1 U15822 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15823 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12599) );
  NAND4_X1 U15824 ( .A1(n12602), .A2(n12601), .A3(n12600), .A4(n12599), .ZN(
        n12603) );
  OR2_X1 U15825 ( .A1(n12604), .A2(n12603), .ZN(n16053) );
  AOI22_X1 U15826 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12608) );
  AOI22_X1 U15827 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12607) );
  AOI22_X1 U15828 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12606) );
  AOI22_X1 U15829 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12605) );
  NAND4_X1 U15830 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        n12614) );
  AOI22_X1 U15831 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12612) );
  AOI22_X1 U15832 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15833 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15834 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12609) );
  NAND4_X1 U15835 ( .A1(n12612), .A2(n12611), .A3(n12610), .A4(n12609), .ZN(
        n12613) );
  OR2_X1 U15836 ( .A1(n12614), .A2(n12613), .ZN(n16047) );
  AOI22_X1 U15837 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11909), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15838 ( .A1(n12583), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15839 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12616) );
  AOI22_X1 U15840 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12615) );
  NAND4_X1 U15841 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12624) );
  AOI22_X1 U15842 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12622) );
  AOI22_X1 U15843 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15844 ( .A1(n11559), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11560), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15845 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12619) );
  NAND4_X1 U15846 ( .A1(n12622), .A2(n12621), .A3(n12620), .A4(n12619), .ZN(
        n12623) );
  NOR2_X1 U15847 ( .A1(n12624), .A2(n12623), .ZN(n16043) );
  AOI22_X1 U15848 ( .A1(n11909), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12583), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12631) );
  AOI22_X1 U15849 ( .A1(n12625), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11637), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12630) );
  AOI22_X1 U15850 ( .A1(n11567), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11568), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12629) );
  AOI22_X1 U15851 ( .A1(n11641), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12628) );
  NAND4_X1 U15852 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        n12638) );
  AOI22_X1 U15853 ( .A1(n11596), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11573), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15854 ( .A1(n12588), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11630), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15855 ( .A1(n11560), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11574), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15856 ( .A1(n12632), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11559), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12633) );
  NAND4_X1 U15857 ( .A1(n12636), .A2(n12635), .A3(n12634), .A4(n12633), .ZN(
        n12637) );
  AOI22_X1 U15858 ( .A1(n12639), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15859 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9739), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12650) );
  INV_X1 U15860 ( .A(n12641), .ZN(n16818) );
  AOI22_X1 U15861 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12649) );
  AND2_X1 U15862 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12643) );
  OR2_X1 U15863 ( .A1(n12643), .A2(n12642), .ZN(n12780) );
  INV_X1 U15864 ( .A(n12780), .ZN(n12753) );
  NAND2_X1 U15865 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12647) );
  INV_X1 U15866 ( .A(n12645), .ZN(n12777) );
  NAND2_X1 U15867 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12646) );
  AND3_X1 U15868 ( .A1(n12753), .A2(n12647), .A3(n12646), .ZN(n12648) );
  NAND4_X1 U15869 ( .A1(n12651), .A2(n12650), .A3(n12649), .A4(n12648), .ZN(
        n12659) );
  AOI22_X1 U15870 ( .A1(n9732), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12657) );
  NAND2_X1 U15871 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12653) );
  NAND2_X1 U15872 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12652) );
  AND3_X1 U15873 ( .A1(n12653), .A2(n12780), .A3(n12652), .ZN(n12656) );
  AOI22_X1 U15874 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12784), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15875 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12654) );
  NAND4_X1 U15876 ( .A1(n12657), .A2(n12656), .A3(n12655), .A4(n12654), .ZN(
        n12658) );
  AND2_X1 U15877 ( .A1(n12659), .A2(n12658), .ZN(n16028) );
  NAND2_X1 U15878 ( .A1(n12676), .A2(n16028), .ZN(n12680) );
  AOI22_X1 U15879 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15880 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U15881 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12661) );
  NAND2_X1 U15882 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12660) );
  AND3_X1 U15883 ( .A1(n12753), .A2(n12661), .A3(n12660), .ZN(n12663) );
  AOI22_X1 U15884 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12662) );
  NAND4_X1 U15885 ( .A1(n12665), .A2(n12664), .A3(n12663), .A4(n12662), .ZN(
        n12674) );
  AOI22_X1 U15886 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15887 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15888 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12670) );
  NAND2_X1 U15889 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12668) );
  NAND2_X1 U15890 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12667) );
  AND3_X1 U15891 ( .A1(n12668), .A2(n12780), .A3(n12667), .ZN(n12669) );
  NAND4_X1 U15892 ( .A1(n12672), .A2(n12671), .A3(n12670), .A4(n12669), .ZN(
        n12673) );
  NAND2_X1 U15893 ( .A1(n12674), .A2(n12673), .ZN(n12679) );
  XNOR2_X1 U15894 ( .A(n12680), .B(n12679), .ZN(n12675) );
  INV_X1 U15895 ( .A(n13939), .ZN(n12714) );
  NOR2_X1 U15896 ( .A1(n12675), .A2(n12714), .ZN(n16032) );
  NAND2_X1 U15897 ( .A1(n16887), .A2(n16028), .ZN(n12677) );
  XNOR2_X1 U15898 ( .A(n12677), .B(n12676), .ZN(n16030) );
  NOR2_X1 U15899 ( .A1(n16887), .A2(n12679), .ZN(n16031) );
  AOI21_X1 U15900 ( .B1(n16026), .B2(n10737), .A(n10736), .ZN(n12678) );
  NOR2_X1 U15901 ( .A1(n12680), .A2(n12679), .ZN(n12695) );
  AOI22_X1 U15902 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15903 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12685) );
  NAND2_X1 U15904 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12682) );
  NAND2_X1 U15905 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12681) );
  AND3_X1 U15906 ( .A1(n12753), .A2(n12682), .A3(n12681), .ZN(n12684) );
  AOI22_X1 U15907 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12683) );
  NAND4_X1 U15908 ( .A1(n12686), .A2(n12685), .A3(n12684), .A4(n12683), .ZN(
        n12694) );
  AOI22_X1 U15909 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15910 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15911 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12690) );
  NAND2_X1 U15912 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U15913 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12687) );
  AND3_X1 U15914 ( .A1(n12688), .A2(n12780), .A3(n12687), .ZN(n12689) );
  NAND4_X1 U15915 ( .A1(n12692), .A2(n12691), .A3(n12690), .A4(n12689), .ZN(
        n12693) );
  AND2_X1 U15916 ( .A1(n12694), .A2(n12693), .ZN(n12697) );
  NAND2_X1 U15917 ( .A1(n12695), .A2(n12697), .ZN(n12717) );
  OAI211_X1 U15918 ( .C1(n12695), .C2(n12697), .A(n13939), .B(n12717), .ZN(
        n12713) );
  NAND2_X1 U15919 ( .A1(n16029), .A2(n12697), .ZN(n16022) );
  AOI22_X1 U15920 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15921 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12702) );
  NAND2_X1 U15922 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12699) );
  NAND2_X1 U15923 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12698) );
  AND3_X1 U15924 ( .A1(n12753), .A2(n12699), .A3(n12698), .ZN(n12701) );
  AOI22_X1 U15925 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15926 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12711) );
  AOI22_X1 U15927 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12709) );
  AOI22_X1 U15928 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12708) );
  AOI22_X1 U15929 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12707) );
  NAND2_X1 U15930 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12705) );
  NAND2_X1 U15931 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12704) );
  AND3_X1 U15932 ( .A1(n12705), .A2(n12780), .A3(n12704), .ZN(n12706) );
  NAND4_X1 U15933 ( .A1(n12709), .A2(n12708), .A3(n12707), .A4(n12706), .ZN(
        n12710) );
  NAND2_X1 U15934 ( .A1(n12711), .A2(n12710), .ZN(n16014) );
  XNOR2_X1 U15935 ( .A(n12717), .B(n16014), .ZN(n12715) );
  NOR2_X1 U15936 ( .A1(n12715), .A2(n12714), .ZN(n16016) );
  NAND2_X1 U15937 ( .A1(n16013), .A2(n16016), .ZN(n12716) );
  OR2_X1 U15938 ( .A1(n12717), .A2(n16014), .ZN(n12732) );
  INV_X1 U15939 ( .A(n12732), .ZN(n12734) );
  AOI22_X1 U15940 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15941 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12722) );
  AOI22_X1 U15942 ( .A1(n16818), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12721) );
  INV_X1 U15943 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n20381) );
  NAND2_X1 U15944 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12719) );
  NAND2_X1 U15945 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12718) );
  AND3_X1 U15946 ( .A1(n12753), .A2(n12719), .A3(n12718), .ZN(n12720) );
  NAND4_X1 U15947 ( .A1(n12723), .A2(n12722), .A3(n12721), .A4(n12720), .ZN(
        n12731) );
  AOI22_X1 U15948 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15949 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12725) );
  NAND2_X1 U15950 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12724) );
  AND3_X1 U15951 ( .A1(n12725), .A2(n12780), .A3(n12724), .ZN(n12728) );
  AOI22_X1 U15952 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15953 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12726) );
  NAND4_X1 U15954 ( .A1(n12729), .A2(n12728), .A3(n12727), .A4(n12726), .ZN(
        n12730) );
  NAND2_X1 U15955 ( .A1(n12731), .A2(n12730), .ZN(n12736) );
  INV_X1 U15956 ( .A(n12736), .ZN(n12733) );
  OAI211_X1 U15957 ( .C1(n12734), .C2(n12733), .A(n12766), .B(n13939), .ZN(
        n12735) );
  NOR2_X1 U15958 ( .A1(n16887), .A2(n12736), .ZN(n16008) );
  AOI22_X1 U15959 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15960 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U15961 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12738) );
  NAND2_X1 U15962 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12737) );
  AND3_X1 U15963 ( .A1(n12753), .A2(n12738), .A3(n12737), .ZN(n12740) );
  AOI22_X1 U15964 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12739) );
  NAND4_X1 U15965 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12750) );
  AOI22_X1 U15966 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12748) );
  AOI22_X1 U15967 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12747) );
  AOI22_X1 U15968 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15969 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12744) );
  NAND2_X1 U15970 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n12743) );
  AND3_X1 U15971 ( .A1(n12744), .A2(n12780), .A3(n12743), .ZN(n12745) );
  NAND4_X1 U15972 ( .A1(n12748), .A2(n12747), .A3(n12746), .A4(n12745), .ZN(
        n12749) );
  NAND2_X1 U15973 ( .A1(n12750), .A2(n12749), .ZN(n16001) );
  AOI22_X1 U15974 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U15975 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12752) );
  NAND2_X1 U15976 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n12751) );
  AND3_X1 U15977 ( .A1(n12753), .A2(n12752), .A3(n12751), .ZN(n12756) );
  AOI22_X1 U15978 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15979 ( .A1(n16818), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12754) );
  NAND4_X1 U15980 ( .A1(n12757), .A2(n12756), .A3(n12755), .A4(n12754), .ZN(
        n12765) );
  AOI22_X1 U15981 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12666), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U15982 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12762) );
  AOI22_X1 U15983 ( .A1(n16818), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U15984 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12759) );
  NAND2_X1 U15985 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12758) );
  AND3_X1 U15986 ( .A1(n12759), .A2(n12780), .A3(n12758), .ZN(n12760) );
  NAND4_X1 U15987 ( .A1(n12763), .A2(n12762), .A3(n12761), .A4(n12760), .ZN(
        n12764) );
  NAND2_X1 U15988 ( .A1(n12765), .A2(n12764), .ZN(n12770) );
  INV_X1 U15989 ( .A(n12766), .ZN(n15999) );
  INV_X1 U15990 ( .A(n16001), .ZN(n12767) );
  AND2_X1 U15991 ( .A1(n16887), .A2(n12767), .ZN(n12768) );
  NAND2_X1 U15992 ( .A1(n15999), .A2(n12768), .ZN(n12769) );
  NOR2_X1 U15993 ( .A1(n12769), .A2(n12770), .ZN(n12771) );
  AOI21_X1 U15994 ( .B1(n12770), .B2(n12769), .A(n12771), .ZN(n15994) );
  AOI22_X1 U15995 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12774) );
  NAND2_X1 U15996 ( .A1(n12781), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12773) );
  NAND2_X1 U15997 ( .A1(n12777), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12772) );
  NAND4_X1 U15998 ( .A1(n12774), .A2(n12773), .A3(n12772), .A4(n12780), .ZN(
        n12792) );
  AOI22_X1 U15999 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12783), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U16000 ( .A1(n12782), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12775) );
  NAND2_X1 U16001 ( .A1(n12776), .A2(n12775), .ZN(n12791) );
  NOR2_X1 U16002 ( .A1(n12645), .A2(n12778), .ZN(n12779) );
  AOI211_X1 U16003 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n12781), .A(
        n12780), .B(n12779), .ZN(n12789) );
  AOI22_X1 U16004 ( .A1(n12783), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12782), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16005 ( .A1(n12666), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9743), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16006 ( .A1(n12785), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16818), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12786) );
  NAND4_X1 U16007 ( .A1(n12789), .A2(n12788), .A3(n12787), .A4(n12786), .ZN(
        n12790) );
  OAI21_X1 U16008 ( .B1(n12792), .B2(n12791), .A(n12790), .ZN(n12793) );
  INV_X1 U16009 ( .A(n12793), .ZN(n12794) );
  XNOR2_X1 U16010 ( .A(n12795), .B(n12794), .ZN(n14719) );
  INV_X1 U16011 ( .A(n16894), .ZN(n12796) );
  OAI21_X1 U16012 ( .B1(n14719), .B2(n16072), .A(n12800), .ZN(P2_U2857) );
  NOR3_X1 U16013 ( .A1(n10154), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16014 ( .A1(n13629), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11242), .ZN(n12808) );
  NAND2_X1 U16015 ( .A1(n15056), .A2(n20998), .ZN(n12818) );
  NOR2_X1 U16016 ( .A1(n12811), .A2(n21867), .ZN(n12815) );
  INV_X1 U16017 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21548) );
  NOR2_X1 U16018 ( .A1(n20904), .A2(n21548), .ZN(n15162) );
  NOR3_X1 U16019 ( .A1(n12813), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12812), .ZN(n12814) );
  AOI211_X1 U16020 ( .C1(n12816), .C2(n12815), .A(n15162), .B(n12814), .ZN(
        n12817) );
  OAI211_X1 U16021 ( .C1(n15168), .C2(n17559), .A(n12818), .B(n12817), .ZN(
        P1_U3000) );
  NAND2_X1 U16022 ( .A1(n10254), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12855) );
  OAI21_X1 U16023 ( .B1(n21173), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n21578), .ZN(n12821) );
  NAND2_X1 U16024 ( .A1(n13339), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12820) );
  OAI211_X1 U16025 ( .C1(n12855), .C2(n17569), .A(n12821), .B(n12820), .ZN(
        n12824) );
  NOR2_X1 U16026 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12851), .ZN(
        n12822) );
  NOR2_X1 U16027 ( .A1(n12861), .A2(n12822), .ZN(n14205) );
  NAND2_X1 U16028 ( .A1(n14205), .A2(n14232), .ZN(n12823) );
  NAND2_X1 U16029 ( .A1(n12824), .A2(n12823), .ZN(n12825) );
  NAND2_X1 U16030 ( .A1(n12826), .A2(n12993), .ZN(n12830) );
  XNOR2_X1 U16031 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15041) );
  AOI22_X1 U16032 ( .A1(n13339), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n14232), .B2(
        n15041), .ZN(n12829) );
  NAND2_X1 U16033 ( .A1(n12827), .A2(n15602), .ZN(n12828) );
  NAND2_X1 U16034 ( .A1(n12830), .A2(n10718), .ZN(n13933) );
  NAND2_X1 U16035 ( .A1(n21578), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13932) );
  OR2_X1 U16036 ( .A1(n13933), .A2(n13346), .ZN(n12860) );
  XNOR2_X2 U16037 ( .A(n12834), .B(n12833), .ZN(n14113) );
  NAND2_X1 U16038 ( .A1(n14113), .A2(n12993), .ZN(n12838) );
  AOI22_X1 U16039 ( .A1(n13339), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21578), .ZN(n12836) );
  NAND2_X1 U16040 ( .A1(n12827), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12835) );
  AND2_X1 U16041 ( .A1(n12836), .A2(n12835), .ZN(n12837) );
  NAND2_X1 U16042 ( .A1(n12838), .A2(n12837), .ZN(n13643) );
  NAND2_X1 U16043 ( .A1(n14375), .A2(n12819), .ZN(n12841) );
  NAND2_X1 U16044 ( .A1(n12841), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13615) );
  OR2_X1 U16045 ( .A1(n14590), .A2(n13014), .ZN(n12846) );
  AOI22_X1 U16046 ( .A1(n12842), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21578), .ZN(n12844) );
  NAND2_X1 U16047 ( .A1(n12827), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12843) );
  AND2_X1 U16048 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NAND2_X1 U16049 ( .A1(n13616), .A2(n14232), .ZN(n12847) );
  NAND2_X1 U16050 ( .A1(n13617), .A2(n12847), .ZN(n13642) );
  NAND2_X1 U16051 ( .A1(n13643), .A2(n13642), .ZN(n13641) );
  NAND2_X1 U16052 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14097) );
  NAND2_X1 U16053 ( .A1(n13641), .A2(n14097), .ZN(n12859) );
  AND2_X1 U16054 ( .A1(n12848), .A2(n12993), .ZN(n12849) );
  NAND2_X1 U16055 ( .A1(n12850), .A2(n12849), .ZN(n12858) );
  AOI21_X1 U16056 ( .B1(n14264), .B2(n12852), .A(n12851), .ZN(n20920) );
  OAI22_X1 U16057 ( .A1(n20920), .A2(n9867), .B1(n13932), .B2(n14264), .ZN(
        n12853) );
  AOI21_X1 U16058 ( .B1(n13339), .B2(P1_EAX_REG_3__SCAN_IN), .A(n12853), .ZN(
        n12854) );
  OAI21_X1 U16059 ( .B1(n14004), .B2(n12855), .A(n12854), .ZN(n12856) );
  INV_X1 U16060 ( .A(n12856), .ZN(n12857) );
  INV_X1 U16061 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21775) );
  INV_X1 U16062 ( .A(n12870), .ZN(n12872) );
  INV_X1 U16063 ( .A(n12861), .ZN(n12862) );
  NAND2_X1 U16064 ( .A1(n12862), .A2(n21775), .ZN(n12863) );
  NAND2_X1 U16065 ( .A1(n12872), .A2(n12863), .ZN(n20891) );
  NAND2_X1 U16066 ( .A1(n20891), .A2(n14232), .ZN(n12864) );
  OAI21_X1 U16067 ( .B1(n13932), .B2(n21775), .A(n12864), .ZN(n12865) );
  AOI21_X1 U16068 ( .B1(n13339), .B2(P1_EAX_REG_5__SCAN_IN), .A(n12865), .ZN(
        n12866) );
  INV_X1 U16069 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12876) );
  INV_X1 U16070 ( .A(n12868), .ZN(n12869) );
  NAND2_X1 U16071 ( .A1(n12869), .A2(n12993), .ZN(n12875) );
  INV_X1 U16072 ( .A(n12877), .ZN(n12878) );
  INV_X1 U16073 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12871) );
  NAND2_X1 U16074 ( .A1(n12872), .A2(n12871), .ZN(n12873) );
  NAND2_X1 U16075 ( .A1(n12878), .A2(n12873), .ZN(n20873) );
  INV_X2 U16076 ( .A(n9867), .ZN(n14232) );
  AOI22_X1 U16077 ( .A1(n20873), .A2(n14232), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13346), .ZN(n12874) );
  INV_X1 U16078 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12881) );
  INV_X1 U16079 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20862) );
  NAND2_X1 U16080 ( .A1(n12878), .A2(n20862), .ZN(n12879) );
  NAND2_X1 U16081 ( .A1(n12909), .A2(n12879), .ZN(n20863) );
  AOI22_X1 U16082 ( .A1(n20863), .A2(n14232), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n13346), .ZN(n12880) );
  OAI21_X1 U16083 ( .B1(n13047), .B2(n12881), .A(n12880), .ZN(n12882) );
  AOI21_X1 U16084 ( .B1(n12883), .B2(n12993), .A(n12882), .ZN(n14362) );
  AOI22_X1 U16085 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12887) );
  AOI22_X1 U16086 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12886) );
  AOI22_X1 U16087 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n9718), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U16088 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13328), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12884) );
  NAND4_X1 U16089 ( .A1(n12887), .A2(n12886), .A3(n12885), .A4(n12884), .ZN(
        n12893) );
  AOI22_X1 U16090 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n13320), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U16091 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13187), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16092 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13285), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16093 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12888) );
  NAND4_X1 U16094 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12892) );
  OAI21_X1 U16095 ( .B1(n12893), .B2(n12892), .A(n12993), .ZN(n12898) );
  NAND2_X1 U16096 ( .A1(n13339), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12897) );
  INV_X1 U16097 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12894) );
  XNOR2_X1 U16098 ( .A(n12909), .B(n12894), .ZN(n15029) );
  NAND2_X1 U16099 ( .A1(n15029), .A2(n14232), .ZN(n12896) );
  NAND2_X1 U16100 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12895) );
  AOI22_X1 U16101 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16102 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16103 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16104 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12899) );
  NAND4_X1 U16105 ( .A1(n12902), .A2(n12901), .A3(n12900), .A4(n12899), .ZN(
        n12908) );
  AOI22_X1 U16106 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10919), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16107 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16108 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10773), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U16109 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12903) );
  NAND4_X1 U16110 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n12907) );
  OAI21_X1 U16111 ( .B1(n12908), .B2(n12907), .A(n12993), .ZN(n12914) );
  NAND2_X1 U16112 ( .A1(n13339), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U16113 ( .A1(n12926), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12910) );
  INV_X1 U16114 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20847) );
  XNOR2_X1 U16115 ( .A(n12910), .B(n20847), .ZN(n20850) );
  NAND2_X1 U16116 ( .A1(n20850), .A2(n14232), .ZN(n12912) );
  NAND2_X1 U16117 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12911) );
  NAND4_X1 U16118 ( .A1(n12914), .A2(n12913), .A3(n12912), .A4(n12911), .ZN(
        n14403) );
  AOI22_X1 U16119 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16120 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16121 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16122 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12915) );
  NAND4_X1 U16123 ( .A1(n12918), .A2(n12917), .A3(n12916), .A4(n12915), .ZN(
        n12924) );
  AOI22_X1 U16124 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U16125 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13995), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16126 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16127 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12919) );
  NAND4_X1 U16128 ( .A1(n12922), .A2(n12921), .A3(n12920), .A4(n12919), .ZN(
        n12923) );
  OAI21_X1 U16129 ( .B1(n12924), .B2(n12923), .A(n12993), .ZN(n12931) );
  NAND2_X1 U16130 ( .A1(n13339), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12930) );
  INV_X1 U16131 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12927) );
  XNOR2_X1 U16132 ( .A(n12932), .B(n12927), .ZN(n15359) );
  NAND2_X1 U16133 ( .A1(n15359), .A2(n14232), .ZN(n12929) );
  NAND2_X1 U16134 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12928) );
  NAND2_X1 U16135 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12934) );
  INV_X1 U16136 ( .A(n12950), .ZN(n12935) );
  INV_X1 U16137 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n14951) );
  XNOR2_X1 U16138 ( .A(n12935), .B(n14951), .ZN(n15319) );
  AOI22_X1 U16139 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13320), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16140 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U16141 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12937) );
  AOI22_X1 U16142 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12936) );
  NAND4_X1 U16143 ( .A1(n12939), .A2(n12938), .A3(n12937), .A4(n12936), .ZN(
        n12945) );
  AOI22_X1 U16144 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16145 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16146 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16147 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12940) );
  NAND4_X1 U16148 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12944) );
  OAI21_X1 U16149 ( .B1(n12945), .B2(n12944), .A(n12993), .ZN(n12948) );
  NAND2_X1 U16150 ( .A1(n13339), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12947) );
  NAND2_X1 U16151 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12946) );
  NAND3_X1 U16152 ( .A1(n12948), .A2(n12947), .A3(n12946), .ZN(n12949) );
  AOI21_X1 U16153 ( .B1(n15319), .B2(n14232), .A(n12949), .ZN(n14947) );
  INV_X1 U16154 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12951) );
  XNOR2_X1 U16155 ( .A(n13017), .B(n12951), .ZN(n15308) );
  AOI22_X1 U16156 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U16157 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16158 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U16159 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12952) );
  NAND4_X1 U16160 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        n12961) );
  AOI22_X1 U16161 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12959) );
  AOI22_X1 U16162 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U16163 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16164 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12956) );
  NAND4_X1 U16165 ( .A1(n12959), .A2(n12958), .A3(n12957), .A4(n12956), .ZN(
        n12960) );
  OAI21_X1 U16166 ( .B1(n12961), .B2(n12960), .A(n12993), .ZN(n12964) );
  NAND2_X1 U16167 ( .A1(n13339), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12963) );
  NAND2_X1 U16168 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12962) );
  NAND3_X1 U16169 ( .A1(n12964), .A2(n12963), .A3(n12962), .ZN(n12965) );
  AOI21_X1 U16170 ( .B1(n15308), .B2(n14232), .A(n12965), .ZN(n14936) );
  AOI22_X1 U16171 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U16172 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16173 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U16174 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U16175 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12975) );
  AOI22_X1 U16176 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16177 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13291), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16178 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16179 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12970) );
  NAND4_X1 U16180 ( .A1(n12973), .A2(n12972), .A3(n12971), .A4(n12970), .ZN(
        n12974) );
  OR2_X1 U16181 ( .A1(n12975), .A2(n12974), .ZN(n12976) );
  AND2_X1 U16182 ( .A1(n12993), .A2(n12976), .ZN(n14961) );
  NAND2_X1 U16183 ( .A1(n13339), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12980) );
  NAND2_X1 U16184 ( .A1(n12977), .A2(n12981), .ZN(n12978) );
  NAND2_X1 U16185 ( .A1(n13011), .A2(n12978), .ZN(n15347) );
  NAND2_X1 U16186 ( .A1(n15347), .A2(n14232), .ZN(n12979) );
  OAI211_X1 U16187 ( .C1(n13932), .C2(n12981), .A(n12980), .B(n12979), .ZN(
        n14935) );
  INV_X1 U16188 ( .A(n13011), .ZN(n12982) );
  NAND2_X1 U16189 ( .A1(n12982), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12984) );
  INV_X1 U16190 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12983) );
  XNOR2_X1 U16191 ( .A(n12984), .B(n12983), .ZN(n15330) );
  NAND2_X1 U16192 ( .A1(n15330), .A2(n14232), .ZN(n12999) );
  AOI22_X1 U16193 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13291), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16194 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16195 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16196 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12985) );
  NAND4_X1 U16197 ( .A1(n12988), .A2(n12987), .A3(n12986), .A4(n12985), .ZN(
        n12995) );
  AOI22_X1 U16198 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16199 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13995), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16200 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12990) );
  AOI22_X1 U16201 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12989) );
  NAND4_X1 U16202 ( .A1(n12992), .A2(n12991), .A3(n12990), .A4(n12989), .ZN(
        n12994) );
  OAI21_X1 U16203 ( .B1(n12995), .B2(n12994), .A(n12993), .ZN(n12998) );
  NAND2_X1 U16204 ( .A1(n13339), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12997) );
  NAND2_X1 U16205 ( .A1(n13346), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12996) );
  NAND2_X1 U16206 ( .A1(n12999), .A2(n10727), .ZN(n14964) );
  AOI22_X1 U16207 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10919), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U16208 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U16209 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U16210 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13000) );
  NAND4_X1 U16211 ( .A1(n13003), .A2(n13002), .A3(n13001), .A4(n13000), .ZN(
        n13009) );
  AOI22_X1 U16212 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16213 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16214 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13005) );
  AOI22_X1 U16215 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13004) );
  NAND4_X1 U16216 ( .A1(n13007), .A2(n13006), .A3(n13005), .A4(n13004), .ZN(
        n13008) );
  NOR2_X1 U16217 ( .A1(n13009), .A2(n13008), .ZN(n13015) );
  INV_X1 U16218 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n13010) );
  XNOR2_X1 U16219 ( .A(n13011), .B(n13010), .ZN(n15336) );
  NAND2_X1 U16220 ( .A1(n15336), .A2(n14232), .ZN(n13013) );
  AOI22_X1 U16221 ( .A1(n13339), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13346), .ZN(n13012) );
  OAI211_X1 U16222 ( .C1(n13015), .C2(n13014), .A(n13013), .B(n13012), .ZN(
        n14962) );
  OAI211_X1 U16223 ( .C1(n14961), .C2(n14935), .A(n14964), .B(n14962), .ZN(
        n13016) );
  NAND2_X1 U16224 ( .A1(n13019), .A2(n15295), .ZN(n13020) );
  AND2_X1 U16225 ( .A1(n13052), .A2(n13020), .ZN(n15297) );
  AOI22_X1 U16226 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13320), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U16227 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n13319), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13023) );
  AOI22_X1 U16228 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13022) );
  AOI22_X1 U16229 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13021) );
  NAND4_X1 U16230 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13021), .ZN(
        n13030) );
  AOI22_X1 U16231 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13995), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13028) );
  AOI22_X1 U16232 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n13293), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13027) );
  AOI22_X1 U16233 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n13138), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13026) );
  AOI22_X1 U16234 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13025) );
  NAND4_X1 U16235 ( .A1(n13028), .A2(n13027), .A3(n13026), .A4(n13025), .ZN(
        n13029) );
  OR2_X1 U16236 ( .A1(n13030), .A2(n13029), .ZN(n13033) );
  INV_X1 U16237 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15137) );
  OAI21_X1 U16238 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n21173), .A(
        n21578), .ZN(n13031) );
  OAI21_X1 U16239 ( .B1(n13047), .B2(n15137), .A(n13031), .ZN(n13032) );
  AOI21_X1 U16240 ( .B1(n13300), .B2(n13033), .A(n13032), .ZN(n13034) );
  AOI21_X1 U16241 ( .B1(n15297), .B2(n14232), .A(n13034), .ZN(n14917) );
  XNOR2_X1 U16242 ( .A(n13052), .B(n14907), .ZN(n15287) );
  NAND2_X1 U16243 ( .A1(n15287), .A2(n14232), .ZN(n13051) );
  AOI22_X1 U16244 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13039) );
  AOI22_X1 U16245 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13038) );
  AOI22_X1 U16246 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U16247 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13036) );
  NAND4_X1 U16248 ( .A1(n13039), .A2(n13038), .A3(n13037), .A4(n13036), .ZN(
        n13046) );
  AOI22_X1 U16249 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13044) );
  AOI22_X1 U16250 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10773), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13043) );
  AOI22_X1 U16251 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13042) );
  AOI22_X1 U16252 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13040), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13041) );
  NAND4_X1 U16253 ( .A1(n13044), .A2(n13043), .A3(n13042), .A4(n13041), .ZN(
        n13045) );
  OR2_X1 U16254 ( .A1(n13046), .A2(n13045), .ZN(n13049) );
  INV_X1 U16255 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15132) );
  OAI22_X1 U16256 ( .A1(n13047), .A2(n15132), .B1(n14907), .B2(n13932), .ZN(
        n13048) );
  AOI21_X1 U16257 ( .B1(n13300), .B2(n13049), .A(n13048), .ZN(n13050) );
  NAND2_X1 U16258 ( .A1(n13051), .A2(n13050), .ZN(n14904) );
  INV_X1 U16259 ( .A(n13053), .ZN(n13055) );
  INV_X1 U16260 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U16261 ( .A1(n13055), .A2(n13054), .ZN(n13056) );
  NAND2_X1 U16262 ( .A1(n13090), .A2(n13056), .ZN(n15271) );
  AOI22_X1 U16263 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13060) );
  AOI22_X1 U16264 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13059) );
  AOI22_X1 U16265 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13058) );
  AOI22_X1 U16266 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13057) );
  NAND4_X1 U16267 ( .A1(n13060), .A2(n13059), .A3(n13058), .A4(n13057), .ZN(
        n13066) );
  AOI22_X1 U16268 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13995), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13064) );
  AOI22_X1 U16269 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13063) );
  AOI22_X1 U16270 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13062) );
  AOI22_X1 U16271 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13061) );
  NAND4_X1 U16272 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        n13065) );
  NOR2_X1 U16273 ( .A1(n13066), .A2(n13065), .ZN(n13070) );
  NAND2_X1 U16274 ( .A1(n21578), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13067) );
  NAND2_X1 U16275 ( .A1(n9867), .A2(n13067), .ZN(n13068) );
  AOI21_X1 U16276 ( .B1(n13339), .B2(P1_EAX_REG_18__SCAN_IN), .A(n13068), .ZN(
        n13069) );
  OAI21_X1 U16277 ( .B1(n13342), .B2(n13070), .A(n13069), .ZN(n13071) );
  XNOR2_X1 U16278 ( .A(n13090), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15265) );
  NAND2_X1 U16279 ( .A1(n15265), .A2(n14232), .ZN(n13088) );
  AOI22_X1 U16280 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13320), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16281 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13075) );
  AOI22_X1 U16282 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13074) );
  AOI22_X1 U16283 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13073) );
  NAND4_X1 U16284 ( .A1(n13076), .A2(n13075), .A3(n13074), .A4(n13073), .ZN(
        n13082) );
  AOI22_X1 U16285 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U16286 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13079) );
  AOI22_X1 U16287 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13078) );
  AOI22_X1 U16288 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13077) );
  NAND4_X1 U16289 ( .A1(n13080), .A2(n13079), .A3(n13078), .A4(n13077), .ZN(
        n13081) );
  NOR2_X1 U16290 ( .A1(n13082), .A2(n13081), .ZN(n13086) );
  NAND2_X1 U16291 ( .A1(n21578), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13083) );
  NAND2_X1 U16292 ( .A1(n9867), .A2(n13083), .ZN(n13084) );
  AOI21_X1 U16293 ( .B1(n13339), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13084), .ZN(
        n13085) );
  OAI21_X1 U16294 ( .B1(n13342), .B2(n13086), .A(n13085), .ZN(n13087) );
  NAND2_X1 U16295 ( .A1(n13088), .A2(n13087), .ZN(n14876) );
  AND2_X2 U16296 ( .A1(n13091), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13092) );
  INV_X1 U16297 ( .A(n13092), .ZN(n13094) );
  INV_X1 U16298 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U16299 ( .A1(n13094), .A2(n13093), .ZN(n13095) );
  NAND2_X1 U16300 ( .A1(n13126), .A2(n13095), .ZN(n15254) );
  AOI22_X1 U16301 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U16302 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16303 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13097) );
  AOI22_X1 U16304 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13096) );
  NAND4_X1 U16305 ( .A1(n13099), .A2(n13098), .A3(n13097), .A4(n13096), .ZN(
        n13105) );
  AOI22_X1 U16306 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13995), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U16307 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13102) );
  AOI22_X1 U16308 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U16309 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13100) );
  NAND4_X1 U16310 ( .A1(n13103), .A2(n13102), .A3(n13101), .A4(n13100), .ZN(
        n13104) );
  NOR2_X1 U16311 ( .A1(n13105), .A2(n13104), .ZN(n13109) );
  NAND2_X1 U16312 ( .A1(n21578), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13106) );
  NAND2_X1 U16313 ( .A1(n9867), .A2(n13106), .ZN(n13107) );
  AOI21_X1 U16314 ( .B1(n13339), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13107), .ZN(
        n13108) );
  OAI21_X1 U16315 ( .B1(n13342), .B2(n13109), .A(n13108), .ZN(n13110) );
  XNOR2_X1 U16316 ( .A(n13126), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15247) );
  INV_X1 U16317 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15249) );
  AOI21_X1 U16318 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15249), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13113) );
  AOI21_X1 U16319 ( .B1(n13339), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13113), .ZN(
        n13125) );
  AOI22_X1 U16320 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13117) );
  AOI22_X1 U16321 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13293), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16322 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U16323 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13114) );
  NAND4_X1 U16324 ( .A1(n13117), .A2(n13116), .A3(n13115), .A4(n13114), .ZN(
        n13123) );
  AOI22_X1 U16325 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16326 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U16327 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U16328 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13118) );
  NAND4_X1 U16329 ( .A1(n13121), .A2(n13120), .A3(n13119), .A4(n13118), .ZN(
        n13122) );
  OAI21_X1 U16330 ( .B1(n13123), .B2(n13122), .A(n13300), .ZN(n13124) );
  AOI22_X1 U16331 ( .A1(n15247), .A2(n14232), .B1(n13125), .B2(n13124), .ZN(
        n14854) );
  INV_X1 U16332 ( .A(n13128), .ZN(n13130) );
  INV_X1 U16333 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16334 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  NAND2_X1 U16335 ( .A1(n13179), .A2(n13131), .ZN(n15237) );
  AOI22_X1 U16336 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16337 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13293), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16338 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16339 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U16340 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13144) );
  AOI22_X1 U16341 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13142) );
  AOI22_X1 U16342 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U16343 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U16344 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13139) );
  NAND4_X1 U16345 ( .A1(n13142), .A2(n13141), .A3(n13140), .A4(n13139), .ZN(
        n13143) );
  NOR2_X1 U16346 ( .A1(n13144), .A2(n13143), .ZN(n13148) );
  NAND2_X1 U16347 ( .A1(n21578), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13145) );
  NAND2_X1 U16348 ( .A1(n9867), .A2(n13145), .ZN(n13146) );
  AOI21_X1 U16349 ( .B1(n13339), .B2(P1_EAX_REG_22__SCAN_IN), .A(n13146), .ZN(
        n13147) );
  OAI21_X1 U16350 ( .B1(n13342), .B2(n13148), .A(n13147), .ZN(n13149) );
  NAND2_X1 U16351 ( .A1(n13150), .A2(n13149), .ZN(n14834) );
  XNOR2_X1 U16352 ( .A(n13179), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15227) );
  NAND2_X1 U16353 ( .A1(n15227), .A2(n14232), .ZN(n13178) );
  AOI22_X1 U16354 ( .A1(n13132), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13154) );
  AOI22_X1 U16355 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13138), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16356 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U16357 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13151) );
  NAND4_X1 U16358 ( .A1(n13154), .A2(n13153), .A3(n13152), .A4(n13151), .ZN(
        n13160) );
  AOI22_X1 U16359 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13158) );
  AOI22_X1 U16360 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13157) );
  AOI22_X1 U16361 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16362 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13155) );
  NAND4_X1 U16363 ( .A1(n13158), .A2(n13157), .A3(n13156), .A4(n13155), .ZN(
        n13159) );
  NOR2_X1 U16364 ( .A1(n13160), .A2(n13159), .ZN(n13184) );
  AOI22_X1 U16365 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13164) );
  AOI22_X1 U16366 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16367 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13162) );
  AOI22_X1 U16368 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13161) );
  NAND4_X1 U16369 ( .A1(n13164), .A2(n13163), .A3(n13162), .A4(n13161), .ZN(
        n13171) );
  AOI22_X1 U16370 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U16371 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n13320), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16372 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n13165), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U16373 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13166) );
  NAND4_X1 U16374 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13170) );
  NOR2_X1 U16375 ( .A1(n13171), .A2(n13170), .ZN(n13185) );
  XOR2_X1 U16376 ( .A(n13184), .B(n13185), .Z(n13172) );
  NAND2_X1 U16377 ( .A1(n13172), .A2(n13300), .ZN(n13176) );
  NAND2_X1 U16378 ( .A1(n21578), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13173) );
  NAND2_X1 U16379 ( .A1(n9867), .A2(n13173), .ZN(n13174) );
  AOI21_X1 U16380 ( .B1(n13339), .B2(P1_EAX_REG_23__SCAN_IN), .A(n13174), .ZN(
        n13175) );
  NAND2_X1 U16381 ( .A1(n13176), .A2(n13175), .ZN(n13177) );
  NAND2_X1 U16382 ( .A1(n13178), .A2(n13177), .ZN(n14824) );
  AND2_X2 U16383 ( .A1(n13180), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13181) );
  INV_X1 U16384 ( .A(n13181), .ZN(n13182) );
  INV_X1 U16385 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16386 ( .A1(n13182), .A2(n13198), .ZN(n13183) );
  NAND2_X1 U16387 ( .A1(n13221), .A2(n13183), .ZN(n15222) );
  NOR2_X1 U16388 ( .A1(n13185), .A2(n13184), .ZN(n13206) );
  AOI22_X1 U16389 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13211), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13191) );
  AOI22_X1 U16390 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13190) );
  AOI22_X1 U16391 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13189) );
  AOI22_X1 U16392 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13188) );
  NAND4_X1 U16393 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13197) );
  AOI22_X1 U16394 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13195) );
  AOI22_X1 U16395 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13194) );
  AOI22_X1 U16396 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13193) );
  AOI22_X1 U16397 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13192) );
  NAND4_X1 U16398 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13196) );
  OR2_X1 U16399 ( .A1(n13197), .A2(n13196), .ZN(n13205) );
  XNOR2_X1 U16400 ( .A(n13206), .B(n13205), .ZN(n13201) );
  AOI21_X1 U16401 ( .B1(n13198), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13199) );
  AOI21_X1 U16402 ( .B1(n13339), .B2(P1_EAX_REG_24__SCAN_IN), .A(n13199), .ZN(
        n13200) );
  OAI21_X1 U16403 ( .B1(n13201), .B2(n13342), .A(n13200), .ZN(n13202) );
  XNOR2_X1 U16404 ( .A(n13221), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15208) );
  INV_X1 U16405 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15206) );
  NOR2_X1 U16406 ( .A1(n15206), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13204) );
  AOI211_X1 U16407 ( .C1(n13339), .C2(P1_EAX_REG_25__SCAN_IN), .A(n14232), .B(
        n13204), .ZN(n13220) );
  NAND2_X1 U16408 ( .A1(n13206), .A2(n13205), .ZN(n13227) );
  AOI22_X1 U16409 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13293), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U16410 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U16411 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13208) );
  AOI22_X1 U16412 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13207) );
  NAND4_X1 U16413 ( .A1(n13210), .A2(n13209), .A3(n13208), .A4(n13207), .ZN(
        n13217) );
  AOI22_X1 U16414 ( .A1(n13211), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13215) );
  AOI22_X1 U16415 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13214) );
  AOI22_X1 U16416 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13213) );
  AOI22_X1 U16417 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13212) );
  NAND4_X1 U16418 ( .A1(n13215), .A2(n13214), .A3(n13213), .A4(n13212), .ZN(
        n13216) );
  NOR2_X1 U16419 ( .A1(n13217), .A2(n13216), .ZN(n13228) );
  XOR2_X1 U16420 ( .A(n13227), .B(n13228), .Z(n13218) );
  NAND2_X1 U16421 ( .A1(n13218), .A2(n13300), .ZN(n13219) );
  AOI22_X1 U16422 ( .A1(n15208), .A2(n14232), .B1(n13220), .B2(n13219), .ZN(
        n14796) );
  AND2_X2 U16423 ( .A1(n13222), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13223) );
  INV_X1 U16424 ( .A(n13223), .ZN(n13225) );
  INV_X1 U16425 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13224) );
  NAND2_X1 U16426 ( .A1(n13225), .A2(n13224), .ZN(n13226) );
  NAND2_X1 U16427 ( .A1(n13259), .A2(n13226), .ZN(n15202) );
  NOR2_X1 U16428 ( .A1(n13228), .A2(n13227), .ZN(n13245) );
  AOI22_X1 U16429 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13232) );
  INV_X1 U16430 ( .A(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n21726) );
  AOI22_X1 U16431 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13231) );
  AOI22_X1 U16432 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13230) );
  AOI22_X1 U16433 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13229) );
  NAND4_X1 U16434 ( .A1(n13232), .A2(n13231), .A3(n13230), .A4(n13229), .ZN(
        n13238) );
  AOI22_X1 U16435 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13236) );
  AOI22_X1 U16436 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13235) );
  AOI22_X1 U16437 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13234) );
  AOI22_X1 U16438 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13233) );
  NAND4_X1 U16439 ( .A1(n13236), .A2(n13235), .A3(n13234), .A4(n13233), .ZN(
        n13237) );
  OR2_X1 U16440 ( .A1(n13238), .A2(n13237), .ZN(n13244) );
  XNOR2_X1 U16441 ( .A(n13245), .B(n13244), .ZN(n13241) );
  AOI21_X1 U16442 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21578), .A(
        n14232), .ZN(n13240) );
  NAND2_X1 U16443 ( .A1(n13339), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13239) );
  OAI211_X1 U16444 ( .C1(n13241), .C2(n13342), .A(n13240), .B(n13239), .ZN(
        n13242) );
  XNOR2_X1 U16445 ( .A(n13259), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15189) );
  INV_X1 U16446 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15187) );
  AOI21_X1 U16447 ( .B1(n15187), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13243) );
  AOI21_X1 U16448 ( .B1(n13339), .B2(P1_EAX_REG_27__SCAN_IN), .A(n13243), .ZN(
        n13258) );
  NAND2_X1 U16449 ( .A1(n13245), .A2(n13244), .ZN(n13263) );
  AOI22_X1 U16450 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U16451 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U16452 ( .A1(n13138), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U16453 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13246) );
  NAND4_X1 U16454 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        n13255) );
  AOI22_X1 U16455 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13320), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13253) );
  AOI22_X1 U16456 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13252) );
  AOI22_X1 U16457 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10773), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13251) );
  AOI22_X1 U16458 ( .A1(n13186), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13250) );
  NAND4_X1 U16459 ( .A1(n13253), .A2(n13252), .A3(n13251), .A4(n13250), .ZN(
        n13254) );
  NOR2_X1 U16460 ( .A1(n13255), .A2(n13254), .ZN(n13264) );
  XOR2_X1 U16461 ( .A(n13263), .B(n13264), .Z(n13256) );
  NAND2_X1 U16462 ( .A1(n13256), .A2(n13300), .ZN(n13257) );
  AOI22_X1 U16463 ( .A1(n15189), .A2(n14232), .B1(n13258), .B2(n13257), .ZN(
        n14770) );
  OR2_X2 U16464 ( .A1(n13259), .A2(n15187), .ZN(n13261) );
  INV_X1 U16465 ( .A(n13261), .ZN(n13262) );
  INV_X1 U16466 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13260) );
  OR2_X2 U16467 ( .A1(n13261), .A2(n13260), .ZN(n13280) );
  OAI21_X1 U16468 ( .B1(n13262), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n13280), .ZN(n15183) );
  NOR2_X1 U16469 ( .A1(n13264), .A2(n13263), .ZN(n13283) );
  AOI22_X1 U16470 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13268) );
  AOI22_X1 U16471 ( .A1(n13319), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13267) );
  AOI22_X1 U16472 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13266) );
  AOI22_X1 U16473 ( .A1(n10919), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13265) );
  NAND4_X1 U16474 ( .A1(n13268), .A2(n13267), .A3(n13266), .A4(n13265), .ZN(
        n13275) );
  AOI22_X1 U16475 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9718), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13273) );
  AOI22_X1 U16476 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13272) );
  AOI22_X1 U16477 ( .A1(n10773), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13271) );
  AOI22_X1 U16478 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13270) );
  NAND4_X1 U16479 ( .A1(n13273), .A2(n13272), .A3(n13271), .A4(n13270), .ZN(
        n13274) );
  OR2_X1 U16480 ( .A1(n13275), .A2(n13274), .ZN(n13282) );
  XNOR2_X1 U16481 ( .A(n13283), .B(n13282), .ZN(n13278) );
  AOI21_X1 U16482 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21578), .A(
        n14232), .ZN(n13277) );
  NAND2_X1 U16483 ( .A1(n12842), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13276) );
  OAI211_X1 U16484 ( .C1(n13278), .C2(n13342), .A(n13277), .B(n13276), .ZN(
        n13279) );
  OAI21_X1 U16485 ( .B1(n15183), .B2(n9867), .A(n13279), .ZN(n14758) );
  XOR2_X1 U16486 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B(n13318), .Z(
        n14727) );
  INV_X1 U16487 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13315) );
  NOR2_X1 U16488 ( .A1(n13315), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13281) );
  AOI211_X1 U16489 ( .C1(n12842), .C2(P1_EAX_REG_29__SCAN_IN), .A(n14232), .B(
        n13281), .ZN(n13303) );
  NAND2_X1 U16490 ( .A1(n13283), .A2(n13282), .ZN(n13335) );
  AOI22_X1 U16491 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13328), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U16492 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U16493 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U16494 ( .A1(n13285), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13286) );
  NAND4_X1 U16495 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13299) );
  AOI22_X1 U16496 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16497 ( .A1(n13291), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13296) );
  AOI22_X1 U16498 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9754), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16499 ( .A1(n13293), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13292), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13294) );
  NAND4_X1 U16500 ( .A1(n13297), .A2(n13296), .A3(n13295), .A4(n13294), .ZN(
        n13298) );
  NOR2_X1 U16501 ( .A1(n13299), .A2(n13298), .ZN(n13336) );
  XOR2_X1 U16502 ( .A(n13335), .B(n13336), .Z(n13301) );
  NAND2_X1 U16503 ( .A1(n13301), .A2(n13300), .ZN(n13302) );
  NAND2_X1 U16504 ( .A1(n13304), .A2(n13305), .ZN(n13345) );
  NAND3_X1 U16505 ( .A1(n20825), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n17572) );
  INV_X1 U16506 ( .A(n17572), .ZN(n13307) );
  NOR2_X2 U16507 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21420) );
  NOR2_X1 U16508 ( .A1(n9885), .A2(n13308), .ZN(n13309) );
  OR2_X1 U16509 ( .A1(n10868), .A2(n20822), .ZN(n13310) );
  NOR2_X1 U16510 ( .A1(n17482), .A2(n13310), .ZN(n13311) );
  NAND2_X1 U16511 ( .A1(n21418), .A2(n13312), .ZN(n21573) );
  NAND2_X1 U16512 ( .A1(n21573), .A2(n20825), .ZN(n13313) );
  NAND2_X1 U16513 ( .A1(n20825), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17494) );
  NAND2_X1 U16514 ( .A1(n21173), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U16515 ( .A1(n17494), .A2(n13314), .ZN(n13624) );
  NAND2_X1 U16516 ( .A1(n17539), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n15373) );
  OAI21_X1 U16517 ( .B1(n17533), .B2(n13315), .A(n15373), .ZN(n13316) );
  AOI21_X1 U16518 ( .B1(n14727), .B2(n17528), .A(n13316), .ZN(n13317) );
  XOR2_X1 U16519 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n14227), .Z(
        n15169) );
  AOI22_X1 U16520 ( .A1(n9718), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13325) );
  AOI22_X1 U16521 ( .A1(n13320), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13319), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13324) );
  AOI22_X1 U16522 ( .A1(n13995), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n13284), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13323) );
  AOI22_X1 U16523 ( .A1(n13321), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10955), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13322) );
  NAND4_X1 U16524 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13334) );
  AOI22_X1 U16525 ( .A1(n13327), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13326), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13332) );
  AOI22_X1 U16526 ( .A1(n13328), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13133), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13331) );
  AOI22_X1 U16527 ( .A1(n13187), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n13186), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13330) );
  AOI22_X1 U16528 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13269), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13329) );
  NAND4_X1 U16529 ( .A1(n13332), .A2(n13331), .A3(n13330), .A4(n13329), .ZN(
        n13333) );
  NOR2_X1 U16530 ( .A1(n13334), .A2(n13333), .ZN(n13338) );
  NOR2_X1 U16531 ( .A1(n13336), .A2(n13335), .ZN(n13337) );
  XOR2_X1 U16532 ( .A(n13338), .B(n13337), .Z(n13343) );
  AOI21_X1 U16533 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21578), .A(
        n14232), .ZN(n13341) );
  NAND2_X1 U16534 ( .A1(n13339), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13340) );
  OAI211_X1 U16535 ( .C1(n13343), .C2(n13342), .A(n13341), .B(n13340), .ZN(
        n13344) );
  OAI21_X1 U16536 ( .B1(n15169), .B2(n9867), .A(n13344), .ZN(n14749) );
  NAND2_X1 U16537 ( .A1(n13348), .A2(n13545), .ZN(n13979) );
  NAND3_X1 U16538 ( .A1(n11324), .A2(n11217), .A3(n21574), .ZN(n13349) );
  NAND2_X1 U16539 ( .A1(n13979), .A2(n13349), .ZN(n13350) );
  NAND2_X1 U16540 ( .A1(n17503), .A2(n13350), .ZN(n13354) );
  INV_X1 U16541 ( .A(n13351), .ZN(n17566) );
  NAND2_X1 U16542 ( .A1(n17566), .A2(n13352), .ZN(n13353) );
  INV_X1 U16543 ( .A(n10872), .ZN(n14730) );
  AND4_X1 U16544 ( .A1(n10866), .A2(n14730), .A3(n13550), .A4(n10858), .ZN(
        n13355) );
  NAND2_X1 U16545 ( .A1(n13356), .A2(n13355), .ZN(n13630) );
  AND2_X1 U16546 ( .A1(n15151), .A2(n14730), .ZN(n13359) );
  NAND2_X1 U16547 ( .A1(n15166), .A2(n13359), .ZN(n13378) );
  NOR4_X1 U16548 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13363) );
  NOR4_X1 U16549 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13362) );
  NOR4_X1 U16550 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13361) );
  NOR4_X1 U16551 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13360) );
  AND4_X1 U16552 ( .A1(n13363), .A2(n13362), .A3(n13361), .A4(n13360), .ZN(
        n13368) );
  NOR4_X1 U16553 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_7__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13366) );
  NOR4_X1 U16554 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13365) );
  NOR4_X1 U16555 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13364) );
  INV_X1 U16556 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21499) );
  AND4_X1 U16557 ( .A1(n13366), .A2(n13365), .A3(n13364), .A4(n21499), .ZN(
        n13367) );
  NAND2_X1 U16558 ( .A1(n13368), .A2(n13367), .ZN(n13369) );
  NOR2_X1 U16559 ( .A1(n13372), .A2(n14274), .ZN(n13370) );
  NAND2_X1 U16560 ( .A1(n15151), .A2(n13370), .ZN(n15138) );
  NOR2_X1 U16561 ( .A1(n15138), .A2(n13371), .ZN(n13376) );
  NOR3_X1 U16562 ( .A1(n15156), .A2(n15096), .A3(n13372), .ZN(n13373) );
  AOI22_X1 U16563 ( .A1(n15140), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15156), .ZN(n13374) );
  INV_X1 U16564 ( .A(n13374), .ZN(n13375) );
  NOR2_X1 U16565 ( .A1(n13376), .A2(n13375), .ZN(n13377) );
  NAND2_X1 U16566 ( .A1(n13378), .A2(n13377), .ZN(P1_U2873) );
  NOR2_X1 U16567 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13380) );
  NOR4_X1 U16568 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13379) );
  NAND4_X1 U16569 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13380), .A4(n13379), .ZN(n13383) );
  INV_X1 U16570 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21571) );
  NOR3_X1 U16571 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21571), .ZN(n13382) );
  NOR4_X1 U16572 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13381) );
  NAND4_X1 U16573 ( .A1(n15096), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13382), .A4(
        n13381), .ZN(U214) );
  INV_X2 U16574 ( .A(n16847), .ZN(n16849) );
  NOR2_X1 U16575 ( .A1(n16849), .A2(n13383), .ZN(n17618) );
  NAND2_X1 U16576 ( .A1(n17618), .A2(U214), .ZN(U212) );
  NAND2_X1 U16577 ( .A1(n15951), .A2(n15825), .ZN(n15828) );
  AOI21_X1 U16578 ( .B1(n10339), .B2(n10340), .A(n15828), .ZN(n13402) );
  INV_X1 U16579 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U16580 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  NOR2_X1 U16581 ( .A1(n13427), .A2(n13386), .ZN(n13387) );
  OR2_X2 U16582 ( .A1(n13388), .A2(n13387), .ZN(n19980) );
  AOI22_X1 U16583 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19980), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19981), .ZN(n13389) );
  OAI211_X1 U16584 ( .C1(n11973), .C2(n15970), .A(n13389), .B(n16464), .ZN(
        n13401) );
  OAI22_X1 U16585 ( .A1(n15969), .A2(n16370), .B1(n13390), .B2(n12363), .ZN(
        n13400) );
  AND2_X1 U16586 ( .A1(n13392), .A2(n13393), .ZN(n13394) );
  NOR2_X1 U16587 ( .A1(n13391), .A2(n13394), .ZN(n16636) );
  INV_X1 U16588 ( .A(n16636), .ZN(n14214) );
  NAND2_X1 U16589 ( .A1(n13396), .A2(n13397), .ZN(n13398) );
  NAND2_X1 U16590 ( .A1(n13395), .A2(n13398), .ZN(n16632) );
  OAI22_X1 U16591 ( .A1(n14214), .A2(n19983), .B1(n16632), .B2(n19987), .ZN(
        n13399) );
  OR4_X1 U16592 ( .A1(n13402), .A2(n13401), .A3(n13400), .A4(n13399), .ZN(
        P2_U2842) );
  INV_X1 U16593 ( .A(n14234), .ZN(n13590) );
  INV_X1 U16594 ( .A(HOLD), .ZN(n21491) );
  INV_X1 U16595 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n21494) );
  NAND2_X1 U16596 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n13403) );
  OAI21_X1 U16597 ( .B1(n21491), .B2(n21483), .A(n13403), .ZN(n13404) );
  OAI21_X1 U16598 ( .B1(n21491), .B2(n21494), .A(n13404), .ZN(n13405) );
  OAI211_X1 U16599 ( .C1(n21483), .C2(n21574), .A(n13590), .B(n13405), .ZN(
        P1_U3195) );
  AND2_X1 U16600 ( .A1(n20812), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16944) );
  OAI21_X1 U16601 ( .B1(n20395), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n20489), 
        .ZN(n13409) );
  INV_X1 U16602 ( .A(n13406), .ZN(n13408) );
  NAND2_X1 U16603 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20778) );
  INV_X1 U16604 ( .A(n20778), .ZN(n13407) );
  NAND2_X1 U16605 ( .A1(n13407), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n17507) );
  OAI211_X1 U16606 ( .C1(n16944), .C2(n13409), .A(n13408), .B(n17507), .ZN(
        n13410) );
  INV_X1 U16607 ( .A(n13410), .ZN(P2_U3178) );
  INV_X1 U16608 ( .A(n13411), .ZN(n13412) );
  INV_X1 U16609 ( .A(n13529), .ZN(n20027) );
  NAND2_X1 U16610 ( .A1(n13412), .A2(n20027), .ZN(n19988) );
  INV_X1 U16611 ( .A(n19988), .ZN(n15988) );
  INV_X1 U16612 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n20820) );
  AND2_X1 U16613 ( .A1(n13427), .A2(n13413), .ZN(n13417) );
  OAI21_X1 U16614 ( .B1(n15988), .B2(n20820), .A(n13417), .ZN(P2_U2814) );
  INV_X1 U16615 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n13414) );
  OAI22_X1 U16616 ( .A1(n13415), .A2(n13414), .B1(n20808), .B2(n13413), .ZN(
        P2_U2816) );
  INV_X1 U16617 ( .A(P2_READREQUEST_REG_SCAN_IN), .ZN(n13416) );
  NAND3_X1 U16618 ( .A1(n13417), .A2(n19988), .A3(n13416), .ZN(n13418) );
  OAI21_X1 U16619 ( .B1(n20805), .B2(n20810), .A(n13418), .ZN(n13419) );
  INV_X1 U16620 ( .A(n13419), .ZN(P2_U3612) );
  NOR2_X1 U16621 ( .A1(n13420), .A2(n13527), .ZN(n13421) );
  AND2_X1 U16622 ( .A1(n13422), .A2(n13421), .ZN(n16922) );
  NOR2_X1 U16623 ( .A1(n16922), .A2(n13423), .ZN(n20797) );
  INV_X1 U16624 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13536) );
  OAI21_X1 U16625 ( .B1(n20797), .B2(n13536), .A(n13424), .ZN(P2_U2819) );
  INV_X1 U16626 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n20062) );
  NOR3_X4 U16627 ( .A1(n13427), .A2(n16029), .A3(n20686), .ZN(n13512) );
  INV_X1 U16628 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17661) );
  OR2_X1 U16629 ( .A1(n16849), .A2(n17661), .ZN(n13426) );
  NAND2_X1 U16630 ( .A1(n16849), .A2(BUF2_REG_0__SCAN_IN), .ZN(n13425) );
  NAND2_X1 U16631 ( .A1(n13426), .A2(n13425), .ZN(n16192) );
  NAND2_X1 U16632 ( .A1(n13512), .A2(n16192), .ZN(n13503) );
  INV_X1 U16633 ( .A(n13427), .ZN(n13428) );
  NAND2_X1 U16634 ( .A1(n13452), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13429) );
  OAI211_X1 U16635 ( .C1(n20062), .C2(n20028), .A(n13503), .B(n13429), .ZN(
        P2_U2952) );
  INV_X1 U16636 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n20066) );
  INV_X1 U16637 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13430) );
  OR2_X1 U16638 ( .A1(n16849), .A2(n13430), .ZN(n13432) );
  NAND2_X1 U16639 ( .A1(n16849), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13431) );
  NAND2_X1 U16640 ( .A1(n13432), .A2(n13431), .ZN(n14708) );
  NAND2_X1 U16641 ( .A1(n13512), .A2(n14708), .ZN(n13525) );
  NAND2_X1 U16642 ( .A1(n13452), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13433) );
  OAI211_X1 U16643 ( .C1(n20066), .C2(n20028), .A(n13525), .B(n13433), .ZN(
        P2_U2981) );
  INV_X1 U16644 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n20040) );
  INV_X1 U16645 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n21784) );
  OR2_X1 U16646 ( .A1(n16849), .A2(n21784), .ZN(n13435) );
  NAND2_X1 U16647 ( .A1(n16849), .A2(BUF2_REG_12__SCAN_IN), .ZN(n13434) );
  NAND2_X1 U16648 ( .A1(n13435), .A2(n13434), .ZN(n16100) );
  NAND2_X1 U16649 ( .A1(n13512), .A2(n16100), .ZN(n13441) );
  NAND2_X1 U16650 ( .A1(n13452), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13436) );
  OAI211_X1 U16651 ( .C1(n20040), .C2(n20028), .A(n13441), .B(n13436), .ZN(
        P2_U2964) );
  INV_X1 U16652 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20073) );
  INV_X1 U16653 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n17644) );
  OR2_X1 U16654 ( .A1(n16849), .A2(n17644), .ZN(n13438) );
  NAND2_X1 U16655 ( .A1(n16849), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13437) );
  NAND2_X1 U16656 ( .A1(n13438), .A2(n13437), .ZN(n16116) );
  NAND2_X1 U16657 ( .A1(n13512), .A2(n16116), .ZN(n13443) );
  NAND2_X1 U16658 ( .A1(n13452), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13439) );
  OAI211_X1 U16659 ( .C1(n20073), .C2(n20028), .A(n13443), .B(n13439), .ZN(
        P2_U2977) );
  INV_X1 U16660 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n20069) );
  NAND2_X1 U16661 ( .A1(n13452), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13440) );
  OAI211_X1 U16662 ( .C1(n20069), .C2(n20028), .A(n13441), .B(n13440), .ZN(
        P2_U2979) );
  INV_X1 U16663 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20043) );
  NAND2_X1 U16664 ( .A1(n13452), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13442) );
  OAI211_X1 U16665 ( .C1(n20043), .C2(n20028), .A(n13443), .B(n13442), .ZN(
        P2_U2962) );
  AND2_X1 U16666 ( .A1(n11324), .A2(n13550), .ZN(n13444) );
  INV_X1 U16667 ( .A(n13555), .ZN(n13445) );
  NOR2_X1 U16668 ( .A1(n13556), .A2(n13445), .ZN(n13546) );
  NAND2_X1 U16669 ( .A1(n13546), .A2(n13550), .ZN(n14225) );
  NAND2_X1 U16670 ( .A1(n21420), .A2(n13446), .ZN(n20826) );
  INV_X1 U16671 ( .A(n20826), .ZN(n14744) );
  AOI21_X1 U16672 ( .B1(n14225), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14744), 
        .ZN(n13447) );
  NAND2_X1 U16673 ( .A1(n14226), .A2(n13447), .ZN(P1_U2801) );
  INV_X1 U16674 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13448) );
  OR2_X1 U16675 ( .A1(n16849), .A2(n13448), .ZN(n13450) );
  NAND2_X1 U16676 ( .A1(n16849), .A2(BUF2_REG_15__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U16677 ( .A1(n13450), .A2(n13449), .ZN(n14357) );
  AOI222_X1 U16678 ( .A1(n14357), .A2(n13512), .B1(n13520), .B2(
        P2_EAX_REG_15__SCAN_IN), .C1(n13452), .C2(P2_LWORD_REG_15__SCAN_IN), 
        .ZN(n13451) );
  INV_X1 U16679 ( .A(n13451), .ZN(P2_U2982) );
  AOI22_X1 U16680 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n13452), .B1(n13520), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n13455) );
  INV_X1 U16681 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17647) );
  OR2_X1 U16682 ( .A1(n16849), .A2(n17647), .ZN(n13454) );
  NAND2_X1 U16683 ( .A1(n16849), .A2(BUF2_REG_8__SCAN_IN), .ZN(n13453) );
  NAND2_X1 U16684 ( .A1(n13454), .A2(n13453), .ZN(n16130) );
  NAND2_X1 U16685 ( .A1(n13512), .A2(n16130), .ZN(n13493) );
  NAND2_X1 U16686 ( .A1(n13455), .A2(n13493), .ZN(P2_U2960) );
  AOI22_X1 U16687 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n13460) );
  INV_X1 U16688 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n13456) );
  OR2_X1 U16689 ( .A1(n16849), .A2(n13456), .ZN(n13458) );
  NAND2_X1 U16690 ( .A1(n16849), .A2(BUF2_REG_1__SCAN_IN), .ZN(n13457) );
  AND2_X1 U16691 ( .A1(n13458), .A2(n13457), .ZN(n20025) );
  INV_X1 U16692 ( .A(n20025), .ZN(n13459) );
  NAND2_X1 U16693 ( .A1(n13512), .A2(n13459), .ZN(n13505) );
  NAND2_X1 U16694 ( .A1(n13460), .A2(n13505), .ZN(P2_U2953) );
  AOI22_X1 U16695 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n13463) );
  INV_X1 U16696 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17654) );
  OR2_X1 U16697 ( .A1(n16849), .A2(n17654), .ZN(n13462) );
  NAND2_X1 U16698 ( .A1(n16849), .A2(BUF2_REG_2__SCAN_IN), .ZN(n13461) );
  NAND2_X1 U16699 ( .A1(n13462), .A2(n13461), .ZN(n16174) );
  NAND2_X1 U16700 ( .A1(n13512), .A2(n16174), .ZN(n13485) );
  NAND2_X1 U16701 ( .A1(n13463), .A2(n13485), .ZN(P2_U2969) );
  AOI22_X1 U16702 ( .A1(P2_LWORD_REG_11__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n13467) );
  INV_X1 U16703 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n13464) );
  OR2_X1 U16704 ( .A1(n16849), .A2(n13464), .ZN(n13466) );
  NAND2_X1 U16705 ( .A1(n16849), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U16706 ( .A1(n13466), .A2(n13465), .ZN(n16108) );
  NAND2_X1 U16707 ( .A1(n13512), .A2(n16108), .ZN(n13487) );
  NAND2_X1 U16708 ( .A1(n13467), .A2(n13487), .ZN(P2_U2978) );
  AOI22_X1 U16709 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n13471) );
  INV_X1 U16710 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n13468) );
  NOR2_X1 U16711 ( .A1(n16849), .A2(n13468), .ZN(n13469) );
  AOI21_X1 U16712 ( .B1(BUF2_REG_3__SCAN_IN), .B2(n16849), .A(n13469), .ZN(
        n20120) );
  INV_X1 U16713 ( .A(n20120), .ZN(n13470) );
  NAND2_X1 U16714 ( .A1(n13512), .A2(n13470), .ZN(n13489) );
  NAND2_X1 U16715 ( .A1(n13471), .A2(n13489), .ZN(P2_U2955) );
  AOI22_X1 U16716 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n13476) );
  INV_X1 U16717 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n13472) );
  OR2_X1 U16718 ( .A1(n16849), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U16719 ( .A1(n16849), .A2(BUF2_REG_4__SCAN_IN), .ZN(n13473) );
  AND2_X1 U16720 ( .A1(n13474), .A2(n13473), .ZN(n20124) );
  INV_X1 U16721 ( .A(n20124), .ZN(n13475) );
  NAND2_X1 U16722 ( .A1(n13512), .A2(n13475), .ZN(n13491) );
  NAND2_X1 U16723 ( .A1(n13476), .A2(n13491), .ZN(P2_U2956) );
  AOI22_X1 U16724 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n13480) );
  INV_X1 U16725 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n13477) );
  OR2_X1 U16726 ( .A1(n16849), .A2(n13477), .ZN(n13479) );
  NAND2_X1 U16727 ( .A1(n16849), .A2(BUF2_REG_5__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U16728 ( .A1(n13479), .A2(n13478), .ZN(n20129) );
  NAND2_X1 U16729 ( .A1(n13512), .A2(n20129), .ZN(n13521) );
  NAND2_X1 U16730 ( .A1(n13480), .A2(n13521), .ZN(P2_U2957) );
  AOI22_X1 U16731 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n13484) );
  INV_X1 U16732 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n13481) );
  OR2_X1 U16733 ( .A1(n16849), .A2(n13481), .ZN(n13483) );
  NAND2_X1 U16734 ( .A1(n16849), .A2(BUF2_REG_6__SCAN_IN), .ZN(n13482) );
  NAND2_X1 U16735 ( .A1(n13483), .A2(n13482), .ZN(n16145) );
  NAND2_X1 U16736 ( .A1(n13512), .A2(n16145), .ZN(n13518) );
  NAND2_X1 U16737 ( .A1(n13484), .A2(n13518), .ZN(P2_U2958) );
  AOI22_X1 U16738 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n13486) );
  NAND2_X1 U16739 ( .A1(n13486), .A2(n13485), .ZN(P2_U2954) );
  AOI22_X1 U16740 ( .A1(P2_UWORD_REG_11__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n13488) );
  NAND2_X1 U16741 ( .A1(n13488), .A2(n13487), .ZN(P2_U2963) );
  AOI22_X1 U16742 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n13490) );
  NAND2_X1 U16743 ( .A1(n13490), .A2(n13489), .ZN(P2_U2970) );
  AOI22_X1 U16744 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n13492) );
  NAND2_X1 U16745 ( .A1(n13492), .A2(n13491), .ZN(P2_U2971) );
  AOI22_X1 U16746 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n13494) );
  NAND2_X1 U16747 ( .A1(n13494), .A2(n13493), .ZN(P2_U2975) );
  AOI22_X1 U16748 ( .A1(P2_UWORD_REG_13__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n13498) );
  INV_X1 U16749 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13495) );
  OR2_X1 U16750 ( .A1(n16849), .A2(n13495), .ZN(n13497) );
  NAND2_X1 U16751 ( .A1(n16849), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13496) );
  NAND2_X1 U16752 ( .A1(n13497), .A2(n13496), .ZN(n16093) );
  NAND2_X1 U16753 ( .A1(n13512), .A2(n16093), .ZN(n13514) );
  NAND2_X1 U16754 ( .A1(n13498), .A2(n13514), .ZN(P2_U2965) );
  AOI22_X1 U16755 ( .A1(P2_LWORD_REG_9__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n13502) );
  INV_X1 U16756 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13499) );
  OR2_X1 U16757 ( .A1(n16849), .A2(n13499), .ZN(n13501) );
  NAND2_X1 U16758 ( .A1(n16849), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13500) );
  NAND2_X1 U16759 ( .A1(n13501), .A2(n13500), .ZN(n16124) );
  NAND2_X1 U16760 ( .A1(n13512), .A2(n16124), .ZN(n13507) );
  NAND2_X1 U16761 ( .A1(n13502), .A2(n13507), .ZN(P2_U2976) );
  AOI22_X1 U16762 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n13504) );
  NAND2_X1 U16763 ( .A1(n13504), .A2(n13503), .ZN(P2_U2967) );
  AOI22_X1 U16764 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n13506) );
  NAND2_X1 U16765 ( .A1(n13506), .A2(n13505), .ZN(P2_U2968) );
  AOI22_X1 U16766 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n13508) );
  NAND2_X1 U16767 ( .A1(n13508), .A2(n13507), .ZN(P2_U2961) );
  AOI22_X1 U16768 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n13513) );
  INV_X1 U16769 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13509) );
  OR2_X1 U16770 ( .A1(n16849), .A2(n13509), .ZN(n13511) );
  NAND2_X1 U16771 ( .A1(n16849), .A2(BUF2_REG_7__SCAN_IN), .ZN(n13510) );
  NAND2_X1 U16772 ( .A1(n13511), .A2(n13510), .ZN(n16138) );
  NAND2_X1 U16773 ( .A1(n13512), .A2(n16138), .ZN(n13516) );
  NAND2_X1 U16774 ( .A1(n13513), .A2(n13516), .ZN(P2_U2959) );
  AOI22_X1 U16775 ( .A1(P2_LWORD_REG_13__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n13515) );
  NAND2_X1 U16776 ( .A1(n13515), .A2(n13514), .ZN(P2_U2980) );
  AOI22_X1 U16777 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U16778 ( .A1(n13517), .A2(n13516), .ZN(P2_U2974) );
  AOI22_X1 U16779 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n13519) );
  NAND2_X1 U16780 ( .A1(n13519), .A2(n13518), .ZN(P2_U2973) );
  AOI22_X1 U16781 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n13523), .B1(n13520), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n13522) );
  NAND2_X1 U16782 ( .A1(n13522), .A2(n13521), .ZN(P2_U2972) );
  INV_X1 U16783 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n20036) );
  NAND2_X1 U16784 ( .A1(n13523), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13524) );
  OAI211_X1 U16785 ( .C1(n20036), .C2(n20028), .A(n13525), .B(n13524), .ZN(
        P2_U2966) );
  INV_X1 U16786 ( .A(n13526), .ZN(n13535) );
  INV_X1 U16787 ( .A(n20030), .ZN(n13531) );
  INV_X1 U16788 ( .A(n13527), .ZN(n13528) );
  NOR2_X1 U16789 ( .A1(n13529), .A2(n13528), .ZN(n13530) );
  NAND2_X1 U16790 ( .A1(n13531), .A2(n13530), .ZN(n13534) );
  NAND4_X1 U16791 ( .A1(n13535), .A2(n13534), .A3(n13533), .A4(n13532), .ZN(
        n16925) );
  OAI22_X1 U16792 ( .A1(n17507), .A2(n13536), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n20800), .ZN(n13537) );
  INV_X1 U16793 ( .A(n16833), .ZN(n13544) );
  INV_X1 U16794 ( .A(n13538), .ZN(n13542) );
  INV_X1 U16795 ( .A(n13539), .ZN(n13540) );
  AND2_X1 U16796 ( .A1(n11465), .A2(n13540), .ZN(n13541) );
  NAND2_X1 U16797 ( .A1(n13542), .A2(n13541), .ZN(n16918) );
  OR3_X1 U16798 ( .A1(n16833), .A2(n20747), .A3(n16918), .ZN(n13543) );
  OAI21_X1 U16799 ( .B1(n13544), .B2(n16924), .A(n13543), .ZN(P2_U3595) );
  INV_X1 U16800 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13562) );
  OR2_X1 U16801 ( .A1(n17503), .A2(n13545), .ZN(n13548) );
  OR2_X1 U16802 ( .A1(n13546), .A2(n11324), .ZN(n13547) );
  NAND2_X1 U16803 ( .A1(n13548), .A2(n13547), .ZN(n20823) );
  NAND3_X1 U16804 ( .A1(n11242), .A2(n10888), .A3(n13590), .ZN(n13549) );
  AND2_X1 U16805 ( .A1(n13549), .A2(n21574), .ZN(n21576) );
  OR2_X1 U16806 ( .A1(n20823), .A2(n21576), .ZN(n17484) );
  AND2_X1 U16807 ( .A1(n17484), .A2(n13550), .ZN(n20831) );
  NAND2_X1 U16808 ( .A1(n11017), .A2(n11218), .ZN(n13552) );
  OAI21_X1 U16809 ( .B1(n11195), .B2(n13552), .A(n13551), .ZN(n13554) );
  MUX2_X1 U16810 ( .A(n13554), .B(n13553), .S(n17503), .Z(n13558) );
  NOR2_X1 U16811 ( .A1(n13556), .A2(n13555), .ZN(n13557) );
  OR2_X1 U16812 ( .A1(n13558), .A2(n13557), .ZN(n13559) );
  NAND2_X1 U16813 ( .A1(n13559), .A2(n10872), .ZN(n17486) );
  INV_X1 U16814 ( .A(n17486), .ZN(n13560) );
  NAND2_X1 U16815 ( .A1(n13560), .A2(n20831), .ZN(n13561) );
  OAI21_X1 U16816 ( .B1(n13562), .B2(n20831), .A(n13561), .ZN(P1_U3484) );
  XNOR2_X1 U16817 ( .A(n13563), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17605) );
  OAI21_X1 U16818 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15983), .A(
        n13573), .ZN(n17600) );
  NAND2_X1 U16819 ( .A1(n16754), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n17611) );
  OAI21_X1 U16820 ( .B1(n16472), .B2(n17600), .A(n17611), .ZN(n13564) );
  AOI21_X1 U16821 ( .B1(n16470), .B2(n17605), .A(n13564), .ZN(n13567) );
  OAI21_X1 U16822 ( .B1(n16445), .B2(n13565), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13566) );
  OAI211_X1 U16823 ( .C1(n17589), .C2(n10204), .A(n13567), .B(n13566), .ZN(
        P2_U3014) );
  XNOR2_X1 U16824 ( .A(n13568), .B(n13580), .ZN(n13576) );
  NAND2_X1 U16825 ( .A1(n16470), .A2(n13576), .ZN(n13569) );
  NAND2_X1 U16826 ( .A1(n16754), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13577) );
  OAI211_X1 U16827 ( .C1(n17599), .C2(n13570), .A(n13569), .B(n13577), .ZN(
        n13571) );
  INV_X1 U16828 ( .A(n13571), .ZN(n13575) );
  XNOR2_X1 U16829 ( .A(n15971), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13572) );
  XNOR2_X1 U16830 ( .A(n13573), .B(n13572), .ZN(n13583) );
  AOI22_X1 U16831 ( .A1(n17586), .A2(n13570), .B1(n17587), .B2(n13583), .ZN(
        n13574) );
  OAI211_X1 U16832 ( .C1(n15977), .C2(n17589), .A(n13575), .B(n13574), .ZN(
        P2_U3013) );
  NAND2_X1 U16833 ( .A1(n17606), .A2(n13576), .ZN(n13578) );
  NAND2_X1 U16834 ( .A1(n13578), .A2(n13577), .ZN(n13582) );
  AOI211_X1 U16835 ( .C1(n12067), .C2(n13580), .A(n13579), .B(n17615), .ZN(
        n13581) );
  AOI211_X1 U16836 ( .C1(n17602), .C2(n13583), .A(n13582), .B(n13581), .ZN(
        n13589) );
  OR2_X1 U16837 ( .A1(n13585), .A2(n13584), .ZN(n13586) );
  NAND2_X1 U16838 ( .A1(n13587), .A2(n13586), .ZN(n20772) );
  AOI22_X1 U16839 ( .A1(n17603), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n17608), .B2(n20772), .ZN(n13588) );
  OAI211_X1 U16840 ( .C1(n15977), .C2(n16764), .A(n13589), .B(n13588), .ZN(
        P2_U3045) );
  INV_X1 U16841 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13594) );
  OR3_X1 U16842 ( .A1(n14226), .A2(n11217), .A3(n13590), .ZN(n13592) );
  NAND2_X1 U16843 ( .A1(n17503), .A2(n14234), .ZN(n17497) );
  INV_X1 U16844 ( .A(n17468), .ZN(n14003) );
  NAND2_X1 U16845 ( .A1(n20940), .A2(n11218), .ZN(n13930) );
  NOR2_X1 U16846 ( .A1(n21578), .A2(n13446), .ZN(n17579) );
  NAND2_X1 U16847 ( .A1(n20825), .A2(n17579), .ZN(n20938) );
  INV_X2 U16848 ( .A(n20938), .ZN(n20967) );
  NOR2_X4 U16849 ( .A1(n20940), .A2(n20967), .ZN(n20966) );
  AOI22_X1 U16850 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13593) );
  OAI21_X1 U16851 ( .B1(n13594), .B2(n13930), .A(n13593), .ZN(P1_U2909) );
  INV_X1 U16852 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U16853 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U16854 ( .B1(n13596), .B2(n13930), .A(n13595), .ZN(P1_U2912) );
  INV_X1 U16855 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U16856 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13597) );
  OAI21_X1 U16857 ( .B1(n13598), .B2(n13930), .A(n13597), .ZN(P1_U2911) );
  INV_X1 U16858 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13600) );
  AOI22_X1 U16859 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U16860 ( .B1(n13600), .B2(n13930), .A(n13599), .ZN(P1_U2907) );
  INV_X1 U16861 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13602) );
  AOI22_X1 U16862 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U16863 ( .B1(n13602), .B2(n13930), .A(n13601), .ZN(P1_U2908) );
  INV_X1 U16864 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21638) );
  AOI22_X1 U16865 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13603) );
  OAI21_X1 U16866 ( .B1(n21638), .B2(n13930), .A(n13603), .ZN(P1_U2910) );
  INV_X1 U16867 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13605) );
  AOI22_X1 U16868 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13604) );
  OAI21_X1 U16869 ( .B1(n13605), .B2(n13930), .A(n13604), .ZN(P1_U2906) );
  NAND2_X1 U16870 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  INV_X1 U16871 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15972) );
  MUX2_X1 U16872 ( .A(n15972), .B(n15977), .S(n16080), .Z(n13610) );
  OAI21_X1 U16873 ( .B1(n20750), .B2(n16072), .A(n13610), .ZN(P2_U2886) );
  NAND2_X1 U16874 ( .A1(n16887), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13611) );
  INV_X1 U16875 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13613) );
  MUX2_X1 U16876 ( .A(n10204), .B(n13613), .S(n16078), .Z(n13614) );
  OAI21_X1 U16877 ( .B1(n20781), .B2(n16072), .A(n13614), .ZN(P2_U2887) );
  INV_X1 U16878 ( .A(n13615), .ZN(n13619) );
  INV_X1 U16879 ( .A(n13616), .ZN(n13618) );
  OAI21_X1 U16880 ( .B1(n13619), .B2(n13618), .A(n13617), .ZN(n14253) );
  INV_X1 U16881 ( .A(n14375), .ZN(n21287) );
  AOI211_X1 U16882 ( .C1(n21287), .C2(n13621), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n13620), .ZN(n13623) );
  NOR2_X1 U16883 ( .A1(n13623), .A2(n13622), .ZN(n21000) );
  OAI21_X1 U16884 ( .B1(n17517), .B2(n13624), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U16885 ( .A1(n17539), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n21005) );
  NAND2_X1 U16886 ( .A1(n13625), .A2(n21005), .ZN(n13626) );
  AOI21_X1 U16887 ( .B1(n21000), .B2(n17531), .A(n13626), .ZN(n13627) );
  OAI21_X1 U16888 ( .B1(n15370), .B2(n14253), .A(n13627), .ZN(P1_U2999) );
  OAI21_X1 U16889 ( .B1(n13629), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13628), .ZN(n20996) );
  OR2_X1 U16890 ( .A1(n13630), .A2(n11242), .ZN(n13631) );
  INV_X2 U16891 ( .A(n20932), .ZN(n15079) );
  OAI222_X1 U16892 ( .A1(n20996), .A2(n20925), .B1(n20936), .B2(n14246), .C1(
        n14253), .C2(n15079), .ZN(P1_U2872) );
  XNOR2_X1 U16893 ( .A(n13633), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13646) );
  OAI21_X1 U16894 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n15533), .A(
        n14464), .ZN(n21002) );
  INV_X1 U16895 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21495) );
  NOR2_X1 U16896 ( .A1(n20904), .A2(n21495), .ZN(n13648) );
  OR2_X1 U16897 ( .A1(n13635), .A2(n13634), .ZN(n13636) );
  AND2_X1 U16898 ( .A1(n13637), .A2(n13636), .ZN(n15048) );
  NOR2_X1 U16899 ( .A1(n15048), .A2(n15576), .ZN(n13638) );
  AOI211_X1 U16900 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n21002), .A(
        n13648), .B(n13638), .ZN(n13640) );
  OAI211_X1 U16901 ( .C1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n21003), .A(
        n15477), .B(n11219), .ZN(n13639) );
  OAI211_X1 U16902 ( .C1(n13646), .C2(n17559), .A(n13640), .B(n13639), .ZN(
        P1_U3030) );
  OAI21_X1 U16903 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(n15055) );
  INV_X1 U16904 ( .A(n15048), .ZN(n13644) );
  AOI22_X1 U16905 ( .A1(n20931), .A2(n13644), .B1(n15075), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13645) );
  OAI21_X1 U16906 ( .B1(n15055), .B2(n15079), .A(n13645), .ZN(P1_U2871) );
  INV_X1 U16907 ( .A(n13646), .ZN(n13649) );
  MUX2_X1 U16908 ( .A(n17528), .B(n17517), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13647) );
  AOI211_X1 U16909 ( .C1(n13649), .C2(n17531), .A(n13648), .B(n13647), .ZN(
        n13650) );
  OAI21_X1 U16910 ( .B1(n15370), .B2(n15055), .A(n13650), .ZN(P1_U2998) );
  AND2_X2 U16911 ( .A1(n13910), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13912) );
  INV_X1 U16912 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13652) );
  AND2_X4 U16913 ( .A1(n13654), .A2(n17415), .ZN(n18419) );
  AOI22_X1 U16914 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13651) );
  OAI21_X1 U16915 ( .B1(n10740), .B2(n13652), .A(n13651), .ZN(n13653) );
  AOI21_X1 U16916 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n13653), .ZN(n13658) );
  AND2_X2 U16917 ( .A1(n17403), .A2(n13665), .ZN(n14524) );
  INV_X4 U16918 ( .A(n18285), .ZN(n18457) );
  AOI22_X1 U16919 ( .A1(n14578), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13657) );
  AND2_X4 U16920 ( .A1(n13910), .A2(n13655), .ZN(n18459) );
  AOI22_X1 U16921 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13656) );
  NAND3_X1 U16922 ( .A1(n13658), .A2(n13657), .A3(n13656), .ZN(n13671) );
  NAND2_X4 U16923 ( .A1(n14479), .A2(n17398), .ZN(n18455) );
  INV_X1 U16924 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U16925 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13661) );
  OAI21_X1 U16926 ( .B1(n18330), .B2(n17440), .A(n13661), .ZN(n13662) );
  AOI21_X1 U16927 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n13662), .ZN(n13669) );
  AOI22_X1 U16928 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13684), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13668) );
  INV_X2 U16929 ( .A(n13705), .ZN(n17006) );
  AOI22_X1 U16930 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13667) );
  NAND3_X1 U16931 ( .A1(n13669), .A2(n13668), .A3(n13667), .ZN(n13670) );
  INV_X1 U16932 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14555) );
  AOI22_X1 U16933 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18419), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U16934 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13672) );
  OAI211_X1 U16935 ( .C1(n14555), .C2(n18301), .A(n13673), .B(n13672), .ZN(
        n13676) );
  INV_X1 U16936 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18132) );
  INV_X1 U16937 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18327) );
  OAI22_X1 U16938 ( .A1(n14490), .A2(n18132), .B1(n18285), .B2(n18327), .ZN(
        n13675) );
  INV_X1 U16939 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n18131) );
  OAI22_X1 U16940 ( .A1(n18328), .A2(n18445), .B1(n9724), .B2(n18131), .ZN(
        n13674) );
  INV_X1 U16941 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18326) );
  INV_X2 U16942 ( .A(n9712), .ZN(n18432) );
  INV_X2 U16943 ( .A(n13703), .ZN(n18237) );
  AOI22_X1 U16944 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13677) );
  OAI21_X1 U16945 ( .B1(n10740), .B2(n18326), .A(n13677), .ZN(n13678) );
  AOI21_X1 U16946 ( .B1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9717), .A(
        n13678), .ZN(n13681) );
  AOI22_X1 U16947 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n17006), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13680) );
  AOI22_X1 U16948 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13679) );
  NAND3_X1 U16949 ( .A1(n13681), .A2(n13680), .A3(n13679), .ZN(n13682) );
  AOI22_X1 U16950 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13688) );
  AOI22_X1 U16951 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13687) );
  AOI22_X1 U16952 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18450), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13686) );
  AOI22_X1 U16953 ( .A1(n14578), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13685) );
  NAND4_X1 U16954 ( .A1(n13688), .A2(n13687), .A3(n13686), .A4(n13685), .ZN(
        n13695) );
  INV_X1 U16955 ( .A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14507) );
  INV_X1 U16956 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14506) );
  INV_X1 U16957 ( .A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18382) );
  OAI22_X1 U16958 ( .A1(n9712), .A2(n14506), .B1(n18402), .B2(n18382), .ZN(
        n13691) );
  INV_X1 U16959 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18379) );
  INV_X1 U16960 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13689) );
  OAI22_X1 U16961 ( .A1(n18443), .A2(n18379), .B1(n13729), .B2(n13689), .ZN(
        n13690) );
  AOI22_X1 U16962 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13692) );
  OAI211_X1 U16963 ( .C1(n18455), .C2(n14507), .A(n13693), .B(n13692), .ZN(
        n13694) );
  INV_X1 U16964 ( .A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13697) );
  INV_X1 U16965 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13696) );
  OAI22_X1 U16966 ( .A1(n18301), .A2(n13697), .B1(n18402), .B2(n13696), .ZN(
        n13702) );
  INV_X1 U16967 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n18400) );
  OAI22_X1 U16968 ( .A1(n18285), .A2(n18400), .B1(n10740), .B2(n18401), .ZN(
        n13701) );
  INV_X1 U16969 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n18404) );
  AOI22_X1 U16970 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U16971 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13698) );
  OAI211_X1 U16972 ( .C1(n18404), .C2(n10739), .A(n13699), .B(n13698), .ZN(
        n13700) );
  AOI22_X1 U16973 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18432), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13709) );
  AOI22_X1 U16974 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13708) );
  AOI22_X1 U16975 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13704) );
  OAI21_X1 U16976 ( .B1(n13705), .B2(n18272), .A(n13704), .ZN(n13706) );
  AOI21_X1 U16977 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n13706), .ZN(n13707) );
  NAND3_X1 U16978 ( .A1(n13709), .A2(n13708), .A3(n13707), .ZN(n13710) );
  NAND2_X1 U16979 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n13713) );
  NAND2_X1 U16980 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13712) );
  OAI211_X1 U16981 ( .C1(n18455), .C2(n21743), .A(n13713), .B(n13712), .ZN(
        n13714) );
  INV_X1 U16982 ( .A(n13714), .ZN(n13718) );
  INV_X2 U16983 ( .A(n18301), .ZN(n18425) );
  AOI22_X1 U16984 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13717) );
  AOI22_X1 U16985 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U16986 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13715) );
  NAND4_X1 U16987 ( .A1(n13718), .A2(n13717), .A3(n13716), .A4(n13715), .ZN(
        n13724) );
  AOI22_X1 U16988 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13722) );
  AOI22_X1 U16989 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13721) );
  INV_X2 U16990 ( .A(n13729), .ZN(n18456) );
  AOI22_X1 U16991 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13720) );
  AOI22_X1 U16992 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13719) );
  NAND4_X1 U16993 ( .A1(n13722), .A2(n13721), .A3(n13720), .A4(n13719), .ZN(
        n13723) );
  INV_X1 U16994 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13727) );
  NAND2_X1 U16995 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13726) );
  NAND2_X1 U16996 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n13725) );
  OAI211_X1 U16997 ( .C1(n18455), .C2(n13727), .A(n13726), .B(n13725), .ZN(
        n13728) );
  INV_X1 U16998 ( .A(n13728), .ZN(n13733) );
  AOI22_X1 U16999 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13732) );
  AOI22_X1 U17000 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13731) );
  NAND2_X1 U17001 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13730) );
  NAND4_X1 U17002 ( .A1(n13733), .A2(n13732), .A3(n13731), .A4(n13730), .ZN(
        n13739) );
  AOI22_X1 U17003 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13737) );
  AOI22_X1 U17004 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13736) );
  AOI22_X1 U17005 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13735) );
  AOI22_X1 U17006 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13734) );
  NAND4_X1 U17007 ( .A1(n13737), .A2(n13736), .A3(n13735), .A4(n13734), .ZN(
        n13738) );
  NAND2_X1 U17008 ( .A1(n19373), .A2(n18502), .ZN(n13767) );
  NAND3_X1 U17009 ( .A1(n13766), .A2(n13898), .A3(n13767), .ZN(n13778) );
  NAND2_X1 U17010 ( .A1(n13766), .A2(n18509), .ZN(n13816) );
  INV_X1 U17011 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13742) );
  NAND2_X1 U17012 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13741) );
  OAI211_X1 U17013 ( .C1(n18455), .C2(n13742), .A(n13741), .B(n13740), .ZN(
        n13743) );
  INV_X1 U17014 ( .A(n13743), .ZN(n13747) );
  AOI22_X1 U17015 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13746) );
  AOI22_X1 U17016 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U17017 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13744) );
  INV_X2 U17018 ( .A(n13748), .ZN(n18153) );
  AOI22_X1 U17019 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13752) );
  AOI22_X1 U17020 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13751) );
  AOI22_X1 U17021 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13750) );
  AOI22_X1 U17022 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13749) );
  INV_X1 U17023 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U17024 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13754) );
  NAND2_X1 U17025 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13753) );
  OAI211_X1 U17026 ( .C1(n18455), .C2(n14527), .A(n13754), .B(n13753), .ZN(
        n13755) );
  INV_X1 U17027 ( .A(n13755), .ZN(n13759) );
  AOI22_X1 U17028 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13758) );
  AOI22_X1 U17029 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13757) );
  NAND2_X1 U17030 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13756) );
  NAND4_X1 U17031 ( .A1(n13759), .A2(n13758), .A3(n13757), .A4(n13756), .ZN(
        n13765) );
  AOI22_X1 U17032 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18269), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17033 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13762) );
  AOI22_X1 U17034 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U17035 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13760) );
  NAND4_X1 U17036 ( .A1(n13763), .A2(n13762), .A3(n13761), .A4(n13760), .ZN(
        n13764) );
  NOR2_X1 U17037 ( .A1(n18651), .A2(n9733), .ZN(n13768) );
  NAND4_X1 U17038 ( .A1(n19369), .A2(n19365), .A3(n13768), .A4(n13771), .ZN(
        n13781) );
  NOR2_X2 U17039 ( .A1(n13766), .A2(n13781), .ZN(n17708) );
  NAND2_X1 U17040 ( .A1(n13766), .A2(n19365), .ZN(n13897) );
  NOR2_X1 U17041 ( .A1(n13767), .A2(n13897), .ZN(n14483) );
  NAND2_X1 U17042 ( .A1(n19943), .A2(n13768), .ZN(n13775) );
  INV_X1 U17043 ( .A(n13775), .ZN(n13769) );
  NOR2_X1 U17044 ( .A1(n18707), .A2(n19355), .ZN(n13787) );
  OAI21_X1 U17045 ( .B1(n9734), .B2(n17397), .A(n13787), .ZN(n13795) );
  INV_X1 U17046 ( .A(n13788), .ZN(n13789) );
  AOI21_X1 U17047 ( .B1(n13766), .B2(n13789), .A(n13771), .ZN(n13774) );
  NOR2_X1 U17048 ( .A1(n9734), .A2(n13771), .ZN(n13772) );
  NOR2_X1 U17049 ( .A1(n13772), .A2(n19369), .ZN(n13773) );
  AOI211_X1 U17050 ( .C1(n19369), .C2(n17397), .A(n13774), .B(n13773), .ZN(
        n13777) );
  NAND3_X1 U17051 ( .A1(n19365), .A2(n13789), .A3(n13775), .ZN(n13776) );
  OAI211_X1 U17052 ( .C1(n13778), .C2(n18651), .A(n13777), .B(n13776), .ZN(
        n13794) );
  INV_X1 U17053 ( .A(n13794), .ZN(n13779) );
  INV_X1 U17054 ( .A(n13782), .ZN(n13784) );
  INV_X1 U17055 ( .A(n17723), .ZN(n13783) );
  NAND3_X1 U17056 ( .A1(n13784), .A2(n18707), .A3(n13783), .ZN(n13785) );
  NOR2_X1 U17057 ( .A1(n13788), .A2(n13787), .ZN(n19951) );
  OAI21_X1 U17058 ( .B1(n19377), .B2(n19369), .A(n13789), .ZN(n13790) );
  NOR2_X1 U17059 ( .A1(n13791), .A2(n13790), .ZN(n13852) );
  INV_X1 U17060 ( .A(n13852), .ZN(n13793) );
  INV_X1 U17061 ( .A(n17708), .ZN(n13792) );
  OAI21_X1 U17062 ( .B1(n13794), .B2(n13793), .A(n13792), .ZN(n13796) );
  AND2_X1 U17063 ( .A1(n13796), .A2(n13795), .ZN(n13907) );
  MUX2_X1 U17064 ( .A(n19806), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n17414), .Z(n13811) );
  NAND2_X1 U17065 ( .A1(n19587), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13812) );
  INV_X1 U17066 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13797) );
  MUX2_X1 U17067 ( .A(n13797), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        n10426), .Z(n13803) );
  OAI22_X1 U17068 ( .A1(n13802), .A2(n13803), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10426), .ZN(n13798) );
  OAI22_X1 U17069 ( .A1(n13798), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19814), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13806) );
  NOR2_X1 U17070 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19814), .ZN(
        n13799) );
  NAND2_X1 U17071 ( .A1(n13798), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13804) );
  AOI22_X1 U17072 ( .A1(n13806), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        n13799), .B2(n13804), .ZN(n13807) );
  INV_X1 U17073 ( .A(n13811), .ZN(n13801) );
  OAI21_X1 U17074 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19587), .A(
        n13812), .ZN(n13819) );
  INV_X1 U17075 ( .A(n13819), .ZN(n13800) );
  NAND3_X1 U17076 ( .A1(n13807), .A2(n13801), .A3(n13800), .ZN(n13809) );
  XOR2_X1 U17077 ( .A(n13803), .B(n13802), .Z(n13808) );
  AND2_X1 U17078 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13804), .ZN(
        n13805) );
  AOI21_X1 U17079 ( .B1(n13812), .B2(n13811), .A(n13810), .ZN(n13813) );
  NOR2_X1 U17080 ( .A1(n13814), .A2(n13813), .ZN(n13820) );
  NAND2_X1 U17081 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19944) );
  NAND2_X1 U17082 ( .A1(n18707), .A2(n13766), .ZN(n13821) );
  OAI211_X1 U17083 ( .C1(n13766), .C2(n18707), .A(n13821), .B(n19941), .ZN(
        n13815) );
  NAND2_X1 U17084 ( .A1(n19944), .A2(n13815), .ZN(n17707) );
  NOR2_X1 U17085 ( .A1(n13902), .A2(n17707), .ZN(n13817) );
  MUX2_X1 U17086 ( .A(n9870), .B(n13817), .S(n13816), .Z(n13824) );
  AOI21_X1 U17087 ( .B1(n13820), .B2(n13819), .A(n13818), .ZN(n19785) );
  INV_X1 U17088 ( .A(n13851), .ZN(n13822) );
  NOR2_X1 U17089 ( .A1(n19785), .A2(n13822), .ZN(n13823) );
  NOR2_X1 U17090 ( .A1(n13824), .A2(n13823), .ZN(n13825) );
  NAND2_X1 U17091 ( .A1(n13907), .A2(n13825), .ZN(n13826) );
  INV_X1 U17092 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14535) );
  NAND2_X1 U17093 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13827) );
  AOI22_X1 U17094 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13830) );
  AOI22_X1 U17095 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U17096 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13828) );
  NAND4_X1 U17097 ( .A1(n9850), .A2(n13830), .A3(n13829), .A4(n13828), .ZN(
        n13837) );
  INV_X2 U17098 ( .A(n9712), .ZN(n18458) );
  AOI22_X1 U17099 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13835) );
  AOI22_X1 U17100 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13834) );
  AOI22_X1 U17101 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13833) );
  AOI22_X1 U17102 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13832) );
  NAND4_X1 U17103 ( .A1(n13835), .A2(n13834), .A3(n13833), .A4(n13832), .ZN(
        n13836) );
  NOR2_X1 U17104 ( .A1(n17127), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17272) );
  INV_X1 U17105 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18284) );
  NAND2_X1 U17106 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13839) );
  NAND2_X1 U17107 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13838) );
  OAI211_X1 U17108 ( .C1(n18455), .C2(n18284), .A(n13839), .B(n13838), .ZN(
        n13840) );
  INV_X1 U17109 ( .A(n13840), .ZN(n13844) );
  AOI22_X1 U17110 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17111 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13842) );
  NAND2_X1 U17112 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13841) );
  AOI22_X1 U17113 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13848) );
  AOI22_X1 U17114 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13847) );
  AOI22_X1 U17115 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13846) );
  AOI22_X1 U17116 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13845) );
  XOR2_X1 U17117 ( .A(n17272), .B(n13849), .Z(n19047) );
  INV_X1 U17118 ( .A(n19047), .ZN(n13857) );
  OAI21_X1 U17119 ( .B1(n13849), .B2(n9808), .A(n17050), .ZN(n13850) );
  INV_X1 U17120 ( .A(n13850), .ZN(n19050) );
  NAND2_X1 U17121 ( .A1(n18649), .A2(n19923), .ZN(n18117) );
  AND2_X2 U17122 ( .A1(n19955), .A2(n17725), .ZN(n19268) );
  INV_X1 U17123 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19924) );
  NOR2_X1 U17124 ( .A1(n19183), .A2(n19336), .ZN(n19291) );
  INV_X1 U17125 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17408) );
  OAI211_X1 U17126 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n19337), .A(
        n19291), .B(n17408), .ZN(n13853) );
  OAI21_X1 U17127 ( .B1(n19156), .B2(n19924), .A(n13853), .ZN(n13855) );
  INV_X1 U17128 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n17406) );
  NAND3_X1 U17129 ( .A1(n19323), .A2(n19121), .A3(n17406), .ZN(n19339) );
  AOI21_X1 U17130 ( .B1(n19329), .B2(n19339), .A(n17408), .ZN(n13854) );
  AOI211_X1 U17131 ( .C1(n19050), .C2(n19331), .A(n13855), .B(n13854), .ZN(
        n13856) );
  OAI21_X1 U17132 ( .B1(n19285), .B2(n13857), .A(n13856), .ZN(P3_U2861) );
  NAND2_X1 U17133 ( .A1(n10889), .A2(n10872), .ZN(n13858) );
  INV_X1 U17134 ( .A(DATAI_1_), .ZN(n13860) );
  NAND2_X1 U17135 ( .A1(n15086), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13859) );
  OAI21_X1 U17136 ( .B1(n15086), .B2(n13860), .A(n13859), .ZN(n15134) );
  INV_X1 U17137 ( .A(n15134), .ZN(n13861) );
  INV_X1 U17138 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20965) );
  OAI222_X1 U17139 ( .A1(n15055), .A2(n15160), .B1(n15153), .B2(n13861), .C1(
        n15151), .C2(n20965), .ZN(P1_U2903) );
  INV_X1 U17140 ( .A(DATAI_0_), .ZN(n13863) );
  NAND2_X1 U17141 ( .A1(n15096), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13862) );
  OAI21_X1 U17142 ( .B1(n15086), .B2(n13863), .A(n13862), .ZN(n15141) );
  INV_X1 U17143 ( .A(n15141), .ZN(n13864) );
  INV_X1 U17144 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20970) );
  OAI222_X1 U17145 ( .A1(n14253), .A2(n15160), .B1(n15153), .B2(n13864), .C1(
        n15151), .C2(n20970), .ZN(P1_U2904) );
  NAND2_X1 U17146 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  MUX2_X1 U17147 ( .A(n13869), .B(n15955), .S(n16070), .Z(n13870) );
  OAI21_X1 U17148 ( .B1(n16856), .B2(n16072), .A(n13870), .ZN(P2_U2885) );
  XNOR2_X1 U17149 ( .A(n13872), .B(n13871), .ZN(n13971) );
  INV_X1 U17150 ( .A(n17547), .ZN(n14129) );
  NAND3_X1 U17151 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n13873), .ZN(n13874) );
  OAI211_X1 U17152 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n14129), .A(
        n14464), .B(n13874), .ZN(n13881) );
  NOR2_X1 U17153 ( .A1(n15533), .A2(n14133), .ZN(n13880) );
  INV_X1 U17154 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21498) );
  NAND2_X1 U17155 ( .A1(n13877), .A2(n13876), .ZN(n13878) );
  NAND2_X1 U17156 ( .A1(n13875), .A2(n13878), .ZN(n13936) );
  OAI22_X1 U17157 ( .A1(n20904), .A2(n21498), .B1(n15576), .B2(n13936), .ZN(
        n13879) );
  AOI211_X1 U17158 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13881), .A(
        n13880), .B(n13879), .ZN(n13888) );
  INV_X1 U17159 ( .A(n21003), .ZN(n13884) );
  NAND2_X1 U17160 ( .A1(n13882), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13883) );
  INV_X1 U17161 ( .A(n15535), .ZN(n13886) );
  NAND3_X1 U17162 ( .A1(n13886), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13885), .ZN(n13887) );
  OAI211_X1 U17163 ( .C1(n13971), .C2(n17559), .A(n13888), .B(n13887), .ZN(
        P1_U3029) );
  NOR2_X1 U17164 ( .A1(n16817), .A2(n16070), .ZN(n13894) );
  AOI21_X1 U17165 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n16070), .A(n13894), .ZN(
        n13895) );
  OAI21_X1 U17166 ( .B1(n20751), .B2(n16072), .A(n13895), .ZN(P2_U2884) );
  INV_X1 U17167 ( .A(n18117), .ZN(n17437) );
  INV_X1 U17168 ( .A(n19337), .ZN(n17359) );
  OAI21_X1 U17169 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n17418) );
  INV_X1 U17170 ( .A(n13912), .ZN(n17427) );
  NAND2_X1 U17171 ( .A1(n17418), .A2(n17427), .ZN(n13899) );
  INV_X1 U17172 ( .A(n17415), .ZN(n17416) );
  NAND2_X1 U17173 ( .A1(n17416), .A2(n10426), .ZN(n17426) );
  OAI211_X1 U17174 ( .C1(n13910), .C2(n17359), .A(n13899), .B(n17426), .ZN(
        n19795) );
  NOR2_X1 U17175 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19923), .ZN(n19354) );
  NAND2_X1 U17176 ( .A1(n19943), .A2(n18704), .ZN(n19824) );
  AOI21_X1 U17177 ( .B1(n13900), .B2(n19824), .A(n19941), .ZN(n13901) );
  NAND2_X1 U17178 ( .A1(n19789), .A2(n19944), .ZN(n13908) );
  AOI21_X1 U17179 ( .B1(n14484), .B2(n9870), .A(n16954), .ZN(n13906) );
  OAI211_X1 U17180 ( .C1(n18650), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        n19798) );
  INV_X1 U17181 ( .A(n19798), .ZN(n19809) );
  INV_X1 U17182 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n19342) );
  NAND3_X1 U17183 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19921)
         );
  OAI22_X1 U17184 ( .A1(n19809), .A2(n19830), .B1(n19342), .B2(n19921), .ZN(
        n13909) );
  AOI21_X1 U17185 ( .B1(n17437), .B2(n19795), .A(n17439), .ZN(n13916) );
  NAND2_X1 U17186 ( .A1(n17359), .A2(n17398), .ZN(n17404) );
  AOI22_X1 U17187 ( .A1(n17404), .A2(n13910), .B1(n19787), .B2(n17426), .ZN(
        n13911) );
  NOR2_X1 U17188 ( .A1(n13911), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n19797) );
  NOR2_X1 U17189 ( .A1(n13912), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13913) );
  NOR2_X1 U17190 ( .A1(n9717), .A2(n13913), .ZN(n18070) );
  AOI22_X1 U17191 ( .A1(n19797), .A2(n17437), .B1(n18070), .B2(n19821), .ZN(
        n13914) );
  OAI22_X1 U17192 ( .A1(n13916), .A2(n13915), .B1(n17439), .B2(n13914), .ZN(
        P3_U3285) );
  INV_X1 U17193 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13918) );
  AOI22_X1 U17194 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13917) );
  OAI21_X1 U17195 ( .B1(n13918), .B2(n13930), .A(n13917), .ZN(P1_U2915) );
  AOI22_X1 U17196 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13919) );
  OAI21_X1 U17197 ( .B1(n15132), .B2(n13930), .A(n13919), .ZN(P1_U2919) );
  INV_X1 U17198 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13921) );
  AOI22_X1 U17199 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13920) );
  OAI21_X1 U17200 ( .B1(n13921), .B2(n13930), .A(n13920), .ZN(P1_U2916) );
  INV_X1 U17201 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13923) );
  AOI22_X1 U17202 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13922) );
  OAI21_X1 U17203 ( .B1(n13923), .B2(n13930), .A(n13922), .ZN(P1_U2918) );
  INV_X1 U17204 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U17205 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13924) );
  OAI21_X1 U17206 ( .B1(n13925), .B2(n13930), .A(n13924), .ZN(P1_U2917) );
  AOI22_X1 U17207 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13926) );
  OAI21_X1 U17208 ( .B1(n15137), .B2(n13930), .A(n13926), .ZN(P1_U2920) );
  INV_X1 U17209 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13928) );
  AOI22_X1 U17210 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13927) );
  OAI21_X1 U17211 ( .B1(n13928), .B2(n13930), .A(n13927), .ZN(P1_U2913) );
  INV_X1 U17212 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U17213 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13929) );
  OAI21_X1 U17214 ( .B1(n13931), .B2(n13930), .A(n13929), .ZN(P1_U2914) );
  INV_X1 U17215 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13966) );
  MUX2_X1 U17216 ( .A(n13966), .B(n13933), .S(n13932), .Z(n13935) );
  INV_X1 U17217 ( .A(n13641), .ZN(n13934) );
  NAND2_X1 U17218 ( .A1(n13935), .A2(n13934), .ZN(n14098) );
  OAI21_X1 U17219 ( .B1(n13935), .B2(n13934), .A(n14098), .ZN(n15046) );
  INV_X1 U17220 ( .A(n13936), .ZN(n15044) );
  AOI22_X1 U17221 ( .A1(n20931), .A2(n15044), .B1(n15075), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13937) );
  OAI21_X1 U17222 ( .B1(n15046), .B2(n15079), .A(n13937), .ZN(P1_U2870) );
  AND2_X1 U17223 ( .A1(n13939), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13940) );
  NAND2_X1 U17224 ( .A1(n13938), .A2(n13940), .ZN(n14090) );
  OR2_X1 U17225 ( .A1(n13938), .A2(n13940), .ZN(n13941) );
  NAND2_X1 U17226 ( .A1(n14090), .A2(n13941), .ZN(n20005) );
  OR2_X1 U17227 ( .A1(n13944), .A2(n13943), .ZN(n13945) );
  NAND2_X1 U17228 ( .A1(n13942), .A2(n13945), .ZN(n19986) );
  INV_X1 U17229 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n13946) );
  MUX2_X1 U17230 ( .A(n19986), .B(n13946), .S(n16070), .Z(n13947) );
  OAI21_X1 U17231 ( .B1(n20005), .B2(n16072), .A(n13947), .ZN(P2_U2883) );
  INV_X1 U17232 ( .A(DATAI_2_), .ZN(n13949) );
  NAND2_X1 U17233 ( .A1(n15086), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13948) );
  OAI21_X1 U17234 ( .B1(n15086), .B2(n13949), .A(n13948), .ZN(n15129) );
  INV_X1 U17235 ( .A(n15129), .ZN(n13950) );
  INV_X1 U17236 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20963) );
  OAI222_X1 U17237 ( .A1(n15046), .A2(n15160), .B1(n15153), .B2(n13950), .C1(
        n15151), .C2(n20963), .ZN(P1_U2902) );
  INV_X1 U17238 ( .A(n16192), .ZN(n16851) );
  OR2_X1 U17239 ( .A1(n13954), .A2(n13953), .ZN(n13956) );
  AND2_X1 U17240 ( .A1(n13956), .A2(n13955), .ZN(n17607) );
  NAND2_X1 U17241 ( .A1(n16855), .A2(n17607), .ZN(n20018) );
  OAI211_X1 U17242 ( .C1(n16855), .C2(n17607), .A(n20018), .B(n20020), .ZN(
        n13958) );
  AOI22_X1 U17243 ( .A1(n20016), .A2(n17607), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n16191), .ZN(n13957) );
  OAI211_X1 U17244 ( .C1(n16851), .C2(n20024), .A(n13958), .B(n13957), .ZN(
        P2_U2919) );
  XOR2_X1 U17245 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n14090), .Z(n13964)
         );
  NAND2_X1 U17246 ( .A1(n13942), .A2(n13960), .ZN(n13961) );
  NAND2_X1 U17247 ( .A1(n13959), .A2(n13961), .ZN(n17590) );
  MUX2_X1 U17248 ( .A(n17590), .B(n13962), .S(n16070), .Z(n13963) );
  OAI21_X1 U17249 ( .B1(n13964), .B2(n16072), .A(n13963), .ZN(P2_U2882) );
  INV_X1 U17250 ( .A(n15046), .ZN(n13965) );
  NAND2_X1 U17251 ( .A1(n13965), .A2(n17530), .ZN(n13970) );
  INV_X1 U17252 ( .A(n15041), .ZN(n13968) );
  OAI22_X1 U17253 ( .A1(n17533), .A2(n13966), .B1(n20904), .B2(n21498), .ZN(
        n13967) );
  AOI21_X1 U17254 ( .B1(n17528), .B2(n13968), .A(n13967), .ZN(n13969) );
  OAI211_X1 U17255 ( .C1(n20829), .C2(n13971), .A(n13970), .B(n13969), .ZN(
        P1_U2997) );
  NOR2_X1 U17256 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13446), .ZN(n14016) );
  AND3_X1 U17257 ( .A1(n13351), .A2(n13973), .A3(n13972), .ZN(n13974) );
  NAND2_X1 U17258 ( .A1(n13975), .A2(n13974), .ZN(n15588) );
  INV_X1 U17259 ( .A(n15588), .ZN(n14589) );
  OR2_X1 U17260 ( .A1(n21291), .A2(n14589), .ZN(n13985) );
  NAND2_X1 U17261 ( .A1(n17468), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13976) );
  NAND2_X1 U17262 ( .A1(n17468), .A2(n10880), .ZN(n15585) );
  MUX2_X1 U17263 ( .A(n13976), .B(n15585), .S(n15602), .Z(n13983) );
  NOR2_X1 U17264 ( .A1(n13977), .A2(n15602), .ZN(n14000) );
  NAND2_X1 U17265 ( .A1(n13977), .A2(n15602), .ZN(n13996) );
  INV_X1 U17266 ( .A(n13996), .ZN(n13978) );
  NOR2_X1 U17267 ( .A1(n14000), .A2(n13978), .ZN(n15597) );
  NAND2_X1 U17268 ( .A1(n10871), .A2(n15597), .ZN(n13980) );
  AND2_X1 U17269 ( .A1(n13979), .A2(n13990), .ZN(n14001) );
  OAI22_X1 U17270 ( .A1(n15588), .A2(n13980), .B1(n14001), .B2(n15597), .ZN(
        n13981) );
  INV_X1 U17271 ( .A(n13981), .ZN(n13982) );
  AND2_X1 U17272 ( .A1(n13983), .A2(n13982), .ZN(n13984) );
  NAND2_X1 U17273 ( .A1(n13985), .A2(n13984), .ZN(n15594) );
  OAI21_X1 U17274 ( .B1(n17468), .B2(n13986), .A(n21574), .ZN(n13987) );
  NOR2_X1 U17275 ( .A1(n17497), .A2(n13987), .ZN(n13993) );
  OR2_X1 U17276 ( .A1(n14239), .A2(n14290), .ZN(n13989) );
  OAI211_X1 U17277 ( .C1(n17503), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n13991) );
  MUX2_X1 U17278 ( .A(n15602), .B(n15594), .S(n14595), .Z(n17477) );
  AOI22_X1 U17279 ( .A1(n14016), .A2(n15602), .B1(n17477), .B2(n13446), .ZN(
        n14011) );
  AOI21_X1 U17280 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13996), .A(
        n13995), .ZN(n15605) );
  NOR3_X1 U17281 ( .A1(n15588), .A2(n15605), .A3(n13997), .ZN(n14008) );
  INV_X1 U17282 ( .A(n14000), .ZN(n13999) );
  NAND2_X1 U17283 ( .A1(n17468), .A2(n10746), .ZN(n13998) );
  OAI211_X1 U17284 ( .C1(n14001), .C2(n13999), .A(n15585), .B(n13998), .ZN(
        n14006) );
  NAND2_X1 U17285 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n15602), .ZN(
        n14002) );
  OAI22_X1 U17286 ( .A1(n14003), .A2(n14002), .B1(n14001), .B2(n14000), .ZN(
        n14005) );
  MUX2_X1 U17287 ( .A(n14006), .B(n14005), .S(n14004), .Z(n14007) );
  AOI211_X1 U17288 ( .C1(n21167), .C2(n15588), .A(n14008), .B(n14007), .ZN(
        n15607) );
  INV_X1 U17289 ( .A(n15607), .ZN(n14009) );
  MUX2_X1 U17290 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14009), .S(
        n14595), .Z(n17480) );
  AOI22_X1 U17291 ( .A1(n14016), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n13446), .B2(n17480), .ZN(n14010) );
  NOR2_X1 U17292 ( .A1(n14011), .A2(n14010), .ZN(n17491) );
  INV_X1 U17293 ( .A(n14012), .ZN(n15584) );
  NAND2_X1 U17294 ( .A1(n17491), .A2(n15584), .ZN(n14023) );
  INV_X1 U17295 ( .A(n14275), .ZN(n21290) );
  OR2_X1 U17296 ( .A1(n14013), .A2(n21290), .ZN(n14014) );
  XNOR2_X1 U17297 ( .A(n14014), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20892) );
  NAND2_X1 U17298 ( .A1(n20892), .A2(n17566), .ZN(n14015) );
  MUX2_X1 U17299 ( .A(n17569), .B(n14015), .S(n14595), .Z(n14018) );
  INV_X1 U17300 ( .A(n14016), .ZN(n14017) );
  OAI22_X1 U17301 ( .A1(n14018), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n14017), 
        .B2(n17569), .ZN(n17490) );
  NOR2_X1 U17302 ( .A1(n17490), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14019) );
  NAND2_X1 U17303 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17579), .ZN(n17581) );
  AOI21_X1 U17304 ( .B1(n14023), .B2(n14019), .A(n17581), .ZN(n14020) );
  INV_X1 U17305 ( .A(n17579), .ZN(n14021) );
  NOR2_X1 U17306 ( .A1(n17490), .A2(n14021), .ZN(n14022) );
  NAND2_X1 U17307 ( .A1(n14023), .A2(n14022), .ZN(n17499) );
  INV_X1 U17308 ( .A(n17499), .ZN(n14026) );
  INV_X1 U17309 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21706) );
  NAND2_X1 U17310 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21706), .ZN(n14112) );
  INV_X1 U17311 ( .A(n14112), .ZN(n14024) );
  OAI22_X1 U17312 ( .A1(n14375), .A2(n21418), .B1(n14590), .B2(n14024), .ZN(
        n14025) );
  OAI21_X1 U17313 ( .B1(n14026), .B2(n14025), .A(n21007), .ZN(n14027) );
  OAI21_X1 U17314 ( .B1(n21007), .B2(n21329), .A(n14027), .ZN(P1_U3478) );
  INV_X1 U17315 ( .A(n14028), .ZN(n14029) );
  NAND2_X1 U17316 ( .A1(n13938), .A2(n14029), .ZN(n14217) );
  INV_X1 U17317 ( .A(n14217), .ZN(n14033) );
  INV_X1 U17318 ( .A(n14032), .ZN(n14030) );
  NOR2_X1 U17319 ( .A1(n14217), .A2(n14030), .ZN(n14152) );
  INV_X1 U17320 ( .A(n14152), .ZN(n14031) );
  OAI211_X1 U17321 ( .C1(n14033), .C2(n14032), .A(n14031), .B(n16086), .ZN(
        n14039) );
  INV_X1 U17322 ( .A(n14035), .ZN(n14222) );
  NAND2_X1 U17323 ( .A1(n14222), .A2(n14036), .ZN(n14037) );
  AND2_X1 U17324 ( .A1(n14034), .A2(n14037), .ZN(n16676) );
  NAND2_X1 U17325 ( .A1(n16676), .A2(n16080), .ZN(n14038) );
  OAI211_X1 U17326 ( .C1(n16080), .C2(n14040), .A(n14039), .B(n14038), .ZN(
        P2_U2877) );
  NAND2_X1 U17327 ( .A1(n14042), .A2(n14043), .ZN(n14044) );
  NAND2_X1 U17328 ( .A1(n14041), .A2(n14044), .ZN(n16691) );
  INV_X1 U17329 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n20075) );
  INV_X1 U17330 ( .A(n16124), .ZN(n14045) );
  OAI222_X1 U17331 ( .A1(n16691), .A2(n16213), .B1(n20001), .B2(n20075), .C1(
        n20024), .C2(n14045), .ZN(P2_U2910) );
  NAND2_X1 U17332 ( .A1(n14047), .A2(n14048), .ZN(n14049) );
  AND2_X1 U17333 ( .A1(n14042), .A2(n14049), .ZN(n16704) );
  INV_X1 U17334 ( .A(n16704), .ZN(n15900) );
  INV_X1 U17335 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n20077) );
  INV_X1 U17336 ( .A(n16130), .ZN(n14050) );
  OAI222_X1 U17337 ( .A1(n15900), .A2(n16213), .B1(n20001), .B2(n20077), .C1(
        n20024), .C2(n14050), .ZN(P2_U2911) );
  OR2_X1 U17338 ( .A1(n14052), .A2(n14053), .ZN(n14054) );
  NAND2_X1 U17339 ( .A1(n14085), .A2(n14054), .ZN(n16661) );
  INV_X1 U17340 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n20071) );
  INV_X1 U17341 ( .A(n16108), .ZN(n14055) );
  OAI222_X1 U17342 ( .A1(n16661), .A2(n16213), .B1(n20001), .B2(n20071), .C1(
        n20024), .C2(n14055), .ZN(P2_U2908) );
  OR2_X1 U17343 ( .A1(n14057), .A2(n14056), .ZN(n14058) );
  NAND2_X1 U17344 ( .A1(n14047), .A2(n14058), .ZN(n16715) );
  INV_X1 U17345 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n20079) );
  INV_X1 U17346 ( .A(n16138), .ZN(n16872) );
  OAI222_X1 U17347 ( .A1(n16715), .A2(n16213), .B1(n20079), .B2(n20001), .C1(
        n20024), .C2(n16872), .ZN(P2_U2912) );
  XOR2_X1 U17348 ( .A(n14059), .B(n14060), .Z(n16735) );
  INV_X1 U17349 ( .A(n16735), .ZN(n15922) );
  INV_X1 U17350 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n20081) );
  INV_X1 U17351 ( .A(n16145), .ZN(n20138) );
  OAI222_X1 U17352 ( .A1(n15922), .A2(n16213), .B1(n20081), .B2(n20001), .C1(
        n20024), .C2(n20138), .ZN(P2_U2913) );
  AND2_X1 U17353 ( .A1(n14041), .A2(n14061), .ZN(n14062) );
  NOR2_X1 U17354 ( .A1(n14052), .A2(n14062), .ZN(n16677) );
  INV_X1 U17355 ( .A(n16677), .ZN(n14064) );
  INV_X1 U17356 ( .A(n20024), .ZN(n16210) );
  AOI22_X1 U17357 ( .A1(n16210), .A2(n16116), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n16191), .ZN(n14063) );
  OAI21_X1 U17358 ( .B1(n14064), .B2(n16213), .A(n14063), .ZN(P2_U2909) );
  NOR2_X1 U17359 ( .A1(n14090), .A2(n14065), .ZN(n14215) );
  XNOR2_X1 U17360 ( .A(n14215), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14071) );
  AND2_X1 U17361 ( .A1(n14066), .A2(n14067), .ZN(n14069) );
  OR2_X1 U17362 ( .A1(n14069), .A2(n14068), .ZN(n16719) );
  MUX2_X1 U17363 ( .A(n16719), .B(n11708), .S(n16070), .Z(n14070) );
  OAI21_X1 U17364 ( .B1(n14071), .B2(n16072), .A(n14070), .ZN(P2_U2880) );
  OR2_X1 U17365 ( .A1(n14073), .A2(n14072), .ZN(n14074) );
  NAND2_X1 U17366 ( .A1(n14075), .A2(n14074), .ZN(n20760) );
  XNOR2_X1 U17367 ( .A(n16856), .B(n20760), .ZN(n14079) );
  NOR2_X1 U17368 ( .A1(n20769), .A2(n20772), .ZN(n14076) );
  AOI21_X1 U17369 ( .B1(n20769), .B2(n20772), .A(n14076), .ZN(n20019) );
  NAND2_X1 U17370 ( .A1(n20019), .A2(n20018), .ZN(n20017) );
  INV_X1 U17371 ( .A(n14076), .ZN(n14077) );
  NAND2_X1 U17372 ( .A1(n20017), .A2(n14077), .ZN(n14078) );
  NAND2_X1 U17373 ( .A1(n14079), .A2(n14078), .ZN(n16204) );
  OAI21_X1 U17374 ( .B1(n14079), .B2(n14078), .A(n16204), .ZN(n14080) );
  NAND2_X1 U17375 ( .A1(n14080), .A2(n20020), .ZN(n14083) );
  INV_X1 U17376 ( .A(n16174), .ZN(n20115) );
  INV_X1 U17377 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20090) );
  OAI22_X1 U17378 ( .A1(n20024), .A2(n20115), .B1(n20001), .B2(n20090), .ZN(
        n14081) );
  AOI21_X1 U17379 ( .B1(n20016), .B2(n20760), .A(n14081), .ZN(n14082) );
  NAND2_X1 U17380 ( .A1(n14083), .A2(n14082), .ZN(P2_U2917) );
  NAND2_X1 U17381 ( .A1(n14085), .A2(n14084), .ZN(n14086) );
  AND2_X1 U17382 ( .A1(n13392), .A2(n14086), .ZN(n16651) );
  INV_X1 U17383 ( .A(n16651), .ZN(n14088) );
  AOI22_X1 U17384 ( .A1(n16210), .A2(n16100), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n16191), .ZN(n14087) );
  OAI21_X1 U17385 ( .B1(n14088), .B2(n16213), .A(n14087), .ZN(P2_U2907) );
  NOR2_X1 U17386 ( .A1(n14090), .A2(n14089), .ZN(n14092) );
  INV_X1 U17387 ( .A(n14215), .ZN(n14091) );
  OAI211_X1 U17388 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n14092), .A(
        n14091), .B(n16086), .ZN(n14096) );
  INV_X1 U17389 ( .A(n14066), .ZN(n14093) );
  AOI21_X1 U17390 ( .B1(n14094), .B2(n13959), .A(n14093), .ZN(n16727) );
  NAND2_X1 U17391 ( .A1(n16727), .A2(n16080), .ZN(n14095) );
  OAI211_X1 U17392 ( .C1(n16080), .C2(n11706), .A(n14096), .B(n14095), .ZN(
        P2_U2881) );
  NAND2_X1 U17393 ( .A1(n14098), .A2(n14097), .ZN(n14100) );
  NAND2_X1 U17394 ( .A1(n14100), .A2(n14099), .ZN(n14108) );
  OAI21_X1 U17395 ( .B1(n14100), .B2(n14099), .A(n14108), .ZN(n20916) );
  AOI21_X1 U17396 ( .B1(n13875), .B2(n14102), .A(n14101), .ZN(n20908) );
  AOI22_X1 U17397 ( .A1(n20931), .A2(n20908), .B1(n15075), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n14103) );
  OAI21_X1 U17398 ( .B1(n20916), .B2(n15079), .A(n14103), .ZN(P1_U2869) );
  INV_X1 U17399 ( .A(n14104), .ZN(n14107) );
  AOI21_X1 U17400 ( .B1(n14108), .B2(n14107), .A(n14106), .ZN(n14208) );
  INV_X1 U17401 ( .A(n14208), .ZN(n20899) );
  INV_X1 U17402 ( .A(DATAI_4_), .ZN(n14110) );
  NAND2_X1 U17403 ( .A1(n15086), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14109) );
  OAI21_X1 U17404 ( .B1(n15086), .B2(n14110), .A(n14109), .ZN(n15121) );
  INV_X1 U17405 ( .A(n15121), .ZN(n14111) );
  INV_X1 U17406 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20959) );
  OAI222_X1 U17407 ( .A1(n20899), .A2(n15160), .B1(n15153), .B2(n14111), .C1(
        n20959), .C2(n15151), .ZN(P1_U2900) );
  NAND2_X1 U17408 ( .A1(n21007), .A2(n14112), .ZN(n14740) );
  INV_X1 U17409 ( .A(n21167), .ZN(n14120) );
  INV_X1 U17410 ( .A(n21007), .ZN(n14736) );
  NAND2_X1 U17411 ( .A1(n14736), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14119) );
  AOI21_X1 U17412 ( .B1(n21264), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n14373), 
        .ZN(n14117) );
  OR2_X1 U17413 ( .A1(n14113), .A2(n21173), .ZN(n21201) );
  NAND2_X1 U17414 ( .A1(n14113), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21414) );
  INV_X1 U17415 ( .A(n21414), .ZN(n21075) );
  NAND2_X1 U17416 ( .A1(n21139), .A2(n21075), .ZN(n14280) );
  OAI21_X1 U17417 ( .B1(n21201), .B2(n21415), .A(n14280), .ZN(n14116) );
  OAI211_X1 U17418 ( .C1(n14117), .C2(n14116), .A(n21007), .B(n21420), .ZN(
        n14118) );
  OAI211_X1 U17419 ( .C1(n14740), .C2(n14120), .A(n14119), .B(n14118), .ZN(
        P1_U3475) );
  NOR2_X1 U17420 ( .A1(n14106), .A2(n14122), .ZN(n14123) );
  OR2_X1 U17421 ( .A1(n14121), .A2(n14123), .ZN(n17527) );
  INV_X1 U17422 ( .A(DATAI_5_), .ZN(n14125) );
  NAND2_X1 U17423 ( .A1(n15086), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14124) );
  OAI21_X1 U17424 ( .B1(n15086), .B2(n14125), .A(n14124), .ZN(n15116) );
  INV_X1 U17425 ( .A(n15116), .ZN(n14126) );
  INV_X1 U17426 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20957) );
  OAI222_X1 U17427 ( .A1(n17527), .A2(n15160), .B1(n15153), .B2(n14126), .C1(
        n15151), .C2(n20957), .ZN(P1_U2899) );
  XNOR2_X1 U17428 ( .A(n14200), .B(n14128), .ZN(n14201) );
  OAI21_X1 U17429 ( .B1(n14129), .B2(n14131), .A(n14464), .ZN(n17545) );
  INV_X1 U17430 ( .A(n17545), .ZN(n14130) );
  OAI21_X1 U17431 ( .B1(n15533), .B2(n14133), .A(n14130), .ZN(n14259) );
  INV_X1 U17432 ( .A(n14131), .ZN(n14132) );
  OR2_X1 U17433 ( .A1(n15535), .A2(n14132), .ZN(n14136) );
  INV_X1 U17434 ( .A(n14133), .ZN(n14134) );
  AOI22_X1 U17435 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14259), .B1(
        n17555), .B2(n14128), .ZN(n14139) );
  INV_X1 U17436 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14137) );
  NOR2_X1 U17437 ( .A1(n20904), .A2(n14137), .ZN(n14266) );
  AOI21_X1 U17438 ( .B1(n20998), .B2(n20908), .A(n14266), .ZN(n14138) );
  OAI211_X1 U17439 ( .C1(n17559), .C2(n14269), .A(n14139), .B(n14138), .ZN(
        P1_U3028) );
  OR2_X1 U17440 ( .A1(n14140), .A2(n14141), .ZN(n14142) );
  NAND2_X1 U17441 ( .A1(n13396), .A2(n14142), .ZN(n16648) );
  NAND2_X1 U17442 ( .A1(n14152), .A2(n14151), .ZN(n14150) );
  INV_X1 U17443 ( .A(n14150), .ZN(n14145) );
  OAI211_X1 U17444 ( .C1(n14145), .C2(n14144), .A(n16086), .B(n14143), .ZN(
        n14147) );
  NAND2_X1 U17445 ( .A1(n16078), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n14146) );
  OAI211_X1 U17446 ( .C1(n16648), .C2(n16078), .A(n14147), .B(n14146), .ZN(
        P2_U2875) );
  AND2_X1 U17447 ( .A1(n14034), .A2(n14148), .ZN(n14149) );
  NOR2_X1 U17448 ( .A1(n14140), .A2(n14149), .ZN(n16664) );
  INV_X1 U17449 ( .A(n16664), .ZN(n14155) );
  OAI211_X1 U17450 ( .C1(n14152), .C2(n14151), .A(n14150), .B(n16086), .ZN(
        n14154) );
  NAND2_X1 U17451 ( .A1(n16078), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n14153) );
  OAI211_X1 U17452 ( .C1(n14155), .C2(n16078), .A(n14154), .B(n14153), .ZN(
        P2_U2876) );
  AND2_X1 U17453 ( .A1(n17492), .A2(n21478), .ZN(n14156) );
  INV_X2 U17454 ( .A(n14169), .ZN(n20988) );
  OR2_X1 U17455 ( .A1(n20988), .A2(n11217), .ZN(n14256) );
  INV_X1 U17456 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14162) );
  INV_X1 U17457 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20939) );
  INV_X1 U17458 ( .A(n20980), .ZN(n14161) );
  INV_X1 U17459 ( .A(DATAI_15_), .ZN(n14159) );
  NAND2_X1 U17460 ( .A1(n15096), .A2(BUF1_REG_15__SCAN_IN), .ZN(n14158) );
  OAI21_X1 U17461 ( .B1(n15086), .B2(n14159), .A(n14158), .ZN(n15145) );
  INV_X1 U17462 ( .A(n15145), .ZN(n14160) );
  OAI222_X1 U17463 ( .A1(n14256), .A2(n14162), .B1(n14169), .B2(n20939), .C1(
        n14161), .C2(n14160), .ZN(P1_U2967) );
  INV_X1 U17464 ( .A(DATAI_3_), .ZN(n14164) );
  NAND2_X1 U17465 ( .A1(n15086), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14163) );
  OAI21_X1 U17466 ( .B1(n15086), .B2(n14164), .A(n14163), .ZN(n15124) );
  INV_X1 U17467 ( .A(n15124), .ZN(n14165) );
  INV_X1 U17468 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20961) );
  OAI222_X1 U17469 ( .A1(n20916), .A2(n15160), .B1(n15153), .B2(n14165), .C1(
        n15151), .C2(n20961), .ZN(P1_U2901) );
  INV_X1 U17470 ( .A(DATAI_10_), .ZN(n14167) );
  NAND2_X1 U17471 ( .A1(n15096), .A2(BUF1_REG_10__SCAN_IN), .ZN(n14166) );
  OAI21_X1 U17472 ( .B1(n15086), .B2(n14167), .A(n14166), .ZN(n15157) );
  NAND2_X1 U17473 ( .A1(n20980), .A2(n15157), .ZN(n20984) );
  NAND2_X1 U17474 ( .A1(n20988), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n14168) );
  OAI211_X1 U17475 ( .C1(n21638), .C2(n14256), .A(n20984), .B(n14168), .ZN(
        P1_U2947) );
  AOI22_X1 U17476 ( .A1(n20993), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20988), .ZN(n14170) );
  NAND2_X1 U17477 ( .A1(n20980), .A2(n15124), .ZN(n14184) );
  NAND2_X1 U17478 ( .A1(n14170), .A2(n14184), .ZN(P1_U2955) );
  AOI22_X1 U17479 ( .A1(n20993), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20988), .ZN(n14171) );
  NAND2_X1 U17480 ( .A1(n20980), .A2(n15129), .ZN(n14182) );
  NAND2_X1 U17481 ( .A1(n14171), .A2(n14182), .ZN(P1_U2954) );
  AOI22_X1 U17482 ( .A1(n20993), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20988), .ZN(n14174) );
  INV_X1 U17483 ( .A(DATAI_7_), .ZN(n14173) );
  NAND2_X1 U17484 ( .A1(n15096), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14172) );
  OAI21_X1 U17485 ( .B1(n15086), .B2(n14173), .A(n14172), .ZN(n15108) );
  NAND2_X1 U17486 ( .A1(n20980), .A2(n15108), .ZN(n14196) );
  NAND2_X1 U17487 ( .A1(n14174), .A2(n14196), .ZN(P1_U2944) );
  AOI22_X1 U17488 ( .A1(n20993), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20988), .ZN(n14177) );
  INV_X1 U17489 ( .A(DATAI_6_), .ZN(n14176) );
  NAND2_X1 U17490 ( .A1(n15096), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14175) );
  OAI21_X1 U17491 ( .B1(n15086), .B2(n14176), .A(n14175), .ZN(n15112) );
  NAND2_X1 U17492 ( .A1(n20980), .A2(n15112), .ZN(n14180) );
  NAND2_X1 U17493 ( .A1(n14177), .A2(n14180), .ZN(P1_U2958) );
  AOI22_X1 U17494 ( .A1(n20993), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20988), .ZN(n14178) );
  NAND2_X1 U17495 ( .A1(n20980), .A2(n15121), .ZN(n14192) );
  NAND2_X1 U17496 ( .A1(n14178), .A2(n14192), .ZN(P1_U2956) );
  AOI22_X1 U17497 ( .A1(n20993), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20988), .ZN(n14179) );
  NAND2_X1 U17498 ( .A1(n20980), .A2(n15116), .ZN(n14186) );
  NAND2_X1 U17499 ( .A1(n14179), .A2(n14186), .ZN(P1_U2942) );
  AOI22_X1 U17500 ( .A1(n20993), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20988), .ZN(n14181) );
  NAND2_X1 U17501 ( .A1(n14181), .A2(n14180), .ZN(P1_U2943) );
  AOI22_X1 U17502 ( .A1(n20993), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20988), .ZN(n14183) );
  NAND2_X1 U17503 ( .A1(n14183), .A2(n14182), .ZN(P1_U2939) );
  AOI22_X1 U17504 ( .A1(n20993), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20988), .ZN(n14185) );
  NAND2_X1 U17505 ( .A1(n14185), .A2(n14184), .ZN(P1_U2940) );
  AOI22_X1 U17506 ( .A1(n20993), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20988), .ZN(n14187) );
  NAND2_X1 U17507 ( .A1(n14187), .A2(n14186), .ZN(P1_U2957) );
  AOI22_X1 U17508 ( .A1(n20993), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20988), .ZN(n14188) );
  NAND2_X1 U17509 ( .A1(n20980), .A2(n15134), .ZN(n14194) );
  NAND2_X1 U17510 ( .A1(n14188), .A2(n14194), .ZN(P1_U2938) );
  AOI22_X1 U17511 ( .A1(n20993), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20988), .ZN(n14189) );
  NAND2_X1 U17512 ( .A1(n20980), .A2(n15141), .ZN(n14190) );
  NAND2_X1 U17513 ( .A1(n14189), .A2(n14190), .ZN(P1_U2952) );
  AOI22_X1 U17514 ( .A1(n20993), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20988), .ZN(n14191) );
  NAND2_X1 U17515 ( .A1(n14191), .A2(n14190), .ZN(P1_U2937) );
  AOI22_X1 U17516 ( .A1(n20993), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20988), .ZN(n14193) );
  NAND2_X1 U17517 ( .A1(n14193), .A2(n14192), .ZN(P1_U2941) );
  AOI22_X1 U17518 ( .A1(n20993), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20988), .ZN(n14195) );
  NAND2_X1 U17519 ( .A1(n14195), .A2(n14194), .ZN(P1_U2953) );
  AOI22_X1 U17520 ( .A1(n20993), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20988), .ZN(n14197) );
  NAND2_X1 U17521 ( .A1(n14197), .A2(n14196), .ZN(P1_U2959) );
  AOI22_X1 U17522 ( .A1(n20993), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20988), .ZN(n14199) );
  INV_X1 U17523 ( .A(DATAI_8_), .ZN(n21845) );
  NAND2_X1 U17524 ( .A1(n15096), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14198) );
  OAI21_X1 U17525 ( .B1(n15086), .B2(n21845), .A(n14198), .ZN(n15104) );
  NAND2_X1 U17526 ( .A1(n20980), .A2(n15104), .ZN(n14255) );
  NAND2_X1 U17527 ( .A1(n14199), .A2(n14255), .ZN(P1_U2945) );
  XNOR2_X1 U17528 ( .A(n14202), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n14203) );
  XNOR2_X1 U17529 ( .A(n14204), .B(n14203), .ZN(n14262) );
  INV_X1 U17530 ( .A(n14205), .ZN(n20898) );
  INV_X1 U17531 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21500) );
  NOR2_X1 U17532 ( .A1(n20904), .A2(n21500), .ZN(n14258) );
  AOI21_X1 U17533 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n14258), .ZN(n14206) );
  OAI21_X1 U17534 ( .B1(n20898), .B2(n17524), .A(n14206), .ZN(n14207) );
  AOI21_X1 U17535 ( .B1(n14208), .B2(n17530), .A(n14207), .ZN(n14209) );
  OAI21_X1 U17536 ( .B1(n14262), .B2(n20829), .A(n14209), .ZN(P1_U2995) );
  OR2_X1 U17537 ( .A1(n14101), .A2(n14211), .ZN(n14212) );
  NAND2_X1 U17538 ( .A1(n14210), .A2(n14212), .ZN(n20893) );
  OAI222_X1 U17539 ( .A1(n20893), .A2(n20925), .B1(n20936), .B2(n11238), .C1(
        n15079), .C2(n20899), .ZN(P1_U2868) );
  INV_X1 U17540 ( .A(n16093), .ZN(n14213) );
  INV_X1 U17541 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n21804) );
  OAI222_X1 U17542 ( .A1(n14214), .A2(n16213), .B1(n14213), .B2(n20024), .C1(
        n21804), .C2(n20001), .ZN(P2_U2906) );
  NAND2_X1 U17543 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14342) );
  INV_X1 U17544 ( .A(n14216), .ZN(n14343) );
  NOR2_X1 U17545 ( .A1(n14342), .A2(n14343), .ZN(n14341) );
  OAI211_X1 U17546 ( .C1(n14341), .C2(n14218), .A(n16086), .B(n14217), .ZN(
        n14224) );
  NAND2_X1 U17547 ( .A1(n14219), .A2(n14220), .ZN(n14221) );
  AND2_X1 U17548 ( .A1(n14222), .A2(n14221), .ZN(n16689) );
  NAND2_X1 U17549 ( .A1(n16689), .A2(n16080), .ZN(n14223) );
  OAI211_X1 U17550 ( .C1(n16080), .C2(n11735), .A(n14224), .B(n14223), .ZN(
        P2_U2878) );
  INV_X1 U17551 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14229) );
  AND2_X1 U17552 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20825), .ZN(n14231) );
  NAND2_X1 U17553 ( .A1(n14232), .A2(n14231), .ZN(n14249) );
  OR2_X4 U17554 ( .A1(n15164), .A2(n14249), .ZN(n20851) );
  OAI21_X1 U17555 ( .B1(n10888), .B2(n14240), .A(n20851), .ZN(n20889) );
  NAND2_X1 U17556 ( .A1(n21574), .A2(n21173), .ZN(n14237) );
  INV_X1 U17557 ( .A(n14237), .ZN(n14233) );
  OAI21_X1 U17558 ( .B1(n11217), .B2(n14234), .A(n14233), .ZN(n14243) );
  NOR3_X1 U17559 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(n21706), .ZN(n17573) );
  NAND2_X1 U17560 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17573), .ZN(n14235) );
  NAND2_X1 U17561 ( .A1(n14249), .A2(n14235), .ZN(n14236) );
  NAND2_X1 U17562 ( .A1(n15047), .A2(n15008), .ZN(n20860) );
  AND2_X1 U17563 ( .A1(n11217), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n14241) );
  NAND2_X1 U17564 ( .A1(n14241), .A2(n14237), .ZN(n14238) );
  NOR2_X1 U17565 ( .A1(n20894), .A2(n20996), .ZN(n14248) );
  NOR2_X1 U17566 ( .A1(n14240), .A2(n14239), .ZN(n20913) );
  INV_X1 U17567 ( .A(n20913), .ZN(n20895) );
  INV_X1 U17568 ( .A(n14241), .ZN(n14242) );
  NAND2_X1 U17569 ( .A1(n14243), .A2(n14242), .ZN(n14244) );
  OAI22_X1 U17570 ( .A1(n20895), .A2(n14590), .B1(n20883), .B2(n14246), .ZN(
        n14247) );
  AOI211_X1 U17571 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n20860), .A(n14248), .B(
        n14247), .ZN(n14252) );
  INV_X1 U17572 ( .A(n14249), .ZN(n14250) );
  AND2_X2 U17573 ( .A1(n15164), .A2(n14250), .ZN(n20919) );
  AND2_X2 U17574 ( .A1(n15008), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20912) );
  OAI21_X1 U17575 ( .B1(n20919), .B2(n20912), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14251) );
  OAI211_X1 U17576 ( .C1(n20917), .C2(n14253), .A(n14252), .B(n14251), .ZN(
        P1_U2840) );
  INV_X1 U17577 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20953) );
  NAND2_X1 U17578 ( .A1(n20988), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14254) );
  OAI211_X1 U17579 ( .C1(n20953), .C2(n14256), .A(n14255), .B(n14254), .ZN(
        P1_U2960) );
  NOR2_X1 U17580 ( .A1(n15576), .A2(n20893), .ZN(n14257) );
  AOI211_X1 U17581 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n14259), .A(
        n14258), .B(n14257), .ZN(n14261) );
  OAI211_X1 U17582 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n17555), .B(n17556), .ZN(n14260) );
  OAI211_X1 U17583 ( .C1(n17559), .C2(n14262), .A(n14261), .B(n14260), .ZN(
        P1_U3027) );
  INV_X1 U17584 ( .A(n20916), .ZN(n14263) );
  NAND2_X1 U17585 ( .A1(n14263), .A2(n17530), .ZN(n14268) );
  NOR2_X1 U17586 ( .A1(n17533), .A2(n14264), .ZN(n14265) );
  AOI211_X1 U17587 ( .C1(n17528), .C2(n20920), .A(n14266), .B(n14265), .ZN(
        n14267) );
  OAI211_X1 U17588 ( .C1(n14269), .C2(n20829), .A(n14268), .B(n14267), .ZN(
        P1_U2996) );
  NOR2_X1 U17589 ( .A1(n13391), .A2(n14271), .ZN(n14272) );
  OR2_X1 U17590 ( .A1(n14270), .A2(n14272), .ZN(n16624) );
  AOI22_X1 U17591 ( .A1(n16210), .A2(n14708), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n16191), .ZN(n14273) );
  OAI21_X1 U17592 ( .B1(n16624), .B2(n16213), .A(n14273), .ZN(P2_U2905) );
  NOR2_X2 U17593 ( .A1(n15096), .A2(n15370), .ZN(n14303) );
  AOI22_X1 U17594 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n14304), .B1(DATAI_21_), 
        .B2(n14303), .ZN(n21456) );
  AOI22_X1 U17595 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14304), .B1(DATAI_29_), 
        .B2(n14303), .ZN(n21355) );
  INV_X1 U17596 ( .A(n21355), .ZN(n21453) );
  INV_X1 U17597 ( .A(n21451), .ZN(n21318) );
  OR2_X1 U17598 ( .A1(n21291), .A2(n14275), .ZN(n21110) );
  OR2_X1 U17599 ( .A1(n14590), .A2(n10970), .ZN(n21260) );
  OAI21_X1 U17600 ( .B1(n21110), .B2(n21260), .A(n14308), .ZN(n14278) );
  NOR2_X1 U17601 ( .A1(n21409), .A2(n21136), .ZN(n14412) );
  AOI22_X1 U17602 ( .A1(n14278), .A2(n21420), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14412), .ZN(n14309) );
  NAND2_X1 U17603 ( .A1(n14307), .A2(n14729), .ZN(n14432) );
  OAI22_X1 U17604 ( .A1(n21318), .A2(n14309), .B1(n14308), .B2(n14432), .ZN(
        n14277) );
  AOI21_X1 U17605 ( .B1(n14311), .B2(n21453), .A(n14277), .ZN(n14283) );
  INV_X1 U17606 ( .A(n14278), .ZN(n14279) );
  NAND3_X1 U17607 ( .A1(n14280), .A2(n21420), .A3(n14279), .ZN(n14281) );
  NAND2_X1 U17608 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14282) );
  OAI211_X1 U17609 ( .C1(n21456), .C2(n21178), .A(n14283), .B(n14282), .ZN(
        P1_U3094) );
  AOI22_X1 U17610 ( .A1(DATAI_16_), .A2(n14303), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n14304), .ZN(n21381) );
  AOI22_X1 U17611 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n14304), .B1(DATAI_24_), 
        .B2(n14303), .ZN(n21424) );
  INV_X1 U17612 ( .A(n21424), .ZN(n21378) );
  INV_X1 U17613 ( .A(n21411), .ZN(n21303) );
  NAND2_X1 U17614 ( .A1(n14307), .A2(n11218), .ZN(n14443) );
  OAI22_X1 U17615 ( .A1(n21303), .A2(n14309), .B1(n14308), .B2(n14443), .ZN(
        n14284) );
  AOI21_X1 U17616 ( .B1(n14311), .B2(n21378), .A(n14284), .ZN(n14286) );
  NAND2_X1 U17617 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n14285) );
  OAI211_X1 U17618 ( .C1(n21381), .C2(n21178), .A(n14286), .B(n14285), .ZN(
        P1_U3089) );
  AOI22_X1 U17619 ( .A1(DATAI_17_), .A2(n14303), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n14304), .ZN(n21385) );
  AOI22_X1 U17620 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14304), .B1(DATAI_25_), 
        .B2(n14303), .ZN(n21430) );
  INV_X1 U17621 ( .A(n21430), .ZN(n21382) );
  INV_X1 U17622 ( .A(n21425), .ZN(n21306) );
  NAND2_X1 U17623 ( .A1(n14307), .A2(n11217), .ZN(n14439) );
  OAI22_X1 U17624 ( .A1(n21306), .A2(n14309), .B1(n14308), .B2(n14439), .ZN(
        n14287) );
  AOI21_X1 U17625 ( .B1(n14311), .B2(n21382), .A(n14287), .ZN(n14289) );
  NAND2_X1 U17626 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n14288) );
  OAI211_X1 U17627 ( .C1(n21385), .C2(n21178), .A(n14289), .B(n14288), .ZN(
        P1_U3090) );
  AOI22_X1 U17628 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n14304), .B1(DATAI_18_), 
        .B2(n14303), .ZN(n21436) );
  AOI22_X1 U17629 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14304), .B1(DATAI_26_), 
        .B2(n14303), .ZN(n21347) );
  INV_X1 U17630 ( .A(n21347), .ZN(n21433) );
  INV_X1 U17631 ( .A(n21431), .ZN(n21309) );
  NAND2_X1 U17632 ( .A1(n14307), .A2(n14290), .ZN(n21019) );
  OAI22_X1 U17633 ( .A1(n21309), .A2(n14309), .B1(n14308), .B2(n21019), .ZN(
        n14291) );
  AOI21_X1 U17634 ( .B1(n14311), .B2(n21433), .A(n14291), .ZN(n14293) );
  NAND2_X1 U17635 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14292) );
  OAI211_X1 U17636 ( .C1(n21436), .C2(n21178), .A(n14293), .B(n14292), .ZN(
        P1_U3091) );
  AOI22_X1 U17637 ( .A1(DATAI_22_), .A2(n14303), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n14304), .ZN(n21462) );
  AOI22_X1 U17638 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14304), .B1(DATAI_30_), 
        .B2(n14303), .ZN(n21359) );
  INV_X1 U17639 ( .A(n21359), .ZN(n21459) );
  INV_X1 U17640 ( .A(n21457), .ZN(n21321) );
  NAND2_X1 U17641 ( .A1(n14307), .A2(n10858), .ZN(n21029) );
  OAI22_X1 U17642 ( .A1(n21321), .A2(n14309), .B1(n14308), .B2(n21029), .ZN(
        n14294) );
  AOI21_X1 U17643 ( .B1(n14311), .B2(n21459), .A(n14294), .ZN(n14296) );
  NAND2_X1 U17644 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n14295) );
  OAI211_X1 U17645 ( .C1(n21462), .C2(n21178), .A(n14296), .B(n14295), .ZN(
        P1_U3095) );
  AOI22_X1 U17646 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n14304), .B1(DATAI_23_), 
        .B2(n14303), .ZN(n21473) );
  AOI22_X1 U17647 ( .A1(DATAI_31_), .A2(n14303), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n14304), .ZN(n21367) );
  INV_X1 U17648 ( .A(n21464), .ZN(n21327) );
  NAND2_X1 U17649 ( .A1(n14307), .A2(n10872), .ZN(n14421) );
  OAI22_X1 U17650 ( .A1(n21327), .A2(n14309), .B1(n14308), .B2(n14421), .ZN(
        n14297) );
  AOI21_X1 U17651 ( .B1(n14311), .B2(n21467), .A(n14297), .ZN(n14299) );
  NAND2_X1 U17652 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14298) );
  OAI211_X1 U17653 ( .C1(n21473), .C2(n21178), .A(n14299), .B(n14298), .ZN(
        P1_U3096) );
  AOI22_X1 U17654 ( .A1(DATAI_19_), .A2(n14303), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n14304), .ZN(n21391) );
  AOI22_X1 U17655 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n14304), .B1(DATAI_27_), 
        .B2(n14303), .ZN(n21442) );
  INV_X1 U17656 ( .A(n21442), .ZN(n21388) );
  OAI22_X1 U17657 ( .A1(n21312), .A2(n14309), .B1(n14308), .B2(n21022), .ZN(
        n14300) );
  AOI21_X1 U17658 ( .B1(n14311), .B2(n21388), .A(n14300), .ZN(n14302) );
  NAND2_X1 U17659 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14301) );
  OAI211_X1 U17660 ( .C1(n21391), .C2(n21178), .A(n14302), .B(n14301), .ZN(
        P1_U3092) );
  AOI22_X1 U17661 ( .A1(DATAI_20_), .A2(n14303), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n14304), .ZN(n21395) );
  AOI22_X1 U17662 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n14304), .B1(DATAI_28_), 
        .B2(n14303), .ZN(n21450) );
  INV_X1 U17663 ( .A(n21450), .ZN(n21392) );
  INV_X1 U17664 ( .A(n21443), .ZN(n21315) );
  NAND2_X1 U17665 ( .A1(n14307), .A2(n14306), .ZN(n14428) );
  OAI22_X1 U17666 ( .A1(n21315), .A2(n14309), .B1(n14308), .B2(n14428), .ZN(
        n14310) );
  AOI21_X1 U17667 ( .B1(n14311), .B2(n21392), .A(n14310), .ZN(n14314) );
  NAND2_X1 U17668 ( .A1(n14312), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14313) );
  OAI211_X1 U17669 ( .C1(n21395), .C2(n21178), .A(n14314), .B(n14313), .ZN(
        P1_U3093) );
  INV_X1 U17670 ( .A(n14316), .ZN(n14324) );
  OR2_X1 U17671 ( .A1(n14317), .A2(n14318), .ZN(n16206) );
  NAND2_X1 U17672 ( .A1(n14317), .A2(n14318), .ZN(n14319) );
  NAND2_X1 U17673 ( .A1(n16206), .A2(n14319), .ZN(n16203) );
  NOR2_X1 U17674 ( .A1(n11505), .A2(n16464), .ZN(n14320) );
  AOI21_X1 U17675 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14321), .A(
        n14320), .ZN(n14322) );
  OAI21_X1 U17676 ( .B1(n16763), .B2(n16203), .A(n14322), .ZN(n14323) );
  AOI21_X1 U17677 ( .B1(n14325), .B2(n14324), .A(n14323), .ZN(n14326) );
  OAI21_X1 U17678 ( .B1(n16817), .B2(n16764), .A(n14326), .ZN(n14327) );
  AOI21_X1 U17679 ( .B1(n14332), .B2(n17606), .A(n14327), .ZN(n14328) );
  OAI21_X1 U17680 ( .B1(n10442), .B2(n14334), .A(n14328), .ZN(P2_U3043) );
  AOI22_X1 U17681 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n16754), .ZN(n14329) );
  OAI211_X1 U17682 ( .C1(n15940), .C2(n16448), .A(n14330), .B(n14329), .ZN(
        n14331) );
  AOI21_X1 U17683 ( .B1(n14332), .B2(n16470), .A(n14331), .ZN(n14333) );
  OAI21_X1 U17684 ( .B1(n16472), .B2(n14334), .A(n14333), .ZN(P2_U3011) );
  XOR2_X1 U17685 ( .A(n14121), .B(n14335), .Z(n20878) );
  INV_X1 U17686 ( .A(n20878), .ZN(n14348) );
  XOR2_X1 U17687 ( .A(n17552), .B(n14337), .Z(n20871) );
  AOI22_X1 U17688 ( .A1(n20871), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U17689 ( .B1(n14348), .B2(n15079), .A(n14338), .ZN(P1_U2866) );
  OR2_X1 U17690 ( .A1(n14068), .A2(n14339), .ZN(n14340) );
  NAND2_X1 U17691 ( .A1(n14219), .A2(n14340), .ZN(n16707) );
  NOR2_X1 U17692 ( .A1(n16707), .A2(n16070), .ZN(n14345) );
  AOI211_X1 U17693 ( .C1(n14343), .C2(n14342), .A(n16072), .B(n14341), .ZN(
        n14344) );
  AOI211_X1 U17694 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n16078), .A(n14345), .B(
        n14344), .ZN(n14346) );
  INV_X1 U17695 ( .A(n14346), .ZN(P2_U2879) );
  INV_X1 U17696 ( .A(n15112), .ZN(n14347) );
  OAI222_X1 U17697 ( .A1(n15160), .A2(n14348), .B1(n15153), .B2(n14347), .C1(
        n15151), .C2(n12876), .ZN(P1_U2898) );
  INV_X1 U17698 ( .A(n16632), .ZN(n14349) );
  NAND2_X1 U17699 ( .A1(n14349), .A2(n16080), .ZN(n14354) );
  INV_X1 U17700 ( .A(n14143), .ZN(n14352) );
  OAI211_X1 U17701 ( .C1(n14352), .C2(n10675), .A(n14351), .B(n16086), .ZN(
        n14353) );
  OAI211_X1 U17702 ( .C1(n16080), .C2(n11756), .A(n14354), .B(n14353), .ZN(
        P2_U2874) );
  OAI21_X1 U17703 ( .B1(n14270), .B2(n14356), .A(n14355), .ZN(n16607) );
  INV_X1 U17704 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n20064) );
  INV_X1 U17705 ( .A(n14357), .ZN(n14358) );
  OAI222_X1 U17706 ( .A1(n16607), .A2(n16213), .B1(n20001), .B2(n20064), .C1(
        n14358), .C2(n20024), .ZN(P2_U2904) );
  INV_X1 U17707 ( .A(n14360), .ZN(n14361) );
  AOI21_X1 U17708 ( .B1(n14362), .B2(n14359), .A(n14361), .ZN(n20868) );
  INV_X1 U17709 ( .A(n20868), .ZN(n14372) );
  AOI21_X1 U17710 ( .B1(n14365), .B2(n14364), .A(n14363), .ZN(n20866) );
  AOI22_X1 U17711 ( .A1(n20866), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n14366) );
  OAI21_X1 U17712 ( .B1(n14372), .B2(n15079), .A(n14366), .ZN(P1_U2865) );
  AND2_X1 U17713 ( .A1(n14360), .A2(n14367), .ZN(n14369) );
  OR2_X1 U17714 ( .A1(n14369), .A2(n14368), .ZN(n15036) );
  AOI22_X1 U17715 ( .A1(n15158), .A2(n15104), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15156), .ZN(n14370) );
  OAI21_X1 U17716 ( .B1(n15036), .B2(n15160), .A(n14370), .ZN(P1_U2896) );
  INV_X1 U17717 ( .A(n15108), .ZN(n14371) );
  OAI222_X1 U17718 ( .A1(n14372), .A2(n15160), .B1(n15153), .B2(n14371), .C1(
        n15151), .C2(n12881), .ZN(P1_U2897) );
  INV_X1 U17719 ( .A(n21082), .ZN(n21076) );
  OAI21_X1 U17720 ( .B1(n21055), .B2(n21104), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14376) );
  NAND2_X1 U17721 ( .A1(n14376), .A2(n21420), .ZN(n14385) );
  INV_X1 U17722 ( .A(n21291), .ZN(n14377) );
  OR2_X1 U17723 ( .A1(n21167), .A2(n14377), .ZN(n21079) );
  INV_X1 U17724 ( .A(n21079), .ZN(n21038) );
  NAND2_X1 U17725 ( .A1(n21037), .A2(n10971), .ZN(n14378) );
  NAND2_X1 U17726 ( .A1(n21038), .A2(n21369), .ZN(n14379) );
  OR2_X1 U17727 ( .A1(n21233), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n14410) );
  OR2_X1 U17728 ( .A1(n14380), .A2(n21578), .ZN(n21171) );
  INV_X1 U17729 ( .A(n14379), .ZN(n14384) );
  INV_X1 U17730 ( .A(n14380), .ZN(n14381) );
  NOR2_X1 U17731 ( .A1(n14381), .A2(n21578), .ZN(n21293) );
  NAND2_X1 U17732 ( .A1(n21234), .A2(n21166), .ZN(n21085) );
  NOR3_X2 U17733 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21409), .A3(
        n21085), .ZN(n21069) );
  INV_X1 U17734 ( .A(n21069), .ZN(n14382) );
  AND2_X1 U17735 ( .A1(n14410), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14416) );
  AOI21_X1 U17736 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n14382), .A(n14416), 
        .ZN(n14383) );
  INV_X1 U17737 ( .A(n21395), .ZN(n21445) );
  AOI22_X1 U17738 ( .A1(n21104), .A2(n21445), .B1(n21444), .B2(n21069), .ZN(
        n14386) );
  OAI21_X1 U17739 ( .B1(n21450), .B2(n21074), .A(n14386), .ZN(n14387) );
  AOI21_X1 U17740 ( .B1(n21071), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n14387), .ZN(n14388) );
  OAI21_X1 U17741 ( .B1(n14401), .B2(n21315), .A(n14388), .ZN(P1_U3053) );
  INV_X1 U17742 ( .A(n21473), .ZN(n21362) );
  AOI22_X1 U17743 ( .A1(n21104), .A2(n21362), .B1(n21466), .B2(n21069), .ZN(
        n14389) );
  OAI21_X1 U17744 ( .B1(n21367), .B2(n21074), .A(n14389), .ZN(n14390) );
  AOI21_X1 U17745 ( .B1(n21071), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n14390), .ZN(n14391) );
  OAI21_X1 U17746 ( .B1(n14401), .B2(n21327), .A(n14391), .ZN(P1_U3056) );
  INV_X1 U17747 ( .A(n21456), .ZN(n21352) );
  AOI22_X1 U17748 ( .A1(n21104), .A2(n21352), .B1(n21452), .B2(n21069), .ZN(
        n14392) );
  OAI21_X1 U17749 ( .B1(n21355), .B2(n21074), .A(n14392), .ZN(n14393) );
  AOI21_X1 U17750 ( .B1(n21071), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n14393), .ZN(n14394) );
  OAI21_X1 U17751 ( .B1(n14401), .B2(n21318), .A(n14394), .ZN(P1_U3054) );
  INV_X1 U17752 ( .A(n21381), .ZN(n21421) );
  AOI22_X1 U17753 ( .A1(n21104), .A2(n21421), .B1(n21412), .B2(n21069), .ZN(
        n14395) );
  OAI21_X1 U17754 ( .B1(n21424), .B2(n21074), .A(n14395), .ZN(n14396) );
  AOI21_X1 U17755 ( .B1(n21071), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n14396), .ZN(n14397) );
  OAI21_X1 U17756 ( .B1(n14401), .B2(n21303), .A(n14397), .ZN(P1_U3049) );
  INV_X1 U17757 ( .A(n21385), .ZN(n21427) );
  AOI22_X1 U17758 ( .A1(n21104), .A2(n21427), .B1(n21426), .B2(n21069), .ZN(
        n14398) );
  OAI21_X1 U17759 ( .B1(n21430), .B2(n21074), .A(n14398), .ZN(n14399) );
  AOI21_X1 U17760 ( .B1(n21071), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n14399), .ZN(n14400) );
  OAI21_X1 U17761 ( .B1(n14401), .B2(n21306), .A(n14400), .ZN(P1_U3050) );
  OR2_X1 U17762 ( .A1(n14368), .A2(n14403), .ZN(n14404) );
  NAND2_X1 U17763 ( .A1(n14402), .A2(n14404), .ZN(n20926) );
  INV_X1 U17764 ( .A(DATAI_9_), .ZN(n14406) );
  NAND2_X1 U17765 ( .A1(n15096), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14405) );
  OAI21_X1 U17766 ( .B1(n15096), .B2(n14406), .A(n14405), .ZN(n20971) );
  AOI22_X1 U17767 ( .A1(n15158), .A2(n20971), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15156), .ZN(n14407) );
  OAI21_X1 U17768 ( .B1(n20926), .B2(n15160), .A(n14407), .ZN(P1_U2895) );
  NAND2_X1 U17769 ( .A1(n14449), .A2(n21420), .ZN(n14409) );
  INV_X1 U17770 ( .A(n21339), .ZN(n14408) );
  AND2_X1 U17771 ( .A1(n21420), .A2(n21173), .ZN(n14649) );
  INV_X1 U17772 ( .A(n14649), .ZN(n21288) );
  NOR2_X1 U17773 ( .A1(n21110), .A2(n14378), .ZN(n14415) );
  INV_X1 U17774 ( .A(n14410), .ZN(n14411) );
  INV_X1 U17775 ( .A(n14412), .ZN(n14413) );
  NOR2_X1 U17776 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14413), .ZN(
        n14420) );
  INV_X1 U17777 ( .A(n21171), .ZN(n21228) );
  INV_X1 U17778 ( .A(n14415), .ZN(n14417) );
  AOI21_X1 U17779 ( .B1(n14418), .B2(n14417), .A(n14416), .ZN(n14419) );
  NAND2_X1 U17780 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n14424) );
  INV_X1 U17781 ( .A(n14420), .ZN(n14448) );
  OAI22_X1 U17782 ( .A1(n14449), .A2(n21473), .B1(n14421), .B2(n14448), .ZN(
        n14422) );
  AOI21_X1 U17783 ( .B1(n21160), .B2(n21467), .A(n14422), .ZN(n14423) );
  OAI211_X1 U17784 ( .C1(n14453), .C2(n21327), .A(n14424), .B(n14423), .ZN(
        P1_U3088) );
  NAND2_X1 U17785 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n14427) );
  OAI22_X1 U17786 ( .A1(n14449), .A2(n21391), .B1(n21022), .B2(n14448), .ZN(
        n14425) );
  AOI21_X1 U17787 ( .B1(n21160), .B2(n21388), .A(n14425), .ZN(n14426) );
  OAI211_X1 U17788 ( .C1(n14453), .C2(n21312), .A(n14427), .B(n14426), .ZN(
        P1_U3084) );
  NAND2_X1 U17789 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n14431) );
  OAI22_X1 U17790 ( .A1(n14449), .A2(n21395), .B1(n14428), .B2(n14448), .ZN(
        n14429) );
  AOI21_X1 U17791 ( .B1(n21160), .B2(n21392), .A(n14429), .ZN(n14430) );
  OAI211_X1 U17792 ( .C1(n14453), .C2(n21315), .A(n14431), .B(n14430), .ZN(
        P1_U3085) );
  NAND2_X1 U17793 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n14435) );
  OAI22_X1 U17794 ( .A1(n14449), .A2(n21456), .B1(n14432), .B2(n14448), .ZN(
        n14433) );
  AOI21_X1 U17795 ( .B1(n21160), .B2(n21453), .A(n14433), .ZN(n14434) );
  OAI211_X1 U17796 ( .C1(n14453), .C2(n21318), .A(n14435), .B(n14434), .ZN(
        P1_U3086) );
  NAND2_X1 U17797 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n14438) );
  OAI22_X1 U17798 ( .A1(n14449), .A2(n21462), .B1(n21029), .B2(n14448), .ZN(
        n14436) );
  AOI21_X1 U17799 ( .B1(n21160), .B2(n21459), .A(n14436), .ZN(n14437) );
  OAI211_X1 U17800 ( .C1(n14453), .C2(n21321), .A(n14438), .B(n14437), .ZN(
        P1_U3087) );
  NAND2_X1 U17801 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n14442) );
  OAI22_X1 U17802 ( .A1(n14449), .A2(n21385), .B1(n14439), .B2(n14448), .ZN(
        n14440) );
  AOI21_X1 U17803 ( .B1(n21160), .B2(n21382), .A(n14440), .ZN(n14441) );
  OAI211_X1 U17804 ( .C1(n14453), .C2(n21306), .A(n14442), .B(n14441), .ZN(
        P1_U3082) );
  NAND2_X1 U17805 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n14446) );
  OAI22_X1 U17806 ( .A1(n14449), .A2(n21381), .B1(n14443), .B2(n14448), .ZN(
        n14444) );
  AOI21_X1 U17807 ( .B1(n21160), .B2(n21378), .A(n14444), .ZN(n14445) );
  OAI211_X1 U17808 ( .C1(n14453), .C2(n21303), .A(n14446), .B(n14445), .ZN(
        P1_U3081) );
  NAND2_X1 U17809 ( .A1(n14447), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n14452) );
  OAI22_X1 U17810 ( .A1(n14449), .A2(n21436), .B1(n21019), .B2(n14448), .ZN(
        n14450) );
  AOI21_X1 U17811 ( .B1(n21160), .B2(n21433), .A(n14450), .ZN(n14451) );
  OAI211_X1 U17812 ( .C1(n14453), .C2(n21309), .A(n14452), .B(n14451), .ZN(
        P1_U3083) );
  OR2_X1 U17813 ( .A1(n14363), .A2(n14455), .ZN(n14456) );
  NAND2_X1 U17814 ( .A1(n15574), .A2(n14456), .ZN(n15032) );
  OAI222_X1 U17815 ( .A1(n15032), .A2(n20925), .B1(n20936), .B2(n11256), .C1(
        n15079), .C2(n15036), .ZN(P1_U2864) );
  XNOR2_X1 U17816 ( .A(n14458), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14459) );
  XNOR2_X1 U17817 ( .A(n14457), .B(n14459), .ZN(n14477) );
  NAND2_X1 U17818 ( .A1(n17555), .A2(n14460), .ZN(n17544) );
  INV_X1 U17819 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15558) );
  XNOR2_X1 U17820 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n14461) );
  NOR2_X1 U17821 ( .A1(n17538), .A2(n14461), .ZN(n14471) );
  NAND2_X1 U17822 ( .A1(n17547), .A2(n14462), .ZN(n14463) );
  NAND2_X1 U17823 ( .A1(n14464), .A2(n14463), .ZN(n15560) );
  INV_X1 U17824 ( .A(n15557), .ZN(n14465) );
  NOR2_X1 U17825 ( .A1(n15533), .A2(n14465), .ZN(n17546) );
  INV_X1 U17826 ( .A(n17540), .ZN(n14467) );
  NAND2_X1 U17827 ( .A1(n15477), .A2(n15558), .ZN(n14466) );
  AND2_X1 U17828 ( .A1(n14467), .A2(n14466), .ZN(n17536) );
  INV_X1 U17829 ( .A(n15032), .ZN(n14468) );
  INV_X1 U17830 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21507) );
  NOR2_X1 U17831 ( .A1(n20904), .A2(n21507), .ZN(n14473) );
  AOI21_X1 U17832 ( .B1(n20998), .B2(n14468), .A(n14473), .ZN(n14469) );
  OAI21_X1 U17833 ( .B1(n17536), .B2(n10220), .A(n14469), .ZN(n14470) );
  AOI211_X1 U17834 ( .C1(n14477), .C2(n20999), .A(n14471), .B(n14470), .ZN(
        n14472) );
  INV_X1 U17835 ( .A(n14472), .ZN(P1_U3023) );
  AOI21_X1 U17836 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n14473), .ZN(n14475) );
  OR2_X1 U17837 ( .A1(n17524), .A2(n15029), .ZN(n14474) );
  OAI211_X1 U17838 ( .C1(n15036), .C2(n15370), .A(n14475), .B(n14474), .ZN(
        n14476) );
  AOI21_X1 U17839 ( .B1(n14477), .B2(n17531), .A(n14476), .ZN(n14478) );
  INV_X1 U17840 ( .A(n14478), .ZN(P1_U2991) );
  NOR2_X1 U17841 ( .A1(n14479), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17459) );
  OR2_X1 U17842 ( .A1(n17459), .A2(n17419), .ZN(n19793) );
  NOR2_X1 U17843 ( .A1(n18117), .A2(n19793), .ZN(n14480) );
  MUX2_X1 U17844 ( .A(n14480), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n17439), .Z(P3_U3284) );
  AND2_X1 U17845 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n18122) );
  NAND2_X1 U17846 ( .A1(n9734), .A2(n9725), .ZN(n18495) );
  INV_X1 U17847 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17803) );
  INV_X1 U17848 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17834) );
  INV_X1 U17849 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n18123) );
  INV_X1 U17850 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n21753) );
  INV_X1 U17851 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17906) );
  INV_X1 U17852 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n21674) );
  INV_X1 U17853 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n18067) );
  NAND3_X1 U17854 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18481) );
  NOR3_X1 U17855 ( .A1(n18067), .A2(n18486), .A3(n18481), .ZN(n17457) );
  NAND4_X1 U17856 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n18438) );
  NOR2_X1 U17857 ( .A1(n18375), .A2(n18438), .ZN(n14485) );
  NAND4_X1 U17858 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(n14485), .ZN(n17455) );
  NAND2_X1 U17859 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n18244), .ZN(n18224) );
  NAND2_X1 U17860 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n18181), .ZN(n18172) );
  INV_X1 U17861 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14488) );
  AOI22_X1 U17862 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14487) );
  NAND2_X1 U17863 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n14486) );
  OAI211_X1 U17864 ( .C1(n14488), .C2(n18455), .A(n14487), .B(n14486), .ZN(
        n14494) );
  INV_X1 U17865 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14489) );
  OAI22_X1 U17866 ( .A1(n14490), .A2(n17440), .B1(n10740), .B2(n14489), .ZN(
        n14493) );
  INV_X1 U17867 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n18209) );
  INV_X1 U17868 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14491) );
  OAI22_X1 U17869 ( .A1(n18445), .A2(n18209), .B1(n18285), .B2(n14491), .ZN(
        n14492) );
  OR3_X1 U17870 ( .A1(n14494), .A2(n14493), .A3(n14492), .ZN(n14502) );
  INV_X1 U17871 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14496) );
  AOI22_X1 U17872 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14495) );
  OAI21_X1 U17873 ( .B1(n10739), .B2(n14496), .A(n14495), .ZN(n14497) );
  AOI21_X1 U17874 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(n14497), .ZN(n14500) );
  AOI22_X1 U17875 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14499) );
  AOI22_X1 U17876 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14498) );
  NAND3_X1 U17877 ( .A1(n14500), .A2(n14499), .A3(n14498), .ZN(n14501) );
  NOR2_X1 U17878 ( .A1(n14502), .A2(n14501), .ZN(n14585) );
  INV_X1 U17879 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18380) );
  AOI22_X1 U17880 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14504) );
  NAND2_X1 U17881 ( .A1(n14578), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n14503) );
  OAI211_X1 U17882 ( .C1(n18380), .C2(n18455), .A(n14504), .B(n14503), .ZN(
        n14510) );
  INV_X1 U17883 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14505) );
  INV_X1 U17884 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18387) );
  OAI22_X1 U17885 ( .A1(n14490), .A2(n14505), .B1(n18285), .B2(n18387), .ZN(
        n14509) );
  OAI22_X1 U17886 ( .A1(n10739), .A2(n14507), .B1(n18301), .B2(n14506), .ZN(
        n14508) );
  OR3_X1 U17887 ( .A1(n14510), .A2(n14509), .A3(n14508), .ZN(n14517) );
  INV_X1 U17888 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n18378) );
  INV_X1 U17889 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16978) );
  OAI22_X1 U17890 ( .A1(n9724), .A2(n18378), .B1(n18443), .B2(n16978), .ZN(
        n14511) );
  AOI21_X1 U17891 ( .B1(n18450), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n14511), .ZN(n14515) );
  AOI22_X1 U17892 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14514) );
  AOI22_X1 U17893 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14513) );
  NAND2_X1 U17894 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14512) );
  NAND4_X1 U17895 ( .A1(n14515), .A2(n14514), .A3(n14513), .A4(n14512), .ZN(
        n14516) );
  NOR2_X1 U17896 ( .A1(n14517), .A2(n14516), .ZN(n18174) );
  INV_X1 U17897 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14518) );
  OAI22_X1 U17898 ( .A1(n9724), .A2(n14518), .B1(n18443), .B2(n18284), .ZN(
        n14519) );
  AOI21_X1 U17899 ( .B1(n18450), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n14519), .ZN(n14523) );
  AOI22_X1 U17900 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14522) );
  AOI22_X1 U17901 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U17902 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14520) );
  NAND4_X1 U17903 ( .A1(n14523), .A2(n14522), .A3(n14521), .A4(n14520), .ZN(
        n14534) );
  INV_X1 U17904 ( .A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18422) );
  INV_X1 U17905 ( .A(n14524), .ZN(n18381) );
  AOI22_X1 U17906 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14526) );
  NAND2_X1 U17907 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14525) );
  OAI211_X1 U17908 ( .C1(n18422), .C2(n18381), .A(n14526), .B(n14525), .ZN(
        n14532) );
  INV_X1 U17909 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14528) );
  OAI22_X1 U17910 ( .A1(n9712), .A2(n14528), .B1(n10739), .B2(n14527), .ZN(
        n14531) );
  INV_X1 U17911 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14529) );
  INV_X1 U17912 ( .A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18291) );
  OAI22_X1 U17913 ( .A1(n14490), .A2(n14529), .B1(n18330), .B2(n18291), .ZN(
        n14530) );
  OR3_X1 U17914 ( .A1(n14532), .A2(n14531), .A3(n14530), .ZN(n14533) );
  NOR2_X1 U17915 ( .A1(n14534), .A2(n14533), .ZN(n18183) );
  INV_X1 U17916 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14542) );
  INV_X1 U17917 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n18303) );
  OAI22_X1 U17918 ( .A1(n18443), .A2(n14535), .B1(n13729), .B2(n18303), .ZN(
        n14539) );
  INV_X1 U17919 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14537) );
  INV_X1 U17920 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14536) );
  OAI22_X1 U17921 ( .A1(n9724), .A2(n14537), .B1(n18445), .B2(n14536), .ZN(
        n14538) );
  AOI211_X1 U17922 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n14539), .B(n14538), .ZN(n14541) );
  AOI22_X1 U17923 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14540) );
  OAI211_X1 U17924 ( .C1(n18455), .C2(n14542), .A(n14541), .B(n14540), .ZN(
        n14548) );
  AOI22_X1 U17925 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U17926 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14545) );
  AOI22_X1 U17927 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14544) );
  AOI22_X1 U17928 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14543) );
  NAND4_X1 U17929 ( .A1(n14546), .A2(n14545), .A3(n14544), .A4(n14543), .ZN(
        n14547) );
  OR2_X1 U17930 ( .A1(n14548), .A2(n14547), .ZN(n18188) );
  INV_X1 U17931 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14550) );
  INV_X1 U17932 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14549) );
  OAI22_X1 U17933 ( .A1(n14550), .A2(n18443), .B1(n13729), .B2(n14549), .ZN(
        n14552) );
  INV_X1 U17934 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18319) );
  OAI22_X1 U17935 ( .A1(n18319), .A2(n18445), .B1(n9724), .B2(n18328), .ZN(
        n14551) );
  AOI211_X1 U17936 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n9717), .A(
        n14552), .B(n14551), .ZN(n14554) );
  AOI22_X1 U17937 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14553) );
  OAI211_X1 U17938 ( .C1(n14555), .C2(n18455), .A(n14554), .B(n14553), .ZN(
        n14561) );
  AOI22_X1 U17939 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14559) );
  INV_X1 U17940 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18471) );
  AOI22_X1 U17941 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14558) );
  AOI22_X1 U17942 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18269), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14557) );
  AOI22_X1 U17943 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14556) );
  NAND4_X1 U17944 ( .A1(n14559), .A2(n14558), .A3(n14557), .A4(n14556), .ZN(
        n14560) );
  OR2_X1 U17945 ( .A1(n14561), .A2(n14560), .ZN(n18189) );
  NAND2_X1 U17946 ( .A1(n18188), .A2(n18189), .ZN(n18187) );
  NOR2_X1 U17947 ( .A1(n18183), .A2(n18187), .ZN(n18182) );
  INV_X1 U17948 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16958) );
  INV_X1 U17949 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14562) );
  OAI22_X1 U17950 ( .A1(n18443), .A2(n16958), .B1(n13729), .B2(n14562), .ZN(
        n14564) );
  INV_X1 U17951 ( .A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n18403) );
  OAI22_X1 U17952 ( .A1(n9724), .A2(n18401), .B1(n18445), .B2(n18403), .ZN(
        n14563) );
  AOI211_X1 U17953 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n14564), .B(n14563), .ZN(n14566) );
  AOI22_X1 U17954 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14565) );
  OAI211_X1 U17955 ( .C1(n18455), .C2(n18272), .A(n14566), .B(n14565), .ZN(
        n14572) );
  AOI22_X1 U17956 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14570) );
  AOI22_X1 U17957 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14569) );
  AOI22_X1 U17958 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14568) );
  AOI22_X1 U17959 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14567) );
  NAND4_X1 U17960 ( .A1(n14570), .A2(n14569), .A3(n14568), .A4(n14567), .ZN(
        n14571) );
  OR2_X1 U17961 ( .A1(n14572), .A2(n14571), .ZN(n18179) );
  NAND2_X1 U17962 ( .A1(n18182), .A2(n18179), .ZN(n18178) );
  NOR2_X1 U17963 ( .A1(n18174), .A2(n18178), .ZN(n18173) );
  INV_X1 U17964 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18361) );
  INV_X1 U17965 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16993) );
  INV_X1 U17966 ( .A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n18230) );
  OAI22_X1 U17967 ( .A1(n18443), .A2(n16993), .B1(n13729), .B2(n18230), .ZN(
        n14575) );
  INV_X1 U17968 ( .A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14573) );
  INV_X1 U17969 ( .A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18228) );
  OAI22_X1 U17970 ( .A1(n9724), .A2(n14573), .B1(n18445), .B2(n18228), .ZN(
        n14574) );
  AOI211_X1 U17971 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n14575), .B(n14574), .ZN(n14577) );
  AOI22_X1 U17972 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14576) );
  OAI211_X1 U17973 ( .C1(n18455), .C2(n18361), .A(n14577), .B(n14576), .ZN(
        n14584) );
  AOI22_X1 U17974 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14582) );
  AOI22_X1 U17975 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14581) );
  AOI22_X1 U17976 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14580) );
  AOI22_X1 U17977 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14579) );
  NAND4_X1 U17978 ( .A1(n14582), .A2(n14581), .A3(n14580), .A4(n14579), .ZN(
        n14583) );
  OR2_X1 U17979 ( .A1(n14584), .A2(n14583), .ZN(n18170) );
  NAND2_X1 U17980 ( .A1(n18173), .A2(n18170), .ZN(n18169) );
  NOR2_X1 U17981 ( .A1(n14585), .A2(n18169), .ZN(n18165) );
  AOI21_X1 U17982 ( .B1(n14585), .B2(n18169), .A(n18165), .ZN(n18519) );
  AOI22_X1 U17983 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n18168), .B1(n18519), 
        .B2(n18498), .ZN(n14588) );
  INV_X1 U17984 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14586) );
  NAND3_X1 U17985 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14586), .A3(n10143), 
        .ZN(n14587) );
  NAND2_X1 U17986 ( .A1(n14588), .A2(n14587), .ZN(P3_U2675) );
  OR2_X1 U17987 ( .A1(n14590), .A2(n14589), .ZN(n14593) );
  INV_X1 U17988 ( .A(n15586), .ZN(n14591) );
  NAND2_X1 U17989 ( .A1(n14591), .A2(n10884), .ZN(n14592) );
  NAND2_X1 U17990 ( .A1(n14593), .A2(n14592), .ZN(n17471) );
  OAI22_X1 U17991 ( .A1(n15604), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n13446), .ZN(n14594) );
  AOI21_X1 U17992 ( .B1(n17471), .B2(n17567), .A(n14594), .ZN(n14597) );
  INV_X1 U17993 ( .A(n14595), .ZN(n17473) );
  INV_X1 U17994 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20830) );
  OAI22_X1 U17995 ( .A1(n17473), .A2(n20822), .B1(n17581), .B2(n20830), .ZN(
        n17565) );
  AOI21_X1 U17996 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20825), .A(n17565), 
        .ZN(n15601) );
  AOI21_X1 U17997 ( .B1(n17468), .B2(n17567), .A(n15601), .ZN(n14596) );
  OAI22_X1 U17998 ( .A1(n14597), .A2(n15601), .B1(n14596), .B2(n10884), .ZN(
        P1_U3474) );
  INV_X1 U17999 ( .A(n14601), .ZN(n14602) );
  NAND2_X1 U18000 ( .A1(n14603), .A2(n14602), .ZN(n14604) );
  NAND2_X1 U18001 ( .A1(n14605), .A2(n14604), .ZN(n14609) );
  OR2_X1 U18002 ( .A1(n15626), .A2(n14606), .ZN(n14607) );
  XNOR2_X1 U18003 ( .A(n14607), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14608) );
  XNOR2_X1 U18004 ( .A(n14609), .B(n14608), .ZN(n14640) );
  NAND2_X1 U18005 ( .A1(n14626), .A2(n16470), .ZN(n14617) );
  NAND2_X1 U18006 ( .A1(n12371), .A2(n14610), .ZN(n14611) );
  INV_X1 U18007 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14612) );
  NAND2_X1 U18008 ( .A1(n16754), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U18009 ( .B1(n17599), .B2(n14612), .A(n14631), .ZN(n14613) );
  INV_X1 U18010 ( .A(n14613), .ZN(n14614) );
  OAI21_X1 U18011 ( .B1(n15628), .B2(n16448), .A(n14614), .ZN(n14615) );
  AOI21_X1 U18012 ( .B1(n16003), .B2(n16454), .A(n14615), .ZN(n14616) );
  OAI211_X1 U18013 ( .C1(n14640), .C2(n16472), .A(n14617), .B(n14616), .ZN(
        P2_U2986) );
  NAND2_X1 U18014 ( .A1(n14618), .A2(n16470), .ZN(n14624) );
  NAND2_X1 U18015 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14619) );
  OAI211_X1 U18016 ( .C1(n14621), .C2(n16448), .A(n14620), .B(n14619), .ZN(
        n14622) );
  AOI21_X1 U18017 ( .B1(n15993), .B2(n16454), .A(n14622), .ZN(n14623) );
  OAI211_X1 U18018 ( .C1(n16472), .C2(n14625), .A(n14624), .B(n14623), .ZN(
        P2_U2983) );
  NAND2_X1 U18019 ( .A1(n14626), .A2(n17606), .ZN(n14639) );
  AND2_X1 U18020 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  NOR2_X1 U18021 ( .A1(n15611), .A2(n14629), .ZN(n16105) );
  INV_X1 U18022 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14636) );
  NAND2_X1 U18023 ( .A1(n16003), .A2(n17604), .ZN(n14635) );
  XNOR2_X1 U18024 ( .A(n14630), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14633) );
  INV_X1 U18025 ( .A(n14631), .ZN(n14632) );
  AOI21_X1 U18026 ( .B1(n16486), .B2(n14633), .A(n14632), .ZN(n14634) );
  OAI211_X1 U18027 ( .C1(n16491), .C2(n14636), .A(n14635), .B(n14634), .ZN(
        n14637) );
  AOI21_X1 U18028 ( .B1(n17608), .B2(n16105), .A(n14637), .ZN(n14638) );
  OAI211_X1 U18029 ( .C1(n14640), .C2(n10442), .A(n14639), .B(n14638), .ZN(
        P2_U3018) );
  INV_X1 U18030 ( .A(n15166), .ZN(n14648) );
  AOI22_X1 U18031 ( .A1(n20907), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20912), .ZN(n14645) );
  INV_X1 U18032 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21541) );
  INV_X1 U18033 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21536) );
  INV_X1 U18034 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n21523) );
  NAND4_X1 U18035 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_14__SCAN_IN), .A4(P1_REIP_REG_13__SCAN_IN), .ZN(n14909) );
  NOR2_X1 U18036 ( .A1(n21523), .A2(n14909), .ZN(n14883) );
  NAND4_X1 U18037 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n14883), .A3(
        P1_REIP_REG_19__SCAN_IN), .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n14840) );
  INV_X1 U18038 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21506) );
  NAND4_X1 U18039 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20858)
         );
  NAND2_X1 U18040 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20859) );
  NOR4_X1 U18041 ( .A1(n21507), .A2(n21506), .A3(n20858), .A4(n20859), .ZN(
        n15007) );
  INV_X1 U18042 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21511) );
  INV_X1 U18043 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21509) );
  NOR2_X1 U18044 ( .A1(n21511), .A2(n21509), .ZN(n15011) );
  NAND4_X1 U18045 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(n15007), .A4(n15011), .ZN(n14838) );
  NOR2_X1 U18046 ( .A1(n14840), .A2(n14838), .ZN(n14641) );
  NAND4_X1 U18047 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_21__SCAN_IN), .A4(n14641), .ZN(n14798) );
  NOR2_X1 U18048 ( .A1(n21536), .A2(n14798), .ZN(n14797) );
  NAND2_X1 U18049 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14797), .ZN(n14785) );
  NOR2_X1 U18050 ( .A1(n21541), .A2(n14785), .ZN(n14771) );
  AND2_X1 U18051 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14771), .ZN(n14762) );
  NAND2_X1 U18052 ( .A1(n14762), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14751) );
  INV_X1 U18053 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21546) );
  NOR3_X1 U18054 ( .A1(n14751), .A2(n21550), .A3(n21546), .ZN(n14642) );
  NAND2_X1 U18055 ( .A1(n15008), .A2(n14642), .ZN(n14752) );
  NAND3_X1 U18056 ( .A1(n20860), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14752), 
        .ZN(n14644) );
  NAND3_X1 U18057 ( .A1(n20857), .A2(n14642), .A3(n21548), .ZN(n14643) );
  NAND3_X1 U18058 ( .A1(n14645), .A2(n14644), .A3(n14643), .ZN(n14646) );
  OAI21_X1 U18059 ( .B1(n14648), .B2(n20851), .A(n14647), .ZN(P1_U2809) );
  NAND2_X1 U18060 ( .A1(n14113), .A2(n14649), .ZN(n14650) );
  OAI21_X1 U18061 ( .B1(n21201), .B2(n21418), .A(n14650), .ZN(n21334) );
  NOR2_X1 U18062 ( .A1(n21007), .A2(n21409), .ZN(n14651) );
  AOI21_X1 U18063 ( .B1(n21007), .B2(n21334), .A(n14651), .ZN(n14652) );
  OAI21_X1 U18064 ( .B1(n14378), .B2(n14740), .A(n14652), .ZN(P1_U3477) );
  INV_X1 U18065 ( .A(n14653), .ZN(n14654) );
  XNOR2_X1 U18066 ( .A(n14655), .B(n14654), .ZN(n14675) );
  AND2_X1 U18067 ( .A1(n16754), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14672) );
  AOI21_X1 U18068 ( .B1(n17606), .B2(n14675), .A(n14672), .ZN(n14662) );
  NAND2_X1 U18069 ( .A1(n17608), .A2(n20760), .ZN(n14661) );
  INV_X1 U18070 ( .A(n14656), .ZN(n14659) );
  INV_X1 U18071 ( .A(n14657), .ZN(n14658) );
  NAND2_X1 U18072 ( .A1(n14659), .A2(n14658), .ZN(n14676) );
  NAND3_X1 U18073 ( .A1(n17602), .A2(n14677), .A3(n14676), .ZN(n14660) );
  NAND4_X1 U18074 ( .A1(n14663), .A2(n14662), .A3(n14661), .A4(n14660), .ZN(
        n14669) );
  NAND2_X1 U18075 ( .A1(n14664), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14666) );
  AOI21_X1 U18076 ( .B1(n14667), .B2(n14666), .A(n14665), .ZN(n14668) );
  AOI211_X1 U18077 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n14670), .A(
        n14669), .B(n14668), .ZN(n14671) );
  OAI21_X1 U18078 ( .B1(n13869), .B2(n16764), .A(n14671), .ZN(P2_U3044) );
  AOI21_X1 U18079 ( .B1(n16445), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14672), .ZN(n14673) );
  OAI21_X1 U18080 ( .B1(n16448), .B2(n15952), .A(n14673), .ZN(n14674) );
  AOI21_X1 U18081 ( .B1(n16470), .B2(n14675), .A(n14674), .ZN(n14679) );
  NAND3_X1 U18082 ( .A1(n17587), .A2(n14677), .A3(n14676), .ZN(n14678) );
  OAI211_X1 U18083 ( .C1(n13869), .C2(n17589), .A(n14679), .B(n14678), .ZN(
        P2_U3012) );
  INV_X1 U18084 ( .A(n15609), .ZN(n14680) );
  OAI21_X1 U18085 ( .B1(n15617), .B2(n16221), .A(n19994), .ZN(n14684) );
  NAND2_X1 U18086 ( .A1(n14685), .A2(n15984), .ZN(n14690) );
  INV_X1 U18087 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14687) );
  AOI22_X1 U18088 ( .A1(n19980), .A2(P2_EBX_REG_30__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_30__SCAN_IN), .ZN(n14686) );
  OAI21_X1 U18089 ( .B1(n15968), .B2(n14687), .A(n14686), .ZN(n14688) );
  INV_X1 U18090 ( .A(n14688), .ZN(n14689) );
  NAND2_X1 U18091 ( .A1(n16473), .A2(n12388), .ZN(n14693) );
  OAI211_X1 U18092 ( .C1(n19983), .C2(n16480), .A(n14694), .B(n14693), .ZN(
        P2_U2825) );
  OR2_X1 U18093 ( .A1(n14698), .A2(n14699), .ZN(n14700) );
  NAND2_X1 U18094 ( .A1(n12463), .A2(n14700), .ZN(n16079) );
  INV_X1 U18095 ( .A(n14701), .ZN(n14702) );
  AOI21_X1 U18096 ( .B1(n14703), .B2(n14355), .A(n14702), .ZN(n16199) );
  NAND2_X1 U18097 ( .A1(n16199), .A2(n17608), .ZN(n14704) );
  NAND2_X1 U18098 ( .A1(n16754), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16334) );
  OAI211_X1 U18099 ( .C1(n16764), .C2(n16079), .A(n14704), .B(n16334), .ZN(
        n14705) );
  INV_X1 U18100 ( .A(n16194), .ZN(n14714) );
  INV_X1 U18101 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14713) );
  INV_X1 U18102 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14710) );
  AOI22_X1 U18103 ( .A1(n16193), .A2(n14708), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n16191), .ZN(n14709) );
  OAI21_X1 U18104 ( .B1(n14710), .B2(n16197), .A(n14709), .ZN(n14711) );
  INV_X1 U18105 ( .A(n14711), .ZN(n14712) );
  OAI21_X1 U18106 ( .B1(n14714), .B2(n14713), .A(n14712), .ZN(n14715) );
  INV_X1 U18107 ( .A(n14717), .ZN(n14718) );
  OAI21_X1 U18108 ( .B1(n14719), .B2(n16202), .A(n14718), .ZN(P2_U2889) );
  INV_X1 U18109 ( .A(n15008), .ZN(n20856) );
  OAI21_X1 U18110 ( .B1(n20856), .B2(n14751), .A(n20860), .ZN(n14764) );
  AOI22_X1 U18111 ( .A1(n20907), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20912), .ZN(n14721) );
  OR3_X1 U18112 ( .A1(n15047), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14751), .ZN(
        n14720) );
  OAI211_X1 U18113 ( .C1(n14764), .C2(n21546), .A(n14721), .B(n14720), .ZN(
        n14726) );
  AND2_X1 U18114 ( .A1(n14759), .A2(n14722), .ZN(n14723) );
  NOR2_X1 U18115 ( .A1(n14741), .A2(n20894), .ZN(n14725) );
  OAI21_X1 U18116 ( .B1(n14742), .B2(n20851), .A(n14728), .ZN(P1_U2811) );
  AOI22_X1 U18117 ( .A1(n15128), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n15156), .ZN(n14735) );
  NOR3_X1 U18118 ( .A1(n15156), .A2(n14730), .A3(n14729), .ZN(n14731) );
  INV_X1 U18119 ( .A(DATAI_13_), .ZN(n14733) );
  NAND2_X1 U18120 ( .A1(n15096), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14732) );
  OAI21_X1 U18121 ( .B1(n15096), .B2(n14733), .A(n14732), .ZN(n20977) );
  AOI22_X1 U18122 ( .A1(n15142), .A2(n20977), .B1(n15140), .B2(DATAI_29_), 
        .ZN(n14734) );
  OAI211_X1 U18123 ( .C1(n14742), .C2(n15160), .A(n14735), .B(n14734), .ZN(
        P1_U2875) );
  NAND2_X1 U18124 ( .A1(n14736), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14739) );
  XNOR2_X1 U18125 ( .A(n9746), .B(n21414), .ZN(n14737) );
  NAND3_X1 U18126 ( .A1(n21007), .A2(n21420), .A3(n14737), .ZN(n14738) );
  OAI211_X1 U18127 ( .C1(n14740), .C2(n21291), .A(n14739), .B(n14738), .ZN(
        P1_U3476) );
  OAI222_X1 U18128 ( .A1(n14743), .A2(n20936), .B1(n20925), .B2(n14741), .C1(
        n14742), .C2(n15079), .ZN(P1_U2843) );
  OR2_X1 U18129 ( .A1(n14744), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14747) );
  INV_X1 U18130 ( .A(n14745), .ZN(n14746) );
  MUX2_X1 U18131 ( .A(n14747), .B(n14746), .S(n21572), .Z(P1_U3487) );
  AOI21_X1 U18132 ( .B1(n14749), .B2(n13345), .A(n14748), .ZN(n14750) );
  INV_X1 U18133 ( .A(n14750), .ZN(n15173) );
  AOI22_X1 U18134 ( .A1(n20907), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20912), .ZN(n14755) );
  NOR3_X1 U18135 ( .A1(n15047), .A2(n14751), .A3(n21546), .ZN(n14753) );
  OAI211_X1 U18136 ( .C1(n14753), .C2(P1_REIP_REG_30__SCAN_IN), .A(n20860), 
        .B(n14752), .ZN(n14754) );
  OAI211_X1 U18137 ( .C1(n20897), .C2(n15169), .A(n14755), .B(n14754), .ZN(
        n14756) );
  AOI21_X1 U18138 ( .B1(n15059), .B2(n20909), .A(n14756), .ZN(n14757) );
  OAI21_X1 U18139 ( .B1(n15173), .B2(n20851), .A(n14757), .ZN(P1_U2810) );
  AOI21_X1 U18140 ( .B1(n14758), .B2(n9772), .A(n13304), .ZN(n15185) );
  INV_X1 U18141 ( .A(n15185), .ZN(n15093) );
  INV_X1 U18142 ( .A(n14759), .ZN(n14760) );
  AOI21_X1 U18143 ( .B1(n14761), .B2(n14776), .A(n14760), .ZN(n15384) );
  NOR2_X1 U18144 ( .A1(n20897), .A2(n15183), .ZN(n14767) );
  AOI21_X1 U18145 ( .B1(n20857), .B2(n14762), .A(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14765) );
  AOI22_X1 U18146 ( .A1(n20907), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20912), .ZN(n14763) );
  OAI21_X1 U18147 ( .B1(n14765), .B2(n14764), .A(n14763), .ZN(n14766) );
  AOI211_X1 U18148 ( .C1(n15384), .C2(n20909), .A(n14767), .B(n14766), .ZN(
        n14768) );
  OAI21_X1 U18149 ( .B1(n15093), .B2(n20851), .A(n14768), .ZN(P1_U2812) );
  OAI21_X1 U18150 ( .B1(n14769), .B2(n14770), .A(n9772), .ZN(n15196) );
  NOR2_X1 U18151 ( .A1(n15047), .A2(n14771), .ZN(n14787) );
  NOR2_X1 U18152 ( .A1(n14787), .A2(n20856), .ZN(n14790) );
  INV_X1 U18153 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21542) );
  AOI22_X1 U18154 ( .A1(n20907), .A2(P1_EBX_REG_27__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20912), .ZN(n14773) );
  NAND3_X1 U18155 ( .A1(n20857), .A2(n21542), .A3(n14771), .ZN(n14772) );
  OAI211_X1 U18156 ( .C1(n14790), .C2(n21542), .A(n14773), .B(n14772), .ZN(
        n14774) );
  AOI21_X1 U18157 ( .B1(n20919), .B2(n15189), .A(n14774), .ZN(n14780) );
  INV_X1 U18158 ( .A(n14776), .ZN(n14777) );
  AOI21_X1 U18159 ( .B1(n14778), .B2(n14775), .A(n14777), .ZN(n15388) );
  NAND2_X1 U18160 ( .A1(n15388), .A2(n20909), .ZN(n14779) );
  OAI211_X1 U18161 ( .C1(n15196), .C2(n20851), .A(n14780), .B(n14779), .ZN(
        P1_U2813) );
  OAI21_X1 U18162 ( .B1(n14781), .B2(n14782), .A(n14775), .ZN(n15397) );
  AOI21_X1 U18163 ( .B1(n14784), .B2(n14783), .A(n14769), .ZN(n15204) );
  NAND2_X1 U18164 ( .A1(n15204), .A2(n20879), .ZN(n14794) );
  INV_X1 U18165 ( .A(n15202), .ZN(n14792) );
  AOI22_X1 U18166 ( .A1(n20907), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20912), .ZN(n14789) );
  INV_X1 U18167 ( .A(n14785), .ZN(n14786) );
  NAND2_X1 U18168 ( .A1(n14787), .A2(n14786), .ZN(n14788) );
  OAI211_X1 U18169 ( .C1(n14790), .C2(n21541), .A(n14789), .B(n14788), .ZN(
        n14791) );
  AOI21_X1 U18170 ( .B1(n20919), .B2(n14792), .A(n14791), .ZN(n14793) );
  OAI211_X1 U18171 ( .C1(n15397), .C2(n20894), .A(n14794), .B(n14793), .ZN(
        P1_U2814) );
  OAI21_X1 U18172 ( .B1(n14795), .B2(n14796), .A(n14783), .ZN(n15215) );
  INV_X1 U18173 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21537) );
  AOI22_X1 U18174 ( .A1(n14797), .A2(n21537), .B1(P1_REIP_REG_25__SCAN_IN), 
        .B2(n21536), .ZN(n14801) );
  INV_X1 U18175 ( .A(n14798), .ZN(n14812) );
  OAI21_X1 U18176 ( .B1(n15047), .B2(n14812), .A(n15008), .ZN(n14811) );
  NAND2_X1 U18177 ( .A1(n14811), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U18178 ( .A1(n20907), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20912), .ZN(n14799) );
  OAI211_X1 U18179 ( .C1(n14801), .C2(n15047), .A(n14800), .B(n14799), .ZN(
        n14805) );
  AND2_X1 U18180 ( .A1(n14807), .A2(n14802), .ZN(n14803) );
  OR2_X1 U18181 ( .A1(n14781), .A2(n14803), .ZN(n15415) );
  NOR2_X1 U18182 ( .A1(n15415), .A2(n20894), .ZN(n14804) );
  AOI211_X1 U18183 ( .C1(n20919), .C2(n15208), .A(n14805), .B(n14804), .ZN(
        n14806) );
  OAI21_X1 U18184 ( .B1(n15215), .B2(n20851), .A(n14806), .ZN(P1_U2815) );
  OAI21_X1 U18185 ( .B1(n14821), .B2(n14808), .A(n14807), .ZN(n15416) );
  AOI21_X1 U18186 ( .B1(n14810), .B2(n14809), .A(n14795), .ZN(n15224) );
  NAND2_X1 U18187 ( .A1(n15224), .A2(n20879), .ZN(n14818) );
  INV_X1 U18188 ( .A(n15222), .ZN(n14816) );
  INV_X1 U18189 ( .A(n14811), .ZN(n14826) );
  AOI22_X1 U18190 ( .A1(n20907), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20912), .ZN(n14814) );
  NAND3_X1 U18191 ( .A1(n20857), .A2(n14812), .A3(n21536), .ZN(n14813) );
  OAI211_X1 U18192 ( .C1(n14826), .C2(n21536), .A(n14814), .B(n14813), .ZN(
        n14815) );
  AOI21_X1 U18193 ( .B1(n20919), .B2(n14816), .A(n14815), .ZN(n14817) );
  OAI211_X1 U18194 ( .C1(n15416), .C2(n20894), .A(n14818), .B(n14817), .ZN(
        P1_U2816) );
  NOR2_X1 U18195 ( .A1(n14836), .A2(n14819), .ZN(n14820) );
  OR2_X1 U18196 ( .A1(n14821), .A2(n14820), .ZN(n15431) );
  INV_X1 U18197 ( .A(n14809), .ZN(n14823) );
  AOI21_X1 U18198 ( .B1(n14824), .B2(n10697), .A(n14823), .ZN(n15231) );
  NAND2_X1 U18199 ( .A1(n15231), .A2(n20879), .ZN(n14832) );
  NOR2_X1 U18200 ( .A1(n15047), .A2(n14838), .ZN(n14973) );
  INV_X1 U18201 ( .A(n14840), .ZN(n14855) );
  AND2_X1 U18202 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n14855), .ZN(n14825) );
  NAND2_X1 U18203 ( .A1(n14973), .A2(n14825), .ZN(n14843) );
  INV_X1 U18204 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21532) );
  OR2_X1 U18205 ( .A1(n14843), .A2(n21532), .ZN(n14828) );
  INV_X1 U18206 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14827) );
  AOI21_X1 U18207 ( .B1(n14828), .B2(n14827), .A(n14826), .ZN(n14830) );
  INV_X1 U18208 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15066) );
  INV_X1 U18209 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15229) );
  OAI22_X1 U18210 ( .A1(n20883), .A2(n15066), .B1(n20882), .B2(n15229), .ZN(
        n14829) );
  AOI211_X1 U18211 ( .C1(n20919), .C2(n15227), .A(n14830), .B(n14829), .ZN(
        n14831) );
  OAI211_X1 U18212 ( .C1(n15431), .C2(n20894), .A(n14832), .B(n14831), .ZN(
        P1_U2817) );
  AOI21_X1 U18213 ( .B1(n14834), .B2(n14833), .A(n14822), .ZN(n15239) );
  INV_X1 U18214 ( .A(n15239), .ZN(n15115) );
  AOI21_X1 U18215 ( .B1(n14837), .B2(n14851), .A(n14836), .ZN(n15440) );
  INV_X1 U18216 ( .A(n14838), .ZN(n14839) );
  NAND2_X1 U18217 ( .A1(n15008), .A2(n14839), .ZN(n14920) );
  OR2_X1 U18218 ( .A1(n14920), .A2(n14840), .ZN(n14841) );
  NAND2_X1 U18219 ( .A1(n20860), .A2(n14841), .ZN(n14870) );
  OAI21_X1 U18220 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n15047), .A(n14870), 
        .ZN(n14845) );
  AOI22_X1 U18221 ( .A1(n20907), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20912), .ZN(n14842) );
  OAI21_X1 U18222 ( .B1(n14843), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14842), 
        .ZN(n14844) );
  AOI21_X1 U18223 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n14845), .A(n14844), 
        .ZN(n14846) );
  OAI21_X1 U18224 ( .B1(n20897), .B2(n15237), .A(n14846), .ZN(n14847) );
  AOI21_X1 U18225 ( .B1(n15440), .B2(n20909), .A(n14847), .ZN(n14848) );
  OAI21_X1 U18226 ( .B1(n15115), .B2(n20851), .A(n14848), .ZN(P1_U2818) );
  INV_X1 U18227 ( .A(n14849), .ZN(n14867) );
  INV_X1 U18228 ( .A(n14850), .ZN(n14852) );
  OAI21_X1 U18229 ( .B1(n14867), .B2(n14852), .A(n14851), .ZN(n15444) );
  XOR2_X1 U18230 ( .A(n14854), .B(n14853), .Z(n15251) );
  NAND2_X1 U18231 ( .A1(n15251), .A2(n20879), .ZN(n14861) );
  INV_X1 U18232 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14858) );
  NAND3_X1 U18233 ( .A1(n14973), .A2(n14858), .A3(n14855), .ZN(n14857) );
  AOI22_X1 U18234 ( .A1(n20907), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20912), .ZN(n14856) );
  OAI211_X1 U18235 ( .C1(n14870), .C2(n14858), .A(n14857), .B(n14856), .ZN(
        n14859) );
  AOI21_X1 U18236 ( .B1(n20919), .B2(n15247), .A(n14859), .ZN(n14860) );
  OAI211_X1 U18237 ( .C1(n15444), .C2(n20894), .A(n14861), .B(n14860), .ZN(
        P1_U2819) );
  INV_X1 U18238 ( .A(n14853), .ZN(n14864) );
  OAI21_X1 U18239 ( .B1(n14865), .B2(n14863), .A(n14864), .ZN(n15261) );
  INV_X1 U18240 ( .A(n14866), .ZN(n14869) );
  INV_X1 U18241 ( .A(n14877), .ZN(n14868) );
  AOI21_X1 U18242 ( .B1(n14869), .B2(n14868), .A(n14867), .ZN(n15452) );
  AND2_X1 U18243 ( .A1(n14973), .A2(n14883), .ZN(n14895) );
  INV_X1 U18244 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21771) );
  INV_X1 U18245 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21526) );
  NOR2_X1 U18246 ( .A1(n21771), .A2(n21526), .ZN(n14879) );
  AOI21_X1 U18247 ( .B1(n14895), .B2(n14879), .A(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14871) );
  NOR2_X1 U18248 ( .A1(n14871), .A2(n14870), .ZN(n14874) );
  AOI22_X1 U18249 ( .A1(n20907), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20912), .ZN(n14872) );
  OAI21_X1 U18250 ( .B1(n20897), .B2(n15254), .A(n14872), .ZN(n14873) );
  AOI211_X1 U18251 ( .C1(n15452), .C2(n20909), .A(n14874), .B(n14873), .ZN(
        n14875) );
  OAI21_X1 U18252 ( .B1(n15261), .B2(n20851), .A(n14875), .ZN(P1_U2820) );
  AOI21_X1 U18253 ( .B1(n14876), .B2(n9822), .A(n14863), .ZN(n15269) );
  INV_X1 U18254 ( .A(n15269), .ZN(n15127) );
  AOI21_X1 U18255 ( .B1(n14878), .B2(n14892), .A(n14877), .ZN(n15468) );
  INV_X1 U18256 ( .A(n15265), .ZN(n14886) );
  AOI21_X1 U18257 ( .B1(n21771), .B2(n21526), .A(n14879), .ZN(n14882) );
  INV_X1 U18258 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15267) );
  NAND2_X1 U18259 ( .A1(n20907), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n14880) );
  OAI211_X1 U18260 ( .C1(n20882), .C2(n15267), .A(n14880), .B(n20904), .ZN(
        n14881) );
  AOI21_X1 U18261 ( .B1(n14895), .B2(n14882), .A(n14881), .ZN(n14885) );
  INV_X1 U18262 ( .A(n20860), .ZN(n15012) );
  NAND2_X1 U18263 ( .A1(n20860), .A2(n14920), .ZN(n14970) );
  OAI21_X1 U18264 ( .B1(n15012), .B2(n14883), .A(n14970), .ZN(n14910) );
  NAND2_X1 U18265 ( .A1(n14910), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14884) );
  OAI211_X1 U18266 ( .C1(n20897), .C2(n14886), .A(n14885), .B(n14884), .ZN(
        n14887) );
  AOI21_X1 U18267 ( .B1(n15468), .B2(n20909), .A(n14887), .ZN(n14888) );
  OAI21_X1 U18268 ( .B1(n15127), .B2(n20851), .A(n14888), .ZN(P1_U2821) );
  INV_X1 U18269 ( .A(n14889), .ZN(n14890) );
  OAI21_X1 U18270 ( .B1(n14890), .B2(n9899), .A(n9822), .ZN(n15276) );
  INV_X1 U18271 ( .A(n14892), .ZN(n14893) );
  AOI21_X1 U18272 ( .B1(n14894), .B2(n14891), .A(n14893), .ZN(n15471) );
  INV_X1 U18273 ( .A(n14895), .ZN(n14898) );
  AOI21_X1 U18274 ( .B1(n20912), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17539), .ZN(n14897) );
  NAND2_X1 U18275 ( .A1(n20907), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14896) );
  OAI211_X1 U18276 ( .C1(n14898), .C2(P1_REIP_REG_18__SCAN_IN), .A(n14897), 
        .B(n14896), .ZN(n14899) );
  AOI21_X1 U18277 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n14910), .A(n14899), 
        .ZN(n14900) );
  OAI21_X1 U18278 ( .B1(n20897), .B2(n15271), .A(n14900), .ZN(n14901) );
  AOI21_X1 U18279 ( .B1(n15471), .B2(n20909), .A(n14901), .ZN(n14902) );
  OAI21_X1 U18280 ( .B1(n15276), .B2(n20851), .A(n14902), .ZN(P1_U2822) );
  OAI21_X1 U18281 ( .B1(n14903), .B2(n14904), .A(n14889), .ZN(n15285) );
  INV_X1 U18282 ( .A(n14891), .ZN(n14905) );
  AOI21_X1 U18283 ( .B1(n14906), .B2(n14918), .A(n14905), .ZN(n15494) );
  OAI21_X1 U18284 ( .B1(n20882), .B2(n14907), .A(n20904), .ZN(n14908) );
  AOI21_X1 U18285 ( .B1(n20907), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14908), .ZN(
        n14913) );
  INV_X1 U18286 ( .A(n14973), .ZN(n14953) );
  NOR2_X1 U18287 ( .A1(n14953), .A2(n14909), .ZN(n14911) );
  OAI21_X1 U18288 ( .B1(n14911), .B2(P1_REIP_REG_17__SCAN_IN), .A(n14910), 
        .ZN(n14912) );
  OAI211_X1 U18289 ( .C1(n20897), .C2(n15287), .A(n14913), .B(n14912), .ZN(
        n14914) );
  AOI21_X1 U18290 ( .B1(n15494), .B2(n20909), .A(n14914), .ZN(n14915) );
  OAI21_X1 U18291 ( .B1(n15285), .B2(n20851), .A(n14915), .ZN(P1_U2823) );
  INV_X1 U18292 ( .A(n14903), .ZN(n14916) );
  OAI21_X1 U18293 ( .B1(n14917), .B2(n9798), .A(n14916), .ZN(n15300) );
  OAI21_X1 U18294 ( .B1(n14933), .B2(n14919), .A(n14918), .ZN(n15501) );
  INV_X1 U18295 ( .A(n15501), .ZN(n14929) );
  INV_X1 U18296 ( .A(n15297), .ZN(n14927) );
  NAND3_X1 U18297 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14923) );
  OR2_X1 U18298 ( .A1(n14920), .A2(n14923), .ZN(n14921) );
  AND2_X1 U18299 ( .A1(n20860), .A2(n14921), .ZN(n14942) );
  INV_X1 U18300 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15073) );
  AOI21_X1 U18301 ( .B1(n20912), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17539), .ZN(n14922) );
  OAI21_X1 U18302 ( .B1(n20883), .B2(n15073), .A(n14922), .ZN(n14925) );
  NOR3_X1 U18303 ( .A1(n14953), .A2(P1_REIP_REG_16__SCAN_IN), .A3(n14923), 
        .ZN(n14924) );
  AOI211_X1 U18304 ( .C1(n14942), .C2(P1_REIP_REG_16__SCAN_IN), .A(n14925), 
        .B(n14924), .ZN(n14926) );
  OAI21_X1 U18305 ( .B1(n20897), .B2(n14927), .A(n14926), .ZN(n14928) );
  AOI21_X1 U18306 ( .B1(n20909), .B2(n14929), .A(n14928), .ZN(n14930) );
  OAI21_X1 U18307 ( .B1(n15300), .B2(n20851), .A(n14930), .ZN(P1_U2824) );
  NOR2_X1 U18308 ( .A1(n14948), .A2(n14931), .ZN(n14932) );
  OR2_X1 U18309 ( .A1(n14933), .A2(n14932), .ZN(n15508) );
  INV_X1 U18310 ( .A(n14961), .ZN(n14996) );
  INV_X1 U18311 ( .A(n14935), .ZN(n14959) );
  OR2_X1 U18312 ( .A1(n14963), .A2(n14947), .ZN(n14945) );
  NAND2_X1 U18313 ( .A1(n15310), .A2(n20879), .ZN(n14944) );
  NAND2_X1 U18314 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14937) );
  INV_X1 U18315 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21520) );
  OAI21_X1 U18316 ( .B1(n14953), .B2(n14937), .A(n21520), .ZN(n14941) );
  INV_X1 U18317 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15074) );
  NAND2_X1 U18318 ( .A1(n20912), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14938) );
  OAI211_X1 U18319 ( .C1(n20883), .C2(n15074), .A(n20904), .B(n14938), .ZN(
        n14940) );
  NOR2_X1 U18320 ( .A1(n20897), .A2(n15308), .ZN(n14939) );
  AOI211_X1 U18321 ( .C1(n14942), .C2(n14941), .A(n14940), .B(n14939), .ZN(
        n14943) );
  OAI211_X1 U18322 ( .C1(n15508), .C2(n20894), .A(n14944), .B(n14943), .ZN(
        P1_U2825) );
  INV_X1 U18323 ( .A(n14945), .ZN(n14946) );
  AOI21_X1 U18324 ( .B1(n14947), .B2(n14963), .A(n14946), .ZN(n15321) );
  INV_X1 U18325 ( .A(n15321), .ZN(n15149) );
  AOI21_X1 U18326 ( .B1(n14949), .B2(n14968), .A(n14948), .ZN(n15513) );
  INV_X1 U18327 ( .A(n14970), .ZN(n14987) );
  NAND2_X1 U18328 ( .A1(n20907), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14950) );
  OAI211_X1 U18329 ( .C1(n20882), .C2(n14951), .A(n14950), .B(n20904), .ZN(
        n14952) );
  AOI21_X1 U18330 ( .B1(n14987), .B2(P1_REIP_REG_14__SCAN_IN), .A(n14952), 
        .ZN(n14956) );
  OAI21_X1 U18331 ( .B1(n14953), .B2(P1_REIP_REG_14__SCAN_IN), .A(
        P1_REIP_REG_13__SCAN_IN), .ZN(n14954) );
  OAI211_X1 U18332 ( .C1(P1_REIP_REG_13__SCAN_IN), .C2(P1_REIP_REG_14__SCAN_IN), .A(n14954), .B(n20860), .ZN(n14955) );
  OAI211_X1 U18333 ( .C1(n20897), .C2(n15319), .A(n14956), .B(n14955), .ZN(
        n14957) );
  AOI21_X1 U18334 ( .B1(n20909), .B2(n15513), .A(n14957), .ZN(n14958) );
  OAI21_X1 U18335 ( .B1(n15149), .B2(n20851), .A(n14958), .ZN(P1_U2826) );
  AOI21_X1 U18336 ( .B1(n14959), .B2(n15015), .A(n14960), .ZN(n14997) );
  AOI21_X1 U18337 ( .B1(n14997), .B2(n14961), .A(n14960), .ZN(n14980) );
  INV_X1 U18338 ( .A(n14962), .ZN(n14979) );
  NOR2_X1 U18339 ( .A1(n14980), .A2(n14979), .ZN(n14978) );
  OAI21_X1 U18340 ( .B1(n14978), .B2(n14964), .A(n14963), .ZN(n15334) );
  INV_X1 U18341 ( .A(n15330), .ZN(n14976) );
  NAND2_X1 U18342 ( .A1(n14965), .A2(n14966), .ZN(n14967) );
  NAND2_X1 U18343 ( .A1(n14968), .A2(n14967), .ZN(n15527) );
  INV_X1 U18344 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21516) );
  INV_X1 U18345 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15077) );
  AOI21_X1 U18346 ( .B1(n20912), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17539), .ZN(n14969) );
  OAI21_X1 U18347 ( .B1(n20883), .B2(n15077), .A(n14969), .ZN(n14972) );
  NOR2_X1 U18348 ( .A1(n14970), .A2(n21516), .ZN(n14971) );
  AOI211_X1 U18349 ( .C1(n14973), .C2(n21516), .A(n14972), .B(n14971), .ZN(
        n14974) );
  OAI21_X1 U18350 ( .B1(n20894), .B2(n15527), .A(n14974), .ZN(n14975) );
  AOI21_X1 U18351 ( .B1(n14976), .B2(n20919), .A(n14975), .ZN(n14977) );
  OAI21_X1 U18352 ( .B1(n15334), .B2(n20851), .A(n14977), .ZN(P1_U2827) );
  AOI21_X1 U18353 ( .B1(n14980), .B2(n14979), .A(n14978), .ZN(n14981) );
  INV_X1 U18354 ( .A(n14981), .ZN(n15343) );
  INV_X1 U18355 ( .A(n15336), .ZN(n14994) );
  OR2_X1 U18356 ( .A1(n14982), .A2(n14983), .ZN(n14984) );
  NAND2_X1 U18357 ( .A1(n14965), .A2(n14984), .ZN(n15540) );
  INV_X1 U18358 ( .A(n15007), .ZN(n14985) );
  NOR2_X1 U18359 ( .A1(n15047), .A2(n14985), .ZN(n20845) );
  NAND3_X1 U18360 ( .A1(n20845), .A2(P1_REIP_REG_11__SCAN_IN), .A3(n15011), 
        .ZN(n14986) );
  INV_X1 U18361 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15335) );
  NAND2_X1 U18362 ( .A1(n14986), .A2(n15335), .ZN(n14988) );
  NAND2_X1 U18363 ( .A1(n14988), .A2(n14987), .ZN(n14992) );
  NAND2_X1 U18364 ( .A1(n20912), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14989) );
  OAI211_X1 U18365 ( .C1(n20883), .C2(n15078), .A(n20904), .B(n14989), .ZN(
        n14990) );
  INV_X1 U18366 ( .A(n14990), .ZN(n14991) );
  OAI211_X1 U18367 ( .C1(n15540), .C2(n20894), .A(n14992), .B(n14991), .ZN(
        n14993) );
  AOI21_X1 U18368 ( .B1(n20919), .B2(n14994), .A(n14993), .ZN(n14995) );
  OAI21_X1 U18369 ( .B1(n15343), .B2(n20851), .A(n14995), .ZN(P1_U2828) );
  XNOR2_X1 U18370 ( .A(n14997), .B(n14996), .ZN(n15349) );
  INV_X1 U18371 ( .A(n15347), .ZN(n15006) );
  NOR2_X1 U18372 ( .A1(n14998), .A2(n14999), .ZN(n15000) );
  OR2_X1 U18373 ( .A1(n14982), .A2(n15000), .ZN(n15545) );
  NAND2_X1 U18374 ( .A1(n20912), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15001) );
  NAND2_X1 U18375 ( .A1(n15001), .A2(n20904), .ZN(n15002) );
  AOI21_X1 U18376 ( .B1(n20907), .B2(P1_EBX_REG_11__SCAN_IN), .A(n15002), .ZN(
        n15004) );
  INV_X1 U18377 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n21513) );
  NAND3_X1 U18378 ( .A1(n20845), .A2(n15011), .A3(n21513), .ZN(n15003) );
  OAI211_X1 U18379 ( .C1(n15545), .C2(n20894), .A(n15004), .B(n15003), .ZN(
        n15005) );
  AOI21_X1 U18380 ( .B1(n20919), .B2(n15006), .A(n15005), .ZN(n15014) );
  NAND2_X1 U18381 ( .A1(n15008), .A2(n15007), .ZN(n15009) );
  AND2_X1 U18382 ( .A1(n20860), .A2(n15009), .ZN(n20849) );
  INV_X1 U18383 ( .A(n20849), .ZN(n15010) );
  OAI21_X1 U18384 ( .B1(n15012), .B2(n15011), .A(n15010), .ZN(n15022) );
  NAND2_X1 U18385 ( .A1(n15022), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n15013) );
  OAI211_X1 U18386 ( .C1(n15155), .C2(n20851), .A(n15014), .B(n15013), .ZN(
        P1_U2829) );
  AOI21_X1 U18387 ( .B1(n15016), .B2(n14402), .A(n14934), .ZN(n15361) );
  INV_X1 U18388 ( .A(n15361), .ZN(n15161) );
  INV_X1 U18389 ( .A(n15359), .ZN(n15026) );
  INV_X1 U18390 ( .A(n20845), .ZN(n15018) );
  NAND2_X1 U18391 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n21511), .ZN(n15017) );
  OAI22_X1 U18392 ( .A1(n15018), .A2(n15017), .B1(n15081), .B2(n20883), .ZN(
        n15025) );
  AND2_X1 U18393 ( .A1(n15019), .A2(n15020), .ZN(n15021) );
  OR2_X1 U18394 ( .A1(n15021), .A2(n14998), .ZN(n15566) );
  AOI22_X1 U18395 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20912), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n15022), .ZN(n15023) );
  OAI211_X1 U18396 ( .C1(n15566), .C2(n20894), .A(n15023), .B(n20904), .ZN(
        n15024) );
  AOI211_X1 U18397 ( .C1(n20919), .C2(n15026), .A(n15025), .B(n15024), .ZN(
        n15027) );
  OAI21_X1 U18398 ( .B1(n15161), .B2(n20851), .A(n15027), .ZN(P1_U2830) );
  NOR2_X1 U18399 ( .A1(n15047), .A2(n21495), .ZN(n20911) );
  NAND4_X1 U18400 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .A4(n20911), .ZN(n20887) );
  NOR2_X1 U18401 ( .A1(n20859), .A2(n20887), .ZN(n20867) );
  NAND3_X1 U18402 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20867), .A3(n21507), 
        .ZN(n15028) );
  OAI21_X1 U18403 ( .B1(n15029), .B2(n20897), .A(n15028), .ZN(n15034) );
  AOI21_X1 U18404 ( .B1(n20912), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17539), .ZN(n15031) );
  AOI22_X1 U18405 ( .A1(n20849), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_EBX_REG_8__SCAN_IN), .B2(n20907), .ZN(n15030) );
  OAI211_X1 U18406 ( .C1(n20894), .C2(n15032), .A(n15031), .B(n15030), .ZN(
        n15033) );
  NOR2_X1 U18407 ( .A1(n15034), .A2(n15033), .ZN(n15035) );
  OAI21_X1 U18408 ( .B1(n20851), .B2(n15036), .A(n15035), .ZN(P1_U2832) );
  NAND2_X1 U18409 ( .A1(n20907), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n15040) );
  AOI21_X1 U18410 ( .B1(n20857), .B2(n21495), .A(n20856), .ZN(n20923) );
  NAND2_X1 U18411 ( .A1(n21498), .A2(n20911), .ZN(n15037) );
  OAI21_X1 U18412 ( .B1(n20923), .B2(n21498), .A(n15037), .ZN(n15038) );
  AOI21_X1 U18413 ( .B1(n20912), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15038), .ZN(n15039) );
  OAI211_X1 U18414 ( .C1(n20895), .C2(n21291), .A(n15040), .B(n15039), .ZN(
        n15043) );
  NOR2_X1 U18415 ( .A1(n20897), .A2(n15041), .ZN(n15042) );
  AOI211_X1 U18416 ( .C1(n15044), .C2(n20909), .A(n15043), .B(n15042), .ZN(
        n15045) );
  OAI21_X1 U18417 ( .B1(n20917), .B2(n15046), .A(n15045), .ZN(P1_U2838) );
  MUX2_X1 U18418 ( .A(n20897), .B(n20882), .S(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15053) );
  AOI22_X1 U18419 ( .A1(n20913), .A2(n21369), .B1(n20856), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n15052) );
  OAI22_X1 U18420 ( .A1(n15048), .A2(n20894), .B1(n15047), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n15049) );
  INV_X1 U18421 ( .A(n15049), .ZN(n15051) );
  NAND2_X1 U18422 ( .A1(n20907), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n15050) );
  AND4_X1 U18423 ( .A1(n15053), .A2(n15052), .A3(n15051), .A4(n15050), .ZN(
        n15054) );
  OAI21_X1 U18424 ( .B1(n20917), .B2(n15055), .A(n15054), .ZN(P1_U2839) );
  INV_X1 U18425 ( .A(n15056), .ZN(n15058) );
  INV_X1 U18426 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15057) );
  OAI22_X1 U18427 ( .A1(n15058), .A2(n20925), .B1(n15057), .B2(n20936), .ZN(
        P1_U2841) );
  AOI22_X1 U18428 ( .A1(n15059), .A2(n20931), .B1(P1_EBX_REG_30__SCAN_IN), 
        .B2(n15075), .ZN(n15060) );
  OAI21_X1 U18429 ( .B1(n15173), .B2(n15079), .A(n15060), .ZN(P1_U2842) );
  AOI22_X1 U18430 ( .A1(n15384), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n15061) );
  OAI21_X1 U18431 ( .B1(n15093), .B2(n15079), .A(n15061), .ZN(P1_U2844) );
  AOI22_X1 U18432 ( .A1(n15388), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n15062) );
  OAI21_X1 U18433 ( .B1(n15196), .B2(n15079), .A(n15062), .ZN(P1_U2845) );
  INV_X1 U18434 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15063) );
  INV_X1 U18435 ( .A(n15204), .ZN(n15101) );
  OAI222_X1 U18436 ( .A1(n15397), .A2(n20925), .B1(n15063), .B2(n20936), .C1(
        n15101), .C2(n15079), .ZN(P1_U2846) );
  INV_X1 U18437 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15064) );
  OAI222_X1 U18438 ( .A1(n15415), .A2(n20925), .B1(n15064), .B2(n20936), .C1(
        n15215), .C2(n15079), .ZN(P1_U2847) );
  INV_X1 U18439 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15065) );
  INV_X1 U18440 ( .A(n15224), .ZN(n15107) );
  OAI222_X1 U18441 ( .A1(n15416), .A2(n20925), .B1(n15065), .B2(n20936), .C1(
        n15107), .C2(n15079), .ZN(P1_U2848) );
  INV_X1 U18442 ( .A(n15231), .ZN(n15111) );
  OAI222_X1 U18443 ( .A1(n15431), .A2(n20925), .B1(n15066), .B2(n20936), .C1(
        n15111), .C2(n15079), .ZN(P1_U2849) );
  AOI22_X1 U18444 ( .A1(n15440), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n15067) );
  OAI21_X1 U18445 ( .B1(n15115), .B2(n15079), .A(n15067), .ZN(P1_U2850) );
  INV_X1 U18446 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15068) );
  INV_X1 U18447 ( .A(n15251), .ZN(n15119) );
  OAI222_X1 U18448 ( .A1(n15444), .A2(n20925), .B1(n15068), .B2(n20936), .C1(
        n15119), .C2(n15079), .ZN(P1_U2851) );
  AOI22_X1 U18449 ( .A1(n15452), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n15069) );
  OAI21_X1 U18450 ( .B1(n15261), .B2(n15079), .A(n15069), .ZN(P1_U2852) );
  AOI22_X1 U18451 ( .A1(n15468), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n15070) );
  OAI21_X1 U18452 ( .B1(n15127), .B2(n15079), .A(n15070), .ZN(P1_U2853) );
  AOI22_X1 U18453 ( .A1(n15471), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_18__SCAN_IN), .ZN(n15071) );
  OAI21_X1 U18454 ( .B1(n15276), .B2(n15079), .A(n15071), .ZN(P1_U2854) );
  AOI22_X1 U18455 ( .A1(n15494), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n15072) );
  OAI21_X1 U18456 ( .B1(n15285), .B2(n15079), .A(n15072), .ZN(P1_U2855) );
  OAI222_X1 U18457 ( .A1(n15501), .A2(n20925), .B1(n15073), .B2(n20936), .C1(
        n15300), .C2(n15079), .ZN(P1_U2856) );
  INV_X1 U18458 ( .A(n15310), .ZN(n15147) );
  OAI222_X1 U18459 ( .A1(n15508), .A2(n20925), .B1(n15074), .B2(n20936), .C1(
        n15147), .C2(n15079), .ZN(P1_U2857) );
  AOI22_X1 U18460 ( .A1(n15513), .A2(n20931), .B1(n15075), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n15076) );
  OAI21_X1 U18461 ( .B1(n15149), .B2(n15079), .A(n15076), .ZN(P1_U2858) );
  OAI222_X1 U18462 ( .A1(n15527), .A2(n20925), .B1(n15077), .B2(n20936), .C1(
        n15334), .C2(n15079), .ZN(P1_U2859) );
  OAI222_X1 U18463 ( .A1(n15540), .A2(n20925), .B1(n15078), .B2(n20936), .C1(
        n15343), .C2(n15079), .ZN(P1_U2860) );
  INV_X1 U18464 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15080) );
  OAI222_X1 U18465 ( .A1(n15545), .A2(n20925), .B1(n15080), .B2(n20936), .C1(
        n15155), .C2(n15079), .ZN(P1_U2861) );
  OAI22_X1 U18466 ( .A1(n15566), .A2(n20925), .B1(n15081), .B2(n20936), .ZN(
        n15082) );
  AOI21_X1 U18467 ( .B1(n15361), .B2(n20932), .A(n15082), .ZN(n15083) );
  INV_X1 U18468 ( .A(n15083), .ZN(P1_U2862) );
  AOI22_X1 U18469 ( .A1(n15128), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n15156), .ZN(n15088) );
  INV_X1 U18470 ( .A(DATAI_14_), .ZN(n15085) );
  NAND2_X1 U18471 ( .A1(n15096), .A2(BUF1_REG_14__SCAN_IN), .ZN(n15084) );
  OAI21_X1 U18472 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n20979) );
  AOI22_X1 U18473 ( .A1(n15142), .A2(n20979), .B1(n15140), .B2(DATAI_30_), 
        .ZN(n15087) );
  OAI211_X1 U18474 ( .C1(n15173), .C2(n15160), .A(n15088), .B(n15087), .ZN(
        P1_U2874) );
  AOI22_X1 U18475 ( .A1(n15128), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n15156), .ZN(n15092) );
  INV_X1 U18476 ( .A(DATAI_12_), .ZN(n15090) );
  NAND2_X1 U18477 ( .A1(n15096), .A2(BUF1_REG_12__SCAN_IN), .ZN(n15089) );
  OAI21_X1 U18478 ( .B1(n15096), .B2(n15090), .A(n15089), .ZN(n20975) );
  AOI22_X1 U18479 ( .A1(n15142), .A2(n20975), .B1(n15140), .B2(DATAI_28_), 
        .ZN(n15091) );
  OAI211_X1 U18480 ( .C1(n15093), .C2(n15160), .A(n15092), .B(n15091), .ZN(
        P1_U2876) );
  AOI22_X1 U18481 ( .A1(n15128), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n15156), .ZN(n15098) );
  INV_X1 U18482 ( .A(DATAI_11_), .ZN(n15095) );
  NAND2_X1 U18483 ( .A1(n15096), .A2(BUF1_REG_11__SCAN_IN), .ZN(n15094) );
  OAI21_X1 U18484 ( .B1(n15096), .B2(n15095), .A(n15094), .ZN(n20973) );
  AOI22_X1 U18485 ( .A1(n15142), .A2(n20973), .B1(n15140), .B2(DATAI_27_), 
        .ZN(n15097) );
  OAI211_X1 U18486 ( .C1(n15196), .C2(n15160), .A(n15098), .B(n15097), .ZN(
        P1_U2877) );
  AOI22_X1 U18487 ( .A1(n15128), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n15156), .ZN(n15100) );
  AOI22_X1 U18488 ( .A1(n15142), .A2(n15157), .B1(n15140), .B2(DATAI_26_), 
        .ZN(n15099) );
  OAI211_X1 U18489 ( .C1(n15101), .C2(n15160), .A(n15100), .B(n15099), .ZN(
        P1_U2878) );
  AOI22_X1 U18490 ( .A1(n15128), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n15156), .ZN(n15103) );
  AOI22_X1 U18491 ( .A1(n15142), .A2(n20971), .B1(n15140), .B2(DATAI_25_), 
        .ZN(n15102) );
  OAI211_X1 U18492 ( .C1(n15215), .C2(n15160), .A(n15103), .B(n15102), .ZN(
        P1_U2879) );
  AOI22_X1 U18493 ( .A1(n15128), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n15156), .ZN(n15106) );
  AOI22_X1 U18494 ( .A1(n15142), .A2(n15104), .B1(n15140), .B2(DATAI_24_), 
        .ZN(n15105) );
  OAI211_X1 U18495 ( .C1(n15107), .C2(n15160), .A(n15106), .B(n15105), .ZN(
        P1_U2880) );
  AOI22_X1 U18496 ( .A1(n15128), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n15156), .ZN(n15110) );
  AOI22_X1 U18497 ( .A1(n15142), .A2(n15108), .B1(n15140), .B2(DATAI_23_), 
        .ZN(n15109) );
  OAI211_X1 U18498 ( .C1(n15111), .C2(n15160), .A(n15110), .B(n15109), .ZN(
        P1_U2881) );
  AOI22_X1 U18499 ( .A1(n15128), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n15156), .ZN(n15114) );
  AOI22_X1 U18500 ( .A1(n15142), .A2(n15112), .B1(n15140), .B2(DATAI_22_), 
        .ZN(n15113) );
  OAI211_X1 U18501 ( .C1(n15115), .C2(n15160), .A(n15114), .B(n15113), .ZN(
        P1_U2882) );
  AOI22_X1 U18502 ( .A1(n15128), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n15156), .ZN(n15118) );
  AOI22_X1 U18503 ( .A1(n15142), .A2(n15116), .B1(n15140), .B2(DATAI_21_), 
        .ZN(n15117) );
  OAI211_X1 U18504 ( .C1(n15119), .C2(n15160), .A(n15118), .B(n15117), .ZN(
        P1_U2883) );
  INV_X1 U18505 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n17632) );
  OAI22_X1 U18506 ( .A1(n15138), .A2(n17632), .B1(n13921), .B2(n15151), .ZN(
        n15120) );
  INV_X1 U18507 ( .A(n15120), .ZN(n15123) );
  AOI22_X1 U18508 ( .A1(n15142), .A2(n15121), .B1(n15140), .B2(DATAI_20_), 
        .ZN(n15122) );
  OAI211_X1 U18509 ( .C1(n15261), .C2(n15160), .A(n15123), .B(n15122), .ZN(
        P1_U2884) );
  AOI22_X1 U18510 ( .A1(n15128), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n15156), .ZN(n15126) );
  AOI22_X1 U18511 ( .A1(n15142), .A2(n15124), .B1(n15140), .B2(DATAI_19_), 
        .ZN(n15125) );
  OAI211_X1 U18512 ( .C1(n15127), .C2(n15160), .A(n15126), .B(n15125), .ZN(
        P1_U2885) );
  AOI22_X1 U18513 ( .A1(n15128), .A2(BUF1_REG_18__SCAN_IN), .B1(
        P1_EAX_REG_18__SCAN_IN), .B2(n15156), .ZN(n15131) );
  AOI22_X1 U18514 ( .A1(n15142), .A2(n15129), .B1(n15140), .B2(DATAI_18_), 
        .ZN(n15130) );
  OAI211_X1 U18515 ( .C1(n15276), .C2(n15160), .A(n15131), .B(n15130), .ZN(
        P1_U2886) );
  INV_X1 U18516 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16181) );
  OAI22_X1 U18517 ( .A1(n15138), .A2(n16181), .B1(n15132), .B2(n15151), .ZN(
        n15133) );
  INV_X1 U18518 ( .A(n15133), .ZN(n15136) );
  AOI22_X1 U18519 ( .A1(n15142), .A2(n15134), .B1(n15140), .B2(DATAI_17_), 
        .ZN(n15135) );
  OAI211_X1 U18520 ( .C1(n15285), .C2(n15160), .A(n15136), .B(n15135), .ZN(
        P1_U2887) );
  OAI22_X1 U18521 ( .A1(n15138), .A2(n17638), .B1(n15137), .B2(n15151), .ZN(
        n15139) );
  INV_X1 U18522 ( .A(n15139), .ZN(n15144) );
  AOI22_X1 U18523 ( .A1(n15142), .A2(n15141), .B1(n15140), .B2(DATAI_16_), 
        .ZN(n15143) );
  OAI211_X1 U18524 ( .C1(n15300), .C2(n15160), .A(n15144), .B(n15143), .ZN(
        P1_U2888) );
  AOI22_X1 U18525 ( .A1(n15158), .A2(n15145), .B1(P1_EAX_REG_15__SCAN_IN), 
        .B2(n15156), .ZN(n15146) );
  OAI21_X1 U18526 ( .B1(n15147), .B2(n15160), .A(n15146), .ZN(P1_U2889) );
  AOI22_X1 U18527 ( .A1(n15158), .A2(n20979), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15156), .ZN(n15148) );
  OAI21_X1 U18528 ( .B1(n15149), .B2(n15160), .A(n15148), .ZN(P1_U2890) );
  AOI22_X1 U18529 ( .A1(n15158), .A2(n20977), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15156), .ZN(n15150) );
  OAI21_X1 U18530 ( .B1(n15334), .B2(n15160), .A(n15150), .ZN(P1_U2891) );
  INV_X1 U18531 ( .A(n20975), .ZN(n15152) );
  INV_X1 U18532 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21643) );
  OAI222_X1 U18533 ( .A1(n15343), .A2(n15160), .B1(n15153), .B2(n15152), .C1(
        n21643), .C2(n15151), .ZN(P1_U2892) );
  AOI22_X1 U18534 ( .A1(n15158), .A2(n20973), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15156), .ZN(n15154) );
  OAI21_X1 U18535 ( .B1(n15155), .B2(n15160), .A(n15154), .ZN(P1_U2893) );
  AOI22_X1 U18536 ( .A1(n15158), .A2(n15157), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15156), .ZN(n15159) );
  OAI21_X1 U18537 ( .B1(n15161), .B2(n15160), .A(n15159), .ZN(P1_U2894) );
  AOI21_X1 U18538 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15162), .ZN(n15163) );
  OAI21_X1 U18539 ( .B1(n15164), .B2(n17524), .A(n15163), .ZN(n15165) );
  AOI21_X1 U18540 ( .B1(n15166), .B2(n17530), .A(n15165), .ZN(n15167) );
  OAI21_X1 U18541 ( .B1(n15168), .B2(n20829), .A(n15167), .ZN(P1_U2968) );
  NOR2_X1 U18542 ( .A1(n15169), .A2(n17524), .ZN(n15170) );
  AOI211_X1 U18543 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15171), .B(n15170), .ZN(n15172) );
  NAND2_X1 U18544 ( .A1(n15175), .A2(n15197), .ZN(n15179) );
  OAI21_X1 U18545 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15176), .A(
        n15179), .ZN(n15178) );
  INV_X1 U18546 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15192) );
  MUX2_X1 U18547 ( .A(n15192), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n10154), .Z(n15177) );
  OAI211_X1 U18548 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15179), .A(
        n15178), .B(n15177), .ZN(n15181) );
  XNOR2_X1 U18549 ( .A(n15181), .B(n15180), .ZN(n15387) );
  NAND2_X1 U18550 ( .A1(n17539), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n15380) );
  NAND2_X1 U18551 ( .A1(n17517), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15182) );
  OAI211_X1 U18552 ( .C1(n15183), .C2(n17524), .A(n15380), .B(n15182), .ZN(
        n15184) );
  AOI21_X1 U18553 ( .B1(n15185), .B2(n17530), .A(n15184), .ZN(n15186) );
  OAI21_X1 U18554 ( .B1(n20829), .B2(n15387), .A(n15186), .ZN(P1_U2971) );
  NOR2_X1 U18555 ( .A1(n20904), .A2(n21542), .ZN(n15392) );
  NOR2_X1 U18556 ( .A1(n17533), .A2(n15187), .ZN(n15188) );
  AOI211_X1 U18557 ( .C1(n15189), .C2(n17528), .A(n15392), .B(n15188), .ZN(
        n15195) );
  INV_X1 U18558 ( .A(n15190), .ZN(n15191) );
  XNOR2_X1 U18559 ( .A(n15193), .B(n15192), .ZN(n15389) );
  NAND2_X1 U18560 ( .A1(n15389), .A2(n17531), .ZN(n15194) );
  OAI211_X1 U18561 ( .C1(n15196), .C2(n15370), .A(n15195), .B(n15194), .ZN(
        P1_U2972) );
  NAND3_X1 U18562 ( .A1(n15198), .A2(n15216), .A3(n15197), .ZN(n15200) );
  XNOR2_X1 U18563 ( .A(n15200), .B(n15199), .ZN(n15407) );
  NOR2_X1 U18564 ( .A1(n20904), .A2(n21541), .ZN(n15404) );
  AOI21_X1 U18565 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15404), .ZN(n15201) );
  OAI21_X1 U18566 ( .B1(n15202), .B2(n17524), .A(n15201), .ZN(n15203) );
  AOI21_X1 U18567 ( .B1(n15204), .B2(n17530), .A(n15203), .ZN(n15205) );
  OAI21_X1 U18568 ( .B1(n20829), .B2(n15407), .A(n15205), .ZN(P1_U2973) );
  NOR2_X1 U18569 ( .A1(n20904), .A2(n21537), .ZN(n15411) );
  NOR2_X1 U18570 ( .A1(n17533), .A2(n15206), .ZN(n15207) );
  AOI211_X1 U18571 ( .C1(n15208), .C2(n17528), .A(n15411), .B(n15207), .ZN(
        n15214) );
  NOR2_X1 U18572 ( .A1(n10735), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15217) );
  AOI21_X1 U18573 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n10735), .A(
        n15217), .ZN(n15226) );
  NAND3_X1 U18574 ( .A1(n15175), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15226), .ZN(n15211) );
  NAND2_X1 U18575 ( .A1(n15209), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15422) );
  NAND2_X1 U18576 ( .A1(n10735), .A2(n15422), .ZN(n15210) );
  AOI21_X1 U18577 ( .B1(n10640), .B2(n15209), .A(n11121), .ZN(n15219) );
  AOI21_X1 U18578 ( .B1(n15211), .B2(n15210), .A(n15219), .ZN(n15212) );
  XNOR2_X1 U18579 ( .A(n15212), .B(n15398), .ZN(n15408) );
  NAND2_X1 U18580 ( .A1(n15408), .A2(n17531), .ZN(n15213) );
  OAI211_X1 U18581 ( .C1(n15215), .C2(n15370), .A(n15214), .B(n15213), .ZN(
        P1_U2974) );
  INV_X1 U18582 ( .A(n15216), .ZN(n15218) );
  NOR3_X1 U18583 ( .A1(n15219), .A2(n15218), .A3(n15217), .ZN(n15220) );
  XNOR2_X1 U18584 ( .A(n15220), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15426) );
  NOR2_X1 U18585 ( .A1(n20904), .A2(n21536), .ZN(n15419) );
  AOI21_X1 U18586 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15419), .ZN(n15221) );
  OAI21_X1 U18587 ( .B1(n15222), .B2(n17524), .A(n15221), .ZN(n15223) );
  AOI21_X1 U18588 ( .B1(n15224), .B2(n17530), .A(n15223), .ZN(n15225) );
  OAI21_X1 U18589 ( .B1(n20829), .B2(n15426), .A(n15225), .ZN(P1_U2975) );
  XNOR2_X1 U18590 ( .A(n15175), .B(n15226), .ZN(n15434) );
  NAND2_X1 U18591 ( .A1(n17528), .A2(n15227), .ZN(n15228) );
  NAND2_X1 U18592 ( .A1(n17539), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15430) );
  OAI211_X1 U18593 ( .C1(n17533), .C2(n15229), .A(n15228), .B(n15430), .ZN(
        n15230) );
  AOI21_X1 U18594 ( .B1(n15231), .B2(n17530), .A(n15230), .ZN(n15232) );
  OAI21_X1 U18595 ( .B1(n15434), .B2(n20829), .A(n15232), .ZN(P1_U2976) );
  NAND2_X1 U18596 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  XNOR2_X1 U18597 ( .A(n15235), .B(n15435), .ZN(n15443) );
  NOR2_X1 U18598 ( .A1(n20904), .A2(n21532), .ZN(n15437) );
  AOI21_X1 U18599 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15437), .ZN(n15236) );
  OAI21_X1 U18600 ( .B1(n15237), .B2(n17524), .A(n15236), .ZN(n15238) );
  AOI21_X1 U18601 ( .B1(n15239), .B2(n17530), .A(n15238), .ZN(n15240) );
  OAI21_X1 U18602 ( .B1(n20829), .B2(n15443), .A(n15240), .ZN(P1_U2977) );
  NOR3_X1 U18603 ( .A1(n15241), .A2(n10154), .A3(n15242), .ZN(n15256) );
  NOR3_X1 U18604 ( .A1(n15243), .A2(n10735), .A3(n15244), .ZN(n15245) );
  AOI21_X1 U18605 ( .B1(n15256), .B2(n10642), .A(n15245), .ZN(n15246) );
  XOR2_X1 U18606 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15246), .Z(
        n15451) );
  NAND2_X1 U18607 ( .A1(n17528), .A2(n15247), .ZN(n15248) );
  NAND2_X1 U18608 ( .A1(n17539), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15445) );
  OAI211_X1 U18609 ( .C1(n17533), .C2(n15249), .A(n15248), .B(n15445), .ZN(
        n15250) );
  AOI21_X1 U18610 ( .B1(n15251), .B2(n17530), .A(n15250), .ZN(n15252) );
  OAI21_X1 U18611 ( .B1(n15451), .B2(n20829), .A(n15252), .ZN(P1_U2978) );
  INV_X1 U18612 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15253) );
  NOR2_X1 U18613 ( .A1(n20904), .A2(n15253), .ZN(n15458) );
  NOR2_X1 U18614 ( .A1(n17524), .A2(n15254), .ZN(n15255) );
  AOI211_X1 U18615 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15458), .B(n15255), .ZN(n15260) );
  NOR3_X1 U18616 ( .A1(n15243), .A2(n10735), .A3(n15456), .ZN(n15257) );
  NOR2_X1 U18617 ( .A1(n15257), .A2(n15256), .ZN(n15258) );
  XNOR2_X1 U18618 ( .A(n15258), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15453) );
  NAND2_X1 U18619 ( .A1(n15453), .A2(n17531), .ZN(n15259) );
  OAI211_X1 U18620 ( .C1(n15261), .C2(n15370), .A(n15260), .B(n15259), .ZN(
        P1_U2979) );
  NAND2_X1 U18621 ( .A1(n15243), .A2(n15262), .ZN(n15264) );
  XNOR2_X1 U18622 ( .A(n11121), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15263) );
  XNOR2_X1 U18623 ( .A(n15264), .B(n15263), .ZN(n15470) );
  NAND2_X1 U18624 ( .A1(n17528), .A2(n15265), .ZN(n15266) );
  NAND2_X1 U18625 ( .A1(n17539), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n15464) );
  OAI211_X1 U18626 ( .C1(n17533), .C2(n15267), .A(n15266), .B(n15464), .ZN(
        n15268) );
  AOI21_X1 U18627 ( .B1(n15269), .B2(n17530), .A(n15268), .ZN(n15270) );
  OAI21_X1 U18628 ( .B1(n15470), .B2(n20829), .A(n15270), .ZN(P1_U2980) );
  NOR2_X1 U18629 ( .A1(n20904), .A2(n21526), .ZN(n15484) );
  NOR2_X1 U18630 ( .A1(n17524), .A2(n15271), .ZN(n15272) );
  AOI211_X1 U18631 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15484), .B(n15272), .ZN(n15275) );
  OR2_X1 U18632 ( .A1(n15241), .A2(n15273), .ZN(n15472) );
  NAND3_X1 U18633 ( .A1(n15472), .A2(n15243), .A3(n17531), .ZN(n15274) );
  OAI211_X1 U18634 ( .C1(n15276), .C2(n15370), .A(n15275), .B(n15274), .ZN(
        P1_U2981) );
  NAND2_X1 U18635 ( .A1(n15293), .A2(n15283), .ZN(n15282) );
  NOR2_X1 U18636 ( .A1(n10735), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15364) );
  AOI21_X1 U18637 ( .B1(n15312), .B2(n15281), .A(n15280), .ZN(n15302) );
  NAND2_X1 U18638 ( .A1(n10735), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15303) );
  NAND2_X1 U18639 ( .A1(n15302), .A2(n15303), .ZN(n15301) );
  MUX2_X1 U18640 ( .A(n15283), .B(n15282), .S(n15301), .Z(n15284) );
  XNOR2_X1 U18641 ( .A(n15284), .B(n15491), .ZN(n15496) );
  INV_X1 U18642 ( .A(n15285), .ZN(n15289) );
  NOR2_X1 U18643 ( .A1(n20904), .A2(n21523), .ZN(n15493) );
  AOI21_X1 U18644 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15493), .ZN(n15286) );
  OAI21_X1 U18645 ( .B1(n15287), .B2(n17524), .A(n15286), .ZN(n15288) );
  AOI21_X1 U18646 ( .B1(n15289), .B2(n17530), .A(n15288), .ZN(n15290) );
  OAI21_X1 U18647 ( .B1(n15496), .B2(n20829), .A(n15290), .ZN(P1_U2982) );
  AOI21_X1 U18648 ( .B1(n15301), .B2(n15305), .A(n15291), .ZN(n15294) );
  INV_X1 U18649 ( .A(n15291), .ZN(n15292) );
  OAI22_X1 U18650 ( .A1(n15294), .A2(n15293), .B1(n15292), .B2(n15301), .ZN(
        n15497) );
  NAND2_X1 U18651 ( .A1(n15497), .A2(n17531), .ZN(n15299) );
  NAND2_X1 U18652 ( .A1(n17539), .A2(P1_REIP_REG_16__SCAN_IN), .ZN(n15500) );
  OAI21_X1 U18653 ( .B1(n17533), .B2(n15295), .A(n15500), .ZN(n15296) );
  AOI21_X1 U18654 ( .B1(n17528), .B2(n15297), .A(n15296), .ZN(n15298) );
  OAI211_X1 U18655 ( .C1(n15370), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        P1_U2983) );
  INV_X1 U18656 ( .A(n15301), .ZN(n15306) );
  AOI21_X1 U18657 ( .B1(n15305), .B2(n15303), .A(n15302), .ZN(n15304) );
  NOR2_X1 U18658 ( .A1(n20904), .A2(n21520), .ZN(n15505) );
  AOI21_X1 U18659 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15505), .ZN(n15307) );
  OAI21_X1 U18660 ( .B1(n15308), .B2(n17524), .A(n15307), .ZN(n15309) );
  AOI21_X1 U18661 ( .B1(n15310), .B2(n17530), .A(n15309), .ZN(n15311) );
  INV_X1 U18662 ( .A(n15312), .ZN(n15315) );
  OAI21_X1 U18663 ( .B1(n15315), .B2(n15314), .A(n15313), .ZN(n15317) );
  XNOR2_X1 U18664 ( .A(n10154), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15316) );
  XNOR2_X1 U18665 ( .A(n15317), .B(n15316), .ZN(n15519) );
  INV_X1 U18666 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n21518) );
  NOR2_X1 U18667 ( .A1(n20904), .A2(n21518), .ZN(n15512) );
  AOI21_X1 U18668 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15512), .ZN(n15318) );
  OAI21_X1 U18669 ( .B1(n15319), .B2(n17524), .A(n15318), .ZN(n15320) );
  AOI21_X1 U18670 ( .B1(n15321), .B2(n17530), .A(n15320), .ZN(n15322) );
  OAI21_X1 U18671 ( .B1(n15519), .B2(n20829), .A(n15322), .ZN(P1_U2985) );
  INV_X1 U18672 ( .A(n15323), .ZN(n15324) );
  AOI21_X1 U18673 ( .B1(n15352), .B2(n15325), .A(n15324), .ZN(n15340) );
  AND2_X1 U18674 ( .A1(n15326), .A2(n15327), .ZN(n15339) );
  NAND2_X1 U18675 ( .A1(n15340), .A2(n15339), .ZN(n15338) );
  NAND2_X1 U18676 ( .A1(n15338), .A2(n15327), .ZN(n15328) );
  XOR2_X1 U18677 ( .A(n15329), .B(n15328), .Z(n15530) );
  NAND2_X1 U18678 ( .A1(n15530), .A2(n17531), .ZN(n15333) );
  NOR2_X1 U18679 ( .A1(n20904), .A2(n21516), .ZN(n15523) );
  NOR2_X1 U18680 ( .A1(n17524), .A2(n15330), .ZN(n15331) );
  AOI211_X1 U18681 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15523), .B(n15331), .ZN(n15332) );
  OAI211_X1 U18682 ( .C1(n15370), .C2(n15334), .A(n15333), .B(n15332), .ZN(
        P1_U2986) );
  NOR2_X1 U18683 ( .A1(n20904), .A2(n15335), .ZN(n15537) );
  NOR2_X1 U18684 ( .A1(n17524), .A2(n15336), .ZN(n15337) );
  AOI211_X1 U18685 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15537), .B(n15337), .ZN(n15342) );
  OAI21_X1 U18686 ( .B1(n15340), .B2(n15339), .A(n15338), .ZN(n15532) );
  NAND2_X1 U18687 ( .A1(n15532), .A2(n17531), .ZN(n15341) );
  OAI211_X1 U18688 ( .C1(n15343), .C2(n15370), .A(n15342), .B(n15341), .ZN(
        P1_U2987) );
  NAND3_X1 U18689 ( .A1(n15351), .A2(n10735), .A3(n15556), .ZN(n15355) );
  NAND2_X1 U18690 ( .A1(n15344), .A2(n15355), .ZN(n15345) );
  XNOR2_X1 U18691 ( .A(n15345), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15555) );
  NOR2_X1 U18692 ( .A1(n20904), .A2(n21513), .ZN(n15548) );
  AOI21_X1 U18693 ( .B1(n17517), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15548), .ZN(n15346) );
  OAI21_X1 U18694 ( .B1(n15347), .B2(n17524), .A(n15346), .ZN(n15348) );
  AOI21_X1 U18695 ( .B1(n15349), .B2(n17530), .A(n15348), .ZN(n15350) );
  OAI21_X1 U18696 ( .B1(n15555), .B2(n20829), .A(n15350), .ZN(P1_U2988) );
  NOR2_X1 U18697 ( .A1(n15351), .A2(n15556), .ZN(n15354) );
  XNOR2_X1 U18698 ( .A(n15352), .B(n15556), .ZN(n15353) );
  MUX2_X1 U18699 ( .A(n15354), .B(n15353), .S(n10154), .Z(n15357) );
  INV_X1 U18700 ( .A(n15355), .ZN(n15356) );
  NOR2_X1 U18701 ( .A1(n15357), .A2(n15356), .ZN(n15570) );
  NAND2_X1 U18702 ( .A1(n17539), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15564) );
  NAND2_X1 U18703 ( .A1(n17517), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15358) );
  OAI211_X1 U18704 ( .C1(n17524), .C2(n15359), .A(n15564), .B(n15358), .ZN(
        n15360) );
  AOI21_X1 U18705 ( .B1(n15361), .B2(n17530), .A(n15360), .ZN(n15362) );
  OAI21_X1 U18706 ( .B1(n15570), .B2(n20829), .A(n15362), .ZN(P1_U2989) );
  NOR2_X1 U18707 ( .A1(n15364), .A2(n15363), .ZN(n15366) );
  XOR2_X1 U18708 ( .A(n15366), .B(n15365), .Z(n15572) );
  NAND2_X1 U18709 ( .A1(n15572), .A2(n17531), .ZN(n15369) );
  NOR2_X1 U18710 ( .A1(n20904), .A2(n21509), .ZN(n15578) );
  NOR2_X1 U18711 ( .A1(n17524), .A2(n20850), .ZN(n15367) );
  AOI211_X1 U18712 ( .C1(n17517), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15578), .B(n15367), .ZN(n15368) );
  OAI211_X1 U18713 ( .C1(n15370), .C2(n20926), .A(n15369), .B(n15368), .ZN(
        P1_U2990) );
  INV_X1 U18714 ( .A(n14741), .ZN(n15377) );
  INV_X1 U18715 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15374) );
  NAND3_X1 U18716 ( .A1(n15371), .A2(n10636), .A3(n15374), .ZN(n15372) );
  OAI211_X1 U18717 ( .C1(n15375), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15376) );
  AOI21_X1 U18718 ( .B1(n15377), .B2(n20998), .A(n15376), .ZN(n15378) );
  OAI21_X1 U18719 ( .B1(n15379), .B2(n17559), .A(n15378), .ZN(P1_U3002) );
  INV_X1 U18720 ( .A(n15380), .ZN(n15383) );
  NOR3_X1 U18721 ( .A1(n15390), .A2(n10636), .A3(n15381), .ZN(n15382) );
  AOI211_X1 U18722 ( .C1(n15393), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15383), .B(n15382), .ZN(n15386) );
  NAND2_X1 U18723 ( .A1(n15384), .A2(n20998), .ZN(n15385) );
  OAI211_X1 U18724 ( .C1(n15387), .C2(n17559), .A(n15386), .B(n15385), .ZN(
        P1_U3003) );
  INV_X1 U18725 ( .A(n15388), .ZN(n15396) );
  NAND2_X1 U18726 ( .A1(n15389), .A2(n20999), .ZN(n15395) );
  NOR2_X1 U18727 ( .A1(n15390), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15391) );
  AOI211_X1 U18728 ( .C1(n15393), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15392), .B(n15391), .ZN(n15394) );
  OAI211_X1 U18729 ( .C1(n15576), .C2(n15396), .A(n15395), .B(n15394), .ZN(
        P1_U3004) );
  INV_X1 U18730 ( .A(n15397), .ZN(n15405) );
  INV_X1 U18731 ( .A(n15428), .ZN(n15417) );
  NAND4_X1 U18732 ( .A1(n15417), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(n15398), .ZN(n15409) );
  INV_X1 U18733 ( .A(n15399), .ZN(n15400) );
  AOI21_X1 U18734 ( .B1(n15417), .B2(n15400), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15401) );
  AOI21_X1 U18735 ( .B1(n15402), .B2(n15409), .A(n15401), .ZN(n15403) );
  AOI211_X1 U18736 ( .C1(n15405), .C2(n20998), .A(n15404), .B(n15403), .ZN(
        n15406) );
  OAI21_X1 U18737 ( .B1(n15407), .B2(n17559), .A(n15406), .ZN(P1_U3005) );
  NAND2_X1 U18738 ( .A1(n15408), .A2(n20999), .ZN(n15414) );
  INV_X1 U18739 ( .A(n15409), .ZN(n15410) );
  AOI211_X1 U18740 ( .C1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15412), .A(
        n15411), .B(n15410), .ZN(n15413) );
  OAI211_X1 U18741 ( .C1(n15576), .C2(n15415), .A(n15414), .B(n15413), .ZN(
        P1_U3006) );
  INV_X1 U18742 ( .A(n15416), .ZN(n15424) );
  NAND2_X1 U18743 ( .A1(n15417), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15418) );
  MUX2_X1 U18744 ( .A(n15418), .B(n15427), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n15421) );
  INV_X1 U18745 ( .A(n15419), .ZN(n15420) );
  OAI211_X1 U18746 ( .C1(n15535), .C2(n15422), .A(n15421), .B(n15420), .ZN(
        n15423) );
  AOI21_X1 U18747 ( .B1(n15424), .B2(n20998), .A(n15423), .ZN(n15425) );
  OAI21_X1 U18748 ( .B1(n15426), .B2(n17559), .A(n15425), .ZN(P1_U3007) );
  MUX2_X1 U18749 ( .A(n15428), .B(n15427), .S(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n15429) );
  OAI211_X1 U18750 ( .C1(n15431), .C2(n15576), .A(n15430), .B(n15429), .ZN(
        n15432) );
  INV_X1 U18751 ( .A(n15432), .ZN(n15433) );
  OAI21_X1 U18752 ( .B1(n15434), .B2(n17559), .A(n15433), .ZN(P1_U3008) );
  NOR2_X1 U18753 ( .A1(n10643), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15438) );
  NAND2_X1 U18754 ( .A1(n15439), .A2(n10643), .ZN(n15446) );
  AOI21_X1 U18755 ( .B1(n15447), .B2(n15446), .A(n15435), .ZN(n15436) );
  AOI211_X1 U18756 ( .C1(n15439), .C2(n15438), .A(n15437), .B(n15436), .ZN(
        n15442) );
  NAND2_X1 U18757 ( .A1(n15440), .A2(n20998), .ZN(n15441) );
  OAI211_X1 U18758 ( .C1(n15443), .C2(n17559), .A(n15442), .B(n15441), .ZN(
        P1_U3009) );
  INV_X1 U18759 ( .A(n15444), .ZN(n15449) );
  OAI211_X1 U18760 ( .C1(n15447), .C2(n10643), .A(n15446), .B(n15445), .ZN(
        n15448) );
  AOI21_X1 U18761 ( .B1(n15449), .B2(n20998), .A(n15448), .ZN(n15450) );
  OAI21_X1 U18762 ( .B1(n15451), .B2(n17559), .A(n15450), .ZN(P1_U3010) );
  INV_X1 U18763 ( .A(n15452), .ZN(n15462) );
  NAND2_X1 U18764 ( .A1(n15453), .A2(n20999), .ZN(n15461) );
  INV_X1 U18765 ( .A(n15463), .ZN(n15455) );
  OAI21_X1 U18766 ( .B1(n15520), .B2(n21003), .A(n15456), .ZN(n15454) );
  AOI21_X1 U18767 ( .B1(n15455), .B2(n15454), .A(n10642), .ZN(n15459) );
  NOR3_X1 U18768 ( .A1(n15466), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15456), .ZN(n15457) );
  NOR3_X1 U18769 ( .A1(n15459), .A2(n15458), .A3(n15457), .ZN(n15460) );
  OAI211_X1 U18770 ( .C1(n15576), .C2(n15462), .A(n15461), .B(n15460), .ZN(
        P1_U3011) );
  NAND2_X1 U18771 ( .A1(n15463), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15465) );
  OAI211_X1 U18772 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15466), .A(
        n15465), .B(n15464), .ZN(n15467) );
  AOI21_X1 U18773 ( .B1(n15468), .B2(n20998), .A(n15467), .ZN(n15469) );
  OAI21_X1 U18774 ( .B1(n15470), .B2(n17559), .A(n15469), .ZN(P1_U3012) );
  INV_X1 U18775 ( .A(n15471), .ZN(n15488) );
  NAND3_X1 U18776 ( .A1(n15472), .A2(n15243), .A3(n20999), .ZN(n15487) );
  INV_X1 U18777 ( .A(n15473), .ZN(n15481) );
  OAI21_X1 U18778 ( .B1(n15524), .B2(n15514), .A(n15477), .ZN(n15474) );
  INV_X1 U18779 ( .A(n15474), .ZN(n15475) );
  NOR2_X1 U18780 ( .A1(n17540), .A2(n15475), .ZN(n15522) );
  NAND2_X1 U18781 ( .A1(n15477), .A2(n15515), .ZN(n15476) );
  NAND2_X1 U18782 ( .A1(n15522), .A2(n15476), .ZN(n15510) );
  AOI21_X1 U18783 ( .B1(n15477), .B2(n15481), .A(n15510), .ZN(n15489) );
  INV_X1 U18784 ( .A(n15489), .ZN(n15485) );
  INV_X1 U18785 ( .A(n15478), .ZN(n15479) );
  INV_X1 U18786 ( .A(n15506), .ZN(n15482) );
  NOR3_X1 U18787 ( .A1(n15482), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15481), .ZN(n15483) );
  AOI211_X1 U18788 ( .C1(n15485), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15484), .B(n15483), .ZN(n15486) );
  OAI211_X1 U18789 ( .C1(n15576), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        P1_U3013) );
  NAND3_X1 U18790 ( .A1(n15506), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15490) );
  AOI21_X1 U18791 ( .B1(n15491), .B2(n15490), .A(n15489), .ZN(n15492) );
  AOI211_X1 U18792 ( .C1(n15494), .C2(n20998), .A(n15493), .B(n15492), .ZN(
        n15495) );
  OAI21_X1 U18793 ( .B1(n15496), .B2(n17559), .A(n15495), .ZN(P1_U3014) );
  INV_X1 U18794 ( .A(n15497), .ZN(n15504) );
  XNOR2_X1 U18795 ( .A(n21704), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15498) );
  NAND2_X1 U18796 ( .A1(n15506), .A2(n15498), .ZN(n15499) );
  OAI211_X1 U18797 ( .C1(n15501), .C2(n15576), .A(n15500), .B(n15499), .ZN(
        n15502) );
  AOI21_X1 U18798 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15510), .A(
        n15502), .ZN(n15503) );
  OAI21_X1 U18799 ( .B1(n15504), .B2(n17559), .A(n15503), .ZN(P1_U3015) );
  AOI21_X1 U18800 ( .B1(n15506), .B2(n21704), .A(n15505), .ZN(n15507) );
  OAI21_X1 U18801 ( .B1(n15508), .B2(n15576), .A(n15507), .ZN(n15509) );
  NOR2_X1 U18802 ( .A1(n15522), .A2(n15515), .ZN(n15511) );
  AOI211_X1 U18803 ( .C1(n15513), .C2(n20998), .A(n15512), .B(n15511), .ZN(
        n15518) );
  INV_X1 U18804 ( .A(n17544), .ZN(n15552) );
  INV_X1 U18805 ( .A(n15514), .ZN(n15516) );
  NAND4_X1 U18806 ( .A1(n15552), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15516), .A4(n15515), .ZN(n15517) );
  OAI211_X1 U18807 ( .C1(n15519), .C2(n17559), .A(n15518), .B(n15517), .ZN(
        P1_U3017) );
  NOR2_X1 U18808 ( .A1(n15520), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15521) );
  NOR2_X1 U18809 ( .A1(n15522), .A2(n15521), .ZN(n15529) );
  AOI21_X1 U18810 ( .B1(n15525), .B2(n15524), .A(n15523), .ZN(n15526) );
  OAI21_X1 U18811 ( .B1(n15527), .B2(n15576), .A(n15526), .ZN(n15528) );
  AOI211_X1 U18812 ( .C1(n15530), .C2(n20999), .A(n15529), .B(n15528), .ZN(
        n15531) );
  INV_X1 U18813 ( .A(n15531), .ZN(P1_U3018) );
  INV_X1 U18814 ( .A(n15532), .ZN(n15544) );
  OAI22_X1 U18815 ( .A1(n15563), .A2(n15551), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15533), .ZN(n15534) );
  NOR2_X1 U18816 ( .A1(n15534), .A2(n17540), .ZN(n15546) );
  OAI21_X1 U18817 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15535), .A(
        n15546), .ZN(n15542) );
  NAND4_X1 U18818 ( .A1(n15552), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15551), .A4(n15536), .ZN(n15539) );
  INV_X1 U18819 ( .A(n15537), .ZN(n15538) );
  OAI211_X1 U18820 ( .C1(n15576), .C2(n15540), .A(n15539), .B(n15538), .ZN(
        n15541) );
  AOI21_X1 U18821 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15542), .A(
        n15541), .ZN(n15543) );
  OAI21_X1 U18822 ( .B1(n15544), .B2(n17559), .A(n15543), .ZN(P1_U3019) );
  INV_X1 U18823 ( .A(n15545), .ZN(n15549) );
  INV_X1 U18824 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15550) );
  NOR2_X1 U18825 ( .A1(n15546), .A2(n15550), .ZN(n15547) );
  AOI211_X1 U18826 ( .C1(n20998), .C2(n15549), .A(n15548), .B(n15547), .ZN(
        n15554) );
  NAND3_X1 U18827 ( .A1(n15552), .A2(n15551), .A3(n15550), .ZN(n15553) );
  OAI211_X1 U18828 ( .C1(n15555), .C2(n17559), .A(n15554), .B(n15553), .ZN(
        P1_U3020) );
  NAND2_X1 U18829 ( .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15559) );
  NOR2_X1 U18830 ( .A1(n17538), .A2(n15559), .ZN(n15571) );
  XNOR2_X1 U18831 ( .A(n15556), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15568) );
  NOR3_X1 U18832 ( .A1(n15559), .A2(n15558), .A3(n15557), .ZN(n15562) );
  INV_X1 U18833 ( .A(n15560), .ZN(n15561) );
  OAI21_X1 U18834 ( .B1(n15563), .B2(n15562), .A(n15561), .ZN(n15579) );
  NAND2_X1 U18835 ( .A1(n15579), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15565) );
  OAI211_X1 U18836 ( .C1(n15576), .C2(n15566), .A(n15565), .B(n15564), .ZN(
        n15567) );
  AOI21_X1 U18837 ( .B1(n15571), .B2(n15568), .A(n15567), .ZN(n15569) );
  OAI21_X1 U18838 ( .B1(n15570), .B2(n17559), .A(n15569), .ZN(P1_U3021) );
  INV_X1 U18839 ( .A(n15571), .ZN(n15582) );
  NAND2_X1 U18840 ( .A1(n15572), .A2(n20999), .ZN(n15581) );
  NAND2_X1 U18841 ( .A1(n15574), .A2(n15573), .ZN(n15575) );
  AND2_X1 U18842 ( .A1(n15019), .A2(n15575), .ZN(n20846) );
  INV_X1 U18843 ( .A(n20846), .ZN(n20924) );
  NOR2_X1 U18844 ( .A1(n20924), .A2(n15576), .ZN(n15577) );
  AOI211_X1 U18845 ( .C1(n15579), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15578), .B(n15577), .ZN(n15580) );
  OAI211_X1 U18846 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15582), .A(
        n15581), .B(n15580), .ZN(P1_U3022) );
  INV_X1 U18847 ( .A(n13977), .ZN(n15583) );
  NAND2_X1 U18848 ( .A1(n15584), .A2(n15583), .ZN(n15589) );
  OAI21_X1 U18849 ( .B1(n15586), .B2(n15589), .A(n15585), .ZN(n15587) );
  AOI21_X1 U18850 ( .B1(n21369), .B2(n15588), .A(n15587), .ZN(n17474) );
  INV_X1 U18851 ( .A(n17567), .ZN(n15606) );
  INV_X1 U18852 ( .A(n15604), .ZN(n15598) );
  INV_X1 U18853 ( .A(n15589), .ZN(n15591) );
  NOR2_X1 U18854 ( .A1(n13446), .A2(n21835), .ZN(n15596) );
  INV_X1 U18855 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21867) );
  AOI22_X1 U18856 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n11219), .B2(n21867), .ZN(
        n15595) );
  INV_X1 U18857 ( .A(n15595), .ZN(n15590) );
  AOI22_X1 U18858 ( .A1(n15598), .A2(n15591), .B1(n15596), .B2(n15590), .ZN(
        n15592) );
  OAI21_X1 U18859 ( .B1(n17474), .B2(n15606), .A(n15592), .ZN(n15593) );
  INV_X1 U18860 ( .A(n15601), .ZN(n17570) );
  MUX2_X1 U18861 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15593), .S(
        n17570), .Z(P1_U3473) );
  NAND2_X1 U18862 ( .A1(n15594), .A2(n17567), .ZN(n15600) );
  AOI22_X1 U18863 ( .A1(n15598), .A2(n15597), .B1(n15596), .B2(n15595), .ZN(
        n15599) );
  NAND2_X1 U18864 ( .A1(n15600), .A2(n15599), .ZN(n15603) );
  MUX2_X1 U18865 ( .A(n15603), .B(n15602), .S(n15601), .Z(P1_U3472) );
  OAI22_X1 U18866 ( .A1(n15607), .A2(n15606), .B1(n15605), .B2(n15604), .ZN(
        n15608) );
  MUX2_X1 U18867 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15608), .S(
        n17570), .Z(P1_U3469) );
  OAI21_X1 U18868 ( .B1(n15611), .B2(n15610), .A(n15609), .ZN(n16494) );
  INV_X1 U18869 ( .A(n15613), .ZN(n15614) );
  OAI21_X1 U18870 ( .B1(n9804), .B2(n10334), .A(n19994), .ZN(n15618) );
  INV_X1 U18871 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16232) );
  NAND2_X1 U18872 ( .A1(n15619), .A2(n15984), .ZN(n15621) );
  AOI22_X1 U18873 ( .A1(n19980), .A2(P2_EBX_REG_29__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_29__SCAN_IN), .ZN(n15620) );
  OAI211_X1 U18874 ( .C1(n15968), .C2(n16232), .A(n15621), .B(n15620), .ZN(
        n15622) );
  OAI21_X1 U18875 ( .B1(n16494), .B2(n19983), .A(n15623), .ZN(P2_U2826) );
  INV_X1 U18876 ( .A(n16105), .ZN(n15633) );
  AOI22_X1 U18877 ( .A1(n19980), .A2(P2_EBX_REG_28__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_28__SCAN_IN), .ZN(n15625) );
  NAND2_X1 U18878 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15624) );
  OAI211_X1 U18879 ( .C1(n15626), .C2(n12363), .A(n15625), .B(n15624), .ZN(
        n15631) );
  OAI21_X1 U18880 ( .B1(n15627), .B2(n15628), .A(n19994), .ZN(n15629) );
  AOI21_X1 U18881 ( .B1(n15969), .B2(n15629), .A(n9804), .ZN(n15630) );
  AOI211_X1 U18882 ( .C1(n12388), .C2(n16003), .A(n15631), .B(n15630), .ZN(
        n15632) );
  OAI21_X1 U18883 ( .B1(n15633), .B2(n19983), .A(n15632), .ZN(P2_U2827) );
  INV_X1 U18884 ( .A(n15634), .ZN(n15648) );
  INV_X1 U18885 ( .A(n15635), .ZN(n15636) );
  OAI21_X1 U18886 ( .B1(n15648), .B2(n15636), .A(n19994), .ZN(n15637) );
  AOI21_X1 U18887 ( .B1(n15969), .B2(n15637), .A(n15627), .ZN(n15642) );
  AOI22_X1 U18888 ( .A1(n19980), .A2(P2_EBX_REG_27__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_27__SCAN_IN), .ZN(n15639) );
  NAND2_X1 U18889 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15638) );
  OAI211_X1 U18890 ( .C1(n15640), .C2(n12363), .A(n15639), .B(n15638), .ZN(
        n15641) );
  AOI211_X1 U18891 ( .C1(n16009), .C2(n12388), .A(n15642), .B(n15641), .ZN(
        n15643) );
  OAI21_X1 U18892 ( .B1(n16111), .B2(n19983), .A(n15643), .ZN(P2_U2828) );
  OAI21_X1 U18893 ( .B1(n15644), .B2(n15645), .A(n12248), .ZN(n16504) );
  NOR2_X1 U18894 ( .A1(n15667), .A2(n15646), .ZN(n15647) );
  OR2_X1 U18895 ( .A1(n12019), .A2(n15647), .ZN(n16246) );
  INV_X1 U18896 ( .A(n16246), .ZN(n16502) );
  OAI21_X1 U18897 ( .B1(n15662), .B2(n16241), .A(n19994), .ZN(n15649) );
  AOI21_X1 U18898 ( .B1(n15969), .B2(n15649), .A(n15648), .ZN(n15655) );
  OAI211_X1 U18899 ( .C1(n15650), .C2(n11842), .A(n15651), .B(n15984), .ZN(
        n15653) );
  AOI22_X1 U18900 ( .A1(n19980), .A2(P2_EBX_REG_26__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_26__SCAN_IN), .ZN(n15652) );
  OAI211_X1 U18901 ( .C1(n15968), .C2(n16242), .A(n15653), .B(n15652), .ZN(
        n15654) );
  AOI211_X1 U18902 ( .C1(n16502), .C2(n12388), .A(n15655), .B(n15654), .ZN(
        n15656) );
  OAI21_X1 U18903 ( .B1(n16504), .B2(n19983), .A(n15656), .ZN(P2_U2829) );
  INV_X1 U18904 ( .A(n15644), .ZN(n15658) );
  OAI21_X1 U18905 ( .B1(n15657), .B2(n15659), .A(n15658), .ZN(n16516) );
  INV_X1 U18906 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U18907 ( .A1(n15681), .A2(n16249), .ZN(n15660) );
  AOI21_X1 U18908 ( .B1(n15660), .B2(n19994), .A(n15981), .ZN(n15661) );
  OR2_X1 U18909 ( .A1(n15662), .A2(n15661), .ZN(n15664) );
  AOI22_X1 U18910 ( .A1(n19980), .A2(P2_EBX_REG_25__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_25__SCAN_IN), .ZN(n15663) );
  OAI211_X1 U18911 ( .C1(n15968), .C2(n16251), .A(n15664), .B(n15663), .ZN(
        n15669) );
  AND2_X1 U18912 ( .A1(n15678), .A2(n15665), .ZN(n15666) );
  NOR2_X1 U18913 ( .A1(n15667), .A2(n15666), .ZN(n16519) );
  INV_X1 U18914 ( .A(n16519), .ZN(n16025) );
  NOR2_X1 U18915 ( .A1(n16025), .A2(n19987), .ZN(n15668) );
  AOI211_X1 U18916 ( .C1(n15984), .C2(n15670), .A(n15669), .B(n15668), .ZN(
        n15671) );
  OAI21_X1 U18917 ( .B1(n16516), .B2(n19983), .A(n15671), .ZN(P2_U2830) );
  INV_X1 U18918 ( .A(n15672), .ZN(n15693) );
  AND2_X1 U18919 ( .A1(n15693), .A2(n15673), .ZN(n15674) );
  NOR2_X1 U18920 ( .A1(n15657), .A2(n15674), .ZN(n16529) );
  INV_X1 U18921 ( .A(n16529), .ZN(n15689) );
  NAND2_X1 U18922 ( .A1(n15675), .A2(n15676), .ZN(n15677) );
  AND2_X1 U18923 ( .A1(n15678), .A2(n15677), .ZN(n16528) );
  NOR2_X1 U18924 ( .A1(n15679), .A2(n12363), .ZN(n15687) );
  AOI21_X1 U18925 ( .B1(n15680), .B2(n10316), .A(n16947), .ZN(n15682) );
  OAI21_X1 U18926 ( .B1(n15682), .B2(n15981), .A(n15681), .ZN(n15685) );
  AOI22_X1 U18927 ( .A1(n19980), .A2(P2_EBX_REG_24__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_24__SCAN_IN), .ZN(n15684) );
  NAND2_X1 U18928 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15683) );
  NAND3_X1 U18929 ( .A1(n15685), .A2(n15684), .A3(n15683), .ZN(n15686) );
  AOI211_X1 U18930 ( .C1(n16528), .C2(n12388), .A(n15687), .B(n15686), .ZN(
        n15688) );
  OAI21_X1 U18931 ( .B1(n15689), .B2(n19983), .A(n15688), .ZN(P2_U2831) );
  NAND2_X1 U18932 ( .A1(n15690), .A2(n15691), .ZN(n15692) );
  AND2_X1 U18933 ( .A1(n15693), .A2(n15692), .ZN(n16549) );
  INV_X1 U18934 ( .A(n16549), .ZN(n15706) );
  INV_X1 U18935 ( .A(n15694), .ZN(n16272) );
  AOI21_X1 U18936 ( .B1(n15695), .B2(n16272), .A(n16947), .ZN(n15696) );
  OAI21_X1 U18937 ( .B1(n15696), .B2(n15981), .A(n15680), .ZN(n15699) );
  AOI22_X1 U18938 ( .A1(n19980), .A2(P2_EBX_REG_23__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_23__SCAN_IN), .ZN(n15698) );
  NAND2_X1 U18939 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15697) );
  NAND3_X1 U18940 ( .A1(n15699), .A2(n15698), .A3(n15697), .ZN(n15703) );
  OR2_X1 U18941 ( .A1(n9839), .A2(n15700), .ZN(n15701) );
  NAND2_X1 U18942 ( .A1(n15675), .A2(n15701), .ZN(n16546) );
  NOR2_X1 U18943 ( .A1(n16546), .A2(n19987), .ZN(n15702) );
  AOI211_X1 U18944 ( .C1(n15984), .C2(n15704), .A(n15703), .B(n15702), .ZN(
        n15705) );
  OAI21_X1 U18945 ( .B1(n15706), .B2(n19983), .A(n15705), .ZN(P2_U2832) );
  OAI21_X1 U18946 ( .B1(n12436), .B2(n15707), .A(n15690), .ZN(n16558) );
  NOR2_X1 U18947 ( .A1(n9839), .A2(n10738), .ZN(n16561) );
  XOR2_X1 U18948 ( .A(n16286), .B(n15710), .Z(n15713) );
  AOI22_X1 U18949 ( .A1(n19980), .A2(P2_EBX_REG_22__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_22__SCAN_IN), .ZN(n15711) );
  OAI21_X1 U18950 ( .B1(n15968), .B2(n16283), .A(n15711), .ZN(n15712) );
  AOI21_X1 U18951 ( .B1(n15713), .B2(n19994), .A(n15712), .ZN(n15714) );
  OAI21_X1 U18952 ( .B1(n15715), .B2(n12363), .A(n15714), .ZN(n15716) );
  AOI21_X1 U18953 ( .B1(n16561), .B2(n12388), .A(n15716), .ZN(n15717) );
  OAI21_X1 U18954 ( .B1(n16558), .B2(n19983), .A(n15717), .ZN(P2_U2833) );
  INV_X1 U18955 ( .A(n16157), .ZN(n15728) );
  NAND2_X1 U18956 ( .A1(n15967), .A2(n15718), .ZN(n15741) );
  XOR2_X1 U18957 ( .A(n15719), .B(n15741), .Z(n15724) );
  INV_X1 U18958 ( .A(n19980), .ZN(n15973) );
  OAI22_X1 U18959 ( .A1(n15973), .A2(n10649), .B1(n21847), .B2(n15970), .ZN(
        n15721) );
  NOR2_X1 U18960 ( .A1(n15968), .A2(n10596), .ZN(n15720) );
  AOI211_X1 U18961 ( .C1(n15722), .C2(n15984), .A(n15721), .B(n15720), .ZN(
        n15723) );
  OAI21_X1 U18962 ( .B1(n15724), .B2(n16947), .A(n15723), .ZN(n15725) );
  AOI21_X1 U18963 ( .B1(n15726), .B2(n12388), .A(n15725), .ZN(n15727) );
  OAI21_X1 U18964 ( .B1(n15728), .B2(n19983), .A(n15727), .ZN(P2_U2834) );
  NAND2_X1 U18965 ( .A1(n15729), .A2(n15730), .ZN(n15731) );
  AND2_X1 U18966 ( .A1(n12437), .A2(n15731), .ZN(n16577) );
  INV_X1 U18967 ( .A(n16577), .ZN(n15747) );
  AOI21_X1 U18968 ( .B1(n15734), .B2(n15732), .A(n12440), .ZN(n16566) );
  INV_X1 U18969 ( .A(n16566), .ZN(n15735) );
  NOR2_X1 U18970 ( .A1(n15735), .A2(n19987), .ZN(n15745) );
  NOR2_X1 U18971 ( .A1(n15736), .A2(n12363), .ZN(n15744) );
  NOR2_X1 U18972 ( .A1(n15969), .A2(n16297), .ZN(n15743) );
  OAI21_X1 U18973 ( .B1(n15737), .B2(n16297), .A(n19994), .ZN(n15740) );
  AOI22_X1 U18974 ( .A1(n19980), .A2(P2_EBX_REG_20__SCAN_IN), .B1(n19985), 
        .B2(P2_REIP_REG_20__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U18975 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15738) );
  OAI211_X1 U18976 ( .C1(n15741), .C2(n15740), .A(n15739), .B(n15738), .ZN(
        n15742) );
  NOR4_X1 U18977 ( .A1(n15745), .A2(n15744), .A3(n15743), .A4(n15742), .ZN(
        n15746) );
  OAI21_X1 U18978 ( .B1(n15747), .B2(n19983), .A(n15746), .ZN(P2_U2835) );
  INV_X1 U18979 ( .A(n15729), .ZN(n15750) );
  AOI21_X1 U18980 ( .B1(n15751), .B2(n15749), .A(n15750), .ZN(n16580) );
  INV_X1 U18981 ( .A(n16580), .ZN(n16173) );
  OAI21_X1 U18982 ( .B1(n15752), .B2(n15753), .A(n15732), .ZN(n16587) );
  INV_X1 U18983 ( .A(n16587), .ZN(n15765) );
  INV_X1 U18984 ( .A(n15755), .ZN(n15754) );
  NOR2_X1 U18985 ( .A1(n15991), .A2(n15754), .ZN(n15757) );
  OAI21_X1 U18986 ( .B1(n15755), .B2(n16947), .A(n15969), .ZN(n15756) );
  MUX2_X1 U18987 ( .A(n15757), .B(n15756), .S(n16308), .Z(n15764) );
  NAND2_X1 U18988 ( .A1(n15758), .A2(n15984), .ZN(n15762) );
  NAND2_X1 U18989 ( .A1(n19980), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15759) );
  OAI211_X1 U18990 ( .C1(n20718), .C2(n15970), .A(n15759), .B(n16464), .ZN(
        n15760) );
  INV_X1 U18991 ( .A(n15760), .ZN(n15761) );
  OAI211_X1 U18992 ( .C1(n15968), .C2(n16306), .A(n15762), .B(n15761), .ZN(
        n15763) );
  AOI211_X1 U18993 ( .C1(n15765), .C2(n12388), .A(n15764), .B(n15763), .ZN(
        n15766) );
  OAI21_X1 U18994 ( .B1(n16173), .B2(n19983), .A(n15766), .ZN(P2_U2836) );
  OR2_X1 U18995 ( .A1(n15768), .A2(n15767), .ZN(n15769) );
  AND2_X1 U18996 ( .A1(n15749), .A2(n15769), .ZN(n16599) );
  INV_X1 U18997 ( .A(n16599), .ZN(n15786) );
  AND2_X1 U18998 ( .A1(n15771), .A2(n15770), .ZN(n15772) );
  OR2_X1 U18999 ( .A1(n15772), .A2(n15752), .ZN(n16602) );
  INV_X1 U19000 ( .A(n16602), .ZN(n15784) );
  NAND2_X1 U19001 ( .A1(n15773), .A2(n15984), .ZN(n15777) );
  NAND2_X1 U19002 ( .A1(n19980), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n15774) );
  OAI211_X1 U19003 ( .C1(n12228), .C2(n15970), .A(n15774), .B(n16464), .ZN(
        n15775) );
  INV_X1 U19004 ( .A(n15775), .ZN(n15776) );
  OAI211_X1 U19005 ( .C1(n15968), .C2(n16316), .A(n15777), .B(n15776), .ZN(
        n15783) );
  INV_X1 U19006 ( .A(n15779), .ZN(n15778) );
  NOR2_X1 U19007 ( .A1(n15991), .A2(n15778), .ZN(n15781) );
  OAI21_X1 U19008 ( .B1(n15779), .B2(n16947), .A(n15969), .ZN(n15780) );
  MUX2_X1 U19009 ( .A(n15781), .B(n15780), .S(n16318), .Z(n15782) );
  AOI211_X1 U19010 ( .C1(n15784), .C2(n12388), .A(n15783), .B(n15782), .ZN(
        n15785) );
  OAI21_X1 U19011 ( .B1(n15786), .B2(n19983), .A(n15785), .ZN(P2_U2837) );
  INV_X1 U19012 ( .A(n16324), .ZN(n16068) );
  AOI21_X1 U19013 ( .B1(n19980), .B2(P2_EBX_REG_17__SCAN_IN), .A(n16754), .ZN(
        n15788) );
  NAND2_X1 U19014 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15787) );
  OAI211_X1 U19015 ( .C1(n15970), .C2(n20715), .A(n15788), .B(n15787), .ZN(
        n15793) );
  NOR2_X1 U19016 ( .A1(n10319), .A2(n15789), .ZN(n15790) );
  XOR2_X1 U19017 ( .A(n16328), .B(n15790), .Z(n15791) );
  NOR2_X1 U19018 ( .A1(n15791), .A2(n16947), .ZN(n15792) );
  AOI211_X1 U19019 ( .C1(n15984), .C2(n15794), .A(n15793), .B(n15792), .ZN(
        n15796) );
  NAND2_X1 U19020 ( .A1(n16187), .A2(n15982), .ZN(n15795) );
  OAI211_X1 U19021 ( .C1(n19987), .C2(n16068), .A(n15796), .B(n15795), .ZN(
        P2_U2838) );
  INV_X1 U19022 ( .A(n16199), .ZN(n15810) );
  INV_X1 U19023 ( .A(n16079), .ZN(n16337) );
  AOI21_X1 U19024 ( .B1(n19980), .B2(P2_EBX_REG_16__SCAN_IN), .A(n16754), .ZN(
        n15797) );
  OAI21_X1 U19025 ( .B1(n15798), .B2(n15970), .A(n15797), .ZN(n15799) );
  AOI21_X1 U19026 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19981), .A(
        n15799), .ZN(n15800) );
  OAI21_X1 U19027 ( .B1(n15801), .B2(n12363), .A(n15800), .ZN(n15808) );
  INV_X1 U19028 ( .A(n15803), .ZN(n15802) );
  NOR2_X1 U19029 ( .A1(n15991), .A2(n15802), .ZN(n15806) );
  OAI21_X1 U19030 ( .B1(n15803), .B2(n16947), .A(n15969), .ZN(n15805) );
  MUX2_X1 U19031 ( .A(n15806), .B(n15805), .S(n15804), .Z(n15807) );
  AOI211_X1 U19032 ( .C1(n12388), .C2(n16337), .A(n15808), .B(n15807), .ZN(
        n15809) );
  OAI21_X1 U19033 ( .B1(n15810), .B2(n19983), .A(n15809), .ZN(P2_U2839) );
  NAND2_X1 U19034 ( .A1(n15951), .A2(n15811), .ZN(n15814) );
  INV_X1 U19035 ( .A(n15811), .ZN(n15812) );
  AOI21_X1 U19036 ( .B1(n15812), .B2(n19994), .A(n15981), .ZN(n15813) );
  MUX2_X1 U19037 ( .A(n15814), .B(n15813), .S(n16348), .Z(n15824) );
  NOR2_X1 U19038 ( .A1(n15815), .A2(n15816), .ZN(n15817) );
  OR2_X1 U19039 ( .A1(n14698), .A2(n15817), .ZN(n16611) );
  INV_X1 U19040 ( .A(n16611), .ZN(n16081) );
  OAI21_X1 U19041 ( .B1(n20712), .B2(n15970), .A(n16464), .ZN(n15819) );
  NOR2_X1 U19042 ( .A1(n15973), .A2(n11786), .ZN(n15818) );
  AOI211_X1 U19043 ( .C1(n19981), .C2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15819), .B(n15818), .ZN(n15820) );
  OAI21_X1 U19044 ( .B1(n15821), .B2(n12363), .A(n15820), .ZN(n15822) );
  AOI21_X1 U19045 ( .B1(n16081), .B2(n12388), .A(n15822), .ZN(n15823) );
  OAI211_X1 U19046 ( .C1(n19983), .C2(n16607), .A(n15824), .B(n15823), .ZN(
        P2_U2840) );
  INV_X1 U19047 ( .A(n15825), .ZN(n15826) );
  AOI21_X1 U19048 ( .B1(n15826), .B2(n19994), .A(n15981), .ZN(n15827) );
  MUX2_X1 U19049 ( .A(n15828), .B(n15827), .S(n16357), .Z(n15839) );
  AND2_X1 U19050 ( .A1(n13395), .A2(n15829), .ZN(n15830) );
  NOR2_X1 U19051 ( .A1(n15815), .A2(n15830), .ZN(n16621) );
  NAND2_X1 U19052 ( .A1(n15831), .A2(n15984), .ZN(n15836) );
  NAND2_X1 U19053 ( .A1(n19980), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15832) );
  OAI211_X1 U19054 ( .C1(n15833), .C2(n15970), .A(n15832), .B(n16464), .ZN(
        n15834) );
  INV_X1 U19055 ( .A(n15834), .ZN(n15835) );
  OAI211_X1 U19056 ( .C1(n15968), .C2(n16359), .A(n15836), .B(n15835), .ZN(
        n15837) );
  AOI21_X1 U19057 ( .B1(n16621), .B2(n12388), .A(n15837), .ZN(n15838) );
  OAI211_X1 U19058 ( .C1(n19983), .C2(n16624), .A(n15839), .B(n15838), .ZN(
        P2_U2841) );
  OAI22_X1 U19059 ( .A1(n15840), .A2(n12363), .B1(n15973), .B2(n21785), .ZN(
        n15841) );
  INV_X1 U19060 ( .A(n15841), .ZN(n15842) );
  OAI211_X1 U19061 ( .C1(n20708), .C2(n15970), .A(n15842), .B(n16464), .ZN(
        n15843) );
  AOI21_X1 U19062 ( .B1(n19981), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15843), .ZN(n15844) );
  OAI21_X1 U19063 ( .B1(n16648), .B2(n19987), .A(n15844), .ZN(n15850) );
  INV_X1 U19064 ( .A(n15846), .ZN(n15845) );
  NOR2_X1 U19065 ( .A1(n15991), .A2(n15845), .ZN(n15848) );
  OAI21_X1 U19066 ( .B1(n15846), .B2(n16947), .A(n15969), .ZN(n15847) );
  MUX2_X1 U19067 ( .A(n15848), .B(n15847), .S(n16382), .Z(n15849) );
  AOI211_X1 U19068 ( .C1(n16651), .C2(n15982), .A(n15850), .B(n15849), .ZN(
        n15851) );
  INV_X1 U19069 ( .A(n15851), .ZN(P2_U2843) );
  NAND2_X1 U19070 ( .A1(n15951), .A2(n15852), .ZN(n15855) );
  INV_X1 U19071 ( .A(n15852), .ZN(n15853) );
  AOI21_X1 U19072 ( .B1(n15853), .B2(n19994), .A(n15981), .ZN(n15854) );
  MUX2_X1 U19073 ( .A(n15855), .B(n15854), .S(n16395), .Z(n15862) );
  OAI21_X1 U19074 ( .B1(n21738), .B2(n15970), .A(n16464), .ZN(n15857) );
  NOR2_X1 U19075 ( .A1(n15968), .A2(n16397), .ZN(n15856) );
  AOI211_X1 U19076 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19980), .A(n15857), .B(
        n15856), .ZN(n15858) );
  OAI21_X1 U19077 ( .B1(n15859), .B2(n12363), .A(n15858), .ZN(n15860) );
  AOI21_X1 U19078 ( .B1(n16664), .B2(n12388), .A(n15860), .ZN(n15861) );
  OAI211_X1 U19079 ( .C1(n19983), .C2(n16661), .A(n15862), .B(n15861), .ZN(
        P2_U2844) );
  AOI21_X1 U19080 ( .B1(n15863), .B2(n19994), .A(n15981), .ZN(n15866) );
  INV_X1 U19081 ( .A(n15863), .ZN(n15864) );
  NAND2_X1 U19082 ( .A1(n15951), .A2(n15864), .ZN(n15865) );
  MUX2_X1 U19083 ( .A(n15866), .B(n15865), .S(n16404), .Z(n15873) );
  AOI22_X1 U19084 ( .A1(n15867), .A2(n15984), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19981), .ZN(n15868) );
  OAI211_X1 U19085 ( .C1(n20705), .C2(n15970), .A(n15868), .B(n16464), .ZN(
        n15869) );
  AOI21_X1 U19086 ( .B1(n19980), .B2(P2_EBX_REG_10__SCAN_IN), .A(n15869), .ZN(
        n15872) );
  NAND2_X1 U19087 ( .A1(n16677), .A2(n15982), .ZN(n15871) );
  NAND2_X1 U19088 ( .A1(n16676), .A2(n12388), .ZN(n15870) );
  NAND4_X1 U19089 ( .A1(n15873), .A2(n15872), .A3(n15871), .A4(n15870), .ZN(
        P2_U2845) );
  NOR2_X1 U19090 ( .A1(n10319), .A2(n15874), .ZN(n15875) );
  XNOR2_X1 U19091 ( .A(n15875), .B(n16413), .ZN(n15876) );
  NAND2_X1 U19092 ( .A1(n15876), .A2(n19994), .ZN(n15885) );
  INV_X1 U19093 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21860) );
  NAND2_X1 U19094 ( .A1(n15877), .A2(n15984), .ZN(n15882) );
  NAND2_X1 U19095 ( .A1(n19980), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n15878) );
  OAI211_X1 U19096 ( .C1(n15879), .C2(n15970), .A(n15878), .B(n16464), .ZN(
        n15880) );
  INV_X1 U19097 ( .A(n15880), .ZN(n15881) );
  OAI211_X1 U19098 ( .C1(n15968), .C2(n21860), .A(n15882), .B(n15881), .ZN(
        n15883) );
  AOI21_X1 U19099 ( .B1(n16689), .B2(n12388), .A(n15883), .ZN(n15884) );
  OAI211_X1 U19100 ( .C1(n16691), .C2(n19983), .A(n15885), .B(n15884), .ZN(
        P2_U2846) );
  NAND2_X1 U19101 ( .A1(n15951), .A2(n15886), .ZN(n15890) );
  INV_X1 U19102 ( .A(n15886), .ZN(n15887) );
  AOI21_X1 U19103 ( .B1(n15887), .B2(n19994), .A(n15981), .ZN(n15889) );
  MUX2_X1 U19104 ( .A(n15890), .B(n15889), .S(n15888), .Z(n15899) );
  INV_X1 U19105 ( .A(n16707), .ZN(n15897) );
  NAND2_X1 U19106 ( .A1(n19980), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n15891) );
  OAI211_X1 U19107 ( .C1(n20702), .C2(n15970), .A(n15891), .B(n16464), .ZN(
        n15892) );
  INV_X1 U19108 ( .A(n15892), .ZN(n15894) );
  NAND2_X1 U19109 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15893) );
  OAI211_X1 U19110 ( .C1(n15895), .C2(n12363), .A(n15894), .B(n15893), .ZN(
        n15896) );
  AOI21_X1 U19111 ( .B1(n15897), .B2(n12388), .A(n15896), .ZN(n15898) );
  OAI211_X1 U19112 ( .C1(n19983), .C2(n15900), .A(n15899), .B(n15898), .ZN(
        P2_U2847) );
  NAND2_X1 U19113 ( .A1(n15951), .A2(n15901), .ZN(n15904) );
  INV_X1 U19114 ( .A(n15901), .ZN(n15902) );
  AOI21_X1 U19115 ( .B1(n15902), .B2(n19994), .A(n15981), .ZN(n15903) );
  MUX2_X1 U19116 ( .A(n15904), .B(n15903), .S(n16440), .Z(n15911) );
  AOI22_X1 U19117 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n15984), .B2(n15905), .ZN(n15906) );
  OAI211_X1 U19118 ( .C1(n20700), .C2(n15970), .A(n15906), .B(n16464), .ZN(
        n15907) );
  AOI21_X1 U19119 ( .B1(n19980), .B2(P2_EBX_REG_7__SCAN_IN), .A(n15907), .ZN(
        n15908) );
  OAI21_X1 U19120 ( .B1(n16719), .B2(n19987), .A(n15908), .ZN(n15909) );
  INV_X1 U19121 ( .A(n15909), .ZN(n15910) );
  OAI211_X1 U19122 ( .C1(n16715), .C2(n19983), .A(n15911), .B(n15910), .ZN(
        P2_U2848) );
  AOI21_X1 U19123 ( .B1(n15912), .B2(n19994), .A(n15981), .ZN(n15914) );
  NAND2_X1 U19124 ( .A1(n15951), .A2(n10345), .ZN(n15913) );
  MUX2_X1 U19125 ( .A(n15914), .B(n15913), .S(n16447), .Z(n15921) );
  OAI21_X1 U19126 ( .B1(n20698), .B2(n15970), .A(n16464), .ZN(n15916) );
  NOR2_X1 U19127 ( .A1(n15973), .A2(n11706), .ZN(n15915) );
  AOI211_X1 U19128 ( .C1(n19981), .C2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15916), .B(n15915), .ZN(n15917) );
  OAI21_X1 U19129 ( .B1(n15918), .B2(n12363), .A(n15917), .ZN(n15919) );
  AOI21_X1 U19130 ( .B1(n16727), .B2(n12388), .A(n15919), .ZN(n15920) );
  OAI211_X1 U19131 ( .C1(n15922), .C2(n19983), .A(n15921), .B(n15920), .ZN(
        P2_U2849) );
  NAND2_X1 U19132 ( .A1(n15967), .A2(n19993), .ZN(n15923) );
  XOR2_X1 U19133 ( .A(n17585), .B(n15923), .Z(n15937) );
  INV_X1 U19134 ( .A(n17590), .ZN(n15931) );
  NAND2_X1 U19135 ( .A1(n19980), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n15924) );
  OAI211_X1 U19136 ( .C1(n15925), .C2(n15970), .A(n15924), .B(n16464), .ZN(
        n15926) );
  INV_X1 U19137 ( .A(n15926), .ZN(n15928) );
  NAND2_X1 U19138 ( .A1(n19981), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15927) );
  OAI211_X1 U19139 ( .C1(n12363), .C2(n15929), .A(n15928), .B(n15927), .ZN(
        n15930) );
  AOI21_X1 U19140 ( .B1(n15931), .B2(n12388), .A(n15930), .ZN(n15936) );
  INV_X1 U19141 ( .A(n15933), .ZN(n15934) );
  XNOR2_X1 U19142 ( .A(n15932), .B(n15934), .ZN(n16753) );
  NAND2_X1 U19143 ( .A1(n16753), .A2(n15982), .ZN(n15935) );
  OAI211_X1 U19144 ( .C1(n15937), .C2(n16947), .A(n15936), .B(n15935), .ZN(
        P2_U2850) );
  AOI21_X1 U19145 ( .B1(n15938), .B2(n19994), .A(n15981), .ZN(n15942) );
  INV_X1 U19146 ( .A(n15938), .ZN(n15939) );
  NAND2_X1 U19147 ( .A1(n15951), .A2(n15939), .ZN(n15941) );
  MUX2_X1 U19148 ( .A(n15942), .B(n15941), .S(n15940), .Z(n15950) );
  NOR2_X1 U19149 ( .A1(n12363), .A2(n15943), .ZN(n15946) );
  OAI22_X1 U19150 ( .A1(n15973), .A2(n15944), .B1(n11505), .B2(n15970), .ZN(
        n15945) );
  AOI211_X1 U19151 ( .C1(n19981), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15946), .B(n15945), .ZN(n15947) );
  OAI21_X1 U19152 ( .B1(n19983), .B2(n16203), .A(n15947), .ZN(n15948) );
  OAI211_X1 U19153 ( .C1(n20751), .C2(n19988), .A(n15950), .B(n15949), .ZN(
        P2_U2852) );
  AOI21_X1 U19154 ( .B1(n15965), .B2(n19994), .A(n15981), .ZN(n15954) );
  NAND2_X1 U19155 ( .A1(n15951), .A2(n10320), .ZN(n15953) );
  MUX2_X1 U19156 ( .A(n15954), .B(n15953), .S(n15952), .Z(n15962) );
  NAND2_X1 U19157 ( .A1(n20760), .A2(n15982), .ZN(n15958) );
  OAI22_X1 U19158 ( .A1(n15973), .A2(n15955), .B1(n20694), .B2(n15970), .ZN(
        n15956) );
  AOI21_X1 U19159 ( .B1(n19981), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n15956), .ZN(n15957) );
  OAI211_X1 U19160 ( .C1(n12363), .C2(n15959), .A(n15958), .B(n15957), .ZN(
        n15960) );
  AOI21_X1 U19161 ( .B1(n10215), .B2(n12388), .A(n15960), .ZN(n15961) );
  OAI211_X1 U19162 ( .C1(n19988), .C2(n16856), .A(n15962), .B(n15961), .ZN(
        P2_U2853) );
  AND2_X1 U19163 ( .A1(n15963), .A2(n16778), .ZN(n15964) );
  NOR2_X1 U19164 ( .A1(n15965), .A2(n15964), .ZN(n15966) );
  NAND2_X1 U19165 ( .A1(n15967), .A2(n15966), .ZN(n16785) );
  MUX2_X1 U19166 ( .A(n15969), .B(n15968), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n15980) );
  NOR2_X1 U19167 ( .A1(n15970), .A2(n20692), .ZN(n15975) );
  OAI22_X1 U19168 ( .A1(n15973), .A2(n15972), .B1(n12363), .B2(n15971), .ZN(
        n15974) );
  AOI211_X1 U19169 ( .C1(n15982), .C2(n20772), .A(n15975), .B(n15974), .ZN(
        n15976) );
  OAI21_X1 U19170 ( .B1(n15977), .B2(n19987), .A(n15976), .ZN(n15978) );
  AOI21_X1 U19171 ( .B1(n20769), .B2(n15988), .A(n15978), .ZN(n15979) );
  OAI211_X1 U19172 ( .C1(n16785), .C2(n16947), .A(n15980), .B(n15979), .ZN(
        P2_U2854) );
  INV_X1 U19173 ( .A(n16778), .ZN(n15992) );
  OAI21_X1 U19174 ( .B1(n15981), .B2(n19981), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15990) );
  AOI22_X1 U19175 ( .A1(n19980), .A2(P2_EBX_REG_0__SCAN_IN), .B1(n15982), .B2(
        n17607), .ZN(n15986) );
  AOI22_X1 U19176 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(n19985), .B1(n15984), 
        .B2(n15983), .ZN(n15985) );
  OAI211_X1 U19177 ( .C1(n10204), .C2(n19987), .A(n15986), .B(n15985), .ZN(
        n15987) );
  AOI21_X1 U19178 ( .B1(n16855), .B2(n15988), .A(n15987), .ZN(n15989) );
  OAI211_X1 U19179 ( .C1(n15992), .C2(n15991), .A(n15990), .B(n15989), .ZN(
        P2_U2855) );
  MUX2_X1 U19180 ( .A(n15993), .B(P2_EBX_REG_31__SCAN_IN), .S(n16078), .Z(
        P2_U2856) );
  INV_X1 U19181 ( .A(n16493), .ZN(n15998) );
  NAND3_X1 U19182 ( .A1(n16092), .A2(n15995), .A3(n16086), .ZN(n15997) );
  NAND2_X1 U19183 ( .A1(n16078), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15996) );
  OAI211_X1 U19184 ( .C1(n16078), .C2(n15998), .A(n15997), .B(n15996), .ZN(
        P2_U2858) );
  NOR2_X1 U19185 ( .A1(n16000), .A2(n15999), .ZN(n16002) );
  XNOR2_X1 U19186 ( .A(n16002), .B(n16001), .ZN(n16107) );
  NAND2_X1 U19187 ( .A1(n16078), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16005) );
  NAND2_X1 U19188 ( .A1(n16003), .A2(n16080), .ZN(n16004) );
  OAI211_X1 U19189 ( .C1(n16107), .C2(n16072), .A(n16005), .B(n16004), .ZN(
        P2_U2859) );
  OAI21_X1 U19190 ( .B1(n16006), .B2(n16008), .A(n16007), .ZN(n16115) );
  NAND2_X1 U19191 ( .A1(n16070), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n16011) );
  NAND2_X1 U19192 ( .A1(n16009), .A2(n16080), .ZN(n16010) );
  OAI211_X1 U19193 ( .C1(n16115), .C2(n16072), .A(n16011), .B(n16010), .ZN(
        P2_U2860) );
  NOR2_X1 U19194 ( .A1(n16012), .A2(n16022), .ZN(n16021) );
  NOR2_X1 U19195 ( .A1(n16021), .A2(n16013), .ZN(n16018) );
  NOR2_X1 U19196 ( .A1(n16887), .A2(n16014), .ZN(n16015) );
  XNOR2_X1 U19197 ( .A(n16016), .B(n16015), .ZN(n16017) );
  XNOR2_X1 U19198 ( .A(n16018), .B(n16017), .ZN(n16122) );
  NOR2_X1 U19199 ( .A1(n16246), .A2(n16070), .ZN(n16019) );
  AOI21_X1 U19200 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16070), .A(n16019), .ZN(
        n16020) );
  OAI21_X1 U19201 ( .B1(n16122), .B2(n16072), .A(n16020), .ZN(P2_U2861) );
  AOI21_X1 U19202 ( .B1(n16012), .B2(n16022), .A(n16021), .ZN(n16123) );
  NAND2_X1 U19203 ( .A1(n16123), .A2(n16086), .ZN(n16024) );
  NAND2_X1 U19204 ( .A1(n16070), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16023) );
  OAI211_X1 U19205 ( .C1(n16025), .C2(n16078), .A(n16024), .B(n16023), .ZN(
        P2_U2862) );
  INV_X1 U19206 ( .A(n16026), .ZN(n16027) );
  XOR2_X1 U19207 ( .A(n16030), .B(n16027), .Z(n16040) );
  NAND2_X1 U19208 ( .A1(n16029), .A2(n16028), .ZN(n16039) );
  NOR2_X1 U19209 ( .A1(n16040), .A2(n16039), .ZN(n16038) );
  AOI21_X1 U19210 ( .B1(n16026), .B2(n16030), .A(n16038), .ZN(n16034) );
  XNOR2_X1 U19211 ( .A(n16032), .B(n16031), .ZN(n16033) );
  XNOR2_X1 U19212 ( .A(n16034), .B(n16033), .ZN(n16136) );
  NOR2_X1 U19213 ( .A1(n16080), .A2(n16035), .ZN(n16036) );
  AOI21_X1 U19214 ( .B1(n16528), .B2(n16080), .A(n16036), .ZN(n16037) );
  OAI21_X1 U19215 ( .B1(n16136), .B2(n16072), .A(n16037), .ZN(P2_U2863) );
  AOI21_X1 U19216 ( .B1(n16040), .B2(n16039), .A(n16038), .ZN(n16137) );
  NAND2_X1 U19217 ( .A1(n16137), .A2(n16086), .ZN(n16042) );
  NAND2_X1 U19218 ( .A1(n16078), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n16041) );
  OAI211_X1 U19219 ( .C1(n16546), .C2(n16078), .A(n16042), .B(n16041), .ZN(
        P2_U2864) );
  NAND2_X1 U19220 ( .A1(n9863), .A2(n16043), .ZN(n16044) );
  NAND2_X1 U19221 ( .A1(n16027), .A2(n16044), .ZN(n16152) );
  NAND2_X1 U19222 ( .A1(n16561), .A2(n16080), .ZN(n16046) );
  NAND2_X1 U19223 ( .A1(n16070), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16045) );
  OAI211_X1 U19224 ( .C1(n16152), .C2(n16072), .A(n16046), .B(n16045), .ZN(
        P2_U2865) );
  OAI21_X1 U19225 ( .B1(n16051), .B2(n16047), .A(n9863), .ZN(n16159) );
  NOR2_X1 U19226 ( .A1(n16048), .A2(n16070), .ZN(n16049) );
  AOI21_X1 U19227 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n16078), .A(n16049), .ZN(
        n16050) );
  OAI21_X1 U19228 ( .B1(n16072), .B2(n16159), .A(n16050), .ZN(P2_U2866) );
  INV_X1 U19229 ( .A(n16051), .ZN(n16052) );
  OAI21_X1 U19230 ( .B1(n16057), .B2(n16053), .A(n16052), .ZN(n16165) );
  NOR2_X1 U19231 ( .A1(n16080), .A2(n11763), .ZN(n16054) );
  AOI21_X1 U19232 ( .B1(n16566), .B2(n16080), .A(n16054), .ZN(n16055) );
  OAI21_X1 U19233 ( .B1(n16072), .B2(n16165), .A(n16055), .ZN(P2_U2867) );
  AOI21_X1 U19234 ( .B1(n16058), .B2(n16056), .A(n16057), .ZN(n16170) );
  NAND2_X1 U19235 ( .A1(n16170), .A2(n16086), .ZN(n16060) );
  NAND2_X1 U19236 ( .A1(n16078), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n16059) );
  OAI211_X1 U19237 ( .C1(n16587), .C2(n16078), .A(n16060), .B(n16059), .ZN(
        P2_U2868) );
  NAND2_X1 U19238 ( .A1(n16061), .A2(n16062), .ZN(n16063) );
  NAND2_X1 U19239 ( .A1(n16056), .A2(n16063), .ZN(n16180) );
  NOR2_X1 U19240 ( .A1(n16602), .A2(n16070), .ZN(n16064) );
  AOI21_X1 U19241 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n16078), .A(n16064), .ZN(
        n16065) );
  OAI21_X1 U19242 ( .B1(n16072), .B2(n16180), .A(n16065), .ZN(P2_U2869) );
  OAI21_X1 U19243 ( .B1(n16066), .B2(n16067), .A(n16061), .ZN(n16189) );
  NOR2_X1 U19244 ( .A1(n16068), .A2(n16070), .ZN(n16069) );
  AOI21_X1 U19245 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16070), .A(n16069), .ZN(
        n16071) );
  OAI21_X1 U19246 ( .B1(n16072), .B2(n16189), .A(n16071), .ZN(P2_U2870) );
  NOR2_X1 U19247 ( .A1(n16073), .A2(n16074), .ZN(n16075) );
  NOR2_X1 U19248 ( .A1(n16066), .A2(n16075), .ZN(n16190) );
  NAND2_X1 U19249 ( .A1(n16190), .A2(n16086), .ZN(n16077) );
  NAND2_X1 U19250 ( .A1(n16078), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n16076) );
  OAI211_X1 U19251 ( .C1(n16079), .C2(n16078), .A(n16077), .B(n16076), .ZN(
        P2_U2871) );
  NAND2_X1 U19252 ( .A1(n16081), .A2(n16080), .ZN(n16084) );
  OAI211_X1 U19253 ( .C1(n16085), .C2(n16082), .A(n10669), .B(n16086), .ZN(
        n16083) );
  OAI211_X1 U19254 ( .C1(n16080), .C2(n11786), .A(n16084), .B(n16083), .ZN(
        P2_U2872) );
  NAND2_X1 U19255 ( .A1(n16621), .A2(n16080), .ZN(n16090) );
  INV_X1 U19256 ( .A(n14351), .ZN(n16088) );
  OAI211_X1 U19257 ( .C1(n16088), .C2(n16087), .A(n10672), .B(n16086), .ZN(
        n16089) );
  OAI211_X1 U19258 ( .C1(n16080), .C2(n16091), .A(n16090), .B(n16089), .ZN(
        P2_U2873) );
  NAND3_X1 U19259 ( .A1(n16092), .A2(n15995), .A3(n20020), .ZN(n16099) );
  INV_X1 U19260 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16095) );
  AOI22_X1 U19261 ( .A1(n16193), .A2(n16093), .B1(P2_EAX_REG_29__SCAN_IN), 
        .B2(n16191), .ZN(n16094) );
  OAI21_X1 U19262 ( .B1(n16197), .B2(n16095), .A(n16094), .ZN(n16097) );
  NOR2_X1 U19263 ( .A1(n16494), .A2(n20002), .ZN(n16096) );
  NAND2_X1 U19264 ( .A1(n16099), .A2(n16098), .ZN(P2_U2890) );
  INV_X1 U19265 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16103) );
  AOI22_X1 U19266 ( .A1(n16193), .A2(n16100), .B1(P2_EAX_REG_28__SCAN_IN), 
        .B2(n16191), .ZN(n16102) );
  NAND2_X1 U19267 ( .A1(n16194), .A2(BUF2_REG_28__SCAN_IN), .ZN(n16101) );
  OAI211_X1 U19268 ( .C1(n16197), .C2(n16103), .A(n16102), .B(n16101), .ZN(
        n16104) );
  AOI21_X1 U19269 ( .B1(n16105), .B2(n20016), .A(n16104), .ZN(n16106) );
  OAI21_X1 U19270 ( .B1(n16107), .B2(n16202), .A(n16106), .ZN(P2_U2891) );
  INV_X1 U19271 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16110) );
  AOI22_X1 U19272 ( .A1(n16193), .A2(n16108), .B1(P2_EAX_REG_27__SCAN_IN), 
        .B2(n16191), .ZN(n16109) );
  OAI21_X1 U19273 ( .B1(n16197), .B2(n16110), .A(n16109), .ZN(n16113) );
  NOR2_X1 U19274 ( .A1(n16111), .A2(n20002), .ZN(n16112) );
  AOI211_X1 U19275 ( .C1(n16194), .C2(BUF2_REG_27__SCAN_IN), .A(n16113), .B(
        n16112), .ZN(n16114) );
  OAI21_X1 U19276 ( .B1(n16115), .B2(n16202), .A(n16114), .ZN(P2_U2892) );
  INV_X1 U19277 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16118) );
  AOI22_X1 U19278 ( .A1(n16193), .A2(n16116), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n16191), .ZN(n16117) );
  OAI21_X1 U19279 ( .B1(n16197), .B2(n16118), .A(n16117), .ZN(n16120) );
  NOR2_X1 U19280 ( .A1(n16504), .A2(n20002), .ZN(n16119) );
  AOI211_X1 U19281 ( .C1(n16194), .C2(BUF2_REG_26__SCAN_IN), .A(n16120), .B(
        n16119), .ZN(n16121) );
  OAI21_X1 U19282 ( .B1(n16122), .B2(n16202), .A(n16121), .ZN(P2_U2893) );
  INV_X1 U19283 ( .A(n16123), .ZN(n16129) );
  AOI22_X1 U19284 ( .A1(n16193), .A2(n16124), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n16191), .ZN(n16125) );
  OAI21_X1 U19285 ( .B1(n16197), .B2(n17626), .A(n16125), .ZN(n16127) );
  NOR2_X1 U19286 ( .A1(n16516), .A2(n20002), .ZN(n16126) );
  AOI211_X1 U19287 ( .C1(n16194), .C2(BUF2_REG_25__SCAN_IN), .A(n16127), .B(
        n16126), .ZN(n16128) );
  OAI21_X1 U19288 ( .B1(n16202), .B2(n16129), .A(n16128), .ZN(P2_U2894) );
  INV_X1 U19289 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U19290 ( .A1(n16193), .A2(n16130), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n16191), .ZN(n16132) );
  NAND2_X1 U19291 ( .A1(n16194), .A2(BUF2_REG_24__SCAN_IN), .ZN(n16131) );
  OAI211_X1 U19292 ( .C1(n16197), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16134) );
  AOI21_X1 U19293 ( .B1(n16529), .B2(n20016), .A(n16134), .ZN(n16135) );
  OAI21_X1 U19294 ( .B1(n16136), .B2(n16202), .A(n16135), .ZN(P2_U2895) );
  INV_X1 U19295 ( .A(n16137), .ZN(n16144) );
  INV_X1 U19296 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16141) );
  NAND2_X1 U19297 ( .A1(n16194), .A2(BUF2_REG_23__SCAN_IN), .ZN(n16140) );
  AOI22_X1 U19298 ( .A1(n16193), .A2(n16138), .B1(P2_EAX_REG_23__SCAN_IN), 
        .B2(n16191), .ZN(n16139) );
  OAI211_X1 U19299 ( .C1(n16141), .C2(n16197), .A(n16140), .B(n16139), .ZN(
        n16142) );
  AOI21_X1 U19300 ( .B1(n16549), .B2(n20016), .A(n16142), .ZN(n16143) );
  OAI21_X1 U19301 ( .B1(n16144), .B2(n16202), .A(n16143), .ZN(P2_U2896) );
  INV_X1 U19302 ( .A(n16558), .ZN(n16150) );
  INV_X1 U19303 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16148) );
  NAND2_X1 U19304 ( .A1(n16194), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U19305 ( .A1(n16193), .A2(n16145), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n16191), .ZN(n16146) );
  OAI211_X1 U19306 ( .C1(n16148), .C2(n16197), .A(n16147), .B(n16146), .ZN(
        n16149) );
  AOI21_X1 U19307 ( .B1(n16150), .B2(n20016), .A(n16149), .ZN(n16151) );
  OAI21_X1 U19308 ( .B1(n16202), .B2(n16152), .A(n16151), .ZN(P2_U2897) );
  INV_X1 U19309 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16155) );
  NAND2_X1 U19310 ( .A1(n16194), .A2(BUF2_REG_21__SCAN_IN), .ZN(n16154) );
  AOI22_X1 U19311 ( .A1(n16193), .A2(n20129), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n16191), .ZN(n16153) );
  OAI211_X1 U19312 ( .C1(n16155), .C2(n16197), .A(n16154), .B(n16153), .ZN(
        n16156) );
  AOI21_X1 U19313 ( .B1(n16157), .B2(n20016), .A(n16156), .ZN(n16158) );
  OAI21_X1 U19314 ( .B1(n16202), .B2(n16159), .A(n16158), .ZN(P2_U2898) );
  NOR2_X1 U19315 ( .A1(n16197), .A2(n17632), .ZN(n16163) );
  NAND2_X1 U19316 ( .A1(n16194), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16161) );
  NAND2_X1 U19317 ( .A1(n16191), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n16160) );
  OAI211_X1 U19318 ( .C1(n20124), .C2(n16184), .A(n16161), .B(n16160), .ZN(
        n16162) );
  AOI211_X1 U19319 ( .C1(n16577), .C2(n20016), .A(n16163), .B(n16162), .ZN(
        n16164) );
  OAI21_X1 U19320 ( .B1(n16202), .B2(n16165), .A(n16164), .ZN(P2_U2899) );
  INV_X1 U19321 ( .A(n16197), .ZN(n16169) );
  INV_X1 U19322 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n20055) );
  OAI22_X1 U19323 ( .A1(n20120), .A2(n16184), .B1(n20001), .B2(n20055), .ZN(
        n16168) );
  INV_X1 U19324 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16166) );
  NOR2_X1 U19325 ( .A1(n14714), .A2(n16166), .ZN(n16167) );
  AOI211_X1 U19326 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n16169), .A(n16168), .B(
        n16167), .ZN(n16172) );
  NAND2_X1 U19327 ( .A1(n16170), .A2(n20020), .ZN(n16171) );
  OAI211_X1 U19328 ( .C1(n16173), .C2(n20002), .A(n16172), .B(n16171), .ZN(
        P2_U2900) );
  INV_X1 U19329 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16177) );
  NAND2_X1 U19330 ( .A1(n16194), .A2(BUF2_REG_18__SCAN_IN), .ZN(n16176) );
  AOI22_X1 U19331 ( .A1(n16193), .A2(n16174), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n16191), .ZN(n16175) );
  OAI211_X1 U19332 ( .C1(n16177), .C2(n16197), .A(n16176), .B(n16175), .ZN(
        n16178) );
  AOI21_X1 U19333 ( .B1(n16599), .B2(n20016), .A(n16178), .ZN(n16179) );
  OAI21_X1 U19334 ( .B1(n16202), .B2(n16180), .A(n16179), .ZN(P2_U2901) );
  NOR2_X1 U19335 ( .A1(n16197), .A2(n16181), .ZN(n16186) );
  NAND2_X1 U19336 ( .A1(n16194), .A2(BUF2_REG_17__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U19337 ( .A1(n16191), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n16182) );
  OAI211_X1 U19338 ( .C1(n20025), .C2(n16184), .A(n16183), .B(n16182), .ZN(
        n16185) );
  AOI211_X1 U19339 ( .C1(n16187), .C2(n20016), .A(n16186), .B(n16185), .ZN(
        n16188) );
  OAI21_X1 U19340 ( .B1(n16202), .B2(n16189), .A(n16188), .ZN(P2_U2902) );
  INV_X1 U19341 ( .A(n16190), .ZN(n16201) );
  AOI22_X1 U19342 ( .A1(n16193), .A2(n16192), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n16191), .ZN(n16196) );
  NAND2_X1 U19343 ( .A1(n16194), .A2(BUF2_REG_16__SCAN_IN), .ZN(n16195) );
  OAI211_X1 U19344 ( .C1(n17638), .C2(n16197), .A(n16196), .B(n16195), .ZN(
        n16198) );
  AOI21_X1 U19345 ( .B1(n16199), .B2(n20016), .A(n16198), .ZN(n16200) );
  OAI21_X1 U19346 ( .B1(n16202), .B2(n16201), .A(n16200), .ZN(P2_U2903) );
  INV_X1 U19347 ( .A(n16753), .ZN(n16214) );
  INV_X1 U19348 ( .A(n16203), .ZN(n20756) );
  INV_X1 U19349 ( .A(n20751), .ZN(n16831) );
  XOR2_X1 U19350 ( .A(n16203), .B(n20751), .Z(n20012) );
  OAI21_X1 U19351 ( .B1(n20762), .B2(n20760), .A(n16204), .ZN(n20011) );
  NAND2_X1 U19352 ( .A1(n20012), .A2(n20011), .ZN(n20010) );
  OAI21_X1 U19353 ( .B1(n20756), .B2(n16831), .A(n20010), .ZN(n16208) );
  NAND2_X1 U19354 ( .A1(n16206), .A2(n16205), .ZN(n16207) );
  NAND2_X1 U19355 ( .A1(n15932), .A2(n16207), .ZN(n20003) );
  NAND2_X1 U19356 ( .A1(n16208), .A2(n20003), .ZN(n20006) );
  INV_X1 U19357 ( .A(n20005), .ZN(n16209) );
  NAND3_X1 U19358 ( .A1(n20006), .A2(n20020), .A3(n16209), .ZN(n16212) );
  AOI22_X1 U19359 ( .A1(n16210), .A2(n20129), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n16191), .ZN(n16211) );
  OAI211_X1 U19360 ( .C1(n16214), .C2(n16213), .A(n16212), .B(n16211), .ZN(
        P2_U2914) );
  NOR2_X1 U19361 ( .A1(n16464), .A2(n16218), .ZN(n16476) );
  AOI21_X1 U19362 ( .B1(n16445), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16476), .ZN(n16219) );
  OAI211_X1 U19363 ( .C1(n16448), .C2(n16221), .A(n16220), .B(n16219), .ZN(
        n16222) );
  AOI21_X1 U19364 ( .B1(n16470), .B2(n16482), .A(n16222), .ZN(n16223) );
  OAI21_X1 U19365 ( .B1(n16484), .B2(n16472), .A(n16223), .ZN(P2_U2984) );
  NAND2_X1 U19366 ( .A1(n16225), .A2(n16224), .ZN(n16227) );
  XOR2_X1 U19367 ( .A(n16227), .B(n16226), .Z(n16496) );
  NAND2_X1 U19368 ( .A1(n16495), .A2(n16470), .ZN(n16235) );
  NAND2_X1 U19369 ( .A1(n16230), .A2(n17586), .ZN(n16231) );
  NAND2_X1 U19370 ( .A1(n16754), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n16489) );
  OAI211_X1 U19371 ( .C1(n16232), .C2(n17599), .A(n16231), .B(n16489), .ZN(
        n16233) );
  AOI21_X1 U19372 ( .B1(n16493), .B2(n16454), .A(n16233), .ZN(n16234) );
  OAI211_X1 U19373 ( .C1(n16496), .C2(n16472), .A(n16235), .B(n16234), .ZN(
        P2_U2985) );
  NAND2_X1 U19374 ( .A1(n16236), .A2(n16252), .ZN(n16237) );
  XOR2_X1 U19375 ( .A(n16238), .B(n16237), .Z(n16508) );
  INV_X1 U19376 ( .A(n16241), .ZN(n16244) );
  NAND2_X1 U19377 ( .A1(n16754), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n16499) );
  OAI21_X1 U19378 ( .B1(n17599), .B2(n16242), .A(n16499), .ZN(n16243) );
  AOI21_X1 U19379 ( .B1(n16244), .B2(n17586), .A(n16243), .ZN(n16245) );
  OAI21_X1 U19380 ( .B1(n16246), .B2(n17589), .A(n16245), .ZN(n16247) );
  AOI21_X1 U19381 ( .B1(n16506), .B2(n16470), .A(n16247), .ZN(n16248) );
  OAI21_X1 U19382 ( .B1(n16508), .B2(n16472), .A(n16248), .ZN(P2_U2988) );
  NAND2_X1 U19383 ( .A1(n16249), .A2(n17586), .ZN(n16250) );
  NAND2_X1 U19384 ( .A1(n16754), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n16513) );
  OAI211_X1 U19385 ( .C1(n16251), .C2(n17599), .A(n16250), .B(n16513), .ZN(
        n16257) );
  INV_X1 U19386 ( .A(n16252), .ZN(n16256) );
  OAI21_X1 U19387 ( .B1(n16254), .B2(n16256), .A(n16253), .ZN(n16255) );
  INV_X1 U19388 ( .A(n16239), .ZN(n16258) );
  NAND2_X1 U19389 ( .A1(n16258), .A2(n16514), .ZN(n16510) );
  NAND3_X1 U19390 ( .A1(n16510), .A2(n16470), .A3(n16509), .ZN(n16259) );
  NAND2_X1 U19391 ( .A1(n16534), .A2(n16470), .ZN(n16269) );
  NAND2_X1 U19392 ( .A1(n16754), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n16523) );
  OAI21_X1 U19393 ( .B1(n17599), .B2(n16263), .A(n16523), .ZN(n16264) );
  INV_X1 U19394 ( .A(n16264), .ZN(n16265) );
  OAI21_X1 U19395 ( .B1(n16266), .B2(n16448), .A(n16265), .ZN(n16267) );
  AOI21_X1 U19396 ( .B1(n16528), .B2(n16454), .A(n16267), .ZN(n16268) );
  OAI211_X1 U19397 ( .C1(n16532), .C2(n16472), .A(n16269), .B(n16268), .ZN(
        P2_U2990) );
  OAI21_X1 U19398 ( .B1(n16270), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16262), .ZN(n16551) );
  NAND2_X1 U19399 ( .A1(n16754), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16541) );
  OAI21_X1 U19400 ( .B1(n17599), .B2(n21644), .A(n16541), .ZN(n16271) );
  AOI21_X1 U19401 ( .B1(n16272), .B2(n17586), .A(n16271), .ZN(n16276) );
  NOR2_X1 U19402 ( .A1(n16274), .A2(n16273), .ZN(n16537) );
  OR3_X1 U19403 ( .A1(n16537), .A2(n16536), .A3(n16472), .ZN(n16275) );
  OAI211_X1 U19404 ( .C1(n16546), .C2(n17589), .A(n16276), .B(n16275), .ZN(
        n16277) );
  INV_X1 U19405 ( .A(n16277), .ZN(n16278) );
  OAI21_X1 U19406 ( .B1(n16551), .B2(n17594), .A(n16278), .ZN(P2_U2991) );
  AND2_X1 U19407 ( .A1(n16281), .A2(n16280), .ZN(n16282) );
  XNOR2_X1 U19408 ( .A(n16279), .B(n16282), .ZN(n16564) );
  INV_X1 U19409 ( .A(n16270), .ZN(n16553) );
  NAND2_X1 U19410 ( .A1(n12432), .A2(n16556), .ZN(n16552) );
  NAND3_X1 U19411 ( .A1(n16553), .A2(n16470), .A3(n16552), .ZN(n16289) );
  NAND2_X1 U19412 ( .A1(n16754), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n16554) );
  OAI21_X1 U19413 ( .B1(n17599), .B2(n16283), .A(n16554), .ZN(n16284) );
  INV_X1 U19414 ( .A(n16284), .ZN(n16285) );
  OAI21_X1 U19415 ( .B1(n16286), .B2(n16448), .A(n16285), .ZN(n16287) );
  AOI21_X1 U19416 ( .B1(n16561), .B2(n16454), .A(n16287), .ZN(n16288) );
  OAI211_X1 U19417 ( .C1(n16564), .C2(n16472), .A(n16289), .B(n16288), .ZN(
        P2_U2992) );
  NAND2_X1 U19418 ( .A1(n16291), .A2(n16290), .ZN(n16295) );
  NAND2_X1 U19419 ( .A1(n16293), .A2(n16292), .ZN(n16294) );
  XNOR2_X1 U19420 ( .A(n16295), .B(n16294), .ZN(n16579) );
  NAND2_X1 U19421 ( .A1(n16754), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U19422 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16296) );
  OAI211_X1 U19423 ( .C1(n16297), .C2(n16448), .A(n16570), .B(n16296), .ZN(
        n16299) );
  OAI21_X1 U19424 ( .B1(n16579), .B2(n16472), .A(n16300), .ZN(P2_U2994) );
  NAND2_X1 U19425 ( .A1(n16302), .A2(n16301), .ZN(n16303) );
  NAND2_X1 U19426 ( .A1(n16754), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n16581) );
  OAI21_X1 U19427 ( .B1(n17599), .B2(n16306), .A(n16581), .ZN(n16307) );
  AOI21_X1 U19428 ( .B1(n16308), .B2(n17586), .A(n16307), .ZN(n16309) );
  OAI21_X1 U19429 ( .B1(n16587), .B2(n17589), .A(n16309), .ZN(n16310) );
  AOI21_X1 U19430 ( .B1(n16589), .B2(n16470), .A(n16310), .ZN(n16311) );
  OAI21_X1 U19431 ( .B1(n16591), .B2(n16472), .A(n16311), .ZN(P2_U2995) );
  AOI21_X1 U19432 ( .B1(n16322), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16315) );
  INV_X1 U19433 ( .A(n16304), .ZN(n16314) );
  NOR2_X2 U19434 ( .A1(n16315), .A2(n16314), .ZN(n16604) );
  NAND2_X1 U19435 ( .A1(n16754), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n16595) );
  OAI21_X1 U19436 ( .B1(n17599), .B2(n16316), .A(n16595), .ZN(n16317) );
  AOI21_X1 U19437 ( .B1(n16318), .B2(n17586), .A(n16317), .ZN(n16319) );
  OAI21_X1 U19438 ( .B1(n16602), .B2(n17589), .A(n16319), .ZN(n16320) );
  AOI21_X1 U19439 ( .B1(n16604), .B2(n16470), .A(n16320), .ZN(n16321) );
  OAI21_X1 U19440 ( .B1(n16606), .B2(n16472), .A(n16321), .ZN(P2_U2996) );
  XNOR2_X1 U19441 ( .A(n16322), .B(n16323), .ZN(n16330) );
  NAND2_X1 U19442 ( .A1(n16324), .A2(n16454), .ZN(n16327) );
  AOI21_X1 U19443 ( .B1(n16445), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n16325), .ZN(n16326) );
  OAI211_X1 U19444 ( .C1(n16448), .C2(n16328), .A(n16327), .B(n16326), .ZN(
        n16329) );
  AOI21_X1 U19445 ( .B1(n16330), .B2(n16470), .A(n16329), .ZN(n16331) );
  OAI21_X1 U19446 ( .B1(n16332), .B2(n16472), .A(n16331), .ZN(P2_U2997) );
  OAI211_X1 U19447 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16345), .A(
        n9944), .B(n16470), .ZN(n16339) );
  NAND2_X1 U19448 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16333) );
  OAI211_X1 U19449 ( .C1(n16335), .C2(n16448), .A(n16334), .B(n16333), .ZN(
        n16336) );
  AOI21_X1 U19450 ( .B1(n16337), .B2(n16454), .A(n16336), .ZN(n16338) );
  OAI211_X1 U19451 ( .C1(n10443), .C2(n16472), .A(n16339), .B(n16338), .ZN(
        P2_U2998) );
  NAND2_X1 U19452 ( .A1(n16341), .A2(n16340), .ZN(n16344) );
  NAND2_X1 U19453 ( .A1(n16342), .A2(n16351), .ZN(n16343) );
  XOR2_X1 U19454 ( .A(n16344), .B(n16343), .Z(n16617) );
  NAND2_X1 U19455 ( .A1(n16754), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16610) );
  OAI21_X1 U19456 ( .B1(n17599), .B2(n16346), .A(n16610), .ZN(n16347) );
  AOI21_X1 U19457 ( .B1(n17586), .B2(n16348), .A(n16347), .ZN(n16349) );
  OAI21_X1 U19458 ( .B1(n16611), .B2(n17589), .A(n16349), .ZN(n16350) );
  NAND2_X1 U19459 ( .A1(n16352), .A2(n16351), .ZN(n16354) );
  XOR2_X1 U19460 ( .A(n16354), .B(n16353), .Z(n16630) );
  AOI21_X1 U19461 ( .B1(n16356), .B2(n16364), .A(n16355), .ZN(n16618) );
  NAND2_X1 U19462 ( .A1(n16618), .A2(n16470), .ZN(n16362) );
  NAND2_X1 U19463 ( .A1(n17586), .A2(n16357), .ZN(n16358) );
  NAND2_X1 U19464 ( .A1(n16754), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n16622) );
  OAI211_X1 U19465 ( .C1(n16359), .C2(n17599), .A(n16358), .B(n16622), .ZN(
        n16360) );
  AOI21_X1 U19466 ( .B1(n16621), .B2(n16454), .A(n16360), .ZN(n16361) );
  OAI211_X1 U19467 ( .C1(n16630), .C2(n16472), .A(n16362), .B(n16361), .ZN(
        P2_U3000) );
  OAI21_X1 U19468 ( .B1(n16378), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16364), .ZN(n16643) );
  NAND2_X1 U19469 ( .A1(n16366), .A2(n16365), .ZN(n16368) );
  XOR2_X1 U19470 ( .A(n16368), .B(n16367), .Z(n16641) );
  NOR2_X1 U19471 ( .A1(n16632), .A2(n17589), .ZN(n16372) );
  NAND2_X1 U19472 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16369) );
  NAND2_X1 U19473 ( .A1(n16754), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16631) );
  OAI211_X1 U19474 ( .C1(n16448), .C2(n16370), .A(n16369), .B(n16631), .ZN(
        n16371) );
  AOI211_X1 U19475 ( .C1(n16641), .C2(n17587), .A(n16372), .B(n16371), .ZN(
        n16373) );
  OAI21_X1 U19476 ( .B1(n16643), .B2(n17594), .A(n16373), .ZN(P2_U3001) );
  XNOR2_X1 U19477 ( .A(n16374), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16375) );
  XNOR2_X1 U19478 ( .A(n16376), .B(n16375), .ZN(n16654) );
  NAND2_X1 U19479 ( .A1(n16644), .A2(n16470), .ZN(n16384) );
  NAND2_X1 U19480 ( .A1(n16754), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n16647) );
  OAI21_X1 U19481 ( .B1(n17599), .B2(n16379), .A(n16647), .ZN(n16381) );
  NOR2_X1 U19482 ( .A1(n16648), .A2(n17589), .ZN(n16380) );
  AOI211_X1 U19483 ( .C1(n16382), .C2(n17586), .A(n16381), .B(n16380), .ZN(
        n16383) );
  OAI211_X1 U19484 ( .C1(n16654), .C2(n16472), .A(n16384), .B(n16383), .ZN(
        P2_U3002) );
  NAND2_X1 U19485 ( .A1(n16386), .A2(n16385), .ZN(n16394) );
  XNOR2_X1 U19486 ( .A(n16388), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16443) );
  OAI21_X1 U19487 ( .B1(n16444), .B2(n16443), .A(n16389), .ZN(n16423) );
  INV_X1 U19488 ( .A(n16400), .ZN(n16393) );
  NAND2_X1 U19489 ( .A1(n17586), .A2(n16395), .ZN(n16396) );
  NAND2_X1 U19490 ( .A1(n16754), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n16659) );
  OAI211_X1 U19491 ( .C1(n16397), .C2(n17599), .A(n16396), .B(n16659), .ZN(
        n16398) );
  NAND2_X1 U19492 ( .A1(n16400), .A2(n16399), .ZN(n16402) );
  XOR2_X1 U19493 ( .A(n16402), .B(n16401), .Z(n16684) );
  NAND2_X1 U19494 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16403) );
  NAND2_X1 U19495 ( .A1(n16754), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n16673) );
  OAI211_X1 U19496 ( .C1(n16448), .C2(n16404), .A(n16403), .B(n16673), .ZN(
        n16406) );
  OAI21_X1 U19497 ( .B1(n16684), .B2(n16472), .A(n16407), .ZN(P2_U3004) );
  NAND2_X1 U19498 ( .A1(n16409), .A2(n16408), .ZN(n16411) );
  XOR2_X1 U19499 ( .A(n16411), .B(n16410), .Z(n16698) );
  NAND2_X1 U19500 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16412) );
  NAND2_X1 U19501 ( .A1(n16754), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n16686) );
  OAI211_X1 U19502 ( .C1(n16448), .C2(n16413), .A(n16412), .B(n16686), .ZN(
        n16414) );
  OAI21_X1 U19503 ( .B1(n16472), .B2(n16698), .A(n16415), .ZN(P2_U3005) );
  XNOR2_X1 U19504 ( .A(n16418), .B(n16701), .ZN(n16419) );
  NAND2_X1 U19505 ( .A1(n16421), .A2(n16420), .ZN(n16425) );
  INV_X1 U19506 ( .A(n16432), .ZN(n16422) );
  AOI21_X1 U19507 ( .B1(n16423), .B2(n16431), .A(n16422), .ZN(n16424) );
  XOR2_X1 U19508 ( .A(n16425), .B(n16424), .Z(n16710) );
  NOR2_X1 U19509 ( .A1(n16707), .A2(n17589), .ZN(n16429) );
  NAND2_X1 U19510 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16426) );
  NAND2_X1 U19511 ( .A1(n16754), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16702) );
  OAI211_X1 U19512 ( .C1(n16448), .C2(n16427), .A(n16426), .B(n16702), .ZN(
        n16428) );
  AOI211_X1 U19513 ( .C1(n16710), .C2(n17587), .A(n16429), .B(n16428), .ZN(
        n16430) );
  OAI21_X1 U19514 ( .B1(n16712), .B2(n17594), .A(n16430), .ZN(P2_U3006) );
  NAND2_X1 U19515 ( .A1(n16432), .A2(n16431), .ZN(n16433) );
  XNOR2_X1 U19516 ( .A(n16434), .B(n16433), .ZN(n16726) );
  INV_X1 U19517 ( .A(n16435), .ZN(n16714) );
  NAND2_X1 U19518 ( .A1(n16436), .A2(n16722), .ZN(n16713) );
  NAND3_X1 U19519 ( .A1(n16714), .A2(n16470), .A3(n16713), .ZN(n16442) );
  NAND2_X1 U19520 ( .A1(n16754), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n16718) );
  OAI21_X1 U19521 ( .B1(n17599), .B2(n16437), .A(n16718), .ZN(n16439) );
  NOR2_X1 U19522 ( .A1(n16719), .A2(n17589), .ZN(n16438) );
  AOI211_X1 U19523 ( .C1(n16440), .C2(n17586), .A(n16439), .B(n16438), .ZN(
        n16441) );
  OAI211_X1 U19524 ( .C1(n16726), .C2(n16472), .A(n16442), .B(n16441), .ZN(
        P2_U3007) );
  XNOR2_X1 U19525 ( .A(n16444), .B(n16443), .ZN(n16736) );
  NAND2_X1 U19526 ( .A1(n16445), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16446) );
  NAND2_X1 U19527 ( .A1(n16754), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16730) );
  OAI211_X1 U19528 ( .C1(n16448), .C2(n16447), .A(n16446), .B(n16730), .ZN(
        n16453) );
  OAI21_X1 U19529 ( .B1(n16450), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16451), .ZN(n16739) );
  NOR2_X1 U19530 ( .A1(n16739), .A2(n17594), .ZN(n16452) );
  AOI211_X1 U19531 ( .C1(n16454), .C2(n16727), .A(n16453), .B(n16452), .ZN(
        n16455) );
  OAI21_X1 U19532 ( .B1(n16472), .B2(n16736), .A(n16455), .ZN(P2_U3008) );
  OAI21_X1 U19533 ( .B1(n16458), .B2(n12032), .A(n16457), .ZN(n16460) );
  XNOR2_X1 U19534 ( .A(n19982), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16459) );
  XNOR2_X1 U19535 ( .A(n16460), .B(n16459), .ZN(n16773) );
  NAND2_X1 U19536 ( .A1(n16462), .A2(n16461), .ZN(n16463) );
  XNOR2_X1 U19537 ( .A(n16463), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n16771) );
  OAI22_X1 U19538 ( .A1(n17599), .A2(n16466), .B1(n16465), .B2(n16464), .ZN(
        n16467) );
  AOI21_X1 U19539 ( .B1(n17586), .B2(n19991), .A(n16467), .ZN(n16468) );
  OAI21_X1 U19540 ( .B1(n19986), .B2(n17589), .A(n16468), .ZN(n16469) );
  AOI21_X1 U19541 ( .B1(n16771), .B2(n16470), .A(n16469), .ZN(n16471) );
  OAI21_X1 U19542 ( .B1(n16773), .B2(n16472), .A(n16471), .ZN(P2_U3010) );
  NAND2_X1 U19543 ( .A1(n16473), .A2(n17604), .ZN(n16479) );
  INV_X1 U19544 ( .A(n16486), .ZN(n16474) );
  NOR3_X1 U19545 ( .A1(n16474), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16485), .ZN(n16475) );
  AOI211_X1 U19546 ( .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n16477), .A(
        n16476), .B(n16475), .ZN(n16478) );
  OAI211_X1 U19547 ( .C1(n16763), .C2(n16480), .A(n16479), .B(n16478), .ZN(
        n16481) );
  AOI21_X1 U19548 ( .B1(n17606), .B2(n16482), .A(n16481), .ZN(n16483) );
  OAI211_X1 U19549 ( .C1(n16487), .C2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16486), .B(n16485), .ZN(n16488) );
  OAI211_X1 U19550 ( .C1(n16491), .C2(n16490), .A(n16489), .B(n16488), .ZN(
        n16492) );
  OAI21_X1 U19551 ( .B1(n16525), .B2(n16514), .A(n16500), .ZN(n16497) );
  NAND3_X1 U19552 ( .A1(n16511), .A2(n10710), .A3(n16497), .ZN(n16498) );
  OAI211_X1 U19553 ( .C1(n16515), .C2(n16500), .A(n16499), .B(n16498), .ZN(
        n16501) );
  AOI21_X1 U19554 ( .B1(n16502), .B2(n17604), .A(n16501), .ZN(n16503) );
  OAI21_X1 U19555 ( .B1(n16763), .B2(n16504), .A(n16503), .ZN(n16505) );
  AOI21_X1 U19556 ( .B1(n16506), .B2(n17606), .A(n16505), .ZN(n16507) );
  OAI21_X1 U19557 ( .B1(n16508), .B2(n10442), .A(n16507), .ZN(P2_U3020) );
  NAND3_X1 U19558 ( .A1(n16510), .A2(n17606), .A3(n16509), .ZN(n16521) );
  NAND3_X1 U19559 ( .A1(n16511), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n16514), .ZN(n16512) );
  OAI211_X1 U19560 ( .C1(n16515), .C2(n16514), .A(n16513), .B(n16512), .ZN(
        n16518) );
  NOR2_X1 U19561 ( .A1(n16516), .A2(n16763), .ZN(n16517) );
  AOI211_X1 U19562 ( .C1(n16519), .C2(n17604), .A(n16518), .B(n16517), .ZN(
        n16520) );
  OAI211_X1 U19563 ( .C1(n16522), .C2(n10442), .A(n16521), .B(n16520), .ZN(
        P2_U3021) );
  OAI211_X1 U19564 ( .C1(n16526), .C2(n16525), .A(n16524), .B(n16523), .ZN(
        n16527) );
  AOI21_X1 U19565 ( .B1(n16528), .B2(n17604), .A(n16527), .ZN(n16531) );
  NAND2_X1 U19566 ( .A1(n16529), .A2(n17608), .ZN(n16530) );
  OAI211_X1 U19567 ( .C1(n16532), .C2(n10442), .A(n16531), .B(n16530), .ZN(
        n16533) );
  AOI21_X1 U19568 ( .B1(n16534), .B2(n17606), .A(n16533), .ZN(n16535) );
  INV_X1 U19569 ( .A(n16535), .ZN(P2_U3022) );
  NOR3_X1 U19570 ( .A1(n16537), .A2(n16536), .A3(n10442), .ZN(n16548) );
  NAND2_X1 U19571 ( .A1(n16540), .A2(n16556), .ZN(n16555) );
  INV_X1 U19572 ( .A(n16538), .ZN(n16557) );
  AOI21_X1 U19573 ( .B1(n16555), .B2(n16557), .A(n16539), .ZN(n16544) );
  NAND3_X1 U19574 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16540), .A3(
        n16539), .ZN(n16542) );
  NAND2_X1 U19575 ( .A1(n16542), .A2(n16541), .ZN(n16543) );
  NOR2_X1 U19576 ( .A1(n16544), .A2(n16543), .ZN(n16545) );
  OAI21_X1 U19577 ( .B1(n16546), .B2(n16764), .A(n16545), .ZN(n16547) );
  AOI211_X1 U19578 ( .C1(n17608), .C2(n16549), .A(n16548), .B(n16547), .ZN(
        n16550) );
  OAI21_X1 U19579 ( .B1(n16551), .B2(n16748), .A(n16550), .ZN(P2_U3023) );
  NAND3_X1 U19580 ( .A1(n16553), .A2(n17606), .A3(n16552), .ZN(n16563) );
  OAI211_X1 U19581 ( .C1(n16557), .C2(n16556), .A(n16555), .B(n16554), .ZN(
        n16560) );
  NOR2_X1 U19582 ( .A1(n16558), .A2(n16763), .ZN(n16559) );
  AOI211_X1 U19583 ( .C1(n16561), .C2(n17604), .A(n16560), .B(n16559), .ZN(
        n16562) );
  OAI211_X1 U19584 ( .C1(n16564), .C2(n10442), .A(n16563), .B(n16562), .ZN(
        P2_U3024) );
  OAI211_X1 U19585 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n16567), .B(n16565), .ZN(
        n16574) );
  NAND2_X1 U19586 ( .A1(n16566), .A2(n17604), .ZN(n16573) );
  NAND2_X1 U19587 ( .A1(n16568), .A2(n10706), .ZN(n16569) );
  NAND2_X1 U19588 ( .A1(n16687), .A2(n16569), .ZN(n16584) );
  INV_X1 U19589 ( .A(n16570), .ZN(n16571) );
  AOI21_X1 U19590 ( .B1(n16584), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16571), .ZN(n16572) );
  OAI211_X1 U19591 ( .C1(n16685), .C2(n16574), .A(n16573), .B(n16572), .ZN(
        n16576) );
  OAI21_X1 U19592 ( .B1(n16579), .B2(n10442), .A(n16578), .ZN(P2_U3026) );
  NAND2_X1 U19593 ( .A1(n16580), .A2(n17608), .ZN(n16586) );
  INV_X1 U19594 ( .A(n16581), .ZN(n16583) );
  NOR3_X1 U19595 ( .A1(n16685), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n10706), .ZN(n16582) );
  AOI211_X1 U19596 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n16584), .A(
        n16583), .B(n16582), .ZN(n16585) );
  OAI211_X1 U19597 ( .C1(n16587), .C2(n16764), .A(n16586), .B(n16585), .ZN(
        n16588) );
  OAI21_X1 U19598 ( .B1(n16591), .B2(n10442), .A(n16590), .ZN(P2_U3027) );
  NOR2_X1 U19599 ( .A1(n16592), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16598) );
  INV_X1 U19600 ( .A(n16592), .ZN(n16593) );
  NOR2_X1 U19601 ( .A1(n17615), .A2(n16593), .ZN(n16594) );
  OAI21_X1 U19602 ( .B1(n16608), .B2(n16594), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16596) );
  NAND2_X1 U19603 ( .A1(n16596), .A2(n16595), .ZN(n16597) );
  AOI21_X1 U19604 ( .B1(n16615), .B2(n16598), .A(n16597), .ZN(n16601) );
  NAND2_X1 U19605 ( .A1(n16599), .A2(n17608), .ZN(n16600) );
  OAI211_X1 U19606 ( .C1(n16602), .C2(n16764), .A(n16601), .B(n16600), .ZN(
        n16603) );
  AOI21_X1 U19607 ( .B1(n16604), .B2(n17606), .A(n16603), .ZN(n16605) );
  OAI21_X1 U19608 ( .B1(n16606), .B2(n10442), .A(n16605), .ZN(P2_U3028) );
  NOR2_X1 U19609 ( .A1(n16607), .A2(n16763), .ZN(n16613) );
  NAND2_X1 U19610 ( .A1(n16608), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16609) );
  OAI211_X1 U19611 ( .C1(n16611), .C2(n16764), .A(n16610), .B(n16609), .ZN(
        n16612) );
  AOI211_X1 U19612 ( .C1(n16615), .C2(n16614), .A(n16613), .B(n16612), .ZN(
        n16616) );
  NAND2_X1 U19613 ( .A1(n16618), .A2(n17606), .ZN(n16629) );
  NOR2_X1 U19614 ( .A1(n16633), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16649) );
  INV_X1 U19615 ( .A(n16656), .ZN(n16619) );
  OAI21_X1 U19616 ( .B1(n16619), .B2(n17615), .A(n16687), .ZN(n16645) );
  NOR2_X1 U19617 ( .A1(n16649), .A2(n16645), .ZN(n16639) );
  OAI21_X1 U19618 ( .B1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16633), .A(
        n16639), .ZN(n16627) );
  NOR2_X1 U19619 ( .A1(n16620), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16626) );
  NAND2_X1 U19620 ( .A1(n16621), .A2(n17604), .ZN(n16623) );
  OAI211_X1 U19621 ( .C1(n16763), .C2(n16624), .A(n16623), .B(n16622), .ZN(
        n16625) );
  AOI211_X1 U19622 ( .C1(n16627), .C2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16626), .B(n16625), .ZN(n16628) );
  OAI211_X1 U19623 ( .C1(n16630), .C2(n10442), .A(n16629), .B(n16628), .ZN(
        P2_U3032) );
  OAI21_X1 U19624 ( .B1(n16632), .B2(n16764), .A(n16631), .ZN(n16635) );
  NOR3_X1 U19625 ( .A1(n16633), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n12416), .ZN(n16634) );
  AOI211_X1 U19626 ( .C1(n17608), .C2(n16636), .A(n16635), .B(n16634), .ZN(
        n16637) );
  OAI21_X1 U19627 ( .B1(n16639), .B2(n16638), .A(n16637), .ZN(n16640) );
  AOI21_X1 U19628 ( .B1(n16641), .B2(n17602), .A(n16640), .ZN(n16642) );
  OAI21_X1 U19629 ( .B1(n16643), .B2(n16748), .A(n16642), .ZN(P2_U3033) );
  NAND2_X1 U19630 ( .A1(n16645), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16646) );
  OAI211_X1 U19631 ( .C1(n16648), .C2(n16764), .A(n16647), .B(n16646), .ZN(
        n16650) );
  AOI211_X1 U19632 ( .C1(n17608), .C2(n16651), .A(n16650), .B(n16649), .ZN(
        n16652) );
  OAI211_X1 U19633 ( .C1(n16654), .C2(n10442), .A(n16653), .B(n16652), .ZN(
        P2_U3034) );
  INV_X1 U19634 ( .A(n16655), .ZN(n16668) );
  NAND2_X1 U19635 ( .A1(n16656), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16658) );
  NAND3_X1 U19636 ( .A1(n10396), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16657) );
  AND2_X1 U19637 ( .A1(n16658), .A2(n16657), .ZN(n16666) );
  OAI21_X1 U19638 ( .B1(n16687), .B2(n16660), .A(n16659), .ZN(n16663) );
  NOR2_X1 U19639 ( .A1(n16661), .A2(n16763), .ZN(n16662) );
  AOI211_X1 U19640 ( .C1(n16664), .C2(n17604), .A(n16663), .B(n16662), .ZN(
        n16665) );
  OAI21_X1 U19641 ( .B1(n16685), .B2(n16666), .A(n16665), .ZN(n16667) );
  AOI21_X1 U19642 ( .B1(n16668), .B2(n17606), .A(n16667), .ZN(n16669) );
  OAI21_X1 U19643 ( .B1(n16670), .B2(n10442), .A(n16669), .ZN(P2_U3035) );
  NOR3_X1 U19644 ( .A1(n16672), .A2(n16671), .A3(n16748), .ZN(n16682) );
  XNOR2_X1 U19645 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16680) );
  OAI21_X1 U19646 ( .B1(n16687), .B2(n16674), .A(n16673), .ZN(n16675) );
  AOI21_X1 U19647 ( .B1(n16676), .B2(n17604), .A(n16675), .ZN(n16679) );
  NAND2_X1 U19648 ( .A1(n16677), .A2(n17608), .ZN(n16678) );
  OAI211_X1 U19649 ( .C1(n16685), .C2(n16680), .A(n16679), .B(n16678), .ZN(
        n16681) );
  NOR2_X1 U19650 ( .A1(n16682), .A2(n16681), .ZN(n16683) );
  OAI21_X1 U19651 ( .B1(n16684), .B2(n10442), .A(n16683), .ZN(P2_U3036) );
  INV_X1 U19652 ( .A(n16685), .ZN(n16696) );
  OAI21_X1 U19653 ( .B1(n16687), .B2(n10209), .A(n16686), .ZN(n16688) );
  AOI21_X1 U19654 ( .B1(n16689), .B2(n17604), .A(n16688), .ZN(n16690) );
  OAI21_X1 U19655 ( .B1(n16763), .B2(n16691), .A(n16690), .ZN(n16695) );
  AOI211_X1 U19656 ( .C1(n16696), .C2(n10209), .A(n16695), .B(n16694), .ZN(
        n16697) );
  OAI21_X1 U19657 ( .B1(n10442), .B2(n16698), .A(n16697), .ZN(P2_U3037) );
  INV_X1 U19658 ( .A(n16723), .ZN(n16699) );
  AOI211_X1 U19659 ( .C1(n16722), .C2(n16701), .A(n16700), .B(n16699), .ZN(
        n16709) );
  INV_X1 U19660 ( .A(n16702), .ZN(n16703) );
  AOI21_X1 U19661 ( .B1(n16716), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n16703), .ZN(n16706) );
  NAND2_X1 U19662 ( .A1(n16704), .A2(n17608), .ZN(n16705) );
  OAI211_X1 U19663 ( .C1(n16707), .C2(n16764), .A(n16706), .B(n16705), .ZN(
        n16708) );
  AOI211_X1 U19664 ( .C1(n16710), .C2(n17602), .A(n16709), .B(n16708), .ZN(
        n16711) );
  OAI21_X1 U19665 ( .B1(n16712), .B2(n16748), .A(n16711), .ZN(P2_U3038) );
  NAND3_X1 U19666 ( .A1(n16714), .A2(n17606), .A3(n16713), .ZN(n16725) );
  NOR2_X1 U19667 ( .A1(n16715), .A2(n16763), .ZN(n16721) );
  NAND2_X1 U19668 ( .A1(n16716), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16717) );
  OAI211_X1 U19669 ( .C1(n16719), .C2(n16764), .A(n16718), .B(n16717), .ZN(
        n16720) );
  AOI211_X1 U19670 ( .C1(n16723), .C2(n16722), .A(n16721), .B(n16720), .ZN(
        n16724) );
  OAI211_X1 U19671 ( .C1(n16726), .C2(n10442), .A(n16725), .B(n16724), .ZN(
        P2_U3039) );
  INV_X1 U19672 ( .A(n16727), .ZN(n16731) );
  NAND2_X1 U19673 ( .A1(n16728), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16729) );
  OAI211_X1 U19674 ( .C1(n16731), .C2(n16764), .A(n16730), .B(n16729), .ZN(
        n16734) );
  NOR3_X1 U19675 ( .A1(n16768), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        n16732), .ZN(n16733) );
  AOI211_X1 U19676 ( .C1(n17608), .C2(n16735), .A(n16734), .B(n16733), .ZN(
        n16738) );
  OR2_X1 U19677 ( .A1(n16736), .A2(n10442), .ZN(n16737) );
  OAI211_X1 U19678 ( .C1(n16739), .C2(n16748), .A(n16738), .B(n16737), .ZN(
        P2_U3040) );
  INV_X1 U19679 ( .A(n16741), .ZN(n16742) );
  XNOR2_X1 U19680 ( .A(n16740), .B(n16742), .ZN(n17588) );
  INV_X1 U19681 ( .A(n17588), .ZN(n16762) );
  NAND2_X1 U19682 ( .A1(n16747), .A2(n16746), .ZN(n17593) );
  NOR2_X1 U19683 ( .A1(n17593), .A2(n16748), .ZN(n16760) );
  INV_X1 U19684 ( .A(n16749), .ZN(n16750) );
  AOI211_X1 U19685 ( .C1(n16752), .C2(n16767), .A(n16751), .B(n16750), .ZN(
        n16759) );
  AND2_X1 U19686 ( .A1(n16753), .A2(n17608), .ZN(n16758) );
  NAND2_X1 U19687 ( .A1(n16754), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n17583) );
  INV_X1 U19688 ( .A(n16766), .ZN(n16755) );
  NAND2_X1 U19689 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n16755), .ZN(
        n16756) );
  OAI211_X1 U19690 ( .C1(n17590), .C2(n16764), .A(n17583), .B(n16756), .ZN(
        n16757) );
  NOR4_X1 U19691 ( .A1(n16760), .A2(n16759), .A3(n16758), .A4(n16757), .ZN(
        n16761) );
  OAI21_X1 U19692 ( .B1(n10442), .B2(n16762), .A(n16761), .ZN(P2_U3041) );
  OAI22_X1 U19693 ( .A1(n19986), .A2(n16764), .B1(n16763), .B2(n20003), .ZN(
        n16770) );
  NAND2_X1 U19694 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n16754), .ZN(n16765) );
  OAI221_X1 U19695 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n16768), .C1(
        n16767), .C2(n16766), .A(n16765), .ZN(n16769) );
  AOI211_X1 U19696 ( .C1(n16771), .C2(n17606), .A(n16770), .B(n16769), .ZN(
        n16772) );
  OAI21_X1 U19697 ( .B1(n10442), .B2(n16773), .A(n16772), .ZN(P2_U3042) );
  INV_X1 U19698 ( .A(n16816), .ZN(n16786) );
  NAND2_X1 U19699 ( .A1(n12527), .A2(n16786), .ZN(n16777) );
  NAND2_X1 U19700 ( .A1(n16775), .A2(n16774), .ZN(n16794) );
  NAND2_X1 U19701 ( .A1(n16794), .A2(n16905), .ZN(n16776) );
  NAND2_X1 U19702 ( .A1(n16777), .A2(n16776), .ZN(n16908) );
  MUX2_X1 U19703 ( .A(n16778), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(
        n10319), .Z(n16783) );
  INV_X1 U19704 ( .A(n16783), .ZN(n16779) );
  AOI222_X1 U19705 ( .A1(n16908), .A2(n16943), .B1(n16780), .B2(n16938), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n16779), .ZN(n16782) );
  AOI21_X1 U19706 ( .B1(n16904), .B2(n16943), .A(n16833), .ZN(n16781) );
  OAI22_X1 U19707 ( .A1(n16782), .A2(n16833), .B1(n16781), .B2(n16905), .ZN(
        P2_U3601) );
  NAND2_X1 U19708 ( .A1(n16783), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n16811) );
  NAND2_X1 U19709 ( .A1(n10319), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16784) );
  NAND2_X1 U19710 ( .A1(n16785), .A2(n16784), .ZN(n16813) );
  NAND2_X1 U19711 ( .A1(n16787), .A2(n16786), .ZN(n16796) );
  INV_X1 U19712 ( .A(n16788), .ZN(n16791) );
  INV_X1 U19713 ( .A(n16789), .ZN(n16790) );
  NAND2_X1 U19714 ( .A1(n16791), .A2(n16790), .ZN(n16793) );
  AOI22_X1 U19715 ( .A1(n16794), .A2(n16793), .B1(n16904), .B2(n16792), .ZN(
        n16795) );
  NAND2_X1 U19716 ( .A1(n16796), .A2(n16795), .ZN(n16909) );
  AOI22_X1 U19717 ( .A1(n20769), .A2(n16938), .B1(n16909), .B2(n16943), .ZN(
        n16797) );
  OAI21_X1 U19718 ( .B1(n16811), .B2(n16813), .A(n16797), .ZN(n16798) );
  MUX2_X1 U19719 ( .A(n16798), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16833), .Z(P2_U3600) );
  OR2_X1 U19720 ( .A1(n13869), .A2(n16816), .ZN(n16810) );
  NAND2_X1 U19721 ( .A1(n16800), .A2(n16799), .ZN(n16801) );
  NAND2_X1 U19722 ( .A1(n16801), .A2(n12641), .ZN(n16825) );
  NOR2_X1 U19723 ( .A1(n11537), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16822) );
  AND2_X1 U19724 ( .A1(n16803), .A2(n16802), .ZN(n16820) );
  OAI21_X1 U19725 ( .B1(n16825), .B2(n16822), .A(n16820), .ZN(n16808) );
  INV_X1 U19726 ( .A(n16822), .ZN(n16804) );
  NAND3_X1 U19727 ( .A1(n16825), .A2(n12641), .A3(n16804), .ZN(n16807) );
  NOR2_X1 U19728 ( .A1(n16805), .A2(n16821), .ZN(n16806) );
  AOI22_X1 U19729 ( .A1(n16808), .A2(n16807), .B1(n16806), .B2(n16904), .ZN(
        n16809) );
  NAND2_X1 U19730 ( .A1(n16810), .A2(n16809), .ZN(n16893) );
  INV_X1 U19731 ( .A(n16811), .ZN(n16812) );
  AOI222_X1 U19732 ( .A1(n16943), .A2(n16893), .B1(n20762), .B2(n16938), .C1(
        n16813), .C2(n16812), .ZN(n16815) );
  NAND2_X1 U19733 ( .A1(n16833), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16814) );
  OAI21_X1 U19734 ( .B1(n16815), .B2(n16833), .A(n16814), .ZN(P2_U3599) );
  OR2_X1 U19735 ( .A1(n16817), .A2(n16816), .ZN(n16830) );
  AOI21_X1 U19736 ( .B1(n16904), .B2(n16821), .A(n16818), .ZN(n16819) );
  OAI21_X1 U19737 ( .B1(n16820), .B2(n16822), .A(n16819), .ZN(n16827) );
  INV_X1 U19738 ( .A(n16821), .ZN(n16823) );
  AOI21_X1 U19739 ( .B1(n16904), .B2(n16823), .A(n16822), .ZN(n16824) );
  NAND2_X1 U19740 ( .A1(n16825), .A2(n16824), .ZN(n16826) );
  MUX2_X1 U19741 ( .A(n16827), .B(n16826), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n16828) );
  INV_X1 U19742 ( .A(n16828), .ZN(n16829) );
  NAND2_X1 U19743 ( .A1(n16830), .A2(n16829), .ZN(n16903) );
  AOI22_X1 U19744 ( .A1(n16831), .A2(n16938), .B1(n16943), .B2(n16903), .ZN(
        n16834) );
  NAND2_X1 U19745 ( .A1(n16833), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16832) );
  OAI21_X1 U19746 ( .B1(n16834), .B2(n16833), .A(n16832), .ZN(P2_U3596) );
  OAI21_X1 U19747 ( .B1(n20312), .B2(n20362), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16836) );
  NAND2_X1 U19748 ( .A1(n20246), .A2(n20276), .ZN(n16835) );
  NAND2_X1 U19749 ( .A1(n16836), .A2(n16835), .ZN(n16846) );
  INV_X1 U19750 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20489) );
  OAI21_X1 U19751 ( .B1(n16837), .B2(n20489), .A(n20800), .ZN(n16844) );
  NAND2_X1 U19752 ( .A1(n20557), .A2(n20758), .ZN(n20338) );
  NOR2_X1 U19753 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20338), .ZN(
        n20327) );
  INV_X1 U19754 ( .A(n20327), .ZN(n16843) );
  INV_X1 U19755 ( .A(n16838), .ZN(n16840) );
  NAND2_X1 U19756 ( .A1(n16840), .A2(n16839), .ZN(n20811) );
  NAND2_X1 U19757 ( .A1(n20811), .A2(n20778), .ZN(n16841) );
  AOI21_X1 U19758 ( .B1(n16844), .B2(n16843), .A(n20494), .ZN(n16845) );
  INV_X1 U19759 ( .A(n20329), .ZN(n20316) );
  INV_X1 U19760 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16854) );
  NOR2_X1 U19761 ( .A1(n20804), .A2(n20395), .ZN(n20767) );
  AOI22_X1 U19762 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n20133), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n20134), .ZN(n20571) );
  AOI22_X1 U19763 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20133), .ZN(n20626) );
  INV_X1 U19764 ( .A(n20626), .ZN(n20558) );
  AOI22_X1 U19765 ( .A1(n20312), .A2(n20621), .B1(n20362), .B2(n20558), .ZN(
        n16853) );
  INV_X1 U19766 ( .A(n20175), .ZN(n16886) );
  OAI21_X1 U19767 ( .B1(n16837), .B2(n20327), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16850) );
  OAI21_X1 U19768 ( .B1(n20274), .B2(n16886), .A(n16850), .ZN(n20328) );
  NOR2_X2 U19769 ( .A1(n20494), .A2(n16851), .ZN(n20614) );
  AND2_X1 U19770 ( .A1(n20136), .A2(n20807), .ZN(n20613) );
  AOI22_X1 U19771 ( .A1(n20328), .A2(n20614), .B1(n20613), .B2(n20327), .ZN(
        n16852) );
  OAI211_X1 U19772 ( .C1(n20316), .C2(n16854), .A(n16853), .B(n16852), .ZN(
        P2_U3096) );
  INV_X1 U19773 ( .A(n20614), .ZN(n16871) );
  NOR2_X4 U19774 ( .A1(n20752), .A2(n20205), .ZN(n20388) );
  OR2_X1 U19775 ( .A1(n20804), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20748) );
  NAND2_X1 U19776 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20766), .ZN(
        n20455) );
  NOR2_X1 U19777 ( .A1(n20247), .A2(n20455), .ZN(n16866) );
  OAI21_X1 U19778 ( .B1(n16862), .B2(n16866), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16860) );
  INV_X1 U19779 ( .A(n16859), .ZN(n20360) );
  NOR2_X1 U19780 ( .A1(n20360), .A2(n16866), .ZN(n16864) );
  INV_X1 U19781 ( .A(n20389), .ZN(n16880) );
  INV_X1 U19782 ( .A(n16861), .ZN(n16865) );
  AOI211_X1 U19783 ( .C1(n16862), .C2(n20800), .A(n20749), .B(n16866), .ZN(
        n16863) );
  INV_X1 U19784 ( .A(n20393), .ZN(n16877) );
  NOR2_X1 U19785 ( .A1(n20626), .A2(n20426), .ZN(n16869) );
  INV_X1 U19786 ( .A(n20388), .ZN(n16874) );
  INV_X1 U19787 ( .A(n20613), .ZN(n16867) );
  INV_X1 U19788 ( .A(n16866), .ZN(n20386) );
  OAI22_X1 U19789 ( .A1(n20571), .A2(n16874), .B1(n16867), .B2(n20386), .ZN(
        n16868) );
  AOI211_X1 U19790 ( .C1(n16877), .C2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n16869), .B(n16868), .ZN(n16870) );
  OAI21_X1 U19791 ( .B1(n16871), .B2(n16880), .A(n16870), .ZN(P2_U3112) );
  NOR2_X2 U19792 ( .A1(n20494), .A2(n16872), .ZN(n20665) );
  INV_X1 U19793 ( .A(n20665), .ZN(n16879) );
  AOI22_X1 U19794 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n20133), .ZN(n20610) );
  NOR2_X1 U19795 ( .A1(n20610), .A2(n20426), .ZN(n16876) );
  AOI22_X2 U19796 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n20133), .ZN(n20673) );
  NAND2_X1 U19797 ( .A1(n20136), .A2(n16873), .ZN(n20602) );
  OAI22_X1 U19798 ( .A1(n20673), .A2(n16874), .B1(n20386), .B2(n20602), .ZN(
        n16875) );
  AOI211_X1 U19799 ( .C1(n16877), .C2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n16876), .B(n16875), .ZN(n16878) );
  OAI21_X1 U19800 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(P2_U3119) );
  NOR2_X1 U19801 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20455), .ZN(
        n20399) );
  NAND2_X1 U19802 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20399), .ZN(
        n20425) );
  OAI221_X1 U19803 ( .B1(n20395), .B2(n20432), .C1(n20395), .C2(n20485), .A(
        n20425), .ZN(n16881) );
  NOR2_X1 U19804 ( .A1(n20776), .A2(n20455), .ZN(n20464) );
  INV_X1 U19805 ( .A(n20464), .ZN(n20454) );
  NOR2_X1 U19806 ( .A1(n20454), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20447) );
  AOI21_X1 U19807 ( .B1(n20749), .B2(n16881), .A(n20447), .ZN(n16882) );
  NAND2_X1 U19808 ( .A1(n16883), .A2(n20619), .ZN(n20450) );
  INV_X1 U19809 ( .A(n20450), .ZN(n20438) );
  OAI21_X1 U19810 ( .B1(n16884), .B2(n20447), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16885) );
  NOR2_X2 U19811 ( .A1(n20494), .A2(n20025), .ZN(n20628) );
  NAND2_X1 U19812 ( .A1(n20136), .A2(n16887), .ZN(n20572) );
  INV_X1 U19813 ( .A(n20447), .ZN(n16889) );
  AOI22_X1 U19814 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20133), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n20134), .ZN(n20632) );
  INV_X1 U19815 ( .A(n20632), .ZN(n20499) );
  AOI22_X1 U19816 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20133), .ZN(n20576) );
  INV_X1 U19817 ( .A(n20576), .ZN(n20629) );
  AOI22_X1 U19818 ( .A1(n20449), .A2(n20499), .B1(n20475), .B2(n20629), .ZN(
        n16888) );
  OAI21_X1 U19819 ( .B1(n20572), .B2(n16889), .A(n16888), .ZN(n16890) );
  AOI21_X1 U19820 ( .B1(n20448), .B2(n20628), .A(n16890), .ZN(n16891) );
  OAI21_X1 U19821 ( .B1(n20438), .B2(n16892), .A(n16891), .ZN(P2_U3129) );
  OR2_X1 U19822 ( .A1(n20801), .A2(n20489), .ZN(n16931) );
  MUX2_X1 U19823 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16903), .S(
        n16925), .Z(n16928) );
  MUX2_X1 U19824 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16893), .S(
        n16925), .Z(n16927) );
  MUX2_X1 U19825 ( .A(n16896), .B(n16895), .S(n16894), .Z(n16901) );
  INV_X1 U19826 ( .A(n16897), .ZN(n16898) );
  AND2_X1 U19827 ( .A1(n16899), .A2(n16898), .ZN(n16900) );
  NOR2_X1 U19828 ( .A1(n16901), .A2(n16900), .ZN(n20796) );
  INV_X1 U19829 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16902) );
  NAND2_X1 U19830 ( .A1(n13536), .A2(n16902), .ZN(n16921) );
  INV_X1 U19831 ( .A(n16903), .ZN(n16912) );
  INV_X1 U19832 ( .A(n16904), .ZN(n16906) );
  OAI21_X1 U19833 ( .B1(n16906), .B2(n16905), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16907) );
  AOI211_X1 U19834 ( .C1(n20776), .C2(n16909), .A(n16908), .B(n16907), .ZN(
        n16911) );
  OAI21_X1 U19835 ( .B1(n20776), .B2(n16909), .A(n16925), .ZN(n16910) );
  AOI211_X1 U19836 ( .C1(n16912), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16911), .B(n16910), .ZN(n16916) );
  INV_X1 U19837 ( .A(n16928), .ZN(n16914) );
  OAI21_X1 U19838 ( .B1(n16916), .B2(n20766), .A(n16927), .ZN(n16913) );
  NAND2_X1 U19839 ( .A1(n16914), .A2(n16913), .ZN(n16915) );
  AOI22_X1 U19840 ( .A1(n16916), .A2(n20766), .B1(n20758), .B2(n16915), .ZN(
        n16919) );
  NAND2_X1 U19841 ( .A1(n11887), .A2(n20807), .ZN(n16917) );
  OAI211_X1 U19842 ( .C1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16919), .A(
        n16918), .B(n16917), .ZN(n16920) );
  AOI21_X1 U19843 ( .B1(n16922), .B2(n16921), .A(n16920), .ZN(n16923) );
  OAI211_X1 U19844 ( .C1(n16925), .C2(n16924), .A(n20796), .B(n16923), .ZN(
        n16926) );
  AOI21_X1 U19845 ( .B1(n16928), .B2(n16927), .A(n16926), .ZN(n16933) );
  INV_X1 U19846 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16929) );
  AOI21_X1 U19847 ( .B1(n16933), .B2(n16929), .A(n20808), .ZN(n16930) );
  AOI211_X2 U19848 ( .C1(n16932), .C2(n11897), .A(n16931), .B(n16930), .ZN(
        n16950) );
  AOI21_X1 U19849 ( .B1(n20489), .B2(n20686), .A(n16950), .ZN(n16942) );
  INV_X1 U19850 ( .A(n16933), .ZN(n16936) );
  OAI21_X1 U19851 ( .B1(n20779), .B2(n17507), .A(n16934), .ZN(n16935) );
  AOI21_X1 U19852 ( .B1(n16936), .B2(n20026), .A(n16935), .ZN(n16941) );
  INV_X1 U19853 ( .A(n16950), .ZN(n16945) );
  INV_X1 U19854 ( .A(n20811), .ZN(n16937) );
  OAI21_X1 U19855 ( .B1(n16938), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16937), 
        .ZN(n16939) );
  OAI21_X1 U19856 ( .B1(n16945), .B2(n20812), .A(n16939), .ZN(n16940) );
  OAI211_X1 U19857 ( .C1(n16942), .C2(n20808), .A(n16941), .B(n16940), .ZN(
        P2_U3176) );
  AOI21_X1 U19858 ( .B1(n16944), .B2(n16943), .A(n20026), .ZN(n16949) );
  OAI21_X1 U19859 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20808), .A(n16945), 
        .ZN(n16946) );
  NAND3_X1 U19860 ( .A1(n16946), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n20686), 
        .ZN(n16948) );
  OAI211_X1 U19861 ( .C1(n16950), .C2(n16949), .A(n16948), .B(n16947), .ZN(
        P2_U3177) );
  OAI21_X1 U19862 ( .B1(n16950), .B2(n20808), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n16951) );
  NAND2_X1 U19863 ( .A1(n16951), .A2(n17507), .ZN(P2_U3593) );
  INV_X1 U19864 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19361) );
  NOR3_X1 U19865 ( .A1(n16952), .A2(n18651), .A3(n18707), .ZN(n16953) );
  NOR2_X1 U19866 ( .A1(n17397), .A2(n18643), .ZN(n18626) );
  NAND2_X1 U19867 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n18504) );
  NAND2_X1 U19868 ( .A1(n9734), .A2(n10427), .ZN(n18505) );
  NOR2_X1 U19869 ( .A1(n18504), .A2(n18505), .ZN(n16955) );
  AOI21_X1 U19870 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n18643), .A(n16955), .ZN(
        n16970) );
  INV_X1 U19871 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18697) );
  NAND2_X1 U19872 ( .A1(n17397), .A2(n10427), .ZN(n18632) );
  NAND2_X1 U19873 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n16957) );
  NAND2_X1 U19874 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n16956) );
  OAI211_X1 U19875 ( .C1(n18455), .C2(n16958), .A(n16957), .B(n16956), .ZN(
        n16959) );
  INV_X1 U19876 ( .A(n16959), .ZN(n16963) );
  AOI22_X1 U19877 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U19878 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16961) );
  NAND2_X1 U19879 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n16960) );
  NAND4_X1 U19880 ( .A1(n16963), .A2(n16962), .A3(n16961), .A4(n16960), .ZN(
        n16969) );
  AOI22_X1 U19881 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U19882 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U19883 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U19884 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16964) );
  NAND4_X1 U19885 ( .A1(n16967), .A2(n16966), .A3(n16965), .A4(n16964), .ZN(
        n16968) );
  INV_X1 U19886 ( .A(n17124), .ZN(n17113) );
  OAI222_X1 U19887 ( .A1(n19361), .A2(n18648), .B1(n16970), .B2(n18642), .C1(
        n18645), .C2(n17113), .ZN(P3_U2733) );
  AOI22_X1 U19888 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18626), .B1(
        P3_EAX_REG_1__SCAN_IN), .B2(n16973), .ZN(n16972) );
  INV_X1 U19889 ( .A(n18505), .ZN(n18628) );
  OAI211_X1 U19890 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n18628), .B(n18504), .ZN(n16971) );
  OAI211_X1 U19891 ( .C1(n17048), .C2(n18645), .A(n16972), .B(n16971), .ZN(
        P3_U2734) );
  NAND2_X1 U19892 ( .A1(n18626), .A2(BUF2_REG_0__SCAN_IN), .ZN(n16975) );
  AOI22_X1 U19893 ( .A1(n16973), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n18625), .B2(
        n17127), .ZN(n16974) );
  OAI211_X1 U19894 ( .C1(P3_EAX_REG_0__SCAN_IN), .C2(n18505), .A(n16975), .B(
        n16974), .ZN(P3_U2735) );
  INV_X1 U19895 ( .A(n17054), .ZN(n16990) );
  NAND2_X1 U19896 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n16977) );
  NAND2_X1 U19897 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n16976) );
  OAI211_X1 U19898 ( .C1(n18455), .C2(n16978), .A(n16977), .B(n16976), .ZN(
        n16979) );
  INV_X1 U19899 ( .A(n16979), .ZN(n16983) );
  AOI22_X1 U19900 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U19901 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16981) );
  NAND2_X1 U19902 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n16980) );
  NAND4_X1 U19903 ( .A1(n16983), .A2(n16982), .A3(n16981), .A4(n16980), .ZN(
        n16989) );
  AOI22_X1 U19904 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U19905 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U19906 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U19907 ( .A1(n14578), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16984) );
  NAND4_X1 U19908 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16988) );
  INV_X1 U19909 ( .A(n17059), .ZN(n17005) );
  NAND2_X1 U19910 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n16992) );
  NAND2_X1 U19911 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n16991) );
  OAI211_X1 U19912 ( .C1(n18455), .C2(n16993), .A(n16992), .B(n16991), .ZN(
        n16994) );
  INV_X1 U19913 ( .A(n16994), .ZN(n16998) );
  AOI22_X1 U19914 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U19915 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16996) );
  NAND2_X1 U19916 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n16995) );
  NAND4_X1 U19917 ( .A1(n16998), .A2(n16997), .A3(n16996), .A4(n16995), .ZN(
        n17004) );
  AOI22_X1 U19918 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U19919 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U19920 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U19921 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16999) );
  NAND4_X1 U19922 ( .A1(n17002), .A2(n17001), .A3(n17000), .A4(n16999), .ZN(
        n17003) );
  NAND2_X1 U19923 ( .A1(n17005), .A2(n17115), .ZN(n17063) );
  INV_X1 U19924 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17448) );
  NAND2_X1 U19925 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n17008) );
  NAND2_X1 U19926 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n17007) );
  OAI211_X1 U19927 ( .C1(n18455), .C2(n17448), .A(n17008), .B(n17007), .ZN(
        n17009) );
  INV_X1 U19928 ( .A(n17009), .ZN(n17013) );
  AOI22_X1 U19929 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U19930 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17011) );
  NAND2_X1 U19931 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n17010) );
  NAND4_X1 U19932 ( .A1(n17013), .A2(n17012), .A3(n17011), .A4(n17010), .ZN(
        n17019) );
  AOI22_X1 U19933 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U19934 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U19935 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U19936 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17014) );
  NAND4_X1 U19937 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n17014), .ZN(
        n17018) );
  INV_X1 U19938 ( .A(n17069), .ZN(n17034) );
  INV_X1 U19939 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18145) );
  NAND2_X1 U19940 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n17021) );
  NAND2_X1 U19941 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n17020) );
  OAI211_X1 U19942 ( .C1(n18455), .C2(n18145), .A(n17021), .B(n17020), .ZN(
        n17022) );
  INV_X1 U19943 ( .A(n17022), .ZN(n17026) );
  AOI22_X1 U19944 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U19945 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17024) );
  NAND2_X1 U19946 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n17023) );
  NAND4_X1 U19947 ( .A1(n17026), .A2(n17025), .A3(n17024), .A4(n17023), .ZN(
        n17033) );
  AOI22_X1 U19948 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17031) );
  INV_X1 U19949 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n21743) );
  AOI22_X1 U19950 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U19951 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U19952 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U19953 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17032) );
  INV_X1 U19954 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18329) );
  NAND2_X1 U19955 ( .A1(n18459), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n17036) );
  NAND2_X1 U19956 ( .A1(n18254), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n17035) );
  OAI211_X1 U19957 ( .C1(n18455), .C2(n18329), .A(n17036), .B(n17035), .ZN(
        n17037) );
  INV_X1 U19958 ( .A(n17037), .ZN(n17041) );
  AOI22_X1 U19959 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U19960 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17039) );
  NAND2_X1 U19961 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n17038) );
  NAND4_X1 U19962 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        n17047) );
  AOI22_X1 U19963 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U19964 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U19965 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U19966 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U19967 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  NAND2_X1 U19968 ( .A1(n17048), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17049) );
  INV_X1 U19969 ( .A(n17051), .ZN(n17052) );
  NAND2_X1 U19970 ( .A1(n17052), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17053) );
  INV_X1 U19971 ( .A(n17114), .ZN(n18644) );
  NAND2_X1 U19972 ( .A1(n18644), .A2(n17054), .ZN(n17055) );
  NAND2_X1 U19973 ( .A1(n17059), .A2(n17055), .ZN(n17056) );
  INV_X1 U19974 ( .A(n17056), .ZN(n17057) );
  INV_X1 U19975 ( .A(n17115), .ZN(n18639) );
  XNOR2_X1 U19976 ( .A(n17059), .B(n18639), .ZN(n17060) );
  XNOR2_X1 U19977 ( .A(n17060), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19015) );
  INV_X1 U19978 ( .A(n17060), .ZN(n17061) );
  NAND2_X1 U19979 ( .A1(n17061), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17062) );
  NAND2_X1 U19980 ( .A1(n17063), .A2(n18635), .ZN(n17064) );
  NAND2_X1 U19981 ( .A1(n17069), .A2(n17064), .ZN(n17065) );
  XNOR2_X1 U19982 ( .A(n17067), .B(n17065), .ZN(n18999) );
  INV_X1 U19983 ( .A(n17065), .ZN(n17066) );
  NAND2_X1 U19984 ( .A1(n17067), .A2(n17066), .ZN(n17068) );
  INV_X1 U19985 ( .A(n17116), .ZN(n18631) );
  NAND2_X1 U19986 ( .A1(n17069), .A2(n18631), .ZN(n17070) );
  NAND2_X1 U19987 ( .A1(n17333), .A2(n17070), .ZN(n17071) );
  XNOR2_X1 U19988 ( .A(n17071), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18986) );
  INV_X1 U19989 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n19270) );
  NAND2_X1 U19990 ( .A1(n17333), .A2(n17330), .ZN(n17073) );
  NAND2_X1 U19991 ( .A1(n18830), .A2(n17073), .ZN(n17074) );
  XNOR2_X1 U19992 ( .A(n17076), .B(n17074), .ZN(n18977) );
  INV_X1 U19993 ( .A(n17074), .ZN(n17075) );
  NAND2_X1 U19994 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n19235) );
  NOR2_X1 U19995 ( .A1(n19235), .A2(n17241), .ZN(n19213) );
  NAND2_X1 U19996 ( .A1(n19210), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n19184) );
  INV_X1 U19997 ( .A(n19184), .ZN(n17078) );
  NAND2_X1 U19998 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17078), .ZN(
        n19163) );
  INV_X1 U19999 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17081) );
  NOR2_X1 U20000 ( .A1(n19163), .A2(n17081), .ZN(n17342) );
  INV_X1 U20001 ( .A(n17342), .ZN(n19147) );
  INV_X1 U20002 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17080) );
  INV_X1 U20003 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17259) );
  INV_X1 U20004 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20005 ( .A1(n17080), .A2(n17259), .A3(n17079), .A4(n17241), .ZN(
        n18907) );
  INV_X1 U20006 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n19187) );
  INV_X1 U20007 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17224) );
  NAND3_X1 U20008 ( .A1(n19187), .A2(n17224), .A3(n17081), .ZN(n17082) );
  INV_X1 U20009 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19143) );
  AND2_X1 U20010 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n19108) );
  INV_X1 U20011 ( .A(n19108), .ZN(n19140) );
  INV_X1 U20012 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19136) );
  INV_X1 U20013 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n19093) );
  NOR2_X1 U20014 ( .A1(n19136), .A2(n19093), .ZN(n19095) );
  AND3_X1 U20015 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n19095), .ZN(n18818) );
  AND2_X1 U20016 ( .A1(n18818), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17284) );
  AND2_X1 U20017 ( .A1(n17284), .A2(n19108), .ZN(n17283) );
  NAND2_X1 U20018 ( .A1(n17283), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18782) );
  AND2_X1 U20019 ( .A1(n18830), .A2(n19105), .ZN(n18871) );
  NAND2_X1 U20020 ( .A1(n18871), .A2(n19136), .ZN(n17083) );
  NOR2_X1 U20021 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17083), .ZN(
        n18833) );
  INV_X1 U20022 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n19114) );
  NAND2_X1 U20023 ( .A1(n18833), .A2(n19114), .ZN(n18806) );
  INV_X1 U20024 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18799) );
  INV_X1 U20025 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n19089) );
  NAND2_X1 U20026 ( .A1(n18799), .A2(n19089), .ZN(n17084) );
  OAI22_X1 U20027 ( .A1(n18889), .A2(n18782), .B1(n18806), .B2(n17084), .ZN(
        n17085) );
  INV_X1 U20028 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17374) );
  NAND2_X1 U20029 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17361) );
  NAND2_X1 U20030 ( .A1(n18910), .A2(n17361), .ZN(n17086) );
  INV_X1 U20031 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17355) );
  NAND2_X1 U20032 ( .A1(n17091), .A2(n17355), .ZN(n17337) );
  INV_X1 U20033 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17338) );
  NAND2_X1 U20034 ( .A1(n18830), .A2(n17338), .ZN(n17087) );
  INV_X1 U20035 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17303) );
  NAND2_X1 U20036 ( .A1(n17162), .A2(n17303), .ZN(n17146) );
  INV_X1 U20037 ( .A(n17146), .ZN(n17090) );
  OAI21_X1 U20038 ( .B1(n18910), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17089) );
  INV_X1 U20039 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17407) );
  AND2_X1 U20040 ( .A1(n18830), .A2(n17407), .ZN(n17093) );
  INV_X1 U20041 ( .A(n17093), .ZN(n17088) );
  OAI211_X1 U20042 ( .C1(n17090), .C2(n18910), .A(n17089), .B(n17088), .ZN(
        n17098) );
  NAND2_X1 U20043 ( .A1(n18910), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17092) );
  NOR2_X2 U20044 ( .A1(n17350), .A2(n17092), .ZN(n17161) );
  NAND2_X1 U20045 ( .A1(n17161), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17164) );
  INV_X1 U20046 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21756) );
  NOR2_X1 U20047 ( .A1(n17164), .A2(n21756), .ZN(n17097) );
  OAI21_X1 U20048 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n21756), .A(
        n17164), .ZN(n17094) );
  OAI21_X1 U20049 ( .B1(n17094), .B2(n17146), .A(n17093), .ZN(n17096) );
  NAND3_X1 U20050 ( .A1(n17094), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n17095) );
  OAI211_X1 U20051 ( .C1(n17098), .C2(n17097), .A(n17096), .B(n17095), .ZN(
        n17300) );
  NOR2_X4 U20052 ( .A1(n17710), .A2(n19943), .ZN(n19051) );
  NAND2_X1 U20053 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19341) );
  NAND2_X1 U20054 ( .A1(n19923), .A2(n19341), .ZN(n19937) );
  INV_X1 U20055 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19832) );
  NOR2_X1 U20056 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19832), .ZN(n18811) );
  NAND2_X1 U20057 ( .A1(n19000), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18989) );
  NAND2_X1 U20058 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n18925), .ZN(
        n18895) );
  NAND2_X1 U20059 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18897) );
  INV_X1 U20060 ( .A(n18897), .ZN(n17099) );
  NAND2_X1 U20061 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18767) );
  INV_X1 U20062 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17215) );
  NAND2_X1 U20063 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17182) );
  NAND2_X1 U20064 ( .A1(n18649), .A2(n19832), .ZN(n19842) );
  INV_X1 U20065 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19942) );
  INV_X1 U20066 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17763) );
  AND2_X1 U20067 ( .A1(n17213), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17202) );
  NAND3_X1 U20068 ( .A1(n17202), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17170) );
  NOR2_X1 U20069 ( .A1(n17763), .A2(n17170), .ZN(n17109) );
  OR2_X1 U20070 ( .A1(n19690), .A2(n17109), .ZN(n17171) );
  INV_X1 U20071 ( .A(n17171), .ZN(n17101) );
  AOI21_X1 U20072 ( .B1(n18811), .B2(n17187), .A(n17101), .ZN(n17102) );
  NAND2_X1 U20073 ( .A1(n9715), .A2(n17102), .ZN(n17175) );
  NOR2_X1 U20074 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18809), .ZN(
        n17167) );
  OR2_X1 U20075 ( .A1(n17175), .A2(n17167), .ZN(n17153) );
  NAND2_X1 U20076 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n17166), .ZN(
        n17103) );
  NAND2_X1 U20077 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18813) );
  NAND2_X2 U20078 ( .A1(n9714), .A2(n18813), .ZN(n19049) );
  AND2_X2 U20079 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17104), .ZN(n18858) );
  INV_X2 U20080 ( .A(n18858), .ZN(n18937) );
  AND2_X2 U20081 ( .A1(n19051), .A2(n17330), .ZN(n18934) );
  INV_X1 U20082 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n19070) );
  NAND2_X1 U20083 ( .A1(n18931), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19170) );
  NOR2_X1 U20084 ( .A1(n19170), .A2(n18782), .ZN(n19072) );
  NAND2_X1 U20085 ( .A1(n19072), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18772) );
  NOR2_X1 U20086 ( .A1(n19070), .A2(n18772), .ZN(n18771) );
  AND2_X1 U20087 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17278) );
  NAND2_X1 U20088 ( .A1(n17278), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17288) );
  INV_X1 U20089 ( .A(n17288), .ZN(n17142) );
  AND2_X1 U20090 ( .A1(n17363), .A2(n17142), .ZN(n17306) );
  NAND2_X1 U20091 ( .A1(n17306), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17106) );
  XNOR2_X1 U20092 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n17106), .ZN(
        n17292) );
  NAND2_X1 U20093 ( .A1(n18934), .A2(n17292), .ZN(n17107) );
  NAND2_X1 U20094 ( .A1(n19268), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n17290) );
  OAI211_X1 U20095 ( .C1(n18098), .C2(n18937), .A(n17107), .B(n17290), .ZN(
        n17112) );
  NOR2_X1 U20096 ( .A1(n18809), .A2(n18110), .ZN(n17108) );
  OR2_X2 U20097 ( .A1(n17108), .A2(n19730), .ZN(n18855) );
  NAND2_X1 U20098 ( .A1(n18855), .A2(n17109), .ZN(n17156) );
  INV_X1 U20099 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17749) );
  XOR2_X1 U20100 ( .A(n17749), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n17110) );
  NOR2_X1 U20101 ( .A1(n17156), .A2(n17110), .ZN(n17111) );
  AOI211_X1 U20102 ( .C1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n17153), .A(
        n17112), .B(n17111), .ZN(n17145) );
  NAND2_X1 U20103 ( .A1(n17125), .A2(n17113), .ZN(n17122) );
  NAND2_X1 U20104 ( .A1(n17121), .A2(n17115), .ZN(n17119) );
  NOR2_X1 U20105 ( .A1(n18635), .A2(n17119), .ZN(n17118) );
  NAND2_X1 U20106 ( .A1(n17118), .A2(n17116), .ZN(n17117) );
  NOR2_X1 U20107 ( .A1(n17330), .A2(n17117), .ZN(n17140) );
  XNOR2_X1 U20108 ( .A(n18624), .B(n17117), .ZN(n18968) );
  XNOR2_X1 U20109 ( .A(n18631), .B(n17118), .ZN(n17134) );
  XOR2_X1 U20110 ( .A(n18635), .B(n17119), .Z(n17120) );
  NAND2_X1 U20111 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17120), .ZN(
        n17133) );
  INV_X1 U20112 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18998) );
  XNOR2_X1 U20113 ( .A(n18998), .B(n17120), .ZN(n18997) );
  INV_X1 U20114 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n21879) );
  XNOR2_X1 U20115 ( .A(n18639), .B(n17121), .ZN(n19010) );
  XNOR2_X1 U20116 ( .A(n17122), .B(n18644), .ZN(n17123) );
  NAND2_X1 U20117 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17123), .ZN(
        n17131) );
  INV_X1 U20118 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21882) );
  XNOR2_X1 U20119 ( .A(n21882), .B(n17123), .ZN(n19025) );
  XNOR2_X1 U20120 ( .A(n17125), .B(n17124), .ZN(n17126) );
  INV_X1 U20121 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n19328) );
  OR2_X1 U20122 ( .A1(n17126), .A2(n19328), .ZN(n17130) );
  XNOR2_X1 U20123 ( .A(n17126), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19034) );
  NOR2_X1 U20124 ( .A1(n17129), .A2(n17128), .ZN(n19033) );
  NAND2_X1 U20125 ( .A1(n19034), .A2(n19033), .ZN(n19032) );
  NAND2_X1 U20126 ( .A1(n17130), .A2(n19032), .ZN(n19024) );
  NAND2_X1 U20127 ( .A1(n19025), .A2(n19024), .ZN(n19023) );
  NAND2_X1 U20128 ( .A1(n17131), .A2(n19023), .ZN(n19011) );
  NAND2_X1 U20129 ( .A1(n19010), .A2(n19011), .ZN(n19009) );
  NOR2_X1 U20130 ( .A1(n19010), .A2(n19011), .ZN(n17132) );
  AOI21_X1 U20131 ( .B1(n21879), .B2(n19009), .A(n17132), .ZN(n18996) );
  NAND2_X1 U20132 ( .A1(n18997), .A2(n18996), .ZN(n18995) );
  NAND2_X1 U20133 ( .A1(n17133), .A2(n18995), .ZN(n17135) );
  NAND2_X1 U20134 ( .A1(n17134), .A2(n17135), .ZN(n17136) );
  NAND2_X1 U20135 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18983), .ZN(
        n18982) );
  INV_X1 U20136 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n19261) );
  NAND2_X1 U20137 ( .A1(n17140), .A2(n17137), .ZN(n17141) );
  NAND2_X1 U20138 ( .A1(n18968), .A2(n18969), .ZN(n18967) );
  NAND2_X1 U20139 ( .A1(n17140), .A2(n17139), .ZN(n17138) );
  OAI211_X1 U20140 ( .C1(n17140), .C2(n17139), .A(n18967), .B(n17138), .ZN(
        n17267) );
  NAND2_X1 U20141 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17267), .ZN(
        n17266) );
  NOR2_X2 U20142 ( .A1(n18782), .A2(n19171), .ZN(n19071) );
  NAND2_X1 U20143 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n19071), .ZN(
        n18774) );
  NOR2_X2 U20144 ( .A1(n18774), .A2(n17361), .ZN(n17356) );
  NAND2_X1 U20145 ( .A1(n17356), .A2(n17278), .ZN(n17276) );
  NAND3_X1 U20146 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n17407), .ZN(n17281) );
  NOR2_X1 U20147 ( .A1(n17276), .A2(n17281), .ZN(n17143) );
  AND2_X1 U20148 ( .A1(n17356), .A2(n17142), .ZN(n17304) );
  AOI21_X1 U20149 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17304), .A(
        n17407), .ZN(n17293) );
  NOR2_X2 U20150 ( .A1(n17710), .A2(n18707), .ZN(n19048) );
  OAI21_X1 U20151 ( .B1(n17143), .B2(n17293), .A(n19048), .ZN(n17144) );
  OAI211_X1 U20152 ( .C1(n17300), .C2(n18966), .A(n17145), .B(n17144), .ZN(
        P3_U2799) );
  NAND2_X1 U20153 ( .A1(n17164), .A2(n17146), .ZN(n17147) );
  XNOR2_X1 U20154 ( .A(n17147), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17315) );
  NOR2_X1 U20155 ( .A1(n17304), .A2(n19040), .ZN(n17176) );
  INV_X1 U20156 ( .A(n17176), .ZN(n17149) );
  INV_X1 U20157 ( .A(n17306), .ZN(n17148) );
  NAND2_X1 U20158 ( .A1(n17148), .A2(n18934), .ZN(n17172) );
  AOI21_X1 U20159 ( .B1(n17149), .B2(n17172), .A(n21756), .ZN(n17159) );
  NAND2_X1 U20160 ( .A1(n18934), .A2(n10313), .ZN(n17151) );
  NAND2_X1 U20161 ( .A1(n17339), .A2(n19048), .ZN(n17150) );
  NAND2_X2 U20162 ( .A1(n17151), .A2(n17150), .ZN(n18960) );
  AND2_X2 U20163 ( .A1(n18960), .A2(n17342), .ZN(n18901) );
  NAND2_X1 U20164 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n19060) );
  NOR2_X1 U20165 ( .A1(n17361), .A2(n19060), .ZN(n17366) );
  INV_X1 U20166 ( .A(n17366), .ZN(n17152) );
  NOR4_X1 U20167 ( .A1(n18798), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17152), .A4(n17288), .ZN(n17158) );
  INV_X1 U20168 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17753) );
  XNOR2_X1 U20169 ( .A(n17166), .B(n17753), .ZN(n17752) );
  INV_X2 U20170 ( .A(n19268), .ZN(n19156) );
  INV_X1 U20171 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19908) );
  NOR2_X1 U20172 ( .A1(n19156), .A2(n19908), .ZN(n17312) );
  AOI21_X1 U20173 ( .B1(n17752), .B2(n18858), .A(n17312), .ZN(n17155) );
  NAND2_X1 U20174 ( .A1(n17153), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17154) );
  OAI211_X1 U20175 ( .C1(n17156), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n17155), .B(n17154), .ZN(n17157) );
  NOR3_X1 U20176 ( .A1(n17159), .A2(n17158), .A3(n17157), .ZN(n17160) );
  OAI21_X1 U20177 ( .B1(n17315), .B2(n18966), .A(n17160), .ZN(P3_U2800) );
  NOR2_X1 U20178 ( .A1(n17161), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17163) );
  INV_X1 U20179 ( .A(n17164), .ZN(n17165) );
  INV_X1 U20180 ( .A(n17316), .ZN(n17179) );
  AOI21_X1 U20181 ( .B1(n17187), .B2(n17763), .A(n17166), .ZN(n17762) );
  OAI21_X1 U20182 ( .B1(n17167), .B2(n18858), .A(n17762), .ZN(n17169) );
  AND2_X1 U20183 ( .A1(n19268), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n17322) );
  INV_X1 U20184 ( .A(n17322), .ZN(n17168) );
  OAI211_X1 U20185 ( .C1(n17171), .C2(n17170), .A(n17169), .B(n17168), .ZN(
        n17174) );
  NAND2_X1 U20186 ( .A1(n17363), .A2(n17278), .ZN(n17329) );
  AOI21_X1 U20187 ( .B1(n17303), .B2(n17329), .A(n17172), .ZN(n17173) );
  AOI211_X1 U20188 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n17175), .A(
        n17174), .B(n17173), .ZN(n17178) );
  INV_X1 U20189 ( .A(n17276), .ZN(n17326) );
  OAI21_X1 U20190 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n17326), .A(
        n17176), .ZN(n17177) );
  OAI211_X1 U20191 ( .C1(n17179), .C2(n18966), .A(n17178), .B(n17177), .ZN(
        P3_U2801) );
  INV_X1 U20192 ( .A(n18934), .ZN(n18820) );
  OR2_X1 U20193 ( .A1(n17356), .A2(n19040), .ZN(n17181) );
  OR2_X1 U20194 ( .A1(n17363), .A2(n18820), .ZN(n17180) );
  NAND2_X1 U20195 ( .A1(n17181), .A2(n17180), .ZN(n17221) );
  NOR2_X1 U20196 ( .A1(n17221), .A2(n17355), .ZN(n17210) );
  AOI211_X1 U20197 ( .C1(n18820), .C2(n19040), .A(n17338), .B(n17210), .ZN(
        n17193) );
  OAI211_X1 U20198 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17202), .B(n17182), .ZN(n17191) );
  NAND2_X1 U20199 ( .A1(n17366), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17282) );
  NOR2_X1 U20200 ( .A1(n17282), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17346) );
  INV_X1 U20201 ( .A(n17346), .ZN(n17183) );
  OR2_X1 U20202 ( .A1(n18798), .A2(n17183), .ZN(n17190) );
  INV_X1 U20203 ( .A(n18811), .ZN(n18892) );
  INV_X1 U20204 ( .A(n17734), .ZN(n17184) );
  OAI22_X1 U20205 ( .A1(n17202), .A2(n18813), .B1(n18892), .B2(n17184), .ZN(
        n17185) );
  INV_X1 U20206 ( .A(n17185), .ZN(n17186) );
  AND2_X1 U20207 ( .A1(n9716), .A2(n17186), .ZN(n17219) );
  OAI21_X1 U20208 ( .B1(n18809), .B2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n17219), .ZN(n17206) );
  INV_X1 U20209 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17784) );
  NOR2_X1 U20210 ( .A1(n10503), .A2(n17784), .ZN(n17199) );
  OAI21_X1 U20211 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17199), .A(
        n17187), .ZN(n17731) );
  NAND2_X1 U20212 ( .A1(n19268), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17348) );
  OAI21_X1 U20213 ( .B1(n18937), .B2(n17731), .A(n17348), .ZN(n17188) );
  AOI21_X1 U20214 ( .B1(n17206), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n17188), .ZN(n17189) );
  OAI211_X1 U20215 ( .C1(n18896), .C2(n17191), .A(n17190), .B(n17189), .ZN(
        n17192) );
  NOR2_X1 U20216 ( .A1(n17193), .A2(n17192), .ZN(n17196) );
  XNOR2_X1 U20217 ( .A(n18830), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17336) );
  OAI211_X1 U20218 ( .C1(n17194), .C2(n17336), .A(n17332), .B(n18946), .ZN(
        n17195) );
  NAND2_X1 U20219 ( .A1(n17196), .A2(n17195), .ZN(P3_U2802) );
  INV_X1 U20220 ( .A(n18798), .ZN(n17197) );
  AOI21_X1 U20221 ( .B1(n17197), .B2(n17366), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17209) );
  NAND2_X1 U20222 ( .A1(n17350), .A2(n17337), .ZN(n17198) );
  XNOR2_X1 U20223 ( .A(n17198), .B(n18830), .ZN(n17370) );
  NAND2_X1 U20224 ( .A1(n17370), .A2(n18946), .ZN(n17208) );
  OR2_X1 U20225 ( .A1(n17214), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17201) );
  INV_X1 U20226 ( .A(n17199), .ZN(n17200) );
  NAND2_X1 U20227 ( .A1(n17201), .A2(n17200), .ZN(n17732) );
  NAND2_X1 U20228 ( .A1(n19268), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20229 ( .B1(n17732), .B2(n18937), .A(n17354), .ZN(n17205) );
  INV_X1 U20230 ( .A(n17202), .ZN(n17203) );
  NOR3_X1 U20231 ( .A1(n18896), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17203), .ZN(n17204) );
  AOI211_X1 U20232 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17206), .A(
        n17205), .B(n17204), .ZN(n17207) );
  OAI211_X1 U20233 ( .C1(n17210), .C2(n17209), .A(n17208), .B(n17207), .ZN(
        P3_U2803) );
  INV_X1 U20234 ( .A(n17211), .ZN(n17212) );
  AOI21_X1 U20235 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n9836), .A(
        n17212), .ZN(n17379) );
  NAND2_X1 U20236 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18773) );
  AOI21_X1 U20237 ( .B1(n17213), .B2(n19730), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17218) );
  INV_X1 U20238 ( .A(n18809), .ZN(n17216) );
  AOI21_X1 U20239 ( .B1(n17734), .B2(n17215), .A(n17214), .ZN(n17796) );
  OAI21_X1 U20240 ( .B1(n18858), .B2(n17216), .A(n17796), .ZN(n17217) );
  NAND2_X1 U20241 ( .A1(n19268), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17373) );
  OAI211_X1 U20242 ( .C1(n17219), .C2(n17218), .A(n17217), .B(n17373), .ZN(
        n17220) );
  NOR2_X1 U20243 ( .A1(n17222), .A2(n18910), .ZN(n18951) );
  NOR2_X1 U20244 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18958) );
  NAND2_X1 U20245 ( .A1(n18951), .A2(n18958), .ZN(n17236) );
  NOR2_X1 U20246 ( .A1(n17236), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18942) );
  NOR3_X1 U20247 ( .A1(n18906), .A2(n18830), .A3(n17224), .ZN(n17223) );
  AOI21_X1 U20248 ( .B1(n18942), .B2(n17224), .A(n17223), .ZN(n17225) );
  XOR2_X1 U20249 ( .A(n17079), .B(n17225), .Z(n19198) );
  INV_X1 U20250 ( .A(n19198), .ZN(n17235) );
  INV_X1 U20251 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18973) );
  NOR2_X1 U20252 ( .A1(n18110), .A2(n18989), .ZN(n18030) );
  NAND2_X1 U20253 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n18030), .ZN(
        n18029) );
  NOR2_X1 U20254 ( .A1(n18973), .A2(n18029), .ZN(n18017) );
  NAND2_X1 U20255 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18017), .ZN(
        n17262) );
  INV_X1 U20256 ( .A(n17262), .ZN(n17255) );
  NAND2_X1 U20257 ( .A1(n17244), .A2(n17255), .ZN(n17243) );
  INV_X1 U20258 ( .A(n17243), .ZN(n17958) );
  INV_X1 U20259 ( .A(n18813), .ZN(n19008) );
  AOI21_X1 U20260 ( .B1(n19008), .B2(n18894), .A(n18811), .ZN(n17226) );
  OAI21_X1 U20261 ( .B1(n17958), .B2(n17226), .A(n9716), .ZN(n18941) );
  INV_X1 U20262 ( .A(n18894), .ZN(n17918) );
  NAND2_X1 U20263 ( .A1(n17918), .A2(n18855), .ZN(n18939) );
  AOI211_X1 U20264 ( .C1(n17227), .C2(n17952), .A(n18925), .B(n18939), .ZN(
        n17229) );
  INV_X1 U20265 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n21778) );
  NOR2_X1 U20266 ( .A1(n17227), .A2(n17243), .ZN(n17941) );
  NAND2_X1 U20267 ( .A1(n18925), .A2(n17958), .ZN(n17935) );
  OAI21_X1 U20268 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17941), .A(
        n17935), .ZN(n17943) );
  OAI22_X1 U20269 ( .A1(n19156), .A2(n21778), .B1(n18937), .B2(n17943), .ZN(
        n17228) );
  AOI211_X1 U20270 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18941), .A(
        n17229), .B(n17228), .ZN(n17234) );
  INV_X1 U20271 ( .A(n19210), .ZN(n17230) );
  NOR2_X1 U20272 ( .A1(n17105), .A2(n17230), .ZN(n19201) );
  INV_X1 U20273 ( .A(n19204), .ZN(n17231) );
  OAI22_X1 U20274 ( .A1(n18820), .A2(n19201), .B1(n19040), .B2(n17231), .ZN(
        n18947) );
  NAND2_X1 U20275 ( .A1(n19210), .A2(n17079), .ZN(n19209) );
  INV_X1 U20276 ( .A(n19209), .ZN(n17232) );
  AOI22_X1 U20277 ( .A1(n18947), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n18960), .B2(n17232), .ZN(n17233) );
  OAI211_X1 U20278 ( .C1(n18966), .C2(n17235), .A(n17234), .B(n17233), .ZN(
        P3_U2817) );
  INV_X1 U20279 ( .A(n19235), .ZN(n17238) );
  NAND2_X1 U20280 ( .A1(n17238), .A2(n17241), .ZN(n19241) );
  OAI21_X1 U20281 ( .B1(n17238), .B2(n17241), .A(n19241), .ZN(n17249) );
  INV_X1 U20282 ( .A(n17339), .ZN(n19223) );
  AOI22_X1 U20283 ( .A1(n18934), .A2(n17105), .B1(n19223), .B2(n19048), .ZN(
        n18962) );
  NAND2_X1 U20284 ( .A1(n10313), .A2(n18910), .ZN(n18944) );
  INV_X1 U20285 ( .A(n18944), .ZN(n18952) );
  INV_X1 U20286 ( .A(n17236), .ZN(n17237) );
  AOI21_X1 U20287 ( .B1(n17238), .B2(n18952), .A(n17237), .ZN(n17239) );
  XNOR2_X1 U20288 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17239), .ZN(
        n19221) );
  INV_X1 U20289 ( .A(n19221), .ZN(n17240) );
  OAI22_X1 U20290 ( .A1(n18962), .A2(n17241), .B1(n18966), .B2(n17240), .ZN(
        n17248) );
  NAND2_X2 U20291 ( .A1(n18809), .A2(n18937), .ZN(n19043) );
  INV_X2 U20292 ( .A(n19043), .ZN(n19054) );
  NAND2_X1 U20293 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17242) );
  NOR2_X1 U20294 ( .A1(n17242), .A2(n17262), .ZN(n17982) );
  OAI21_X1 U20295 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17982), .A(
        n17243), .ZN(n17966) );
  NOR3_X1 U20296 ( .A1(n21671), .A2(n18006), .A3(n19690), .ZN(n17254) );
  AND2_X1 U20297 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17254), .ZN(
        n18954) );
  AND2_X1 U20298 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18954), .ZN(
        n18957) );
  NAND2_X1 U20299 ( .A1(n17244), .A2(n17254), .ZN(n18927) );
  OAI211_X1 U20300 ( .C1(n18957), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19049), .B(n18927), .ZN(n17246) );
  NAND2_X1 U20301 ( .A1(n19268), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17245) );
  OAI211_X1 U20302 ( .C1(n19054), .C2(n17966), .A(n17246), .B(n17245), .ZN(
        n17247) );
  AOI211_X1 U20303 ( .C1(n18960), .C2(n17249), .A(n17248), .B(n17247), .ZN(
        n17250) );
  INV_X1 U20304 ( .A(n17250), .ZN(P3_U2819) );
  NOR2_X1 U20305 ( .A1(n18951), .A2(n18952), .ZN(n17251) );
  XNOR2_X1 U20306 ( .A(n17251), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n19254) );
  NOR2_X1 U20307 ( .A1(n19156), .A2(n21816), .ZN(n17252) );
  AOI21_X1 U20308 ( .B1(n18946), .B2(n19254), .A(n17252), .ZN(n17253) );
  OAI21_X1 U20309 ( .B1(n18962), .B2(n17259), .A(n17253), .ZN(n17258) );
  AOI21_X1 U20310 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19049), .A(
        n17254), .ZN(n17256) );
  NAND2_X1 U20311 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17255), .ZN(
        n17984) );
  OAI21_X1 U20312 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17255), .A(
        n17984), .ZN(n17997) );
  OAI22_X1 U20313 ( .A1(n18954), .A2(n17256), .B1(n19054), .B2(n17997), .ZN(
        n17257) );
  AOI211_X1 U20314 ( .C1(n17259), .C2(n18960), .A(n17258), .B(n17257), .ZN(
        n17260) );
  INV_X1 U20315 ( .A(n17260), .ZN(P3_U2821) );
  XNOR2_X1 U20316 ( .A(n17268), .B(n18910), .ZN(n17396) );
  NOR2_X1 U20317 ( .A1(n18006), .A2(n19690), .ZN(n17265) );
  INV_X1 U20318 ( .A(n17261), .ZN(n18972) );
  INV_X1 U20319 ( .A(n9715), .ZN(n19006) );
  AOI21_X1 U20320 ( .B1(n19008), .B2(n18972), .A(n19006), .ZN(n18974) );
  OAI21_X1 U20321 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19690), .A(
        n18974), .ZN(n17264) );
  OAI21_X1 U20322 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18017), .A(
        n17262), .ZN(n18008) );
  INV_X1 U20323 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19870) );
  OAI22_X1 U20324 ( .A1(n19054), .A2(n18008), .B1(n19156), .B2(n19870), .ZN(
        n17263) );
  AOI221_X1 U20325 ( .B1(n17265), .B2(n21671), .C1(n17264), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n17263), .ZN(n17271) );
  OAI21_X1 U20326 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17267), .A(
        n17266), .ZN(n17392) );
  INV_X1 U20327 ( .A(n17392), .ZN(n17269) );
  INV_X1 U20328 ( .A(n17268), .ZN(n17394) );
  AOI22_X1 U20329 ( .A1(n17269), .A2(n19048), .B1(n17394), .B2(n18934), .ZN(
        n17270) );
  OAI211_X1 U20330 ( .C1(n17396), .C2(n18966), .A(n17271), .B(n17270), .ZN(
        P3_U2822) );
  NOR2_X1 U20331 ( .A1(n17272), .A2(n9808), .ZN(n19330) );
  NAND3_X1 U20332 ( .A1(n18649), .A2(n9716), .A3(n18892), .ZN(n17273) );
  AOI22_X1 U20333 ( .A1(n19268), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17273), .ZN(n17275) );
  NAND2_X1 U20334 ( .A1(n19051), .A2(n19330), .ZN(n17274) );
  OAI211_X1 U20335 ( .C1(n19040), .C2(n19330), .A(n17275), .B(n17274), .ZN(
        P3_U2830) );
  OR2_X1 U20336 ( .A1(n17276), .A2(n19285), .ZN(n17280) );
  NOR3_X1 U20337 ( .A1(n21879), .A2(n21882), .A3(n18998), .ZN(n17382) );
  OAI21_X1 U20338 ( .B1(n17408), .B2(n17406), .A(n19328), .ZN(n19313) );
  NAND2_X1 U20339 ( .A1(n17382), .A2(n19313), .ZN(n17384) );
  INV_X1 U20340 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17389) );
  NOR3_X1 U20341 ( .A1(n19270), .A2(n19261), .A3(n17389), .ZN(n19145) );
  INV_X1 U20342 ( .A(n19145), .ZN(n17277) );
  NOR2_X1 U20343 ( .A1(n17384), .A2(n17277), .ZN(n19227) );
  AND3_X1 U20344 ( .A1(n19108), .A2(n17342), .A3(n19227), .ZN(n19142) );
  OAI21_X1 U20345 ( .B1(n19237), .B2(n17406), .A(n17359), .ZN(n19317) );
  NAND2_X1 U20346 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19289) );
  INV_X1 U20347 ( .A(n19289), .ZN(n17380) );
  NAND2_X1 U20348 ( .A1(n17382), .A2(n17380), .ZN(n17383) );
  OR2_X1 U20349 ( .A1(n17277), .A2(n17383), .ZN(n19161) );
  NOR2_X1 U20350 ( .A1(n19147), .A2(n19161), .ZN(n19138) );
  INV_X1 U20351 ( .A(n19138), .ZN(n19091) );
  NOR2_X1 U20352 ( .A1(n19140), .A2(n19091), .ZN(n17358) );
  AOI22_X1 U20353 ( .A1(n19787), .A2(n19142), .B1(n19317), .B2(n17358), .ZN(
        n17343) );
  INV_X1 U20354 ( .A(n17284), .ZN(n17345) );
  NOR2_X1 U20355 ( .A1(n17343), .A2(n17345), .ZN(n19058) );
  NAND4_X1 U20356 ( .A1(n19323), .A2(n17366), .A3(n17278), .A4(n19058), .ZN(
        n17279) );
  NAND2_X1 U20357 ( .A1(n17280), .A2(n17279), .ZN(n17302) );
  INV_X1 U20358 ( .A(n17281), .ZN(n17298) );
  NOR2_X1 U20359 ( .A1(n17406), .A2(n19161), .ZN(n19224) );
  NAND2_X1 U20360 ( .A1(n17342), .A2(n19224), .ZN(n19111) );
  INV_X1 U20361 ( .A(n19111), .ZN(n19160) );
  NAND2_X1 U20362 ( .A1(n17283), .A2(n19160), .ZN(n17357) );
  OAI21_X1 U20363 ( .B1(n17357), .B2(n17282), .A(n19226), .ZN(n17287) );
  NAND3_X1 U20364 ( .A1(n19138), .A2(n17283), .A3(n17366), .ZN(n17285) );
  NAND2_X1 U20365 ( .A1(n17284), .A2(n19142), .ZN(n19055) );
  INV_X1 U20366 ( .A(n19055), .ZN(n19075) );
  AOI21_X1 U20367 ( .B1(n19075), .B2(n17366), .A(n19314), .ZN(n17360) );
  AOI21_X1 U20368 ( .B1(n19337), .B2(n17285), .A(n17360), .ZN(n17286) );
  AND2_X1 U20369 ( .A1(n17287), .A2(n17286), .ZN(n17319) );
  NAND2_X1 U20370 ( .A1(n19291), .A2(n17288), .ZN(n17289) );
  OAI211_X1 U20371 ( .C1(n17319), .C2(n19336), .A(n17289), .B(n19329), .ZN(
        n17309) );
  AOI21_X1 U20372 ( .B1(n19291), .B2(n21756), .A(n17309), .ZN(n17296) );
  OR2_X1 U20373 ( .A1(n19791), .A2(n18624), .ZN(n19200) );
  AND2_X1 U20374 ( .A1(n19323), .A2(n19232), .ZN(n19193) );
  INV_X1 U20375 ( .A(n17290), .ZN(n17291) );
  AOI21_X1 U20376 ( .B1(n19193), .B2(n17292), .A(n17291), .ZN(n17295) );
  NAND2_X1 U20377 ( .A1(n19335), .A2(n17293), .ZN(n17294) );
  OAI211_X1 U20378 ( .C1(n17296), .C2(n17407), .A(n17295), .B(n17294), .ZN(
        n17297) );
  AOI21_X1 U20379 ( .B1(n17302), .B2(n17298), .A(n17297), .ZN(n17299) );
  OAI21_X1 U20380 ( .B1(n17300), .B2(n19249), .A(n17299), .ZN(P3_U2831) );
  INV_X1 U20381 ( .A(n19193), .ZN(n17305) );
  NOR2_X1 U20382 ( .A1(n17329), .A2(n17305), .ZN(n17301) );
  NOR2_X1 U20383 ( .A1(n17302), .A2(n17301), .ZN(n17325) );
  NOR3_X1 U20384 ( .A1(n17325), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n17303), .ZN(n17313) );
  OR2_X1 U20385 ( .A1(n17304), .A2(n19285), .ZN(n17308) );
  OR2_X1 U20386 ( .A1(n17306), .A2(n17305), .ZN(n17307) );
  AND2_X1 U20387 ( .A1(n17308), .A2(n17307), .ZN(n17321) );
  INV_X1 U20388 ( .A(n17309), .ZN(n17310) );
  AOI21_X1 U20389 ( .B1(n17321), .B2(n17310), .A(n21756), .ZN(n17311) );
  NOR3_X1 U20390 ( .A1(n17313), .A2(n17312), .A3(n17311), .ZN(n17314) );
  OAI21_X1 U20391 ( .B1(n17315), .B2(n19249), .A(n17314), .ZN(P3_U2832) );
  NOR2_X1 U20392 ( .A1(n19337), .A2(n19787), .ZN(n19096) );
  AND2_X1 U20393 ( .A1(n19323), .A2(n19096), .ZN(n19242) );
  AND2_X1 U20394 ( .A1(n19323), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17317) );
  OR2_X1 U20395 ( .A1(n19242), .A2(n17317), .ZN(n17318) );
  NAND2_X1 U20396 ( .A1(n17319), .A2(n17318), .ZN(n17328) );
  AOI22_X1 U20397 ( .A1(n17328), .A2(n19156), .B1(n19291), .B2(n17338), .ZN(
        n17320) );
  NAND2_X1 U20398 ( .A1(n17321), .A2(n17320), .ZN(n17323) );
  AOI21_X1 U20399 ( .B1(n17323), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n17322), .ZN(n17324) );
  NOR2_X1 U20400 ( .A1(n17326), .A2(n19321), .ZN(n17327) );
  NOR2_X1 U20401 ( .A1(n19791), .A2(n17330), .ZN(n17331) );
  AOI211_X1 U20402 ( .C1(n17335), .C2(n17334), .A(n19268), .B(n17338), .ZN(
        n17353) );
  NOR3_X1 U20403 ( .A1(n17337), .A2(n17336), .A3(n19249), .ZN(n17352) );
  NAND3_X1 U20404 ( .A1(n19331), .A2(n18910), .A3(n17338), .ZN(n17349) );
  NAND2_X1 U20405 ( .A1(n17339), .A2(n19786), .ZN(n17341) );
  OR2_X1 U20406 ( .A1(n17105), .A2(n19200), .ZN(n17340) );
  NAND2_X1 U20407 ( .A1(n17341), .A2(n17340), .ZN(n19144) );
  NAND3_X1 U20408 ( .A1(n19144), .A2(n19108), .A3(n17342), .ZN(n17344) );
  NOR2_X1 U20409 ( .A1(n19106), .A2(n17345), .ZN(n19083) );
  NAND3_X1 U20410 ( .A1(n19083), .A2(n19323), .A3(n17346), .ZN(n17347) );
  OAI211_X1 U20411 ( .C1(n17350), .C2(n17349), .A(n17348), .B(n17347), .ZN(
        n17351) );
  OAI21_X1 U20412 ( .B1(n19329), .B2(n17355), .A(n17354), .ZN(n17369) );
  INV_X1 U20413 ( .A(n17356), .ZN(n17365) );
  OAI21_X1 U20414 ( .B1(n19089), .B2(n19226), .A(n17357), .ZN(n19097) );
  NAND3_X1 U20415 ( .A1(n17358), .A2(n18818), .A3(n19097), .ZN(n19074) );
  NAND2_X1 U20416 ( .A1(n19237), .A2(n17359), .ZN(n19288) );
  OAI21_X1 U20417 ( .B1(n19060), .B2(n19074), .A(n19288), .ZN(n19057) );
  AOI21_X1 U20418 ( .B1(n17361), .B2(n19288), .A(n17360), .ZN(n17362) );
  OAI211_X1 U20419 ( .C1(n17363), .C2(n19200), .A(n19057), .B(n17362), .ZN(
        n17364) );
  AOI21_X1 U20420 ( .B1(n17365), .B2(n19786), .A(n17364), .ZN(n17372) );
  AOI21_X1 U20421 ( .B1(n19083), .B2(n17366), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17367) );
  AOI211_X1 U20422 ( .C1(n17372), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n17367), .B(n19336), .ZN(n17368) );
  AOI211_X1 U20423 ( .C1(n19255), .C2(n17370), .A(n17369), .B(n17368), .ZN(
        n17371) );
  INV_X1 U20424 ( .A(n17371), .ZN(P3_U2835) );
  INV_X1 U20425 ( .A(n17372), .ZN(n17377) );
  NAND3_X1 U20426 ( .A1(n19083), .A2(n19323), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19079) );
  OAI22_X1 U20427 ( .A1(n17374), .A2(n19336), .B1(n18773), .B2(n19079), .ZN(
        n17376) );
  OAI21_X1 U20428 ( .B1(n19329), .B2(n17374), .A(n17373), .ZN(n17375) );
  AOI21_X1 U20429 ( .B1(n17377), .B2(n17376), .A(n17375), .ZN(n17378) );
  OAI21_X1 U20430 ( .B1(n17379), .B2(n19249), .A(n17378), .ZN(P3_U2836) );
  AOI22_X1 U20431 ( .A1(n19787), .A2(n19313), .B1(n17380), .B2(n19317), .ZN(
        n17381) );
  INV_X1 U20432 ( .A(n17381), .ZN(n19308) );
  NAND2_X1 U20433 ( .A1(n19323), .A2(n19263), .ZN(n19271) );
  NOR3_X1 U20434 ( .A1(n19270), .A2(n19261), .A3(n19271), .ZN(n17390) );
  NOR2_X1 U20435 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n19336), .ZN(
        n17386) );
  AOI22_X1 U20436 ( .A1(n19787), .A2(n17384), .B1(n17383), .B2(n19288), .ZN(
        n17385) );
  NAND2_X1 U20437 ( .A1(n19226), .A2(n17406), .ZN(n19286) );
  AOI21_X1 U20438 ( .B1(n17385), .B2(n19286), .A(n19336), .ZN(n19267) );
  AOI211_X1 U20439 ( .C1(n19291), .C2(n19270), .A(n17386), .B(n19267), .ZN(
        n19260) );
  OAI21_X1 U20440 ( .B1(n19183), .B2(n19260), .A(n19329), .ZN(n17388) );
  NOR2_X1 U20441 ( .A1(n19156), .A2(n19870), .ZN(n17387) );
  AOI221_X1 U20442 ( .B1(n17390), .B2(n17389), .C1(n17388), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17387), .ZN(n17391) );
  OAI21_X1 U20443 ( .B1(n17392), .B2(n19285), .A(n17391), .ZN(n17393) );
  AOI21_X1 U20444 ( .B1(n17394), .B2(n19193), .A(n17393), .ZN(n17395) );
  OAI21_X1 U20445 ( .B1(n17396), .B2(n19249), .A(n17395), .ZN(P3_U2854) );
  NAND2_X1 U20446 ( .A1(n19821), .A2(n17398), .ZN(n17402) );
  INV_X1 U20447 ( .A(n17439), .ZN(n17434) );
  MUX2_X1 U20448 ( .A(n19337), .B(n10721), .S(n17398), .Z(n19805) );
  NAND2_X1 U20449 ( .A1(n19805), .A2(n17437), .ZN(n17399) );
  OAI211_X1 U20450 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18649), .A(
        n17399), .B(n17434), .ZN(n17400) );
  OAI21_X1 U20451 ( .B1(n17434), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n17400), .ZN(n17401) );
  OAI21_X1 U20452 ( .B1(n17439), .B2(n17402), .A(n17401), .ZN(P3_U3290) );
  NOR2_X1 U20453 ( .A1(n17403), .A2(n17415), .ZN(n17405) );
  AOI22_X1 U20454 ( .A1(n17405), .A2(n10721), .B1(n17404), .B2(n17414), .ZN(
        n19801) );
  INV_X1 U20455 ( .A(n19801), .ZN(n17412) );
  INV_X1 U20456 ( .A(n19821), .ZN(n17435) );
  INV_X1 U20457 ( .A(n17405), .ZN(n18104) );
  NOR2_X1 U20458 ( .A1(n18649), .A2(n17406), .ZN(n17432) );
  AOI22_X1 U20459 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n17408), .B2(n17407), .ZN(
        n17431) );
  INV_X1 U20460 ( .A(n17431), .ZN(n17409) );
  NAND2_X1 U20461 ( .A1(n17432), .A2(n17409), .ZN(n17410) );
  OAI211_X1 U20462 ( .C1(n17435), .C2(n18104), .A(n17434), .B(n17410), .ZN(
        n17411) );
  AOI21_X1 U20463 ( .B1(n17412), .B2(n17437), .A(n17411), .ZN(n17413) );
  AOI21_X1 U20464 ( .B1(n17439), .B2(n17414), .A(n17413), .ZN(P3_U3289) );
  NAND2_X1 U20465 ( .A1(n19226), .A2(n17415), .ZN(n17423) );
  NOR2_X1 U20466 ( .A1(n17425), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n17417) );
  OAI21_X1 U20467 ( .B1(n17418), .B2(n17417), .A(n17416), .ZN(n17421) );
  INV_X1 U20468 ( .A(n17419), .ZN(n17724) );
  NAND2_X1 U20469 ( .A1(n17724), .A2(n17420), .ZN(n17424) );
  AND2_X1 U20470 ( .A1(n17421), .A2(n17424), .ZN(n17422) );
  MUX2_X1 U20471 ( .A(n17423), .B(n17422), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n17430) );
  OAI21_X1 U20472 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n17425), .A(
        n17424), .ZN(n17428) );
  NAND2_X1 U20473 ( .A1(n17427), .A2(n17426), .ZN(n18088) );
  AOI22_X1 U20474 ( .A1(n17428), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n19787), .B2(n18088), .ZN(n17429) );
  NAND2_X1 U20475 ( .A1(n17430), .A2(n17429), .ZN(n19799) );
  NAND2_X1 U20476 ( .A1(n17432), .A2(n17431), .ZN(n17433) );
  OAI211_X1 U20477 ( .C1(n18088), .C2(n17435), .A(n17434), .B(n17433), .ZN(
        n17436) );
  AOI21_X1 U20478 ( .B1(n19799), .B2(n17437), .A(n17436), .ZN(n17438) );
  AOI21_X1 U20479 ( .B1(n17439), .B2(n10426), .A(n17438), .ZN(P3_U3288) );
  OAI22_X1 U20480 ( .A1(n14490), .A2(n18209), .B1(n18443), .B2(n17440), .ZN(
        n17441) );
  AOI21_X1 U20481 ( .B1(n18450), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17441), .ZN(n17445) );
  AOI22_X1 U20482 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20483 ( .A1(n14578), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17443) );
  NAND2_X1 U20484 ( .A1(n9717), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n17442) );
  NAND4_X1 U20485 ( .A1(n17445), .A2(n17444), .A3(n17443), .A4(n17442), .ZN(
        n17454) );
  AOI22_X1 U20486 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17446), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U20487 ( .B1(n18330), .B2(n17448), .A(n17447), .ZN(n17449) );
  AOI21_X1 U20488 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n17449), .ZN(n17452) );
  AOI22_X1 U20489 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13684), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U20490 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17450) );
  NAND3_X1 U20491 ( .A1(n17452), .A2(n17451), .A3(n17450), .ZN(n17453) );
  NOR2_X1 U20492 ( .A1(n17454), .A2(n17453), .ZN(n18599) );
  NOR2_X1 U20493 ( .A1(n18498), .A2(n9761), .ZN(n18376) );
  INV_X1 U20494 ( .A(n18495), .ZN(n18497) );
  INV_X1 U20495 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17949) );
  NAND2_X1 U20496 ( .A1(n18497), .A2(n17949), .ZN(n18358) );
  NOR2_X1 U20497 ( .A1(n17455), .A2(n18358), .ZN(n17456) );
  AOI22_X1 U20498 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n18376), .B1(n17457), 
        .B2(n17456), .ZN(n17458) );
  OAI21_X1 U20499 ( .B1(n18599), .B2(n18484), .A(n17458), .ZN(P3_U2690) );
  OR2_X1 U20500 ( .A1(n19937), .A2(n19008), .ZN(n17462) );
  NAND2_X1 U20501 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19350) );
  NAND2_X1 U20502 ( .A1(n17459), .A2(n18330), .ZN(n19343) );
  INV_X1 U20503 ( .A(n19921), .ZN(n17460) );
  OAI21_X1 U20504 ( .B1(n19343), .B2(P3_FLUSH_REG_SCAN_IN), .A(n17460), .ZN(
        n17461) );
  AND2_X1 U20505 ( .A1(n19635), .A2(n17461), .ZN(n17466) );
  AOI21_X1 U20506 ( .B1(n17462), .B2(n19350), .A(n17466), .ZN(n17467) );
  INV_X1 U20507 ( .A(n17467), .ZN(n17464) );
  NOR2_X1 U20508 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19923), .ZN(
        n19428) );
  NOR4_X1 U20509 ( .A1(n19428), .A2(n19407), .A3(n17466), .A4(n19806), .ZN(
        n17463) );
  AOI21_X1 U20510 ( .B1(n19806), .B2(n17464), .A(n17463), .ZN(P3_U2864) );
  NAND2_X1 U20511 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19497) );
  OAI21_X1 U20512 ( .B1(n19008), .B2(n19937), .A(n19923), .ZN(n17465) );
  AOI211_X1 U20513 ( .C1(n19497), .C2(n17465), .A(n19428), .B(n17466), .ZN(
        n19347) );
  INV_X1 U20514 ( .A(n17466), .ZN(n19348) );
  AOI22_X1 U20515 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n17467), .B1(
        n19407), .B2(n19348), .ZN(n19346) );
  AOI22_X1 U20516 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19347), .B1(
        n19346), .B2(n13797), .ZN(P3_U2865) );
  NAND2_X1 U20517 ( .A1(n17468), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n17469) );
  NAND2_X1 U20518 ( .A1(n17469), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n17470) );
  NOR2_X1 U20519 ( .A1(n17471), .A2(n17470), .ZN(n17472) );
  INV_X1 U20520 ( .A(n17472), .ZN(n17476) );
  OAI22_X1 U20521 ( .A1(n17474), .A2(n17473), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n17472), .ZN(n17475) );
  OAI21_X1 U20522 ( .B1(n17476), .B2(n21409), .A(n17475), .ZN(n17479) );
  INV_X1 U20523 ( .A(n17477), .ZN(n17478) );
  AOI222_X1 U20524 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n17479), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17478), .C1(n17479), 
        .C2(n17478), .ZN(n17481) );
  AOI222_X1 U20525 ( .A1(n17481), .A2(n21234), .B1(n17481), .B2(n17480), .C1(
        n21234), .C2(n17480), .ZN(n17488) );
  NOR2_X1 U20526 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(P1_MORE_REG_SCAN_IN), .ZN(
        n17483) );
  OAI22_X1 U20527 ( .A1(n17484), .A2(n17483), .B1(n10868), .B2(n17482), .ZN(
        n17485) );
  INV_X1 U20528 ( .A(n17485), .ZN(n17487) );
  OAI211_X1 U20529 ( .C1(n17488), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n17487), .B(n17486), .ZN(n17489) );
  NOR3_X1 U20530 ( .A1(n17491), .A2(n17490), .A3(n17489), .ZN(n17501) );
  INV_X1 U20531 ( .A(n17501), .ZN(n17498) );
  NOR2_X1 U20532 ( .A1(n17492), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21575) );
  NAND2_X1 U20533 ( .A1(n17493), .A2(n21575), .ZN(n17496) );
  OAI21_X1 U20534 ( .B1(n17494), .B2(n21574), .A(n21475), .ZN(n17495) );
  OAI21_X1 U20535 ( .B1(n17497), .B2(n17496), .A(n17495), .ZN(n17578) );
  AOI21_X1 U20536 ( .B1(n21478), .B2(n21578), .A(n17573), .ZN(n17500) );
  OAI211_X1 U20537 ( .C1(n17501), .C2(n21475), .A(n17500), .B(n17499), .ZN(
        n17502) );
  NOR2_X1 U20538 ( .A1(n17580), .A2(n17502), .ZN(n17506) );
  NAND2_X1 U20539 ( .A1(n17573), .A2(n17503), .ZN(n17504) );
  NAND2_X1 U20540 ( .A1(n20825), .A2(n17504), .ZN(n17505) );
  OAI22_X1 U20541 ( .A1(n17506), .A2(n20825), .B1(n17580), .B2(n17505), .ZN(
        P1_U3161) );
  AND2_X1 U20542 ( .A1(n20966), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U20543 ( .A(n17507), .ZN(n17508) );
  OAI21_X1 U20544 ( .B1(n17509), .B2(P2_FLUSH_REG_SCAN_IN), .A(n17508), .ZN(
        n17510) );
  AND2_X1 U20545 ( .A1(n20494), .A2(n17510), .ZN(n20784) );
  AND2_X1 U20546 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20784), .ZN(
        P2_U3047) );
  AOI22_X1 U20547 ( .A1(n17517), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n17539), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17516) );
  OAI21_X1 U20548 ( .B1(n17513), .B2(n17512), .A(n17511), .ZN(n17514) );
  INV_X1 U20549 ( .A(n17514), .ZN(n17534) );
  AOI22_X1 U20550 ( .A1(n17534), .A2(n17531), .B1(n20868), .B2(n17530), .ZN(
        n17515) );
  OAI211_X1 U20551 ( .C1(n17524), .C2(n20863), .A(n17516), .B(n17515), .ZN(
        P1_U2992) );
  AOI22_X1 U20552 ( .A1(n17517), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n17539), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17523) );
  NAND2_X1 U20553 ( .A1(n17520), .A2(n17519), .ZN(n17521) );
  XNOR2_X1 U20554 ( .A(n17518), .B(n17521), .ZN(n17541) );
  AOI22_X1 U20555 ( .A1(n17530), .A2(n20878), .B1(n17541), .B2(n17531), .ZN(
        n17522) );
  OAI211_X1 U20556 ( .C1(n17524), .C2(n20873), .A(n17523), .B(n17522), .ZN(
        P1_U2993) );
  XOR2_X1 U20557 ( .A(n17526), .B(n17525), .Z(n17554) );
  INV_X1 U20558 ( .A(n20891), .ZN(n17529) );
  AOI222_X1 U20559 ( .A1(n17554), .A2(n17531), .B1(n17530), .B2(n20933), .C1(
        n17529), .C2(n17528), .ZN(n17532) );
  NAND2_X1 U20560 ( .A1(n17539), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n17553) );
  OAI211_X1 U20561 ( .C1(n21775), .C2(n17533), .A(n17532), .B(n17553), .ZN(
        P1_U2994) );
  AOI222_X1 U20562 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n17539), .B1(n20998), 
        .B2(n20866), .C1(n20999), .C2(n17534), .ZN(n17535) );
  OAI221_X1 U20563 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17538), .C1(
        n17537), .C2(n17536), .A(n17535), .ZN(P1_U3024) );
  AOI22_X1 U20564 ( .A1(n17539), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20998), 
        .B2(n20871), .ZN(n17543) );
  AOI22_X1 U20565 ( .A1(n17541), .A2(n20999), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17540), .ZN(n17542) );
  OAI211_X1 U20566 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n17544), .A(
        n17543), .B(n17542), .ZN(P1_U3025) );
  NOR2_X1 U20567 ( .A1(n17546), .A2(n17545), .ZN(n17549) );
  NAND2_X1 U20568 ( .A1(n17547), .A2(n17556), .ZN(n17548) );
  AND2_X1 U20569 ( .A1(n17549), .A2(n17548), .ZN(n17564) );
  NAND2_X1 U20570 ( .A1(n14210), .A2(n17550), .ZN(n17551) );
  AND2_X1 U20571 ( .A1(n17552), .A2(n17551), .ZN(n20930) );
  INV_X1 U20572 ( .A(n17553), .ZN(n17562) );
  INV_X1 U20573 ( .A(n17554), .ZN(n17560) );
  INV_X1 U20574 ( .A(n17555), .ZN(n17558) );
  OR2_X1 U20575 ( .A1(n17556), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17557) );
  OAI22_X1 U20576 ( .A1(n17560), .A2(n17559), .B1(n17558), .B2(n17557), .ZN(
        n17561) );
  AOI211_X1 U20577 ( .C1(n20998), .C2(n20930), .A(n17562), .B(n17561), .ZN(
        n17563) );
  OAI21_X1 U20578 ( .B1(n17564), .B2(n21873), .A(n17563), .ZN(P1_U3026) );
  NAND4_X1 U20579 ( .A1(n20892), .A2(n17567), .A3(n17566), .A4(n17565), .ZN(
        n17568) );
  OAI21_X1 U20580 ( .B1(n17570), .B2(n17569), .A(n17568), .ZN(P1_U3468) );
  NAND4_X1 U20581 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n21578), .A4(n21574), .ZN(n17571) );
  NAND2_X1 U20582 ( .A1(n17572), .A2(n17571), .ZN(n21474) );
  NAND2_X1 U20583 ( .A1(n21478), .A2(n21578), .ZN(n17576) );
  OAI21_X1 U20584 ( .B1(n17580), .B2(n20825), .A(n13446), .ZN(n17575) );
  INV_X1 U20585 ( .A(n17573), .ZN(n17574) );
  OAI211_X1 U20586 ( .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n17576), .A(n17575), 
        .B(n17574), .ZN(n17577) );
  AOI221_X1 U20587 ( .B1(n17579), .B2(n17578), .C1(n21474), .C2(n17578), .A(
        n17577), .ZN(P1_U3162) );
  NOR2_X1 U20588 ( .A1(n17580), .A2(n20825), .ZN(n17582) );
  OAI21_X1 U20589 ( .B1(n17582), .B2(n21706), .A(n17581), .ZN(P1_U3466) );
  INV_X1 U20590 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17598) );
  INV_X1 U20591 ( .A(n17583), .ZN(n17584) );
  AOI21_X1 U20592 ( .B1(n17586), .B2(n17585), .A(n17584), .ZN(n17597) );
  NAND2_X1 U20593 ( .A1(n17588), .A2(n17587), .ZN(n17592) );
  OR2_X1 U20594 ( .A1(n17590), .A2(n17589), .ZN(n17591) );
  OAI211_X1 U20595 ( .C1(n17594), .C2(n17593), .A(n17592), .B(n17591), .ZN(
        n17595) );
  INV_X1 U20596 ( .A(n17595), .ZN(n17596) );
  OAI211_X1 U20597 ( .C1(n17599), .C2(n17598), .A(n17597), .B(n17596), .ZN(
        P2_U3009) );
  INV_X1 U20598 ( .A(n17600), .ZN(n17601) );
  AOI22_X1 U20599 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17603), .B1(
        n17602), .B2(n17601), .ZN(n17614) );
  NAND2_X1 U20600 ( .A1(n17604), .A2(n12527), .ZN(n17612) );
  NAND2_X1 U20601 ( .A1(n17606), .A2(n17605), .ZN(n17610) );
  NAND2_X1 U20602 ( .A1(n17608), .A2(n17607), .ZN(n17609) );
  AND4_X1 U20603 ( .A1(n17612), .A2(n17611), .A3(n17610), .A4(n17609), .ZN(
        n17613) );
  OAI211_X1 U20604 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n17615), .A(
        n17614), .B(n17613), .ZN(P2_U3046) );
  NOR3_X1 U20605 ( .A1(P3_D_C_N_REG_SCAN_IN), .A2(P3_W_R_N_REG_SCAN_IN), .A3(
        P3_BE_N_REG_0__SCAN_IN), .ZN(n17617) );
  NOR4_X1 U20606 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_2__SCAN_IN), 
        .A3(P3_BE_N_REG_3__SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17616) );
  NAND4_X1 U20607 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17617), .A3(n17616), .A4(
        U215), .ZN(U213) );
  AOI222_X1 U20608 ( .A1(n17658), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(n17656), 
        .B2(BUF1_REG_31__SCAN_IN), .C1(n17655), .C2(P1_DATAO_REG_31__SCAN_IN), 
        .ZN(n17619) );
  INV_X1 U20609 ( .A(n17619), .ZN(U216) );
  AOI22_X1 U20610 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n17658), .ZN(n17620) );
  OAI21_X1 U20611 ( .B1(n14710), .B2(n17660), .A(n17620), .ZN(U217) );
  AOI22_X1 U20612 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17658), .ZN(n17621) );
  OAI21_X1 U20613 ( .B1(n16095), .B2(n17660), .A(n17621), .ZN(U218) );
  AOI22_X1 U20614 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17658), .ZN(n17622) );
  OAI21_X1 U20615 ( .B1(n16103), .B2(n17660), .A(n17622), .ZN(U219) );
  AOI22_X1 U20616 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17658), .ZN(n17623) );
  OAI21_X1 U20617 ( .B1(n16110), .B2(n17660), .A(n17623), .ZN(U220) );
  AOI22_X1 U20618 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n17658), .ZN(n17624) );
  OAI21_X1 U20619 ( .B1(n16118), .B2(n17660), .A(n17624), .ZN(U221) );
  INV_X1 U20620 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n17626) );
  AOI22_X1 U20621 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17658), .ZN(n17625) );
  OAI21_X1 U20622 ( .B1(n17626), .B2(n17660), .A(n17625), .ZN(U222) );
  AOI22_X1 U20623 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n17658), .ZN(n17627) );
  OAI21_X1 U20624 ( .B1(n16133), .B2(n17660), .A(n17627), .ZN(U223) );
  INV_X1 U20625 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n21774) );
  AOI22_X1 U20626 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n17655), .ZN(n17628) );
  OAI21_X1 U20627 ( .B1(n21774), .B2(U212), .A(n17628), .ZN(U224) );
  INV_X1 U20628 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n21853) );
  AOI22_X1 U20629 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n17655), .ZN(n17629) );
  OAI21_X1 U20630 ( .B1(n21853), .B2(U212), .A(n17629), .ZN(U225) );
  AOI22_X1 U20631 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17658), .ZN(n17630) );
  OAI21_X1 U20632 ( .B1(n16155), .B2(n17660), .A(n17630), .ZN(U226) );
  AOI22_X1 U20633 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17658), .ZN(n17631) );
  OAI21_X1 U20634 ( .B1(n17632), .B2(n17660), .A(n17631), .ZN(U227) );
  INV_X1 U20635 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n17634) );
  AOI22_X1 U20636 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17658), .ZN(n17633) );
  OAI21_X1 U20637 ( .B1(n17634), .B2(n17660), .A(n17633), .ZN(U228) );
  AOI22_X1 U20638 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17658), .ZN(n17635) );
  OAI21_X1 U20639 ( .B1(n16177), .B2(n17660), .A(n17635), .ZN(U229) );
  AOI22_X1 U20640 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17658), .ZN(n17636) );
  OAI21_X1 U20641 ( .B1(n16181), .B2(n17660), .A(n17636), .ZN(U230) );
  INV_X1 U20642 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17638) );
  AOI22_X1 U20643 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17658), .ZN(n17637) );
  OAI21_X1 U20644 ( .B1(n17638), .B2(n17660), .A(n17637), .ZN(U231) );
  AOI22_X1 U20645 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17658), .ZN(n17639) );
  OAI21_X1 U20646 ( .B1(n13448), .B2(n17660), .A(n17639), .ZN(U232) );
  INV_X1 U20647 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U20648 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n17655), .ZN(n17640) );
  OAI21_X1 U20649 ( .B1(n17678), .B2(U212), .A(n17640), .ZN(U233) );
  INV_X1 U20650 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n17676) );
  AOI22_X1 U20651 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n17655), .ZN(n17641) );
  OAI21_X1 U20652 ( .B1(n17676), .B2(U212), .A(n17641), .ZN(U234) );
  INV_X1 U20653 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17674) );
  INV_X1 U20654 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n21851) );
  OAI222_X1 U20655 ( .A1(U212), .A2(n17674), .B1(n17660), .B2(n21784), .C1(
        U214), .C2(n21851), .ZN(U235) );
  INV_X1 U20656 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U20657 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n17655), .ZN(n17642) );
  OAI21_X1 U20658 ( .B1(n17673), .B2(U212), .A(n17642), .ZN(U236) );
  AOI22_X1 U20659 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17658), .ZN(n17643) );
  OAI21_X1 U20660 ( .B1(n17644), .B2(n17660), .A(n17643), .ZN(U237) );
  INV_X1 U20661 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17671) );
  AOI22_X1 U20662 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n17655), .ZN(n17645) );
  OAI21_X1 U20663 ( .B1(n17671), .B2(U212), .A(n17645), .ZN(U238) );
  AOI22_X1 U20664 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17658), .ZN(n17646) );
  OAI21_X1 U20665 ( .B1(n17647), .B2(n17660), .A(n17646), .ZN(U239) );
  INV_X1 U20666 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17668) );
  AOI22_X1 U20667 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n17655), .ZN(n17648) );
  OAI21_X1 U20668 ( .B1(n17668), .B2(U212), .A(n17648), .ZN(U240) );
  AOI22_X1 U20669 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17658), .ZN(n17649) );
  OAI21_X1 U20670 ( .B1(n13481), .B2(n17660), .A(n17649), .ZN(U241) );
  INV_X1 U20671 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n21807) );
  AOI22_X1 U20672 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n17655), .ZN(n17650) );
  OAI21_X1 U20673 ( .B1(n21807), .B2(U212), .A(n17650), .ZN(U242) );
  AOI22_X1 U20674 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17658), .ZN(n17651) );
  OAI21_X1 U20675 ( .B1(n13472), .B2(n17660), .A(n17651), .ZN(U243) );
  INV_X1 U20676 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U20677 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n17655), .ZN(n17652) );
  OAI21_X1 U20678 ( .B1(n17665), .B2(U212), .A(n17652), .ZN(U244) );
  AOI22_X1 U20679 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17658), .ZN(n17653) );
  OAI21_X1 U20680 ( .B1(n17654), .B2(n17660), .A(n17653), .ZN(U245) );
  INV_X1 U20681 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n17663) );
  AOI22_X1 U20682 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n17656), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n17655), .ZN(n17657) );
  OAI21_X1 U20683 ( .B1(n17663), .B2(U212), .A(n17657), .ZN(U246) );
  AOI22_X1 U20684 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17655), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17658), .ZN(n17659) );
  OAI21_X1 U20685 ( .B1(n17661), .B2(n17660), .A(n17659), .ZN(U247) );
  INV_X1 U20686 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17662) );
  INV_X1 U20687 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n19349) );
  AOI22_X1 U20688 ( .A1(n17693), .A2(n17662), .B1(n19349), .B2(U215), .ZN(U251) );
  INV_X1 U20689 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n19358) );
  AOI22_X1 U20690 ( .A1(n17693), .A2(n17663), .B1(n19358), .B2(U215), .ZN(U252) );
  INV_X1 U20691 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U20692 ( .A1(n17693), .A2(n17664), .B1(n19361), .B2(U215), .ZN(U253) );
  INV_X1 U20693 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19364) );
  AOI22_X1 U20694 ( .A1(n17693), .A2(n17665), .B1(n19364), .B2(U215), .ZN(U254) );
  INV_X1 U20695 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17666) );
  INV_X1 U20696 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19368) );
  AOI22_X1 U20697 ( .A1(n17693), .A2(n17666), .B1(n19368), .B2(U215), .ZN(U255) );
  INV_X1 U20698 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n19372) );
  AOI22_X1 U20699 ( .A1(n17694), .A2(n21807), .B1(n19372), .B2(U215), .ZN(U256) );
  INV_X1 U20700 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17667) );
  INV_X1 U20701 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19376) );
  AOI22_X1 U20702 ( .A1(n17693), .A2(n17667), .B1(n19376), .B2(U215), .ZN(U257) );
  INV_X1 U20703 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n19380) );
  AOI22_X1 U20704 ( .A1(n17694), .A2(n17668), .B1(n19380), .B2(U215), .ZN(U258) );
  OAI22_X1 U20705 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17693), .ZN(n17669) );
  INV_X1 U20706 ( .A(n17669), .ZN(U259) );
  INV_X1 U20707 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17670) );
  AOI22_X1 U20708 ( .A1(n17694), .A2(n17671), .B1(n17670), .B2(U215), .ZN(U260) );
  INV_X1 U20709 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17672) );
  INV_X1 U20710 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n18745) );
  AOI22_X1 U20711 ( .A1(n17693), .A2(n17672), .B1(n18745), .B2(U215), .ZN(U261) );
  INV_X1 U20712 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n18747) );
  AOI22_X1 U20713 ( .A1(n17693), .A2(n17673), .B1(n18747), .B2(U215), .ZN(U262) );
  INV_X1 U20714 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n18751) );
  AOI22_X1 U20715 ( .A1(n17694), .A2(n17674), .B1(n18751), .B2(U215), .ZN(U263) );
  INV_X1 U20716 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17675) );
  AOI22_X1 U20717 ( .A1(n17693), .A2(n17676), .B1(n17675), .B2(U215), .ZN(U264) );
  INV_X1 U20718 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U20719 ( .A1(n17694), .A2(n17678), .B1(n17677), .B2(U215), .ZN(U265) );
  OAI22_X1 U20720 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n17693), .ZN(n17679) );
  INV_X1 U20721 ( .A(n17679), .ZN(U266) );
  OAI22_X1 U20722 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17693), .ZN(n17680) );
  INV_X1 U20723 ( .A(n17680), .ZN(U267) );
  OAI22_X1 U20724 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17693), .ZN(n17681) );
  INV_X1 U20725 ( .A(n17681), .ZN(U268) );
  OAI22_X1 U20726 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17693), .ZN(n17682) );
  INV_X1 U20727 ( .A(n17682), .ZN(U269) );
  OAI22_X1 U20728 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17693), .ZN(n17683) );
  INV_X1 U20729 ( .A(n17683), .ZN(U270) );
  OAI22_X1 U20730 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17694), .ZN(n17684) );
  INV_X1 U20731 ( .A(n17684), .ZN(U271) );
  OAI22_X1 U20732 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17694), .ZN(n17685) );
  INV_X1 U20733 ( .A(n17685), .ZN(U272) );
  INV_X1 U20734 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n21654) );
  AOI22_X1 U20735 ( .A1(n17694), .A2(n21853), .B1(n21654), .B2(U215), .ZN(U273) );
  OAI22_X1 U20736 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17694), .ZN(n17686) );
  INV_X1 U20737 ( .A(n17686), .ZN(U274) );
  INV_X1 U20738 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n17687) );
  INV_X1 U20739 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18543) );
  AOI22_X1 U20740 ( .A1(n17693), .A2(n17687), .B1(n18543), .B2(U215), .ZN(U275) );
  OAI22_X1 U20741 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17693), .ZN(n17688) );
  INV_X1 U20742 ( .A(n17688), .ZN(U276) );
  INV_X1 U20743 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n17689) );
  INV_X1 U20744 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18531) );
  AOI22_X1 U20745 ( .A1(n17693), .A2(n17689), .B1(n18531), .B2(U215), .ZN(U277) );
  OAI22_X1 U20746 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17693), .ZN(n17690) );
  INV_X1 U20747 ( .A(n17690), .ZN(U278) );
  INV_X1 U20748 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17691) );
  INV_X1 U20749 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n21768) );
  AOI22_X1 U20750 ( .A1(n17693), .A2(n17691), .B1(n21768), .B2(U215), .ZN(U279) );
  OAI22_X1 U20751 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17693), .ZN(n17692) );
  INV_X1 U20752 ( .A(n17692), .ZN(U280) );
  INV_X1 U20753 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n17695) );
  AOI22_X1 U20754 ( .A1(n17693), .A2(n17695), .B1(n14713), .B2(U215), .ZN(U281) );
  INV_X1 U20755 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n21787) );
  INV_X1 U20756 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n21701) );
  AOI22_X1 U20757 ( .A1(n17694), .A2(n21787), .B1(n21701), .B2(U215), .ZN(U282) );
  INV_X1 U20758 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n17696) );
  INV_X1 U20759 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n21866) );
  OAI222_X1 U20760 ( .A1(P1_DATAO_REG_31__SCAN_IN), .A2(n17696), .B1(
        P2_DATAO_REG_31__SCAN_IN), .B2(n17695), .C1(P3_DATAO_REG_31__SCAN_IN), 
        .C2(n21866), .ZN(n17698) );
  INV_X2 U20761 ( .A(n17699), .ZN(n17697) );
  INV_X1 U20762 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19874) );
  INV_X1 U20763 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20706) );
  AOI22_X1 U20764 ( .A1(n17697), .A2(n19874), .B1(n20706), .B2(n17699), .ZN(
        U347) );
  INV_X1 U20765 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19872) );
  INV_X1 U20766 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20704) );
  AOI22_X1 U20767 ( .A1(n17697), .A2(n19872), .B1(n20704), .B2(n17699), .ZN(
        U348) );
  INV_X1 U20768 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19871) );
  INV_X1 U20769 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20703) );
  AOI22_X1 U20770 ( .A1(n17697), .A2(n19871), .B1(n20703), .B2(n17699), .ZN(
        U349) );
  INV_X1 U20771 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19869) );
  INV_X1 U20772 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20701) );
  AOI22_X1 U20773 ( .A1(n17697), .A2(n19869), .B1(n20701), .B2(n17699), .ZN(
        U350) );
  INV_X1 U20774 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19867) );
  INV_X1 U20775 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20699) );
  AOI22_X1 U20776 ( .A1(n17697), .A2(n19867), .B1(n20699), .B2(n17699), .ZN(
        U351) );
  INV_X1 U20777 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19865) );
  INV_X1 U20778 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n21790) );
  AOI22_X1 U20779 ( .A1(n17697), .A2(n19865), .B1(n21790), .B2(n17699), .ZN(
        U352) );
  INV_X1 U20780 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19863) );
  INV_X1 U20781 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20697) );
  AOI22_X1 U20782 ( .A1(n17697), .A2(n19863), .B1(n20697), .B2(n17699), .ZN(
        U353) );
  INV_X1 U20783 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U20784 ( .A1(n17697), .A2(n19861), .B1(n20696), .B2(n17699), .ZN(
        U354) );
  INV_X1 U20785 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19907) );
  INV_X1 U20786 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20735) );
  AOI22_X1 U20787 ( .A1(n17697), .A2(n19907), .B1(n20735), .B2(n17698), .ZN(
        U355) );
  INV_X1 U20788 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19905) );
  INV_X1 U20789 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20732) );
  AOI22_X1 U20790 ( .A1(n17697), .A2(n19905), .B1(n20732), .B2(n17699), .ZN(
        U356) );
  INV_X1 U20791 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n21588) );
  INV_X1 U20792 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20730) );
  AOI22_X1 U20793 ( .A1(n17697), .A2(n21588), .B1(n20730), .B2(n17699), .ZN(
        U357) );
  INV_X1 U20794 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19903) );
  INV_X1 U20795 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20728) );
  AOI22_X1 U20796 ( .A1(n17697), .A2(n19903), .B1(n20728), .B2(n17698), .ZN(
        U358) );
  INV_X1 U20797 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19901) );
  INV_X1 U20798 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20727) );
  AOI22_X1 U20799 ( .A1(n17697), .A2(n19901), .B1(n20727), .B2(n17698), .ZN(
        U359) );
  INV_X1 U20800 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19899) );
  INV_X1 U20801 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n21817) );
  AOI22_X1 U20802 ( .A1(n17697), .A2(n19899), .B1(n21817), .B2(n17698), .ZN(
        U360) );
  INV_X1 U20803 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19897) );
  INV_X1 U20804 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20724) );
  AOI22_X1 U20805 ( .A1(n17697), .A2(n19897), .B1(n20724), .B2(n17698), .ZN(
        U361) );
  INV_X1 U20806 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19894) );
  INV_X1 U20807 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20723) );
  AOI22_X1 U20808 ( .A1(n17697), .A2(n19894), .B1(n20723), .B2(n17698), .ZN(
        U362) );
  INV_X1 U20809 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19893) );
  INV_X1 U20810 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20722) );
  AOI22_X1 U20811 ( .A1(n17697), .A2(n19893), .B1(n20722), .B2(n17698), .ZN(
        U363) );
  INV_X1 U20812 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19891) );
  INV_X1 U20813 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20721) );
  AOI22_X1 U20814 ( .A1(n17697), .A2(n19891), .B1(n20721), .B2(n17699), .ZN(
        U364) );
  INV_X1 U20815 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19859) );
  INV_X1 U20816 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20695) );
  AOI22_X1 U20817 ( .A1(n17697), .A2(n19859), .B1(n20695), .B2(n17699), .ZN(
        U365) );
  INV_X1 U20818 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n21850) );
  INV_X1 U20819 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20720) );
  AOI22_X1 U20820 ( .A1(n17697), .A2(n21850), .B1(n20720), .B2(n17699), .ZN(
        U366) );
  INV_X1 U20821 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19888) );
  INV_X1 U20822 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U20823 ( .A1(n17697), .A2(n19888), .B1(n20719), .B2(n17699), .ZN(
        U367) );
  INV_X1 U20824 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19886) );
  INV_X1 U20825 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20717) );
  AOI22_X1 U20826 ( .A1(n17697), .A2(n19886), .B1(n20717), .B2(n17699), .ZN(
        U368) );
  INV_X1 U20827 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n21670) );
  INV_X1 U20828 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20716) );
  AOI22_X1 U20829 ( .A1(n17697), .A2(n21670), .B1(n20716), .B2(n17699), .ZN(
        U369) );
  INV_X1 U20830 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19884) );
  INV_X1 U20831 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20714) );
  AOI22_X1 U20832 ( .A1(n17697), .A2(n19884), .B1(n20714), .B2(n17699), .ZN(
        U370) );
  INV_X1 U20833 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19882) );
  INV_X1 U20834 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20713) );
  AOI22_X1 U20835 ( .A1(n17697), .A2(n19882), .B1(n20713), .B2(n17699), .ZN(
        U371) );
  INV_X1 U20836 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19880) );
  INV_X1 U20837 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U20838 ( .A1(n17697), .A2(n19880), .B1(n20711), .B2(n17699), .ZN(
        U372) );
  INV_X1 U20839 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19879) );
  INV_X1 U20840 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20710) );
  AOI22_X1 U20841 ( .A1(n17697), .A2(n19879), .B1(n20710), .B2(n17699), .ZN(
        U373) );
  INV_X1 U20842 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19877) );
  INV_X1 U20843 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20709) );
  AOI22_X1 U20844 ( .A1(n17697), .A2(n19877), .B1(n20709), .B2(n17699), .ZN(
        U374) );
  INV_X1 U20845 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19876) );
  INV_X1 U20846 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20707) );
  AOI22_X1 U20847 ( .A1(n17697), .A2(n19876), .B1(n20707), .B2(n17698), .ZN(
        U375) );
  INV_X1 U20848 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19857) );
  INV_X1 U20849 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20693) );
  AOI22_X1 U20850 ( .A1(n17697), .A2(n19857), .B1(n20693), .B2(n17699), .ZN(
        U376) );
  INV_X1 U20851 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17701) );
  INV_X1 U20852 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19856) );
  NAND3_X1 U20853 ( .A1(n19856), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n17700) );
  OR2_X1 U20854 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n19845) );
  NAND2_X1 U20855 ( .A1(n17700), .A2(n19845), .ZN(n19920) );
  OAI21_X1 U20856 ( .B1(n19853), .B2(n17701), .A(n19917), .ZN(P3_U2633) );
  INV_X1 U20857 ( .A(n19955), .ZN(n17704) );
  NOR2_X1 U20858 ( .A1(n18704), .A2(n17708), .ZN(n17702) );
  OAI21_X1 U20859 ( .B1(n17702), .B2(n18705), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17703) );
  OAI21_X1 U20860 ( .B1(n17704), .B2(n17725), .A(n17703), .ZN(P3_U2634) );
  AOI21_X1 U20861 ( .B1(n19853), .B2(n19856), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17705) );
  AOI22_X1 U20862 ( .A1(n21589), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17705), 
        .B2(n19933), .ZN(P3_U2635) );
  NOR2_X1 U20863 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n17706) );
  OAI21_X1 U20864 ( .B1(n17706), .B2(BS16), .A(n19920), .ZN(n19918) );
  OAI21_X1 U20865 ( .B1(n19920), .B2(n19942), .A(n19918), .ZN(P3_U2636) );
  OAI211_X1 U20866 ( .C1(n18704), .C2(n17708), .A(n17707), .B(n19789), .ZN(
        n17709) );
  INV_X1 U20867 ( .A(n17709), .ZN(n19792) );
  NOR2_X1 U20868 ( .A1(n19792), .A2(n19830), .ZN(n19935) );
  OAI21_X1 U20869 ( .B1(n19935), .B2(n19342), .A(n17710), .ZN(P3_U2637) );
  INV_X1 U20870 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19919) );
  INV_X1 U20871 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21646) );
  NOR2_X1 U20872 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21596) );
  NOR4_X1 U20873 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n17711) );
  OAI211_X1 U20874 ( .C1(n19919), .C2(n21646), .A(n21596), .B(n17711), .ZN(
        n17719) );
  OR4_X1 U20875 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17718) );
  OR4_X1 U20876 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17717) );
  NOR4_X1 U20877 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17715) );
  NOR4_X1 U20878 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17714) );
  NOR4_X1 U20879 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_27__SCAN_IN), .A3(P3_DATAWIDTH_REG_28__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n17713) );
  NOR4_X1 U20880 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n17712) );
  NAND4_X1 U20881 ( .A1(n17715), .A2(n17714), .A3(n17713), .A4(n17712), .ZN(
        n17716) );
  INV_X1 U20882 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19914) );
  NOR3_X1 U20883 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n17721) );
  OAI21_X1 U20884 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17721), .A(n19928), .ZN(
        n17720) );
  OAI21_X1 U20885 ( .B1(n19928), .B2(n19914), .A(n17720), .ZN(P3_U2638) );
  AOI21_X1 U20886 ( .B1(n19924), .B2(n19919), .A(n17721), .ZN(n17722) );
  INV_X1 U20887 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19911) );
  INV_X1 U20888 ( .A(n19928), .ZN(n19931) );
  AOI22_X1 U20889 ( .A1(n19928), .A2(n17722), .B1(n19911), .B2(n19931), .ZN(
        P3_U2639) );
  NAND3_X1 U20890 ( .A1(n17725), .A2(n19832), .A3(n19942), .ZN(n19841) );
  NOR2_X2 U20891 ( .A1(n18649), .A2(n19841), .ZN(n18101) );
  NAND2_X1 U20892 ( .A1(n19835), .A2(n19688), .ZN(n19828) );
  INV_X1 U20893 ( .A(n19944), .ZN(n19844) );
  AOI211_X1 U20894 ( .C1(n19943), .C2(n19941), .A(n19844), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17728) );
  NAND2_X1 U20895 ( .A1(n18707), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17730) );
  INV_X1 U20896 ( .A(n19956), .ZN(n17726) );
  NAND2_X1 U20897 ( .A1(n17730), .A2(n17726), .ZN(n17727) );
  INV_X1 U20898 ( .A(n17728), .ZN(n19823) );
  INV_X1 U20899 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19896) );
  INV_X1 U20900 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19875) );
  INV_X1 U20901 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19866) );
  INV_X1 U20902 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19862) );
  NAND3_X1 U20903 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n18054) );
  NOR2_X1 U20904 ( .A1(n19862), .A2(n18054), .ZN(n18040) );
  NAND2_X1 U20905 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18040), .ZN(n18034) );
  NOR2_X1 U20906 ( .A1(n19866), .A2(n18034), .ZN(n18011) );
  NAND3_X1 U20907 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(n18011), .ZN(n17981) );
  NOR2_X1 U20908 ( .A1(n21816), .A2(n17981), .ZN(n17980) );
  NAND2_X1 U20909 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17980), .ZN(n17964) );
  NOR2_X1 U20910 ( .A1(n19875), .A2(n17964), .ZN(n17956) );
  NAND2_X1 U20911 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17956), .ZN(n17930) );
  NAND2_X1 U20912 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n17891) );
  NOR2_X1 U20913 ( .A1(n17930), .A2(n17891), .ZN(n17865) );
  NAND4_X1 U20914 ( .A1(n17865), .A2(P3_REIP_REG_17__SCAN_IN), .A3(
        P3_REIP_REG_15__SCAN_IN), .A4(P3_REIP_REG_16__SCAN_IN), .ZN(n17826) );
  NAND3_X1 U20915 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n17827) );
  NOR2_X1 U20916 ( .A1(n17826), .A2(n17827), .ZN(n17838) );
  NAND4_X1 U20917 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17838), .A3(
        P3_REIP_REG_22__SCAN_IN), .A4(P3_REIP_REG_21__SCAN_IN), .ZN(n17825) );
  NOR2_X1 U20918 ( .A1(n19896), .A2(n17825), .ZN(n17808) );
  NAND3_X1 U20919 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(P3_REIP_REG_25__SCAN_IN), 
        .A3(n17808), .ZN(n17743) );
  NOR2_X1 U20920 ( .A1(n18102), .A2(n17743), .ZN(n17787) );
  NAND4_X1 U20921 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n17787), .ZN(n17745) );
  NOR3_X1 U20922 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19908), .A3(n17745), 
        .ZN(n17729) );
  AOI21_X1 U20923 ( .B1(n18091), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17729), .ZN(
        n17748) );
  AOI211_X4 U20924 ( .C1(n19942), .C2(n19944), .A(n19956), .B(n17730), .ZN(
        n18076) );
  NOR3_X2 U20925 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18079) );
  NAND2_X1 U20926 ( .A1(n18079), .A2(n18486), .ZN(n18075) );
  NAND2_X1 U20927 ( .A1(n18053), .A2(n18478), .ZN(n18047) );
  NOR2_X2 U20928 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18047), .ZN(n18027) );
  NAND2_X1 U20929 ( .A1(n18027), .A2(n18020), .ZN(n18019) );
  NOR2_X2 U20930 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18019), .ZN(n17995) );
  INV_X1 U20931 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n18374) );
  NAND2_X1 U20932 ( .A1(n17995), .A2(n18374), .ZN(n17977) );
  NAND2_X1 U20933 ( .A1(n17976), .A2(n18375), .ZN(n17968) );
  NAND2_X1 U20934 ( .A1(n17953), .A2(n17949), .ZN(n17948) );
  NOR2_X2 U20935 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17948), .ZN(n17929) );
  INV_X1 U20936 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17924) );
  NAND2_X1 U20937 ( .A1(n17929), .A2(n17924), .ZN(n17922) );
  NOR2_X2 U20938 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17922), .ZN(n17905) );
  INV_X1 U20939 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n18298) );
  NAND2_X1 U20940 ( .A1(n17905), .A2(n18298), .ZN(n17900) );
  INV_X1 U20941 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17875) );
  NAND2_X1 U20942 ( .A1(n17880), .A2(n17875), .ZN(n17874) );
  NAND2_X1 U20943 ( .A1(n17856), .A2(n18123), .ZN(n17852) );
  NAND2_X1 U20944 ( .A1(n17840), .A2(n17834), .ZN(n17833) );
  NOR2_X2 U20945 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17833), .ZN(n17817) );
  NAND2_X1 U20946 ( .A1(n17817), .A2(n17803), .ZN(n17814) );
  INV_X1 U20947 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17789) );
  NAND2_X1 U20948 ( .A1(n17793), .A2(n17789), .ZN(n17788) );
  NOR2_X1 U20949 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17788), .ZN(n17772) );
  INV_X1 U20950 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n21832) );
  NAND2_X1 U20951 ( .A1(n17772), .A2(n21832), .ZN(n17750) );
  NOR2_X1 U20952 ( .A1(n18112), .A2(n17750), .ZN(n17757) );
  INV_X1 U20953 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n18129) );
  INV_X1 U20954 ( .A(n17731), .ZN(n17775) );
  INV_X1 U20955 ( .A(n17732), .ZN(n17783) );
  INV_X1 U20956 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18780) );
  NOR3_X1 U20957 ( .A1(n18110), .A2(n17733), .A3(n18780), .ZN(n17735) );
  OAI21_X1 U20958 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17735), .A(
        n17734), .ZN(n18769) );
  INV_X1 U20959 ( .A(n18769), .ZN(n17807) );
  NOR2_X1 U20960 ( .A1(n18110), .A2(n17733), .ZN(n17737) );
  INV_X1 U20961 ( .A(n17737), .ZN(n17736) );
  AOI21_X1 U20962 ( .B1(n18780), .B2(n17736), .A(n17735), .ZN(n18778) );
  INV_X1 U20963 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18804) );
  INV_X1 U20964 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n21722) );
  NAND3_X1 U20965 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18814), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17739) );
  NOR2_X1 U20966 ( .A1(n21722), .A2(n17739), .ZN(n18765) );
  INV_X1 U20967 ( .A(n18765), .ZN(n17738) );
  AOI21_X1 U20968 ( .B1(n18804), .B2(n17738), .A(n17737), .ZN(n18791) );
  AOI21_X1 U20969 ( .B1(n21722), .B2(n17739), .A(n18765), .ZN(n18825) );
  INV_X1 U20970 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18828) );
  NAND2_X1 U20971 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18814), .ZN(
        n17741) );
  INV_X1 U20972 ( .A(n17739), .ZN(n17740) );
  AOI21_X1 U20973 ( .B1(n18828), .B2(n17741), .A(n17740), .ZN(n18837) );
  NOR3_X1 U20974 ( .A1(n18110), .A2(n18882), .A3(n18881), .ZN(n18856) );
  NAND3_X1 U20975 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n18856), .ZN(n18810) );
  AOI22_X1 U20976 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18814), .B1(
        n18843), .B2(n18810), .ZN(n18847) );
  NOR2_X1 U20977 ( .A1(n18110), .A2(n18891), .ZN(n18893) );
  NAND2_X1 U20978 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18893), .ZN(
        n17917) );
  NOR2_X1 U20979 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17917), .ZN(
        n17912) );
  INV_X1 U20980 ( .A(n17912), .ZN(n17911) );
  NOR2_X1 U20981 ( .A1(n17828), .A2(n18098), .ZN(n17819) );
  NOR2_X1 U20982 ( .A1(n17773), .A2(n18098), .ZN(n17761) );
  NAND2_X1 U20983 ( .A1(n17742), .A2(n18101), .ZN(n18055) );
  NAND2_X1 U20984 ( .A1(n18116), .A2(n18102), .ZN(n18114) );
  NAND3_X1 U20985 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n17744) );
  INV_X1 U20986 ( .A(n18116), .ZN(n18107) );
  AOI21_X1 U20987 ( .B1(n17743), .B2(n18093), .A(n18107), .ZN(n17792) );
  INV_X1 U20988 ( .A(n17792), .ZN(n17799) );
  AOI21_X1 U20989 ( .B1(n18114), .B2(n17744), .A(n17799), .ZN(n17771) );
  NOR2_X1 U20990 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17745), .ZN(n17755) );
  INV_X1 U20991 ( .A(n17755), .ZN(n17746) );
  INV_X1 U20992 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19906) );
  AOI21_X1 U20993 ( .B1(n17771), .B2(n17746), .A(n19906), .ZN(n17747) );
  NAND2_X1 U20994 ( .A1(n18076), .A2(n17750), .ZN(n17767) );
  XOR2_X1 U20995 ( .A(n17752), .B(n17751), .Z(n17756) );
  OAI22_X1 U20996 ( .A1(n17771), .A2(n19908), .B1(n17753), .B2(n18096), .ZN(
        n17754) );
  OAI21_X1 U20997 ( .B1(n18091), .B2(n17757), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17758) );
  OAI211_X1 U20998 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17767), .A(n17759), .B(
        n17758), .ZN(P3_U2641) );
  INV_X1 U20999 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n21585) );
  AOI211_X1 U21000 ( .C1(n17762), .C2(n17761), .A(n17760), .B(n19839), .ZN(
        n17766) );
  NAND3_X1 U21001 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n17787), .ZN(n17764) );
  OAI22_X1 U21002 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17764), .B1(n17763), 
        .B2(n18096), .ZN(n17765) );
  AOI211_X1 U21003 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n18091), .A(n17766), .B(
        n17765), .ZN(n17770) );
  INV_X1 U21004 ( .A(n17767), .ZN(n17768) );
  OAI21_X1 U21005 ( .B1(n17772), .B2(n21832), .A(n17768), .ZN(n17769) );
  OAI211_X1 U21006 ( .C1(n17771), .C2(n21585), .A(n17770), .B(n17769), .ZN(
        P3_U2642) );
  AOI22_X1 U21007 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17781) );
  AOI211_X1 U21008 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17788), .A(n17772), .B(
        n18112), .ZN(n17777) );
  AOI211_X1 U21009 ( .C1(n17775), .C2(n17774), .A(n17773), .B(n19839), .ZN(
        n17776) );
  AOI211_X1 U21010 ( .C1(n17799), .C2(P3_REIP_REG_28__SCAN_IN), .A(n17777), 
        .B(n17776), .ZN(n17780) );
  NAND2_X1 U21011 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17778) );
  OAI211_X1 U21012 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(P3_REIP_REG_27__SCAN_IN), .A(n17787), .B(n17778), .ZN(n17779) );
  NAND3_X1 U21013 ( .A1(n17781), .A2(n17780), .A3(n17779), .ZN(P3_U2643) );
  INV_X1 U21014 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19902) );
  AOI211_X1 U21015 ( .C1(n17783), .C2(n9875), .A(n17782), .B(n19839), .ZN(
        n17786) );
  OAI22_X1 U21016 ( .A1(n17784), .A2(n18096), .B1(n18113), .B2(n17789), .ZN(
        n17785) );
  AOI211_X1 U21017 ( .C1(n17787), .C2(n19902), .A(n17786), .B(n17785), .ZN(
        n17791) );
  OAI211_X1 U21018 ( .C1(n17793), .C2(n17789), .A(n18076), .B(n17788), .ZN(
        n17790) );
  OAI211_X1 U21019 ( .C1(n17792), .C2(n19902), .A(n17791), .B(n17790), .ZN(
        P3_U2644) );
  NAND3_X1 U21020 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n18093), .A3(n17808), 
        .ZN(n17802) );
  AOI22_X1 U21021 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17801) );
  AOI211_X1 U21022 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17814), .A(n17793), .B(
        n18112), .ZN(n17798) );
  AOI211_X1 U21023 ( .C1(n17796), .C2(n17795), .A(n17794), .B(n19839), .ZN(
        n17797) );
  AOI211_X1 U21024 ( .C1(n17799), .C2(P3_REIP_REG_26__SCAN_IN), .A(n17798), 
        .B(n17797), .ZN(n17800) );
  OAI211_X1 U21025 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17802), .A(n17801), 
        .B(n17800), .ZN(P3_U2645) );
  INV_X1 U21026 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19898) );
  AOI21_X1 U21027 ( .B1(n18093), .B2(n17825), .A(n18107), .ZN(n17816) );
  NAND2_X1 U21028 ( .A1(n18093), .A2(n19896), .ZN(n17824) );
  NOR2_X1 U21029 ( .A1(n17817), .A2(n17803), .ZN(n17804) );
  OAI22_X1 U21030 ( .A1(n18112), .A2(n17804), .B1(n18113), .B2(n17803), .ZN(
        n17813) );
  AOI211_X1 U21031 ( .C1(n17807), .C2(n17806), .A(n17805), .B(n19839), .ZN(
        n17812) );
  NAND2_X1 U21032 ( .A1(n18093), .A2(n17808), .ZN(n17810) );
  INV_X1 U21033 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17809) );
  OAI22_X1 U21034 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17810), .B1(n17809), 
        .B2(n18096), .ZN(n17811) );
  AOI211_X1 U21035 ( .C1(n17814), .C2(n17813), .A(n17812), .B(n17811), .ZN(
        n17815) );
  OAI221_X1 U21036 ( .B1(n19898), .B2(n17816), .C1(n19898), .C2(n17824), .A(
        n17815), .ZN(P3_U2646) );
  AOI22_X1 U21037 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n17823) );
  INV_X1 U21038 ( .A(n17816), .ZN(n17832) );
  AOI211_X1 U21039 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17833), .A(n17817), .B(
        n18112), .ZN(n17821) );
  AOI211_X1 U21040 ( .C1(n18778), .C2(n17819), .A(n17818), .B(n19839), .ZN(
        n17820) );
  AOI211_X1 U21041 ( .C1(n17832), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17821), 
        .B(n17820), .ZN(n17822) );
  OAI211_X1 U21042 ( .C1(n17825), .C2(n17824), .A(n17823), .B(n17822), .ZN(
        P3_U2647) );
  NOR2_X1 U21043 ( .A1(n18102), .A2(n17826), .ZN(n17876) );
  INV_X1 U21044 ( .A(n17876), .ZN(n17890) );
  NOR2_X1 U21045 ( .A1(n17827), .A2(n17890), .ZN(n17850) );
  NAND3_X1 U21046 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .A3(n17850), .ZN(n17837) );
  AOI211_X1 U21047 ( .C1(n18791), .C2(n17829), .A(n17828), .B(n19839), .ZN(
        n17831) );
  OAI22_X1 U21048 ( .A1(n18804), .A2(n18096), .B1(n18113), .B2(n17834), .ZN(
        n17830) );
  AOI211_X1 U21049 ( .C1(n17832), .C2(P3_REIP_REG_23__SCAN_IN), .A(n17831), 
        .B(n17830), .ZN(n17836) );
  OAI211_X1 U21050 ( .C1(n17840), .C2(n17834), .A(n18076), .B(n17833), .ZN(
        n17835) );
  OAI211_X1 U21051 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n17837), .A(n17836), 
        .B(n17835), .ZN(P3_U2648) );
  OAI21_X1 U21052 ( .B1(n18102), .B2(n17838), .A(n18116), .ZN(n17851) );
  INV_X1 U21053 ( .A(n17851), .ZN(n17864) );
  INV_X1 U21054 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19892) );
  AOI211_X1 U21055 ( .C1(n18825), .C2(n9903), .A(n17839), .B(n19839), .ZN(
        n17843) );
  AOI211_X1 U21056 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17852), .A(n17840), .B(
        n18112), .ZN(n17842) );
  OAI22_X1 U21057 ( .A1(n21722), .A2(n18096), .B1(n18113), .B2(n10149), .ZN(
        n17841) );
  NOR3_X1 U21058 ( .A1(n17843), .A2(n17842), .A3(n17841), .ZN(n17846) );
  NAND2_X1 U21059 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(P3_REIP_REG_21__SCAN_IN), 
        .ZN(n17844) );
  OAI211_X1 U21060 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17850), .B(n17844), .ZN(n17845) );
  OAI211_X1 U21061 ( .C1(n17864), .C2(n19892), .A(n17846), .B(n17845), .ZN(
        P3_U2649) );
  AOI22_X1 U21062 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n17855) );
  INV_X1 U21063 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19890) );
  AOI211_X1 U21064 ( .C1(n18837), .C2(n17848), .A(n17847), .B(n19839), .ZN(
        n17849) );
  AOI221_X1 U21065 ( .B1(n17851), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n17850), 
        .C2(n19890), .A(n17849), .ZN(n17854) );
  OAI211_X1 U21066 ( .C1(n17856), .C2(n18123), .A(n18076), .B(n17852), .ZN(
        n17853) );
  NAND3_X1 U21067 ( .A1(n17855), .A2(n17854), .A3(n17853), .ZN(P3_U2650) );
  INV_X1 U21068 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19889) );
  AOI211_X1 U21069 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17874), .A(n17856), .B(
        n18112), .ZN(n17857) );
  AOI21_X1 U21070 ( .B1(n18099), .B2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n17857), .ZN(n17863) );
  AOI211_X1 U21071 ( .C1(n18847), .C2(n17859), .A(n17858), .B(n19839), .ZN(
        n17861) );
  INV_X1 U21072 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19887) );
  INV_X1 U21073 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19885) );
  NOR4_X1 U21074 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n19887), .A3(n19885), 
        .A4(n17890), .ZN(n17860) );
  AOI211_X1 U21075 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n18091), .A(n17861), .B(
        n17860), .ZN(n17862) );
  OAI211_X1 U21076 ( .C1(n19889), .C2(n17864), .A(n17863), .B(n17862), .ZN(
        P3_U2651) );
  NAND3_X1 U21077 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .ZN(n17866) );
  NAND2_X1 U21078 ( .A1(n17865), .A2(n18116), .ZN(n17931) );
  OAI21_X1 U21079 ( .B1(n17866), .B2(n17931), .A(n18114), .ZN(n17897) );
  OAI21_X1 U21080 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17890), .A(n17897), 
        .ZN(n17873) );
  NAND2_X1 U21081 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18856), .ZN(
        n17881) );
  INV_X1 U21082 ( .A(n17881), .ZN(n17867) );
  AOI21_X1 U21083 ( .B1(n17912), .B2(n17867), .A(n18098), .ZN(n17884) );
  OAI21_X1 U21084 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17867), .A(
        n18810), .ZN(n17868) );
  INV_X1 U21085 ( .A(n17868), .ZN(n18857) );
  AOI221_X1 U21086 ( .B1(n17884), .B2(n18857), .C1(n17869), .C2(n17868), .A(
        n19839), .ZN(n17872) );
  INV_X1 U21087 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17870) );
  OAI22_X1 U21088 ( .A1(n17870), .A2(n18096), .B1(n18113), .B2(n17875), .ZN(
        n17871) );
  AOI211_X1 U21089 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n17873), .A(n17872), 
        .B(n17871), .ZN(n17879) );
  OAI211_X1 U21090 ( .C1(n17880), .C2(n17875), .A(n18076), .B(n17874), .ZN(
        n17878) );
  NAND3_X1 U21091 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n17876), .A3(n19887), 
        .ZN(n17877) );
  NAND4_X1 U21092 ( .A1(n17879), .A2(n19156), .A3(n17878), .A4(n17877), .ZN(
        P3_U2652) );
  AOI211_X1 U21093 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17900), .A(n17880), .B(
        n18112), .ZN(n17888) );
  OAI21_X1 U21094 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18856), .A(
        n17881), .ZN(n18866) );
  INV_X1 U21095 ( .A(n18866), .ZN(n17885) );
  INV_X1 U21096 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18869) );
  AOI21_X1 U21097 ( .B1(n17912), .B2(n18869), .A(n18866), .ZN(n17882) );
  AOI21_X1 U21098 ( .B1(n17742), .B2(n17882), .A(n19839), .ZN(n17883) );
  OAI21_X1 U21099 ( .B1(n17885), .B2(n17884), .A(n17883), .ZN(n17886) );
  OAI211_X1 U21100 ( .C1(n18113), .C2(n21753), .A(n19156), .B(n17886), .ZN(
        n17887) );
  AOI211_X1 U21101 ( .C1(n18099), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n17888), .B(n17887), .ZN(n17889) );
  OAI221_X1 U21102 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17890), .C1(n19885), 
        .C2(n17897), .A(n17889), .ZN(P3_U2653) );
  INV_X1 U21103 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n21819) );
  INV_X1 U21104 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19883) );
  NOR2_X1 U21105 ( .A1(n21819), .A2(n19883), .ZN(n17904) );
  NOR3_X1 U21106 ( .A1(n18102), .A2(n17930), .A3(n17891), .ZN(n17903) );
  AOI21_X1 U21107 ( .B1(n17904), .B2(n17903), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n17898) );
  INV_X1 U21108 ( .A(n18882), .ZN(n17892) );
  NAND2_X1 U21109 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17892), .ZN(
        n17893) );
  AOI21_X1 U21110 ( .B1(n18881), .B2(n17893), .A(n18856), .ZN(n18884) );
  INV_X1 U21111 ( .A(n17917), .ZN(n17894) );
  OAI21_X1 U21112 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17894), .A(
        n17893), .ZN(n18899) );
  AOI21_X1 U21113 ( .B1(n17912), .B2(n18899), .A(n18098), .ZN(n17895) );
  XNOR2_X1 U21114 ( .A(n18884), .B(n17895), .ZN(n17896) );
  OAI22_X1 U21115 ( .A1(n17898), .A2(n17897), .B1(n19839), .B2(n17896), .ZN(
        n17899) );
  AOI211_X1 U21116 ( .C1(n18091), .C2(P3_EBX_REG_17__SCAN_IN), .A(n19268), .B(
        n17899), .ZN(n17902) );
  OAI211_X1 U21117 ( .C1(n17905), .C2(n18298), .A(n18076), .B(n17900), .ZN(
        n17901) );
  OAI211_X1 U21118 ( .C1(n18096), .C2(n18881), .A(n17902), .B(n17901), .ZN(
        P3_U2654) );
  NAND2_X1 U21119 ( .A1(n18114), .A2(n17931), .ZN(n17940) );
  INV_X1 U21120 ( .A(n17903), .ZN(n17928) );
  AOI211_X1 U21121 ( .C1(n21819), .C2(n19883), .A(n17904), .B(n17928), .ZN(
        n17910) );
  AOI211_X1 U21122 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17922), .A(n17905), .B(
        n18112), .ZN(n17909) );
  OAI22_X1 U21123 ( .A1(n17907), .A2(n18096), .B1(n18113), .B2(n17906), .ZN(
        n17908) );
  NOR4_X1 U21124 ( .A1(n19268), .A2(n17910), .A3(n17909), .A4(n17908), .ZN(
        n17916) );
  NAND2_X1 U21125 ( .A1(n17742), .A2(n17911), .ZN(n17914) );
  OAI21_X1 U21126 ( .B1(n17912), .B2(n18098), .A(n18899), .ZN(n17913) );
  OAI211_X1 U21127 ( .C1(n18899), .C2(n17914), .A(n18101), .B(n17913), .ZN(
        n17915) );
  OAI211_X1 U21128 ( .C1(n17940), .C2(n19883), .A(n17916), .B(n17915), .ZN(
        P3_U2655) );
  OAI21_X1 U21129 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18893), .A(
        n17917), .ZN(n18917) );
  INV_X1 U21130 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n18097) );
  NAND2_X1 U21131 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18097), .ZN(
        n18018) );
  INV_X1 U21132 ( .A(n18018), .ZN(n18085) );
  NAND2_X1 U21133 ( .A1(n17918), .A2(n18085), .ZN(n17919) );
  OAI21_X1 U21134 ( .B1(n18895), .B2(n17919), .A(n17742), .ZN(n17921) );
  OAI21_X1 U21135 ( .B1(n18917), .B2(n17921), .A(n18101), .ZN(n17920) );
  AOI21_X1 U21136 ( .B1(n18917), .B2(n17921), .A(n17920), .ZN(n17926) );
  OAI211_X1 U21137 ( .C1(n17929), .C2(n17924), .A(n18076), .B(n17922), .ZN(
        n17923) );
  OAI211_X1 U21138 ( .C1(n18113), .C2(n17924), .A(n19156), .B(n17923), .ZN(
        n17925) );
  AOI211_X1 U21139 ( .C1(n18099), .C2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n17926), .B(n17925), .ZN(n17927) );
  OAI221_X1 U21140 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n17928), .C1(n21819), 
        .C2(n17940), .A(n17927), .ZN(P3_U2656) );
  INV_X1 U21141 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19881) );
  AOI211_X1 U21142 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17948), .A(n17929), .B(
        n18112), .ZN(n17934) );
  INV_X1 U21143 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n21689) );
  NOR2_X1 U21144 ( .A1(n18102), .A2(n17930), .ZN(n17944) );
  NAND3_X1 U21145 ( .A1(n17944), .A2(P3_REIP_REG_13__SCAN_IN), .A3(n17931), 
        .ZN(n17932) );
  OAI211_X1 U21146 ( .C1(n21689), .C2(n18096), .A(n19156), .B(n17932), .ZN(
        n17933) );
  AOI211_X1 U21147 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n18091), .A(n17934), .B(
        n17933), .ZN(n17939) );
  AOI21_X1 U21148 ( .B1(n21689), .B2(n17935), .A(n18893), .ZN(n18930) );
  OAI21_X1 U21149 ( .B1(n18894), .B2(n18018), .A(n17742), .ZN(n17959) );
  OAI21_X1 U21150 ( .B1(n18925), .B2(n18098), .A(n17959), .ZN(n17937) );
  AOI21_X1 U21151 ( .B1(n18930), .B2(n17937), .A(n19839), .ZN(n17936) );
  OAI21_X1 U21152 ( .B1(n18930), .B2(n17937), .A(n17936), .ZN(n17938) );
  OAI211_X1 U21153 ( .C1(n17940), .C2(n19881), .A(n17939), .B(n17938), .ZN(
        P3_U2657) );
  OAI21_X1 U21154 ( .B1(n17956), .B2(n18102), .A(n18116), .ZN(n17974) );
  NOR2_X1 U21155 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n18102), .ZN(n17955) );
  INV_X1 U21156 ( .A(n17941), .ZN(n17957) );
  OAI21_X1 U21157 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17957), .A(
        n17742), .ZN(n17942) );
  XNOR2_X1 U21158 ( .A(n17943), .B(n17942), .ZN(n17946) );
  AOI22_X1 U21159 ( .A1(n18091), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17944), 
        .B2(n21778), .ZN(n17945) );
  OAI211_X1 U21160 ( .C1(n19839), .C2(n17946), .A(n17945), .B(n19156), .ZN(
        n17947) );
  AOI221_X1 U21161 ( .B1(n17974), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17955), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17947), .ZN(n17951) );
  OAI211_X1 U21162 ( .C1(n17953), .C2(n17949), .A(n18076), .B(n17948), .ZN(
        n17950) );
  OAI211_X1 U21163 ( .C1(n18096), .C2(n17952), .A(n17951), .B(n17950), .ZN(
        P3_U2658) );
  AOI22_X1 U21164 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n17963) );
  AOI211_X1 U21165 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17968), .A(n17953), .B(
        n18112), .ZN(n17954) );
  AOI211_X1 U21166 ( .C1(n17956), .C2(n17955), .A(n19268), .B(n17954), .ZN(
        n17962) );
  OAI21_X1 U21167 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17958), .A(
        n17957), .ZN(n18938) );
  XOR2_X1 U21168 ( .A(n18938), .B(n17959), .Z(n17960) );
  AOI22_X1 U21169 ( .A1(n18101), .A2(n17960), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17974), .ZN(n17961) );
  NAND3_X1 U21170 ( .A1(n17963), .A2(n17962), .A3(n17961), .ZN(P3_U2659) );
  OAI21_X1 U21171 ( .B1(n18102), .B2(n17964), .A(n19875), .ZN(n17973) );
  INV_X1 U21172 ( .A(n17966), .ZN(n17967) );
  NOR2_X1 U21173 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17984), .ZN(
        n18005) );
  AOI21_X1 U21174 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18005), .A(
        n18098), .ZN(n17986) );
  INV_X1 U21175 ( .A(n17986), .ZN(n17965) );
  OAI221_X1 U21176 ( .B1(n17967), .B2(n17986), .C1(n17966), .C2(n17965), .A(
        n18101), .ZN(n17970) );
  OAI211_X1 U21177 ( .C1(n17976), .C2(n18375), .A(n18076), .B(n17968), .ZN(
        n17969) );
  OAI211_X1 U21178 ( .C1(n18096), .C2(n17971), .A(n17970), .B(n17969), .ZN(
        n17972) );
  AOI21_X1 U21179 ( .B1(n17974), .B2(n17973), .A(n17972), .ZN(n17975) );
  OAI211_X1 U21180 ( .C1(n18113), .C2(n18375), .A(n17975), .B(n19156), .ZN(
        P3_U2660) );
  AOI22_X1 U21181 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18099), .B1(
        n18091), .B2(P3_EBX_REG_10__SCAN_IN), .ZN(n17991) );
  NOR2_X1 U21182 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n18102), .ZN(n17979) );
  AOI211_X1 U21183 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17977), .A(n17976), .B(
        n18112), .ZN(n17978) );
  AOI211_X1 U21184 ( .C1(n17980), .C2(n17979), .A(n19268), .B(n17978), .ZN(
        n17990) );
  AOI21_X1 U21185 ( .B1(n17981), .B2(n18093), .A(n18107), .ZN(n18012) );
  INV_X1 U21186 ( .A(n18012), .ZN(n18001) );
  NOR3_X1 U21187 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n18102), .A3(n17981), .ZN(
        n17994) );
  OAI21_X1 U21188 ( .B1(n18001), .B2(n17994), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n17989) );
  AOI21_X1 U21189 ( .B1(n17983), .B2(n17984), .A(n17982), .ZN(n17987) );
  INV_X1 U21190 ( .A(n17987), .ZN(n18955) );
  OAI21_X1 U21191 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17984), .A(
        n17742), .ZN(n17985) );
  OAI221_X1 U21192 ( .B1(n17987), .B2(n17986), .C1(n18955), .C2(n17985), .A(
        n18101), .ZN(n17988) );
  NAND4_X1 U21193 ( .A1(n17991), .A2(n17990), .A3(n17989), .A4(n17988), .ZN(
        P3_U2661) );
  NOR2_X1 U21194 ( .A1(n19839), .A2(n18018), .ZN(n18057) );
  INV_X1 U21195 ( .A(n18055), .ZN(n17992) );
  AOI22_X1 U21196 ( .A1(n17993), .A2(n18057), .B1(n17992), .B2(n17997), .ZN(
        n18004) );
  NOR2_X1 U21197 ( .A1(n17995), .A2(n18112), .ZN(n18010) );
  AOI211_X1 U21198 ( .C1(n18010), .C2(n18374), .A(n19268), .B(n17994), .ZN(
        n18003) );
  INV_X1 U21199 ( .A(n17995), .ZN(n17996) );
  AOI221_X1 U21200 ( .B1(n18112), .B2(n18113), .C1(n17996), .C2(n18113), .A(
        n18374), .ZN(n18000) );
  NAND2_X1 U21201 ( .A1(n18101), .A2(n18098), .ZN(n18051) );
  OAI22_X1 U21202 ( .A1(n17998), .A2(n18096), .B1(n17997), .B2(n18051), .ZN(
        n17999) );
  AOI211_X1 U21203 ( .C1(n18001), .C2(P3_REIP_REG_9__SCAN_IN), .A(n18000), .B(
        n17999), .ZN(n18002) );
  OAI211_X1 U21204 ( .C1(n18005), .C2(n18004), .A(n18003), .B(n18002), .ZN(
        P3_U2662) );
  OAI21_X1 U21205 ( .B1(n18006), .B2(n18018), .A(n17742), .ZN(n18007) );
  XNOR2_X1 U21206 ( .A(n18008), .B(n18007), .ZN(n18016) );
  NAND2_X1 U21207 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18019), .ZN(n18009) );
  AOI22_X1 U21208 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n18099), .B1(
        n18010), .B2(n18009), .ZN(n18015) );
  INV_X1 U21209 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19868) );
  NAND2_X1 U21210 ( .A1(n18093), .A2(n18011), .ZN(n18022) );
  AOI221_X1 U21211 ( .B1(n19868), .B2(n19870), .C1(n18022), .C2(n19870), .A(
        n18012), .ZN(n18013) );
  AOI211_X1 U21212 ( .C1(n18091), .C2(P3_EBX_REG_8__SCAN_IN), .A(n19268), .B(
        n18013), .ZN(n18014) );
  OAI211_X1 U21213 ( .C1(n19839), .C2(n18016), .A(n18015), .B(n18014), .ZN(
        P3_U2663) );
  AOI21_X1 U21214 ( .B1(n18093), .B2(n18034), .A(n18107), .ZN(n18045) );
  NAND2_X1 U21215 ( .A1(n18093), .A2(n19866), .ZN(n18033) );
  AOI21_X1 U21216 ( .B1(n18973), .B2(n18029), .A(n18017), .ZN(n18979) );
  OAI21_X1 U21217 ( .B1(n18972), .B2(n18018), .A(n17742), .ZN(n18032) );
  XNOR2_X1 U21218 ( .A(n18979), .B(n18032), .ZN(n18025) );
  OAI22_X1 U21219 ( .A1(n18973), .A2(n18096), .B1(n18113), .B2(n18020), .ZN(
        n18024) );
  OAI211_X1 U21220 ( .C1(n18027), .C2(n18020), .A(n18076), .B(n18019), .ZN(
        n18021) );
  OAI211_X1 U21221 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n18022), .A(n19156), .B(
        n18021), .ZN(n18023) );
  AOI211_X1 U21222 ( .C1(n18101), .C2(n18025), .A(n18024), .B(n18023), .ZN(
        n18026) );
  OAI221_X1 U21223 ( .B1(n19868), .B2(n18045), .C1(n19868), .C2(n18033), .A(
        n18026), .ZN(P3_U2664) );
  AOI211_X1 U21224 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n18047), .A(n18027), .B(
        n18112), .ZN(n18028) );
  AOI211_X1 U21225 ( .C1(n18091), .C2(P3_EBX_REG_6__SCAN_IN), .A(n19268), .B(
        n18028), .ZN(n18039) );
  INV_X1 U21226 ( .A(n18045), .ZN(n18037) );
  INV_X1 U21227 ( .A(n18030), .ZN(n18041) );
  OAI21_X1 U21228 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18030), .A(
        n18029), .ZN(n18991) );
  OAI21_X1 U21229 ( .B1(n18098), .B2(n18097), .A(n18101), .ZN(n18111) );
  AOI211_X1 U21230 ( .C1(n17742), .C2(n18041), .A(n18991), .B(n18111), .ZN(
        n18036) );
  NAND2_X1 U21231 ( .A1(n18101), .A2(n18991), .ZN(n18031) );
  OAI22_X1 U21232 ( .A1(n18034), .A2(n18033), .B1(n18032), .B2(n18031), .ZN(
        n18035) );
  AOI211_X1 U21233 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n18037), .A(n18036), .B(
        n18035), .ZN(n18038) );
  OAI211_X1 U21234 ( .C1(n18990), .C2(n18096), .A(n18039), .B(n18038), .ZN(
        P3_U2665) );
  INV_X1 U21235 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18050) );
  AOI21_X1 U21236 ( .B1(n18093), .B2(n18040), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n18044) );
  AND2_X1 U21237 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19000), .ZN(
        n18056) );
  AOI21_X1 U21238 ( .B1(n18056), .B2(n18097), .A(n18098), .ZN(n18042) );
  OAI21_X1 U21239 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18056), .A(
        n18041), .ZN(n19003) );
  XOR2_X1 U21240 ( .A(n18042), .B(n19003), .Z(n18043) );
  OAI22_X1 U21241 ( .A1(n18045), .A2(n18044), .B1(n19839), .B2(n18043), .ZN(
        n18046) );
  AOI211_X1 U21242 ( .C1(n18091), .C2(P3_EBX_REG_5__SCAN_IN), .A(n19268), .B(
        n18046), .ZN(n18049) );
  OAI211_X1 U21243 ( .C1(n18053), .C2(n18478), .A(n18076), .B(n18047), .ZN(
        n18048) );
  OAI211_X1 U21244 ( .C1(n18096), .C2(n18050), .A(n18049), .B(n18048), .ZN(
        P3_U2666) );
  INV_X1 U21245 ( .A(n18051), .ZN(n18082) );
  OR2_X1 U21246 ( .A1(n18110), .A2(n19007), .ZN(n18068) );
  AOI21_X1 U21247 ( .B1(n19022), .B2(n18068), .A(n18056), .ZN(n19019) );
  NOR3_X1 U21248 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n18102), .A3(n18054), .ZN(
        n18052) );
  AOI21_X1 U21249 ( .B1(n18082), .B2(n19019), .A(n18052), .ZN(n18066) );
  AOI211_X1 U21250 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n18075), .A(n18053), .B(
        n18112), .ZN(n18064) );
  AOI21_X1 U21251 ( .B1(n18093), .B2(n18054), .A(n18107), .ZN(n18069) );
  AOI211_X1 U21252 ( .C1(n18056), .C2(n18097), .A(n19019), .B(n18055), .ZN(
        n18061) );
  NAND2_X1 U21253 ( .A1(n19958), .A2(n19355), .ZN(n18120) );
  NOR2_X1 U21254 ( .A1(n9717), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n18059) );
  NOR2_X1 U21255 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19007), .ZN(
        n19014) );
  NAND2_X1 U21256 ( .A1(n18057), .A2(n19014), .ZN(n18058) );
  OAI21_X1 U21257 ( .B1(n18120), .B2(n18059), .A(n18058), .ZN(n18060) );
  NOR2_X1 U21258 ( .A1(n18061), .A2(n18060), .ZN(n18062) );
  OAI211_X1 U21259 ( .C1(n18069), .C2(n19862), .A(n18062), .B(n19156), .ZN(
        n18063) );
  AOI211_X1 U21260 ( .C1(n18099), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n18064), .B(n18063), .ZN(n18065) );
  OAI211_X1 U21261 ( .C1(n18113), .C2(n18067), .A(n18066), .B(n18065), .ZN(
        P3_U2667) );
  INV_X1 U21262 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21676) );
  INV_X1 U21263 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19046) );
  NOR2_X1 U21264 ( .A1(n18110), .A2(n19046), .ZN(n18081) );
  AOI21_X1 U21265 ( .B1(n18081), .B2(n18097), .A(n18098), .ZN(n18083) );
  OAI21_X1 U21266 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n18081), .A(
        n18068), .ZN(n19029) );
  XNOR2_X1 U21267 ( .A(n18083), .B(n19029), .ZN(n18074) );
  INV_X1 U21268 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19860) );
  NAND2_X1 U21269 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n18092) );
  AOI221_X1 U21270 ( .B1(n18102), .B2(n19860), .C1(n18092), .C2(n19860), .A(
        n18069), .ZN(n18073) );
  INV_X1 U21271 ( .A(n18070), .ZN(n18071) );
  OAI22_X1 U21272 ( .A1(n18120), .A2(n18071), .B1(n18486), .B2(n18113), .ZN(
        n18072) );
  AOI211_X1 U21273 ( .C1(n18074), .C2(n18101), .A(n18073), .B(n18072), .ZN(
        n18078) );
  OAI211_X1 U21274 ( .C1(n18079), .C2(n18486), .A(n18076), .B(n18075), .ZN(
        n18077) );
  OAI211_X1 U21275 ( .C1(n18096), .C2(n21676), .A(n18078), .B(n18077), .ZN(
        P3_U2668) );
  INV_X1 U21276 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18500) );
  INV_X1 U21277 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18494) );
  NAND2_X1 U21278 ( .A1(n18500), .A2(n18494), .ZN(n18080) );
  AOI211_X1 U21279 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18080), .A(n18079), .B(
        n18112), .ZN(n18090) );
  AOI21_X1 U21280 ( .B1(n18110), .B2(n19046), .A(n18081), .ZN(n19042) );
  AOI22_X1 U21281 ( .A1(n18107), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19042), 
        .B2(n18082), .ZN(n18087) );
  INV_X1 U21282 ( .A(n19042), .ZN(n18084) );
  OAI211_X1 U21283 ( .C1(n18085), .C2(n18084), .A(n18101), .B(n18083), .ZN(
        n18086) );
  OAI211_X1 U21284 ( .C1(n18120), .C2(n18088), .A(n18087), .B(n18086), .ZN(
        n18089) );
  AOI211_X1 U21285 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n18091), .A(n18090), .B(
        n18089), .ZN(n18095) );
  OAI211_X1 U21286 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n18093), .B(n18092), .ZN(n18094) );
  OAI211_X1 U21287 ( .C1(n18096), .C2(n19046), .A(n18095), .B(n18094), .ZN(
        P3_U2669) );
  NOR2_X1 U21288 ( .A1(n18098), .A2(n18097), .ZN(n18100) );
  AOI21_X1 U21289 ( .B1(n18101), .B2(n18100), .A(n18099), .ZN(n18109) );
  OAI22_X1 U21290 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18102), .B1(n18113), 
        .B2(n18494), .ZN(n18106) );
  NOR2_X1 U21291 ( .A1(n18500), .A2(n18494), .ZN(n18490) );
  INV_X1 U21292 ( .A(n18490), .ZN(n18103) );
  OAI21_X1 U21293 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n18103), .ZN(n18496) );
  OAI22_X1 U21294 ( .A1(n18112), .A2(n18496), .B1(n18120), .B2(n18104), .ZN(
        n18105) );
  AOI211_X1 U21295 ( .C1(n18107), .C2(P3_REIP_REG_1__SCAN_IN), .A(n18106), .B(
        n18105), .ZN(n18108) );
  OAI221_X1 U21296 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18111), .C1(
        n18110), .C2(n18109), .A(n18108), .ZN(P3_U2670) );
  NAND2_X1 U21297 ( .A1(n18113), .A2(n18112), .ZN(n18115) );
  AOI22_X1 U21298 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n18115), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n18114), .ZN(n18119) );
  NAND3_X1 U21299 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18117), .A3(
        n18116), .ZN(n18118) );
  OAI211_X1 U21300 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18120), .A(
        n18119), .B(n18118), .ZN(P3_U2671) );
  INV_X1 U21301 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n18121) );
  NOR2_X1 U21302 ( .A1(n18121), .A2(n18261), .ZN(n18207) );
  INV_X1 U21303 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n18124) );
  NAND3_X1 U21304 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n18122), .ZN(n18166) );
  NOR4_X1 U21305 ( .A1(n21832), .A2(n18124), .A3(n18123), .A4(n18166), .ZN(
        n18125) );
  NAND4_X1 U21306 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n18207), .A4(n18125), .ZN(n18128) );
  NOR2_X1 U21307 ( .A1(n18129), .A2(n18128), .ZN(n18162) );
  NAND2_X1 U21308 ( .A1(n18484), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n18127) );
  NAND2_X1 U21309 ( .A1(n18162), .A2(n9734), .ZN(n18126) );
  OAI22_X1 U21310 ( .A1(n18162), .A2(n18127), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n18126), .ZN(P3_U2672) );
  NAND2_X1 U21311 ( .A1(n18129), .A2(n18128), .ZN(n18130) );
  NAND2_X1 U21312 ( .A1(n18130), .A2(n18484), .ZN(n18161) );
  INV_X1 U21313 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18137) );
  OAI22_X1 U21314 ( .A1(n9712), .A2(n18132), .B1(n18381), .B2(n18131), .ZN(
        n18134) );
  OAI22_X1 U21315 ( .A1(n9724), .A2(n18326), .B1(n18443), .B2(n18329), .ZN(
        n18133) );
  AOI211_X1 U21316 ( .C1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .C2(n9717), .A(
        n18134), .B(n18133), .ZN(n18136) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17006), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18135) );
  OAI211_X1 U21318 ( .C1(n18137), .C2(n18455), .A(n18136), .B(n18135), .ZN(
        n18143) );
  AOI22_X1 U21319 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18141) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18269), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n18140) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18420), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18139) );
  AOI22_X1 U21322 ( .A1(n18457), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n18138) );
  NAND4_X1 U21323 ( .A1(n18141), .A2(n18140), .A3(n18139), .A4(n18138), .ZN(
        n18142) );
  NOR2_X1 U21324 ( .A1(n18143), .A2(n18142), .ZN(n18160) );
  INV_X1 U21325 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18152) );
  INV_X1 U21326 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18144) );
  OAI22_X1 U21327 ( .A1(n18443), .A2(n18145), .B1(n13729), .B2(n18144), .ZN(
        n18149) );
  INV_X1 U21328 ( .A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18147) );
  INV_X1 U21329 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n18146) );
  OAI22_X1 U21330 ( .A1(n9724), .A2(n18147), .B1(n18445), .B2(n18146), .ZN(
        n18148) );
  AOI211_X1 U21331 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n18149), .B(n18148), .ZN(n18151) );
  AOI22_X1 U21332 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18150) );
  OAI211_X1 U21333 ( .C1(n18455), .C2(n18152), .A(n18151), .B(n18150), .ZN(
        n18159) );
  AOI22_X1 U21334 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n18153), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18157) );
  AOI22_X1 U21335 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U21336 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U21337 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18154) );
  NAND4_X1 U21338 ( .A1(n18157), .A2(n18156), .A3(n18155), .A4(n18154), .ZN(
        n18158) );
  OR2_X1 U21339 ( .A1(n18159), .A2(n18158), .ZN(n18164) );
  NAND2_X1 U21340 ( .A1(n18165), .A2(n18164), .ZN(n18163) );
  XNOR2_X1 U21341 ( .A(n18160), .B(n18163), .ZN(n18510) );
  OAI22_X1 U21342 ( .A1(n18162), .A2(n18161), .B1(n18510), .B2(n18484), .ZN(
        P3_U2673) );
  OAI21_X1 U21343 ( .B1(n18165), .B2(n18164), .A(n18163), .ZN(n18518) );
  NOR2_X1 U21344 ( .A1(n18177), .A2(n18166), .ZN(n18167) );
  OAI21_X1 U21345 ( .B1(n18173), .B2(n18170), .A(n18169), .ZN(n18526) );
  NAND3_X1 U21346 ( .A1(n18172), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n18484), 
        .ZN(n18171) );
  OAI221_X1 U21347 ( .B1(n18172), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n18484), 
        .C2(n18526), .A(n18171), .ZN(P3_U2676) );
  AOI21_X1 U21348 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18484), .A(n18181), .ZN(
        n18176) );
  AOI21_X1 U21349 ( .B1(n18174), .B2(n18178), .A(n18173), .ZN(n18527) );
  INV_X1 U21350 ( .A(n18527), .ZN(n18175) );
  OAI22_X1 U21351 ( .A1(n10143), .A2(n18176), .B1(n18484), .B2(n18175), .ZN(
        P3_U2677) );
  INV_X1 U21352 ( .A(n18177), .ZN(n18186) );
  AOI21_X1 U21353 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18484), .A(n18186), .ZN(
        n18180) );
  OAI21_X1 U21354 ( .B1(n18182), .B2(n18179), .A(n18178), .ZN(n18536) );
  OAI22_X1 U21355 ( .A1(n18181), .A2(n18180), .B1(n18484), .B2(n18536), .ZN(
        P3_U2678) );
  AOI21_X1 U21356 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18484), .A(n9802), .ZN(
        n18185) );
  AOI21_X1 U21357 ( .B1(n18183), .B2(n18187), .A(n18182), .ZN(n18537) );
  INV_X1 U21358 ( .A(n18537), .ZN(n18184) );
  OAI22_X1 U21359 ( .A1(n18186), .A2(n18185), .B1(n18484), .B2(n18184), .ZN(
        P3_U2679) );
  AOI21_X1 U21360 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18484), .A(n9803), .ZN(
        n18190) );
  OAI21_X1 U21361 ( .B1(n18189), .B2(n18188), .A(n18187), .ZN(n18549) );
  OAI22_X1 U21362 ( .A1(n9802), .A2(n18190), .B1(n18484), .B2(n18549), .ZN(
        P3_U2680) );
  AOI21_X1 U21363 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18484), .A(n18191), .ZN(
        n18206) );
  INV_X1 U21364 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18199) );
  INV_X1 U21365 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n18192) );
  INV_X1 U21366 ( .A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18343) );
  OAI22_X1 U21367 ( .A1(n18445), .A2(n18192), .B1(n13729), .B2(n18343), .ZN(
        n18196) );
  INV_X1 U21368 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18194) );
  INV_X1 U21369 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18340) );
  OAI22_X1 U21370 ( .A1(n14490), .A2(n18194), .B1(n13705), .B2(n18340), .ZN(
        n18195) );
  AOI211_X1 U21371 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n18196), .B(n18195), .ZN(n18198) );
  AOI22_X1 U21372 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18197) );
  OAI211_X1 U21373 ( .C1(n18455), .C2(n18199), .A(n18198), .B(n18197), .ZN(
        n18205) );
  AOI22_X1 U21374 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18203) );
  AOI22_X1 U21375 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U21376 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18201) );
  AOI22_X1 U21377 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18200) );
  NAND4_X1 U21378 ( .A1(n18203), .A2(n18202), .A3(n18201), .A4(n18200), .ZN(
        n18204) );
  NOR2_X1 U21379 ( .A1(n18205), .A2(n18204), .ZN(n18552) );
  OAI22_X1 U21380 ( .A1(n9803), .A2(n18206), .B1(n18552), .B2(n18484), .ZN(
        P3_U2681) );
  NOR2_X1 U21381 ( .A1(n18498), .A2(n18207), .ZN(n18243) );
  AOI22_X1 U21382 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n18208) );
  OAI21_X1 U21383 ( .B1(n10740), .B2(n18209), .A(n18208), .ZN(n18210) );
  AOI21_X1 U21384 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(n18210), .ZN(n18213) );
  AOI22_X1 U21385 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n18212) );
  AOI22_X1 U21386 ( .A1(n18457), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18211) );
  NAND3_X1 U21387 ( .A1(n18213), .A2(n18212), .A3(n18211), .ZN(n18221) );
  INV_X1 U21388 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U21389 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18420), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n18214) );
  OAI21_X1 U21390 ( .B1(n13705), .B2(n18215), .A(n18214), .ZN(n18216) );
  AOI21_X1 U21391 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A(
        n18216), .ZN(n18219) );
  AOI22_X1 U21392 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n18218) );
  AOI22_X1 U21393 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18217) );
  NAND3_X1 U21394 ( .A1(n18219), .A2(n18218), .A3(n18217), .ZN(n18220) );
  NOR2_X1 U21395 ( .A1(n18221), .A2(n18220), .ZN(n18560) );
  INV_X1 U21396 ( .A(n18560), .ZN(n18222) );
  AOI22_X1 U21397 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n18243), .B1(n18498), 
        .B2(n18222), .ZN(n18223) );
  OAI21_X1 U21398 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n18224), .A(n18223), .ZN(
        P3_U2682) );
  INV_X1 U21399 ( .A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n18227) );
  AOI22_X1 U21400 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18226) );
  NAND2_X1 U21401 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n18225) );
  OAI211_X1 U21402 ( .C1(n18227), .C2(n18381), .A(n18226), .B(n18225), .ZN(
        n18233) );
  INV_X1 U21403 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n18367) );
  OAI22_X1 U21404 ( .A1(n14490), .A2(n18367), .B1(n10740), .B2(n18228), .ZN(
        n18232) );
  INV_X1 U21405 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18229) );
  OAI22_X1 U21406 ( .A1(n9724), .A2(n18230), .B1(n18301), .B2(n18229), .ZN(
        n18231) );
  OR3_X1 U21407 ( .A1(n18233), .A2(n18232), .A3(n18231), .ZN(n18242) );
  AOI22_X1 U21408 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18235) );
  NAND2_X1 U21409 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n18234) );
  OAI211_X1 U21410 ( .C1(n9799), .C2(n18361), .A(n18235), .B(n18234), .ZN(
        n18236) );
  INV_X1 U21411 ( .A(n18236), .ZN(n18240) );
  AOI22_X1 U21412 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18237), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18239) );
  AOI22_X1 U21413 ( .A1(n18153), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18238) );
  NAND3_X1 U21414 ( .A1(n18240), .A2(n18239), .A3(n18238), .ZN(n18241) );
  NOR2_X1 U21415 ( .A1(n18242), .A2(n18241), .ZN(n18565) );
  OAI21_X1 U21416 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n18244), .A(n18243), .ZN(
        n18245) );
  OAI21_X1 U21417 ( .B1(n18565), .B2(n18484), .A(n18245), .ZN(P3_U2683) );
  INV_X1 U21418 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18253) );
  INV_X1 U21419 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n18247) );
  INV_X1 U21420 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18246) );
  OAI22_X1 U21421 ( .A1(n14490), .A2(n18247), .B1(n18402), .B2(n18246), .ZN(
        n18250) );
  INV_X1 U21422 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n18248) );
  OAI22_X1 U21423 ( .A1(n9724), .A2(n18248), .B1(n13729), .B2(n18382), .ZN(
        n18249) );
  AOI211_X1 U21424 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n18250), .B(n18249), .ZN(n18252) );
  AOI22_X1 U21425 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18251) );
  OAI211_X1 U21426 ( .C1(n18455), .C2(n18253), .A(n18252), .B(n18251), .ZN(
        n18260) );
  AOI22_X1 U21427 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18258) );
  AOI22_X1 U21428 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18254), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U21429 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18256) );
  AOI22_X1 U21430 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18255) );
  NAND4_X1 U21431 ( .A1(n18258), .A2(n18257), .A3(n18256), .A4(n18255), .ZN(
        n18259) );
  NOR2_X1 U21432 ( .A1(n18260), .A2(n18259), .ZN(n18569) );
  OAI21_X1 U21433 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n9880), .A(n18261), .ZN(
        n18262) );
  AOI22_X1 U21434 ( .A1(n18498), .A2(n18569), .B1(n18262), .B2(n18484), .ZN(
        P3_U2684) );
  INV_X1 U21435 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18264) );
  AOI22_X1 U21436 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U21437 ( .B1(n18402), .B2(n18264), .A(n18263), .ZN(n18265) );
  AOI21_X1 U21438 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n18265), .ZN(n18268) );
  AOI22_X1 U21439 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18267) );
  AOI22_X1 U21440 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18266) );
  NAND3_X1 U21441 ( .A1(n18268), .A2(n18267), .A3(n18266), .ZN(n18278) );
  AOI22_X1 U21442 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n18271) );
  NAND2_X1 U21443 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n18270) );
  OAI211_X1 U21444 ( .C1(n9799), .C2(n18272), .A(n18271), .B(n18270), .ZN(
        n18276) );
  OAI22_X1 U21445 ( .A1(n9712), .A2(n18401), .B1(n18273), .B2(n18400), .ZN(
        n18275) );
  INV_X1 U21446 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18493) );
  INV_X1 U21447 ( .A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n18405) );
  OAI22_X1 U21448 ( .A1(n18330), .A2(n18493), .B1(n18381), .B2(n18405), .ZN(
        n18274) );
  OR3_X1 U21449 ( .A1(n18276), .A2(n18275), .A3(n18274), .ZN(n18277) );
  NOR2_X1 U21450 ( .A1(n18278), .A2(n18277), .ZN(n18574) );
  INV_X1 U21451 ( .A(n18280), .ZN(n18279) );
  OAI33_X1 U21452 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n18595), .A3(n18280), 
        .B1(n21753), .B2(n18498), .B3(n18279), .ZN(n18281) );
  INV_X1 U21453 ( .A(n18281), .ZN(n18282) );
  OAI21_X1 U21454 ( .B1(n18574), .B2(n18484), .A(n18282), .ZN(P3_U2685) );
  INV_X1 U21455 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n18430) );
  INV_X1 U21456 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18283) );
  OAI22_X1 U21457 ( .A1(n18445), .A2(n18430), .B1(n13729), .B2(n18283), .ZN(
        n18288) );
  INV_X1 U21458 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n18286) );
  OAI22_X1 U21459 ( .A1(n9724), .A2(n18286), .B1(n18285), .B2(n18284), .ZN(
        n18287) );
  AOI211_X1 U21460 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A(
        n18288), .B(n18287), .ZN(n18290) );
  AOI22_X1 U21461 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18289) );
  OAI211_X1 U21462 ( .C1(n18455), .C2(n18291), .A(n18290), .B(n18289), .ZN(
        n18297) );
  AOI22_X1 U21463 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18295) );
  AOI22_X1 U21464 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18294) );
  AOI22_X1 U21465 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n18293) );
  AOI22_X1 U21466 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18292) );
  NAND4_X1 U21467 ( .A1(n18295), .A2(n18294), .A3(n18293), .A4(n18292), .ZN(
        n18296) );
  NOR2_X1 U21468 ( .A1(n18297), .A2(n18296), .ZN(n18579) );
  NOR2_X1 U21469 ( .A1(n18498), .A2(n18299), .ZN(n18315) );
  OAI222_X1 U21470 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n9734), .B1(
        P3_EBX_REG_17__SCAN_IN), .B2(n18299), .C1(n18315), .C2(n18298), .ZN(
        n18300) );
  OAI21_X1 U21471 ( .B1(n18579), .B2(n18484), .A(n18300), .ZN(P3_U2686) );
  INV_X1 U21472 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18308) );
  INV_X1 U21473 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n18442) );
  INV_X1 U21474 ( .A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18446) );
  OAI22_X1 U21475 ( .A1(n10739), .A2(n18442), .B1(n18301), .B2(n18446), .ZN(
        n18305) );
  INV_X1 U21476 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18302) );
  OAI22_X1 U21477 ( .A1(n9724), .A2(n18303), .B1(n13705), .B2(n18302), .ZN(
        n18304) );
  AOI211_X1 U21478 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n18305), .B(n18304), .ZN(n18307) );
  AOI22_X1 U21479 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18306) );
  OAI211_X1 U21480 ( .C1(n18455), .C2(n18308), .A(n18307), .B(n18306), .ZN(
        n18314) );
  AOI22_X1 U21481 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n18312) );
  AOI22_X1 U21482 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18311) );
  AOI22_X1 U21483 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18310) );
  AOI22_X1 U21484 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18309) );
  NAND4_X1 U21485 ( .A1(n18312), .A2(n18311), .A3(n18310), .A4(n18309), .ZN(
        n18313) );
  NOR2_X1 U21486 ( .A1(n18314), .A2(n18313), .ZN(n18585) );
  INV_X1 U21487 ( .A(n18337), .ZN(n18316) );
  OAI21_X1 U21488 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n18316), .A(n18315), .ZN(
        n18317) );
  OAI21_X1 U21489 ( .B1(n18585), .B2(n18484), .A(n18317), .ZN(P3_U2687) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18419), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18318) );
  OAI21_X1 U21491 ( .B1(n18319), .B2(n10740), .A(n18318), .ZN(n18320) );
  AOI21_X1 U21492 ( .B1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9717), .A(n18320), .ZN(n18323) );
  AOI22_X1 U21493 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18322) );
  AOI22_X1 U21494 ( .A1(n18193), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18321) );
  NAND3_X1 U21495 ( .A1(n18323), .A2(n18322), .A3(n18321), .ZN(n18336) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n13684), .B1(
        n18388), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18325) );
  NAND2_X1 U21497 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n18324) );
  OAI211_X1 U21498 ( .C1(n18326), .C2(n18402), .A(n18325), .B(n18324), .ZN(
        n18334) );
  OAI22_X1 U21499 ( .A1(n9712), .A2(n18328), .B1(n10739), .B2(n18327), .ZN(
        n18333) );
  INV_X1 U21500 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18331) );
  OAI22_X1 U21501 ( .A1(n18301), .A2(n18331), .B1(n18330), .B2(n18329), .ZN(
        n18332) );
  OR3_X1 U21502 ( .A1(n18334), .A2(n18333), .A3(n18332), .ZN(n18335) );
  NOR2_X1 U21503 ( .A1(n18336), .A2(n18335), .ZN(n18589) );
  OAI21_X1 U21504 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n18338), .A(n18337), .ZN(
        n18339) );
  AOI22_X1 U21505 ( .A1(n18498), .A2(n18589), .B1(n18339), .B2(n18484), .ZN(
        P3_U2688) );
  INV_X1 U21506 ( .A(n18376), .ZN(n18359) );
  INV_X1 U21507 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18348) );
  INV_X1 U21508 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n18341) );
  OAI22_X1 U21509 ( .A1(n18443), .A2(n18341), .B1(n13729), .B2(n18340), .ZN(
        n18345) );
  INV_X1 U21510 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18342) );
  OAI22_X1 U21511 ( .A1(n9724), .A2(n18343), .B1(n18445), .B2(n18342), .ZN(
        n18344) );
  AOI211_X1 U21512 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n18345), .B(n18344), .ZN(n18347) );
  AOI22_X1 U21513 ( .A1(n18450), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18346) );
  OAI211_X1 U21514 ( .C1(n18455), .C2(n18348), .A(n18347), .B(n18346), .ZN(
        n18354) );
  AOI22_X1 U21515 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17006), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n18352) );
  AOI22_X1 U21516 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n18351) );
  AOI22_X1 U21517 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18350) );
  AOI22_X1 U21518 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18349) );
  NAND4_X1 U21519 ( .A1(n18352), .A2(n18351), .A3(n18350), .A4(n18349), .ZN(
        n18353) );
  OR2_X1 U21520 ( .A1(n18354), .A2(n18353), .ZN(n18590) );
  NOR3_X1 U21521 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n18595), .A3(n18355), .ZN(
        n18356) );
  AOI21_X1 U21522 ( .B1(n18498), .B2(n18590), .A(n18356), .ZN(n18357) );
  OAI221_X1 U21523 ( .B1(n21674), .B2(n18359), .C1(n21674), .C2(n18358), .A(
        n18357), .ZN(P3_U2689) );
  AOI22_X1 U21524 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18360) );
  OAI21_X1 U21525 ( .B1(n18381), .B2(n18361), .A(n18360), .ZN(n18362) );
  AOI21_X1 U21526 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(n18362), .ZN(n18365) );
  AOI22_X1 U21527 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n18364) );
  AOI22_X1 U21528 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18363) );
  NAND3_X1 U21529 ( .A1(n18365), .A2(n18364), .A3(n18363), .ZN(n18373) );
  AOI22_X1 U21530 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n18366) );
  OAI21_X1 U21531 ( .B1(n10739), .B2(n18367), .A(n18366), .ZN(n18368) );
  AOI21_X1 U21532 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n18368), .ZN(n18371) );
  AOI22_X1 U21533 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18370) );
  AOI22_X1 U21534 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n18450), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n18369) );
  NAND3_X1 U21535 ( .A1(n18371), .A2(n18370), .A3(n18369), .ZN(n18372) );
  NOR2_X1 U21536 ( .A1(n18373), .A2(n18372), .ZN(n18601) );
  NOR3_X1 U21537 ( .A1(n18374), .A2(n18477), .A3(n18438), .ZN(n18441) );
  NAND2_X1 U21538 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n18441), .ZN(n18417) );
  NOR2_X1 U21539 ( .A1(n18375), .A2(n18417), .ZN(n18397) );
  OAI21_X1 U21540 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n18397), .A(n18376), .ZN(
        n18377) );
  OAI21_X1 U21541 ( .B1(n18601), .B2(n18484), .A(n18377), .ZN(P3_U2691) );
  OAI22_X1 U21542 ( .A1(n14490), .A2(n18379), .B1(n18402), .B2(n18378), .ZN(
        n18384) );
  OAI22_X1 U21543 ( .A1(n9724), .A2(n18382), .B1(n18381), .B2(n18380), .ZN(
        n18383) );
  AOI211_X1 U21544 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n18384), .B(n18383), .ZN(n18386) );
  AOI22_X1 U21545 ( .A1(n17006), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18450), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n18385) );
  OAI211_X1 U21546 ( .C1(n18455), .C2(n18387), .A(n18386), .B(n18385), .ZN(
        n18394) );
  AOI22_X1 U21547 ( .A1(n18388), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18451), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U21548 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n18391) );
  AOI22_X1 U21549 ( .A1(n18419), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18390) );
  AOI22_X1 U21550 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18389) );
  NAND4_X1 U21551 ( .A1(n18392), .A2(n18391), .A3(n18390), .A4(n18389), .ZN(
        n18393) );
  NOR2_X1 U21552 ( .A1(n18394), .A2(n18393), .ZN(n18605) );
  INV_X1 U21553 ( .A(n18417), .ZN(n18395) );
  OAI21_X1 U21554 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18395), .A(n18484), .ZN(
        n18396) );
  OAI22_X1 U21555 ( .A1(n18605), .A2(n18484), .B1(n18397), .B2(n18396), .ZN(
        P3_U2692) );
  AOI22_X1 U21556 ( .A1(n9738), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18399) );
  NAND2_X1 U21557 ( .A1(n18424), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n18398) );
  OAI211_X1 U21558 ( .C1(n18400), .C2(n10739), .A(n18399), .B(n18398), .ZN(
        n18408) );
  OAI22_X1 U21559 ( .A1(n14490), .A2(n18403), .B1(n18402), .B2(n18401), .ZN(
        n18407) );
  OAI22_X1 U21560 ( .A1(n18301), .A2(n18405), .B1(n10740), .B2(n18404), .ZN(
        n18406) );
  OR3_X1 U21561 ( .A1(n18408), .A2(n18407), .A3(n18406), .ZN(n18416) );
  INV_X1 U21562 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18410) );
  AOI22_X1 U21563 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n18409) );
  OAI21_X1 U21564 ( .B1(n13705), .B2(n18410), .A(n18409), .ZN(n18411) );
  AOI21_X1 U21565 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(n18411), .ZN(n18414) );
  AOI22_X1 U21566 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n18413) );
  AOI22_X1 U21567 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18412) );
  NAND3_X1 U21568 ( .A1(n18414), .A2(n18413), .A3(n18412), .ZN(n18415) );
  NOR2_X1 U21569 ( .A1(n18416), .A2(n18415), .ZN(n18611) );
  OAI21_X1 U21570 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n18441), .A(n18417), .ZN(
        n18418) );
  AOI22_X1 U21571 ( .A1(n18498), .A2(n18611), .B1(n18418), .B2(n18484), .ZN(
        P3_U2693) );
  AOI22_X1 U21572 ( .A1(n18420), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18419), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n18421) );
  OAI21_X1 U21573 ( .B1(n13705), .B2(n18422), .A(n18421), .ZN(n18423) );
  AOI21_X1 U21574 ( .B1(n18424), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n18423), .ZN(n18428) );
  AOI22_X1 U21575 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18427) );
  AOI22_X1 U21576 ( .A1(n18425), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18426) );
  NAND3_X1 U21577 ( .A1(n18428), .A2(n18427), .A3(n18426), .ZN(n18437) );
  AOI22_X1 U21578 ( .A1(n13684), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n18429) );
  OAI21_X1 U21579 ( .B1(n10740), .B2(n18430), .A(n18429), .ZN(n18431) );
  AOI21_X1 U21580 ( .B1(n9717), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(n18431), .ZN(n18435) );
  AOI22_X1 U21581 ( .A1(n18432), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17027), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18434) );
  AOI22_X1 U21582 ( .A1(n18269), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14578), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18433) );
  NAND3_X1 U21583 ( .A1(n18435), .A2(n18434), .A3(n18433), .ZN(n18436) );
  NOR2_X1 U21584 ( .A1(n18437), .A2(n18436), .ZN(n18616) );
  NOR2_X1 U21585 ( .A1(n18477), .A2(n18438), .ZN(n18439) );
  OAI21_X1 U21586 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n18439), .A(n18484), .ZN(
        n18440) );
  OAI22_X1 U21587 ( .A1(n18616), .A2(n18484), .B1(n18441), .B2(n18440), .ZN(
        P3_U2694) );
  INV_X1 U21588 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18454) );
  INV_X1 U21589 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18444) );
  OAI22_X1 U21590 ( .A1(n18445), .A2(n18444), .B1(n18443), .B2(n18442), .ZN(
        n18449) );
  INV_X1 U21591 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18447) );
  OAI22_X1 U21592 ( .A1(n9724), .A2(n18447), .B1(n13705), .B2(n18446), .ZN(
        n18448) );
  AOI211_X1 U21593 ( .C1(n9717), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n18449), .B(n18448), .ZN(n18453) );
  AOI22_X1 U21594 ( .A1(n18451), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n18450), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18452) );
  OAI211_X1 U21595 ( .C1(n18455), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        n18466) );
  AOI22_X1 U21596 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18456), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18464) );
  AOI22_X1 U21597 ( .A1(n17027), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14524), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18463) );
  AOI22_X1 U21598 ( .A1(n18458), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18457), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18462) );
  AOI22_X1 U21599 ( .A1(n18460), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18459), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18461) );
  NAND4_X1 U21600 ( .A1(n18464), .A2(n18463), .A3(n18462), .A4(n18461), .ZN(
        n18465) );
  NOR2_X1 U21601 ( .A1(n18466), .A2(n18465), .ZN(n18622) );
  INV_X1 U21602 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n18476) );
  NOR3_X1 U21603 ( .A1(n18476), .A2(n18478), .A3(n18477), .ZN(n18470) );
  NAND2_X1 U21604 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n18470), .ZN(n18469) );
  INV_X1 U21605 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n21833) );
  OAI21_X1 U21606 ( .B1(n18498), .B2(n21833), .A(n18469), .ZN(n18467) );
  OAI221_X1 U21607 ( .B1(n9734), .B2(n18469), .C1(n18469), .C2(n21833), .A(
        n18467), .ZN(n18468) );
  OAI21_X1 U21608 ( .B1(n18622), .B2(n18484), .A(n18468), .ZN(P3_U2695) );
  INV_X1 U21609 ( .A(n18469), .ZN(n18473) );
  AOI22_X1 U21610 ( .A1(n9734), .A2(n18470), .B1(P3_EBX_REG_7__SCAN_IN), .B2(
        n18484), .ZN(n18472) );
  OAI22_X1 U21611 ( .A1(n18473), .A2(n18472), .B1(n18471), .B2(n18484), .ZN(
        P3_U2696) );
  OAI21_X1 U21612 ( .B1(n18478), .B2(n18477), .A(n18484), .ZN(n18479) );
  NOR4_X1 U21613 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n18595), .A3(n18478), .A4(
        n18477), .ZN(n18474) );
  AOI21_X1 U21614 ( .B1(n18498), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n18474), .ZN(n18475) );
  OAI21_X1 U21615 ( .B1(n18476), .B2(n18479), .A(n18475), .ZN(P3_U2697) );
  AND2_X1 U21616 ( .A1(n18478), .A2(n18477), .ZN(n18480) );
  OAI22_X1 U21617 ( .A1(n18480), .A2(n18479), .B1(n14491), .B2(n18484), .ZN(
        P3_U2698) );
  NOR2_X1 U21618 ( .A1(n18481), .A2(n18495), .ZN(n18491) );
  NAND2_X1 U21619 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n18491), .ZN(n18488) );
  INV_X1 U21620 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18483) );
  NAND3_X1 U21621 ( .A1(n18488), .A2(P3_EBX_REG_4__SCAN_IN), .A3(n18484), .ZN(
        n18482) );
  OAI221_X1 U21622 ( .B1(n18488), .B2(P3_EBX_REG_4__SCAN_IN), .C1(n18484), 
        .C2(n18483), .A(n18482), .ZN(P3_U2699) );
  INV_X1 U21623 ( .A(n18491), .ZN(n18485) );
  OAI21_X1 U21624 ( .B1(n18486), .B2(n18498), .A(n18485), .ZN(n18487) );
  AOI22_X1 U21625 ( .A1(n18488), .A2(n18487), .B1(
        P3_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n18498), .ZN(n18489) );
  INV_X1 U21626 ( .A(n18489), .ZN(P3_U2700) );
  AOI221_X1 U21627 ( .B1(n18490), .B2(n9725), .C1(n18595), .C2(n9725), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n18492) );
  AOI211_X1 U21628 ( .C1(n18498), .C2(n18493), .A(n18492), .B(n18491), .ZN(
        P3_U2701) );
  INV_X1 U21629 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n21641) );
  OAI222_X1 U21630 ( .A1(n18496), .A2(n18495), .B1(n18494), .B2(n9725), .C1(
        n21641), .C2(n18484), .ZN(P3_U2702) );
  AOI22_X1 U21631 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18498), .B1(
        n18497), .B2(n18500), .ZN(n18499) );
  OAI21_X1 U21632 ( .B1(n9725), .B2(n18500), .A(n18499), .ZN(P3_U2703) );
  NAND2_X1 U21633 ( .A1(n18618), .A2(n18502), .ZN(n18551) );
  INV_X1 U21634 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18657) );
  INV_X1 U21635 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18721) );
  INV_X1 U21636 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18719) );
  NAND2_X1 U21637 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n18623) );
  NAND4_X1 U21638 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n18503) );
  NOR3_X1 U21639 ( .A1(n18504), .A2(n18623), .A3(n18503), .ZN(n18629) );
  INV_X1 U21640 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18741) );
  INV_X1 U21641 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18685) );
  INV_X1 U21642 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18743) );
  NOR2_X1 U21643 ( .A1(n18685), .A2(n18743), .ZN(n18600) );
  INV_X1 U21644 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18753) );
  NOR2_X2 U21645 ( .A1(n18596), .A2(n18753), .ZN(n18592) );
  INV_X1 U21646 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n21685) );
  INV_X1 U21647 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18669) );
  NAND2_X1 U21648 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18550), .ZN(n18545) );
  INV_X1 U21649 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18717) );
  NAND2_X1 U21650 ( .A1(n18544), .A2(n19383), .ZN(n18538) );
  NAND2_X1 U21651 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n18515), .ZN(n18514) );
  NOR2_X1 U21652 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n18514), .ZN(n18507) );
  NAND2_X1 U21653 ( .A1(n18643), .A2(n18514), .ZN(n18513) );
  OAI21_X1 U21654 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18505), .A(n18513), .ZN(
        n18506) );
  AOI22_X1 U21655 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18507), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18506), .ZN(n18508) );
  OAI21_X1 U21656 ( .B1(n21701), .B2(n18551), .A(n18508), .ZN(P3_U2704) );
  INV_X1 U21657 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18728) );
  NOR2_X2 U21658 ( .A1(n18509), .A2(n18643), .ZN(n18581) );
  OAI22_X1 U21659 ( .A1(n18510), .A2(n18645), .B1(n14713), .B2(n18551), .ZN(
        n18511) );
  AOI21_X1 U21660 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n18581), .A(n18511), .ZN(
        n18512) );
  OAI221_X1 U21661 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n18514), .C1(n18728), 
        .C2(n18513), .A(n18512), .ZN(P3_U2705) );
  AOI22_X1 U21662 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18580), .ZN(n18517) );
  OAI211_X1 U21663 ( .C1(n18515), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18643), .B(
        n18514), .ZN(n18516) );
  OAI211_X1 U21664 ( .C1(n18518), .C2(n18645), .A(n18517), .B(n18516), .ZN(
        P3_U2706) );
  AOI22_X1 U21665 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18581), .B1(n18625), .B2(
        n18519), .ZN(n18522) );
  OAI211_X1 U21666 ( .C1(n9805), .C2(P3_EAX_REG_28__SCAN_IN), .A(n18643), .B(
        n18520), .ZN(n18521) );
  OAI211_X1 U21667 ( .C1(n18551), .C2(n21768), .A(n18522), .B(n18521), .ZN(
        P3_U2707) );
  AOI22_X1 U21668 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18580), .ZN(n18525) );
  AOI211_X1 U21669 ( .C1(n18657), .C2(n18528), .A(n9805), .B(n18618), .ZN(
        n18523) );
  INV_X1 U21670 ( .A(n18523), .ZN(n18524) );
  OAI211_X1 U21671 ( .C1(n18526), .C2(n18645), .A(n18525), .B(n18524), .ZN(
        P3_U2708) );
  AOI22_X1 U21672 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18581), .B1(n18625), .B2(
        n18527), .ZN(n18530) );
  OAI211_X1 U21673 ( .C1(n18532), .C2(P3_EAX_REG_26__SCAN_IN), .A(n18643), .B(
        n18528), .ZN(n18529) );
  OAI211_X1 U21674 ( .C1(n18551), .C2(n18531), .A(n18530), .B(n18529), .ZN(
        P3_U2709) );
  AOI22_X1 U21675 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18580), .ZN(n18535) );
  AOI211_X1 U21676 ( .C1(n18721), .C2(n18539), .A(n18532), .B(n18618), .ZN(
        n18533) );
  INV_X1 U21677 ( .A(n18533), .ZN(n18534) );
  OAI211_X1 U21678 ( .C1(n18536), .C2(n18645), .A(n18535), .B(n18534), .ZN(
        P3_U2710) );
  AOI22_X1 U21679 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18581), .B1(n18625), .B2(
        n18537), .ZN(n18542) );
  OAI21_X1 U21680 ( .B1(n18719), .B2(n18618), .A(n18538), .ZN(n18540) );
  NAND2_X1 U21681 ( .A1(n18540), .A2(n18539), .ZN(n18541) );
  OAI211_X1 U21682 ( .C1(n18551), .C2(n18543), .A(n18542), .B(n18541), .ZN(
        P3_U2711) );
  AOI211_X1 U21683 ( .C1(n18717), .C2(n18545), .A(n18618), .B(n18544), .ZN(
        n18546) );
  AOI21_X1 U21684 ( .B1(n18580), .B2(BUF2_REG_23__SCAN_IN), .A(n18546), .ZN(
        n18548) );
  NAND2_X1 U21685 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18581), .ZN(n18547) );
  OAI211_X1 U21686 ( .C1(n18549), .C2(n18645), .A(n18548), .B(n18547), .ZN(
        P3_U2712) );
  NAND2_X1 U21687 ( .A1(n19383), .A2(n18550), .ZN(n18557) );
  NAND2_X1 U21688 ( .A1(n18557), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n18555) );
  OAI22_X1 U21689 ( .A1(n18552), .A2(n18645), .B1(n21654), .B2(n18551), .ZN(
        n18553) );
  AOI21_X1 U21690 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n18581), .A(n18553), .ZN(
        n18554) );
  OAI221_X1 U21691 ( .B1(n18557), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n18555), 
        .C2(n18618), .A(n18554), .ZN(P3_U2713) );
  AOI22_X1 U21692 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n18580), .ZN(n18559) );
  INV_X1 U21693 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18667) );
  NAND2_X1 U21694 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .ZN(n18556) );
  NOR2_X1 U21695 ( .A1(n18582), .A2(n18556), .ZN(n18570) );
  NAND2_X1 U21696 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18570), .ZN(n18566) );
  NOR2_X1 U21697 ( .A1(n18667), .A2(n18566), .ZN(n18561) );
  OAI211_X1 U21698 ( .C1(n18561), .C2(P3_EAX_REG_21__SCAN_IN), .A(n18643), .B(
        n18557), .ZN(n18558) );
  OAI211_X1 U21699 ( .C1(n18560), .C2(n18645), .A(n18559), .B(n18558), .ZN(
        P3_U2714) );
  AOI22_X1 U21700 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n18580), .ZN(n18564) );
  AOI211_X1 U21701 ( .C1(n18667), .C2(n18566), .A(n18561), .B(n18618), .ZN(
        n18562) );
  INV_X1 U21702 ( .A(n18562), .ZN(n18563) );
  OAI211_X1 U21703 ( .C1(n18565), .C2(n18645), .A(n18564), .B(n18563), .ZN(
        P3_U2715) );
  AOI22_X1 U21704 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18580), .ZN(n18568) );
  OAI211_X1 U21705 ( .C1(n18570), .C2(P3_EAX_REG_19__SCAN_IN), .A(n18643), .B(
        n18566), .ZN(n18567) );
  OAI211_X1 U21706 ( .C1(n18569), .C2(n18645), .A(n18568), .B(n18567), .ZN(
        P3_U2716) );
  AOI22_X1 U21707 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n18580), .ZN(n18573) );
  INV_X1 U21708 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n21733) );
  INV_X1 U21709 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18710) );
  OR2_X1 U21710 ( .A1(n18710), .A2(n18582), .ZN(n18575) );
  AOI211_X1 U21711 ( .C1(n21733), .C2(n18575), .A(n18570), .B(n18618), .ZN(
        n18571) );
  INV_X1 U21712 ( .A(n18571), .ZN(n18572) );
  OAI211_X1 U21713 ( .C1(n18574), .C2(n18645), .A(n18573), .B(n18572), .ZN(
        P3_U2717) );
  AOI22_X1 U21714 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18580), .ZN(n18578) );
  INV_X1 U21715 ( .A(n18582), .ZN(n18576) );
  OAI211_X1 U21716 ( .C1(n18576), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18643), .B(
        n18575), .ZN(n18577) );
  OAI211_X1 U21717 ( .C1(n18579), .C2(n18645), .A(n18578), .B(n18577), .ZN(
        P3_U2718) );
  AOI22_X1 U21718 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18581), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18580), .ZN(n18584) );
  OAI211_X1 U21719 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18586), .A(n18643), .B(
        n18582), .ZN(n18583) );
  OAI211_X1 U21720 ( .C1(n18585), .C2(n18645), .A(n18584), .B(n18583), .ZN(
        P3_U2719) );
  AOI211_X1 U21721 ( .C1(n21685), .C2(n18591), .A(n18618), .B(n18586), .ZN(
        n18587) );
  AOI21_X1 U21722 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n18626), .A(n18587), .ZN(
        n18588) );
  OAI21_X1 U21723 ( .B1(n18589), .B2(n18645), .A(n18588), .ZN(P3_U2720) );
  AOI22_X1 U21724 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18626), .B1(n18625), .B2(
        n18590), .ZN(n18594) );
  OAI211_X1 U21725 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n18592), .A(n18643), .B(
        n18591), .ZN(n18593) );
  NAND2_X1 U21726 ( .A1(n18594), .A2(n18593), .ZN(P3_U2721) );
  NOR2_X1 U21727 ( .A1(n18595), .A2(n18596), .ZN(n18603) );
  AOI22_X1 U21728 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18626), .B1(n18603), .B2(
        n18753), .ZN(n18598) );
  NAND3_X1 U21729 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18643), .A3(n18596), 
        .ZN(n18597) );
  OAI211_X1 U21730 ( .C1(n18599), .C2(n18645), .A(n18598), .B(n18597), .ZN(
        P3_U2722) );
  INV_X1 U21731 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18683) );
  NAND3_X1 U21732 ( .A1(n9734), .A2(n18617), .A3(n18600), .ZN(n18604) );
  NOR2_X1 U21733 ( .A1(n18683), .A2(n18604), .ZN(n18607) );
  AOI21_X1 U21734 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18643), .A(n18607), .ZN(
        n18602) );
  OAI222_X1 U21735 ( .A1(n18648), .A2(n18751), .B1(n18603), .B2(n18602), .C1(
        n18632), .C2(n18601), .ZN(P3_U2723) );
  INV_X1 U21736 ( .A(n18604), .ZN(n18608) );
  AOI21_X1 U21737 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18643), .A(n18608), .ZN(
        n18606) );
  OAI222_X1 U21738 ( .A1(n18648), .A2(n18747), .B1(n18607), .B2(n18606), .C1(
        n18632), .C2(n18605), .ZN(P3_U2724) );
  NAND2_X1 U21739 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n18617), .ZN(n18614) );
  AOI211_X1 U21740 ( .C1(n18685), .C2(n18614), .A(n18618), .B(n18608), .ZN(
        n18609) );
  AOI21_X1 U21741 ( .B1(n18626), .B2(BUF2_REG_10__SCAN_IN), .A(n18609), .ZN(
        n18610) );
  OAI21_X1 U21742 ( .B1(n18611), .B2(n18645), .A(n18610), .ZN(P3_U2725) );
  NAND2_X1 U21743 ( .A1(n9734), .A2(n18617), .ZN(n18612) );
  OAI21_X1 U21744 ( .B1(n18618), .B2(n18743), .A(n18612), .ZN(n18613) );
  AOI22_X1 U21745 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18626), .B1(n18614), .B2(
        n18613), .ZN(n18615) );
  OAI21_X1 U21746 ( .B1(n18616), .B2(n18645), .A(n18615), .ZN(P3_U2726) );
  AOI211_X1 U21747 ( .C1(n18741), .C2(n18619), .A(n18618), .B(n18617), .ZN(
        n18620) );
  AOI21_X1 U21748 ( .B1(n18626), .B2(BUF2_REG_8__SCAN_IN), .A(n18620), .ZN(
        n18621) );
  OAI21_X1 U21749 ( .B1(n18622), .B2(n18645), .A(n18621), .ZN(P3_U2727) );
  NAND2_X1 U21750 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18642), .ZN(n18638) );
  NOR2_X1 U21751 ( .A1(n18623), .A2(n18638), .ZN(n18637) );
  AOI22_X1 U21752 ( .A1(n18637), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n18643), .ZN(n18630) );
  AOI22_X1 U21753 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18626), .B1(n18625), .B2(
        n18624), .ZN(n18627) );
  OAI221_X1 U21754 ( .B1(n18630), .B2(n18629), .C1(n18630), .C2(n18628), .A(
        n18627), .ZN(P3_U2728) );
  AOI21_X1 U21755 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n18643), .A(n18637), .ZN(
        n18634) );
  AND2_X1 U21756 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18637), .ZN(n18633) );
  OAI222_X1 U21757 ( .A1(n18648), .A2(n19376), .B1(n18634), .B2(n18633), .C1(
        n18632), .C2(n18631), .ZN(P3_U2729) );
  INV_X1 U21758 ( .A(n18638), .ZN(n18647) );
  AOI22_X1 U21759 ( .A1(n18647), .A2(P3_EAX_REG_4__SCAN_IN), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n18643), .ZN(n18636) );
  OAI222_X1 U21760 ( .A1(n19372), .A2(n18648), .B1(n18637), .B2(n18636), .C1(
        n18645), .C2(n18635), .ZN(P3_U2730) );
  INV_X1 U21761 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18693) );
  NOR2_X1 U21762 ( .A1(n18693), .A2(n18638), .ZN(n18641) );
  AOI21_X1 U21763 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18643), .A(n18647), .ZN(
        n18640) );
  OAI222_X1 U21764 ( .A1(n19368), .A2(n18648), .B1(n18641), .B2(n18640), .C1(
        n18645), .C2(n18639), .ZN(P3_U2731) );
  AOI21_X1 U21765 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18643), .A(n18642), .ZN(
        n18646) );
  OAI222_X1 U21766 ( .A1(n19364), .A2(n18648), .B1(n18647), .B2(n18646), .C1(
        n18645), .C2(n18644), .ZN(P3_U2732) );
  NOR2_X2 U21767 ( .A1(n18649), .A2(n18892), .ZN(n19940) );
  NOR2_X4 U21768 ( .A1(n19940), .A2(n18676), .ZN(n18672) );
  AND2_X1 U21769 ( .A1(n18672), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U21770 ( .A1(n18676), .A2(n18651), .ZN(n18674) );
  AOI22_X1 U21771 ( .A1(n19940), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n18672), .ZN(n18652) );
  OAI21_X1 U21772 ( .B1(n18728), .B2(n18674), .A(n18652), .ZN(P3_U2737) );
  INV_X1 U21773 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18726) );
  AOI22_X1 U21774 ( .A1(n19940), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18653) );
  OAI21_X1 U21775 ( .B1(n18726), .B2(n18674), .A(n18653), .ZN(P3_U2738) );
  INV_X1 U21776 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18655) );
  AOI22_X1 U21777 ( .A1(n19940), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18654) );
  OAI21_X1 U21778 ( .B1(n18655), .B2(n18674), .A(n18654), .ZN(P3_U2739) );
  AOI22_X1 U21779 ( .A1(n19940), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18656) );
  OAI21_X1 U21780 ( .B1(n18657), .B2(n18674), .A(n18656), .ZN(P3_U2740) );
  AOI22_X1 U21781 ( .A1(n19940), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18658) );
  OAI21_X1 U21782 ( .B1(n10423), .B2(n18674), .A(n18658), .ZN(P3_U2741) );
  AOI22_X1 U21783 ( .A1(n19940), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18659) );
  OAI21_X1 U21784 ( .B1(n18721), .B2(n18674), .A(n18659), .ZN(P3_U2742) );
  AOI22_X1 U21785 ( .A1(n19940), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18660) );
  OAI21_X1 U21786 ( .B1(n18719), .B2(n18674), .A(n18660), .ZN(P3_U2743) );
  CLKBUF_X1 U21787 ( .A(n19940), .Z(n18699) );
  AOI22_X1 U21788 ( .A1(n18699), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18661) );
  OAI21_X1 U21789 ( .B1(n18717), .B2(n18674), .A(n18661), .ZN(P3_U2744) );
  INV_X1 U21790 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18663) );
  AOI22_X1 U21791 ( .A1(n18699), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18662) );
  OAI21_X1 U21792 ( .B1(n18663), .B2(n18674), .A(n18662), .ZN(P3_U2745) );
  INV_X1 U21793 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18665) );
  AOI22_X1 U21794 ( .A1(n18699), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18664) );
  OAI21_X1 U21795 ( .B1(n18665), .B2(n18674), .A(n18664), .ZN(P3_U2746) );
  AOI22_X1 U21796 ( .A1(n18699), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18666) );
  OAI21_X1 U21797 ( .B1(n18667), .B2(n18674), .A(n18666), .ZN(P3_U2747) );
  AOI22_X1 U21798 ( .A1(n18699), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18668) );
  OAI21_X1 U21799 ( .B1(n18669), .B2(n18674), .A(n18668), .ZN(P3_U2748) );
  AOI22_X1 U21800 ( .A1(n18699), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18670) );
  OAI21_X1 U21801 ( .B1(n21733), .B2(n18674), .A(n18670), .ZN(P3_U2749) );
  AOI22_X1 U21802 ( .A1(n18699), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18671) );
  OAI21_X1 U21803 ( .B1(n18710), .B2(n18674), .A(n18671), .ZN(P3_U2750) );
  INV_X1 U21804 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18675) );
  AOI22_X1 U21805 ( .A1(n18699), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18673) );
  OAI21_X1 U21806 ( .B1(n18675), .B2(n18674), .A(n18673), .ZN(P3_U2751) );
  AOI22_X1 U21807 ( .A1(n18699), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18677) );
  OAI21_X1 U21808 ( .B1(n21685), .B2(n18701), .A(n18677), .ZN(P3_U2752) );
  AOI22_X1 U21809 ( .A1(n18699), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18678) );
  OAI21_X1 U21810 ( .B1(n10425), .B2(n18701), .A(n18678), .ZN(P3_U2753) );
  AOI22_X1 U21811 ( .A1(n18699), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18679) );
  OAI21_X1 U21812 ( .B1(n18753), .B2(n18701), .A(n18679), .ZN(P3_U2754) );
  INV_X1 U21813 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18681) );
  AOI22_X1 U21814 ( .A1(n18699), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18680) );
  OAI21_X1 U21815 ( .B1(n18681), .B2(n18701), .A(n18680), .ZN(P3_U2755) );
  AOI22_X1 U21816 ( .A1(n18699), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18682) );
  OAI21_X1 U21817 ( .B1(n18683), .B2(n18701), .A(n18682), .ZN(P3_U2756) );
  AOI22_X1 U21818 ( .A1(n18699), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18684) );
  OAI21_X1 U21819 ( .B1(n18685), .B2(n18701), .A(n18684), .ZN(P3_U2757) );
  AOI22_X1 U21820 ( .A1(n18699), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18686) );
  OAI21_X1 U21821 ( .B1(n18743), .B2(n18701), .A(n18686), .ZN(P3_U2758) );
  AOI22_X1 U21822 ( .A1(n18699), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18687) );
  OAI21_X1 U21823 ( .B1(n18741), .B2(n18701), .A(n18687), .ZN(P3_U2759) );
  INV_X1 U21824 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18739) );
  AOI22_X1 U21825 ( .A1(n18699), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18688) );
  OAI21_X1 U21826 ( .B1(n18739), .B2(n18701), .A(n18688), .ZN(P3_U2760) );
  INV_X1 U21827 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18690) );
  AOI22_X1 U21828 ( .A1(n18699), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18689) );
  OAI21_X1 U21829 ( .B1(n18690), .B2(n18701), .A(n18689), .ZN(P3_U2761) );
  INV_X1 U21830 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21793) );
  AOI22_X1 U21831 ( .A1(n18699), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18691) );
  OAI21_X1 U21832 ( .B1(n21793), .B2(n18701), .A(n18691), .ZN(P3_U2762) );
  AOI22_X1 U21833 ( .A1(n18699), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18692) );
  OAI21_X1 U21834 ( .B1(n18693), .B2(n18701), .A(n18692), .ZN(P3_U2763) );
  INV_X1 U21835 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18695) );
  AOI22_X1 U21836 ( .A1(n18699), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18694) );
  OAI21_X1 U21837 ( .B1(n18695), .B2(n18701), .A(n18694), .ZN(P3_U2764) );
  AOI22_X1 U21838 ( .A1(n18699), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18696) );
  OAI21_X1 U21839 ( .B1(n18697), .B2(n18701), .A(n18696), .ZN(P3_U2765) );
  INV_X1 U21840 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18731) );
  AOI22_X1 U21841 ( .A1(n18699), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18698) );
  OAI21_X1 U21842 ( .B1(n18731), .B2(n18701), .A(n18698), .ZN(P3_U2766) );
  INV_X1 U21843 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18702) );
  AOI22_X1 U21844 ( .A1(n18699), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18672), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18700) );
  OAI21_X1 U21845 ( .B1(n18702), .B2(n18701), .A(n18700), .ZN(P3_U2767) );
  INV_X1 U21846 ( .A(n18705), .ZN(n18703) );
  NOR3_X4 U21847 ( .A1(n18707), .A2(n18706), .A3(n18705), .ZN(n18748) );
  AOI22_X1 U21848 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18755), .ZN(n18708) );
  OAI21_X1 U21849 ( .B1(n19349), .B2(n18750), .A(n18708), .ZN(P3_U2768) );
  INV_X1 U21850 ( .A(n18748), .ZN(n18758) );
  AOI22_X1 U21851 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18755), .ZN(n18709) );
  OAI21_X1 U21852 ( .B1(n18710), .B2(n18758), .A(n18709), .ZN(P3_U2769) );
  AOI22_X1 U21853 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18755), .ZN(n18711) );
  OAI21_X1 U21854 ( .B1(n19361), .B2(n18750), .A(n18711), .ZN(P3_U2770) );
  AOI22_X1 U21855 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18755), .ZN(n18712) );
  OAI21_X1 U21856 ( .B1(n19364), .B2(n18750), .A(n18712), .ZN(P3_U2771) );
  AOI22_X1 U21857 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18755), .ZN(n18713) );
  OAI21_X1 U21858 ( .B1(n19368), .B2(n18750), .A(n18713), .ZN(P3_U2772) );
  AOI22_X1 U21859 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18755), .ZN(n18714) );
  OAI21_X1 U21860 ( .B1(n19372), .B2(n18750), .A(n18714), .ZN(P3_U2773) );
  AOI22_X1 U21861 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18755), .ZN(n18715) );
  OAI21_X1 U21862 ( .B1(n19376), .B2(n18750), .A(n18715), .ZN(P3_U2774) );
  AOI22_X1 U21863 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18755), .ZN(n18716) );
  OAI21_X1 U21864 ( .B1(n18717), .B2(n18758), .A(n18716), .ZN(P3_U2775) );
  AOI22_X1 U21865 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18755), .ZN(n18718) );
  OAI21_X1 U21866 ( .B1(n18719), .B2(n18758), .A(n18718), .ZN(P3_U2776) );
  AOI22_X1 U21867 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18755), .ZN(n18720) );
  OAI21_X1 U21868 ( .B1(n18721), .B2(n18758), .A(n18720), .ZN(P3_U2777) );
  AOI22_X1 U21869 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18755), .ZN(n18722) );
  OAI21_X1 U21870 ( .B1(n18745), .B2(n18750), .A(n18722), .ZN(P3_U2778) );
  AOI22_X1 U21871 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18734), .ZN(n18723) );
  OAI21_X1 U21872 ( .B1(n18747), .B2(n18750), .A(n18723), .ZN(P3_U2779) );
  AOI22_X1 U21873 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n18748), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18734), .ZN(n18724) );
  OAI21_X1 U21874 ( .B1(n18751), .B2(n18750), .A(n18724), .ZN(P3_U2780) );
  AOI22_X1 U21875 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18734), .ZN(n18725) );
  OAI21_X1 U21876 ( .B1(n18726), .B2(n18758), .A(n18725), .ZN(P3_U2781) );
  AOI22_X1 U21877 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18756), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18734), .ZN(n18727) );
  OAI21_X1 U21878 ( .B1(n18728), .B2(n18758), .A(n18727), .ZN(P3_U2782) );
  AOI22_X1 U21879 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18734), .ZN(n18729) );
  OAI21_X1 U21880 ( .B1(n19349), .B2(n18750), .A(n18729), .ZN(P3_U2783) );
  AOI22_X1 U21881 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18734), .ZN(n18730) );
  OAI21_X1 U21882 ( .B1(n18731), .B2(n18758), .A(n18730), .ZN(P3_U2784) );
  AOI22_X1 U21883 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18734), .ZN(n18732) );
  OAI21_X1 U21884 ( .B1(n19361), .B2(n18750), .A(n18732), .ZN(P3_U2785) );
  AOI22_X1 U21885 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18734), .ZN(n18733) );
  OAI21_X1 U21886 ( .B1(n19364), .B2(n18750), .A(n18733), .ZN(P3_U2786) );
  AOI22_X1 U21887 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18734), .ZN(n18735) );
  OAI21_X1 U21888 ( .B1(n19368), .B2(n18750), .A(n18735), .ZN(P3_U2787) );
  AOI22_X1 U21889 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18755), .ZN(n18736) );
  OAI21_X1 U21890 ( .B1(n19372), .B2(n18750), .A(n18736), .ZN(P3_U2788) );
  AOI22_X1 U21891 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18755), .ZN(n18737) );
  OAI21_X1 U21892 ( .B1(n19376), .B2(n18750), .A(n18737), .ZN(P3_U2789) );
  AOI22_X1 U21893 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18755), .ZN(n18738) );
  OAI21_X1 U21894 ( .B1(n18739), .B2(n18758), .A(n18738), .ZN(P3_U2790) );
  AOI22_X1 U21895 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18755), .ZN(n18740) );
  OAI21_X1 U21896 ( .B1(n18741), .B2(n18758), .A(n18740), .ZN(P3_U2791) );
  AOI22_X1 U21897 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18755), .ZN(n18742) );
  OAI21_X1 U21898 ( .B1(n18743), .B2(n18758), .A(n18742), .ZN(P3_U2792) );
  AOI22_X1 U21899 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18755), .ZN(n18744) );
  OAI21_X1 U21900 ( .B1(n18745), .B2(n18750), .A(n18744), .ZN(P3_U2793) );
  AOI22_X1 U21901 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18755), .ZN(n18746) );
  OAI21_X1 U21902 ( .B1(n18747), .B2(n18750), .A(n18746), .ZN(P3_U2794) );
  AOI22_X1 U21903 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18748), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18755), .ZN(n18749) );
  OAI21_X1 U21904 ( .B1(n18751), .B2(n18750), .A(n18749), .ZN(P3_U2795) );
  AOI22_X1 U21905 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18755), .ZN(n18752) );
  OAI21_X1 U21906 ( .B1(n18753), .B2(n18758), .A(n18752), .ZN(P3_U2796) );
  AOI22_X1 U21907 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18755), .ZN(n18754) );
  OAI21_X1 U21908 ( .B1(n10425), .B2(n18758), .A(n18754), .ZN(P3_U2797) );
  AOI22_X1 U21909 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18756), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18755), .ZN(n18757) );
  OAI21_X1 U21910 ( .B1(n21685), .B2(n18758), .A(n18757), .ZN(P3_U2798) );
  XNOR2_X1 U21911 ( .A(n18783), .B(n19070), .ZN(n18761) );
  NOR2_X1 U21912 ( .A1(n18759), .A2(n19070), .ZN(n18760) );
  MUX2_X1 U21913 ( .A(n18761), .B(n18760), .S(n18910), .Z(n18762) );
  INV_X1 U21914 ( .A(n18762), .ZN(n18763) );
  OAI21_X1 U21915 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n18764), .A(
        n18763), .ZN(n19064) );
  OAI21_X1 U21916 ( .B1(n18765), .B2(n18892), .A(n9716), .ZN(n18766) );
  AOI21_X1 U21917 ( .B1(n19730), .B2(n17733), .A(n18766), .ZN(n18805) );
  OAI21_X1 U21918 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18892), .A(
        n18805), .ZN(n18779) );
  NOR2_X1 U21919 ( .A1(n18896), .A2(n17733), .ZN(n18781) );
  OAI211_X1 U21920 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n18781), .B(n18767), .ZN(n18768) );
  NAND2_X1 U21921 ( .A1(n19268), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n19068) );
  OAI211_X1 U21922 ( .C1(n18937), .C2(n18769), .A(n18768), .B(n19068), .ZN(
        n18770) );
  AOI21_X1 U21923 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18779), .A(
        n18770), .ZN(n18777) );
  AOI21_X1 U21924 ( .B1(n19070), .B2(n18772), .A(n18771), .ZN(n19067) );
  INV_X1 U21925 ( .A(n18773), .ZN(n18775) );
  AOI22_X1 U21926 ( .A1(n18775), .A2(n19071), .B1(n19070), .B2(n18774), .ZN(
        n19063) );
  AOI22_X1 U21927 ( .A1(n18934), .A2(n19067), .B1(n19048), .B2(n19063), .ZN(
        n18776) );
  OAI211_X1 U21928 ( .C1(n18966), .C2(n19064), .A(n18777), .B(n18776), .ZN(
        P3_U2805) );
  INV_X1 U21929 ( .A(n18778), .ZN(n18790) );
  NOR2_X1 U21930 ( .A1(n19156), .A2(n19896), .ZN(n19082) );
  AOI221_X1 U21931 ( .B1(n18781), .B2(n18780), .C1(n18779), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n19082), .ZN(n18789) );
  NOR2_X1 U21932 ( .A1(n18799), .A2(n18798), .ZN(n18787) );
  NAND2_X1 U21933 ( .A1(n19048), .A2(n19171), .ZN(n18921) );
  NAND2_X1 U21934 ( .A1(n18934), .A2(n19170), .ZN(n18912) );
  NAND2_X1 U21935 ( .A1(n18921), .A2(n18912), .ZN(n18902) );
  AOI21_X1 U21936 ( .B1(n18901), .B2(n18782), .A(n18902), .ZN(n18797) );
  INV_X1 U21937 ( .A(n18783), .ZN(n18784) );
  AOI21_X1 U21938 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n18785), .A(
        n18784), .ZN(n19078) );
  OAI22_X1 U21939 ( .A1(n18797), .A2(n10061), .B1(n19078), .B2(n18966), .ZN(
        n18786) );
  AOI21_X1 U21940 ( .B1(n18787), .B2(n10061), .A(n18786), .ZN(n18788) );
  OAI211_X1 U21941 ( .C1(n18937), .C2(n18790), .A(n18789), .B(n18788), .ZN(
        P3_U2806) );
  AOI22_X1 U21942 ( .A1(n19268), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18858), 
        .B2(n18791), .ZN(n18803) );
  INV_X1 U21943 ( .A(n18806), .ZN(n18794) );
  NAND2_X1 U21944 ( .A1(n18830), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18793) );
  OAI211_X1 U21945 ( .C1(n18795), .C2(n18794), .A(n18792), .B(n18793), .ZN(
        n18796) );
  XNOR2_X1 U21946 ( .A(n18796), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n19084) );
  NAND2_X1 U21947 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18815) );
  NAND2_X1 U21948 ( .A1(n18814), .A2(n18855), .ZN(n18829) );
  NOR3_X1 U21949 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18815), .A3(
        n18829), .ZN(n18801) );
  AOI21_X1 U21950 ( .B1(n18799), .B2(n18798), .A(n18797), .ZN(n18800) );
  AOI211_X1 U21951 ( .C1(n18946), .C2(n19084), .A(n18801), .B(n18800), .ZN(
        n18802) );
  OAI211_X1 U21952 ( .C1(n18805), .C2(n18804), .A(n18803), .B(n18802), .ZN(
        P3_U2807) );
  INV_X1 U21953 ( .A(n18818), .ZN(n19088) );
  OAI21_X1 U21954 ( .B1(n18831), .B2(n19088), .A(n18806), .ZN(n18807) );
  NAND2_X1 U21955 ( .A1(n18792), .A2(n18807), .ZN(n18808) );
  XNOR2_X1 U21956 ( .A(n18808), .B(n19089), .ZN(n19104) );
  NAND2_X1 U21957 ( .A1(n18811), .A2(n18810), .ZN(n18812) );
  OAI211_X1 U21958 ( .C1(n18814), .C2(n18813), .A(n9716), .B(n18812), .ZN(
        n18846) );
  AOI21_X1 U21959 ( .B1(n17216), .B2(n18843), .A(n18846), .ZN(n18827) );
  NAND2_X1 U21960 ( .A1(n19268), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n19102) );
  INV_X1 U21961 ( .A(n18829), .ZN(n18816) );
  OAI211_X1 U21962 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18816), .B(n18815), .ZN(n18817) );
  OAI211_X1 U21963 ( .C1(n18827), .C2(n21722), .A(n19102), .B(n18817), .ZN(
        n18824) );
  INV_X1 U21964 ( .A(n18901), .ZN(n18819) );
  NAND2_X1 U21965 ( .A1(n19108), .A2(n18818), .ZN(n19092) );
  NOR2_X1 U21966 ( .A1(n18819), .A2(n19092), .ZN(n18822) );
  NAND2_X1 U21967 ( .A1(n18820), .A2(n19040), .ZN(n18840) );
  AOI21_X1 U21968 ( .B1(n18840), .B2(n19092), .A(n18902), .ZN(n18839) );
  INV_X1 U21969 ( .A(n18839), .ZN(n18821) );
  MUX2_X1 U21970 ( .A(n18822), .B(n18821), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n18823) );
  AOI211_X1 U21971 ( .C1(n18858), .C2(n18825), .A(n18824), .B(n18823), .ZN(
        n18826) );
  OAI21_X1 U21972 ( .B1(n18966), .B2(n19104), .A(n18826), .ZN(P3_U2808) );
  NAND2_X1 U21973 ( .A1(n19268), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n19118) );
  OAI221_X1 U21974 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n18829), .C1(
        n18828), .C2(n18827), .A(n19118), .ZN(n18836) );
  INV_X1 U21975 ( .A(n18873), .ZN(n18852) );
  INV_X1 U21976 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19105) );
  OR3_X1 U21977 ( .A1(n18831), .A2(n19105), .A3(n18830), .ZN(n18853) );
  INV_X1 U21978 ( .A(n18853), .ZN(n18832) );
  AOI22_X1 U21979 ( .A1(n18852), .A2(n18833), .B1(n19095), .B2(n18832), .ZN(
        n18834) );
  XNOR2_X1 U21980 ( .A(n18834), .B(n19114), .ZN(n19120) );
  NAND2_X1 U21981 ( .A1(n19095), .A2(n19114), .ZN(n19107) );
  NAND3_X1 U21982 ( .A1(n19108), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n18901), .ZN(n18864) );
  OAI22_X1 U21983 ( .A1(n19120), .A2(n18966), .B1(n19107), .B2(n18864), .ZN(
        n18835) );
  AOI211_X1 U21984 ( .C1(n18858), .C2(n18837), .A(n18836), .B(n18835), .ZN(
        n18838) );
  OAI21_X1 U21985 ( .B1(n18839), .B2(n19114), .A(n18838), .ZN(P3_U2809) );
  NAND3_X1 U21986 ( .A1(n19108), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n19124) );
  AOI21_X1 U21987 ( .B1(n18840), .B2(n19124), .A(n18902), .ZN(n18863) );
  INV_X1 U21988 ( .A(n18864), .ZN(n18850) );
  NOR2_X1 U21989 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19136), .ZN(
        n19126) );
  NAND2_X1 U21990 ( .A1(n18853), .A2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18841) );
  OAI211_X1 U21991 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18871), .A(
        n18792), .B(n18841), .ZN(n18842) );
  XNOR2_X1 U21992 ( .A(n18842), .B(n19093), .ZN(n19130) );
  OAI21_X1 U21993 ( .B1(n18844), .B2(n19690), .A(n18843), .ZN(n18845) );
  AOI22_X1 U21994 ( .A1(n18847), .A2(n19043), .B1(n18846), .B2(n18845), .ZN(
        n18848) );
  NAND2_X1 U21995 ( .A1(n19268), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n19128) );
  OAI211_X1 U21996 ( .C1(n18966), .C2(n19130), .A(n18848), .B(n19128), .ZN(
        n18849) );
  AOI21_X1 U21997 ( .B1(n18850), .B2(n19126), .A(n18849), .ZN(n18851) );
  OAI21_X1 U21998 ( .B1(n18863), .B2(n19093), .A(n18851), .ZN(P3_U2810) );
  NAND2_X1 U21999 ( .A1(n18852), .A2(n18871), .ZN(n18876) );
  NAND2_X1 U22000 ( .A1(n18876), .A2(n18853), .ZN(n18854) );
  XOR2_X1 U22001 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n18854), .Z(
        n19132) );
  OAI211_X1 U22002 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n9908), .B(n18855), .ZN(n18860)
         );
  INV_X1 U22003 ( .A(n9908), .ZN(n18865) );
  AOI21_X1 U22004 ( .B1(n19008), .B2(n18865), .A(n19006), .ZN(n18880) );
  OAI21_X1 U22005 ( .B1(n18856), .B2(n18892), .A(n18880), .ZN(n18868) );
  AOI22_X1 U22006 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18868), .B1(
        n18858), .B2(n18857), .ZN(n18859) );
  NAND2_X1 U22007 ( .A1(n19268), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n19133) );
  OAI211_X1 U22008 ( .C1(n10730), .C2(n18860), .A(n18859), .B(n19133), .ZN(
        n18861) );
  AOI21_X1 U22009 ( .B1(n18946), .B2(n19132), .A(n18861), .ZN(n18862) );
  OAI221_X1 U22010 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18864), 
        .C1(n19136), .C2(n18863), .A(n18862), .ZN(P3_U2811) );
  AOI21_X1 U22011 ( .B1(n18901), .B2(n19140), .A(n18902), .ZN(n18887) );
  NOR2_X1 U22012 ( .A1(n18896), .A2(n18865), .ZN(n18870) );
  OAI22_X1 U22013 ( .A1(n19156), .A2(n19885), .B1(n18937), .B2(n18866), .ZN(
        n18867) );
  AOI221_X1 U22014 ( .B1(n18870), .B2(n18869), .C1(n18868), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18867), .ZN(n18879) );
  NAND2_X1 U22015 ( .A1(n18910), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18875) );
  INV_X1 U22016 ( .A(n18871), .ZN(n18872) );
  NAND2_X1 U22017 ( .A1(n18872), .A2(n18875), .ZN(n18874) );
  MUX2_X1 U22018 ( .A(n18875), .B(n18874), .S(n18873), .Z(n18877) );
  NAND2_X1 U22019 ( .A1(n18877), .A2(n18876), .ZN(n19149) );
  NOR2_X1 U22020 ( .A1(n19140), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19148) );
  AOI22_X1 U22021 ( .A1(n19149), .A2(n18946), .B1(n18901), .B2(n19148), .ZN(
        n18878) );
  OAI211_X1 U22022 ( .C1(n18887), .C2(n19105), .A(n18879), .B(n18878), .ZN(
        P3_U2812) );
  INV_X1 U22023 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n21717) );
  NOR2_X1 U22024 ( .A1(n19156), .A2(n21717), .ZN(n19154) );
  AOI221_X1 U22025 ( .B1(n18882), .B2(n18881), .C1(n19690), .C2(n18881), .A(
        n18880), .ZN(n18883) );
  AOI211_X1 U22026 ( .C1(n18884), .C2(n19043), .A(n19154), .B(n18883), .ZN(
        n18886) );
  NOR2_X1 U22027 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10542), .ZN(
        n19152) );
  XNOR2_X1 U22028 ( .A(n9884), .B(n19143), .ZN(n19153) );
  AOI22_X1 U22029 ( .A1(n18901), .A2(n19152), .B1(n18946), .B2(n19153), .ZN(
        n18885) );
  OAI211_X1 U22030 ( .C1(n18887), .C2(n19143), .A(n18886), .B(n18885), .ZN(
        P3_U2813) );
  AOI21_X1 U22031 ( .B1(n18889), .B2(n18910), .A(n18888), .ZN(n18890) );
  XNOR2_X1 U22032 ( .A(n18890), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19169) );
  AOI21_X1 U22033 ( .B1(n19008), .B2(n18891), .A(n19006), .ZN(n18926) );
  OAI21_X1 U22034 ( .B1(n18893), .B2(n18892), .A(n18926), .ZN(n18915) );
  NOR3_X1 U22035 ( .A1(n18896), .A2(n18895), .A3(n18894), .ZN(n18914) );
  OAI211_X1 U22036 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18914), .B(n18897), .ZN(n18898) );
  NAND2_X1 U22037 ( .A1(n19268), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n19167) );
  OAI211_X1 U22038 ( .C1(n18937), .C2(n18899), .A(n18898), .B(n19167), .ZN(
        n18900) );
  AOI21_X1 U22039 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18915), .A(
        n18900), .ZN(n18904) );
  AOI22_X1 U22040 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n10542), .ZN(n18903) );
  OAI211_X1 U22041 ( .C1(n18966), .C2(n19169), .A(n18904), .B(n18903), .ZN(
        P3_U2814) );
  NOR2_X1 U22042 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18933), .ZN(
        n19175) );
  NOR2_X1 U22043 ( .A1(n18931), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n19177) );
  NAND2_X1 U22044 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18905) );
  NOR2_X1 U22045 ( .A1(n18906), .A2(n18905), .ZN(n18909) );
  INV_X1 U22046 ( .A(n18951), .ZN(n18908) );
  NOR2_X1 U22047 ( .A1(n18908), .A2(n18907), .ZN(n18922) );
  OAI222_X1 U22048 ( .A1(n19187), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), 
        .B1(n18910), .B2(n17224), .C1(n18909), .C2(n18922), .ZN(n18911) );
  XOR2_X1 U22049 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n18911), .Z(
        n19182) );
  OAI22_X1 U22050 ( .A1(n19177), .A2(n18912), .B1(n18966), .B2(n19182), .ZN(
        n18919) );
  INV_X1 U22051 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18913) );
  AOI22_X1 U22052 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18915), .B1(
        n18914), .B2(n18913), .ZN(n18916) );
  NAND2_X1 U22053 ( .A1(n19268), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n19180) );
  OAI211_X1 U22054 ( .C1(n18937), .C2(n18917), .A(n18916), .B(n19180), .ZN(
        n18918) );
  NOR2_X1 U22055 ( .A1(n18919), .A2(n18918), .ZN(n18920) );
  OAI21_X1 U22056 ( .B1(n19175), .B2(n18921), .A(n18920), .ZN(P3_U2815) );
  INV_X1 U22057 ( .A(n18922), .ZN(n18923) );
  OAI22_X1 U22058 ( .A1(n18923), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n19184), .B2(n18944), .ZN(n18924) );
  XNOR2_X1 U22059 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18924), .ZN(
        n19197) );
  INV_X1 U22060 ( .A(n18925), .ZN(n18928) );
  AOI221_X1 U22061 ( .B1(n18928), .B2(n21689), .C1(n18927), .C2(n21689), .A(
        n18926), .ZN(n18929) );
  NOR2_X1 U22062 ( .A1(n19156), .A2(n19881), .ZN(n19191) );
  AOI211_X1 U22063 ( .C1(n18930), .C2(n19043), .A(n18929), .B(n19191), .ZN(
        n18936) );
  AOI21_X1 U22064 ( .B1(n19201), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18932) );
  NOR2_X1 U22065 ( .A1(n18932), .A2(n18931), .ZN(n19192) );
  AOI221_X1 U22066 ( .B1(n17079), .B2(n19187), .C1(n19204), .C2(n19187), .A(
        n18933), .ZN(n19194) );
  AOI22_X1 U22067 ( .A1(n18934), .A2(n19192), .B1(n19048), .B2(n19194), .ZN(
        n18935) );
  OAI211_X1 U22068 ( .C1(n19197), .C2(n18966), .A(n18936), .B(n18935), .ZN(
        P3_U2816) );
  OAI22_X1 U22069 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18939), .B1(
        n18938), .B2(n18937), .ZN(n18940) );
  AOI21_X1 U22070 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18941), .A(
        n18940), .ZN(n18950) );
  INV_X1 U22071 ( .A(n18942), .ZN(n18943) );
  OAI21_X1 U22072 ( .B1(n10312), .B2(n18944), .A(n18943), .ZN(n18945) );
  XNOR2_X1 U22073 ( .A(n18945), .B(n17224), .ZN(n19218) );
  AOI22_X1 U22074 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18947), .B1(
        n18946), .B2(n19218), .ZN(n18949) );
  NAND2_X1 U22075 ( .A1(n19268), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n19219) );
  NAND3_X1 U22076 ( .A1(n18960), .A2(n19213), .A3(n17224), .ZN(n18948) );
  NAND4_X1 U22077 ( .A1(n18950), .A2(n18949), .A3(n19219), .A4(n18948), .ZN(
        P3_U2818) );
  AOI22_X1 U22078 ( .A1(n18952), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n18951), .B2(n17259), .ZN(n18953) );
  XOR2_X1 U22079 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18953), .Z(
        n19250) );
  AOI21_X1 U22080 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19049), .A(
        n18954), .ZN(n18956) );
  OAI22_X1 U22081 ( .A1(n18957), .A2(n18956), .B1(n19054), .B2(n18955), .ZN(
        n18964) );
  INV_X1 U22082 ( .A(n18958), .ZN(n18959) );
  NAND3_X1 U22083 ( .A1(n18960), .A2(n19235), .A3(n18959), .ZN(n18961) );
  OAI21_X1 U22084 ( .B1(n18962), .B2(n17080), .A(n18961), .ZN(n18963) );
  AOI211_X1 U22085 ( .C1(n19268), .C2(P3_REIP_REG_10__SCAN_IN), .A(n18964), 
        .B(n18963), .ZN(n18965) );
  OAI21_X1 U22086 ( .B1(n19250), .B2(n18966), .A(n18965), .ZN(P3_U2820) );
  OAI21_X1 U22087 ( .B1(n18969), .B2(n18968), .A(n18967), .ZN(n18970) );
  XNOR2_X1 U22088 ( .A(n18970), .B(n19261), .ZN(n19266) );
  NAND2_X1 U22089 ( .A1(n19730), .A2(n18973), .ZN(n18971) );
  OAI22_X1 U22090 ( .A1(n18974), .A2(n18973), .B1(n18972), .B2(n18971), .ZN(
        n18975) );
  AOI21_X1 U22091 ( .B1(n19268), .B2(P3_REIP_REG_7__SCAN_IN), .A(n18975), .ZN(
        n18981) );
  OAI21_X1 U22092 ( .B1(n18977), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18976), .ZN(n18978) );
  INV_X1 U22093 ( .A(n18978), .ZN(n19259) );
  AOI22_X1 U22094 ( .A1(n19043), .A2(n18979), .B1(n19051), .B2(n19259), .ZN(
        n18980) );
  OAI211_X1 U22095 ( .C1(n19040), .C2(n19266), .A(n18981), .B(n18980), .ZN(
        P3_U2823) );
  OAI21_X1 U22096 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18983), .A(
        n18982), .ZN(n19275) );
  NOR2_X1 U22097 ( .A1(n18989), .A2(n19690), .ZN(n18984) );
  AOI22_X1 U22098 ( .A1(n19268), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18984), 
        .B2(n18990), .ZN(n18994) );
  OAI21_X1 U22099 ( .B1(n18987), .B2(n18986), .A(n18985), .ZN(n18988) );
  INV_X1 U22100 ( .A(n18988), .ZN(n19273) );
  OAI21_X1 U22101 ( .B1(n19690), .B2(n18989), .A(n19049), .ZN(n19001) );
  OAI22_X1 U22102 ( .A1(n19054), .A2(n18991), .B1(n18990), .B2(n19001), .ZN(
        n18992) );
  AOI21_X1 U22103 ( .B1(n19051), .B2(n19273), .A(n18992), .ZN(n18993) );
  OAI211_X1 U22104 ( .C1(n19040), .C2(n19275), .A(n18994), .B(n18993), .ZN(
        P3_U2824) );
  OAI21_X1 U22105 ( .B1(n18997), .B2(n18996), .A(n18995), .ZN(n19284) );
  XNOR2_X1 U22106 ( .A(n18999), .B(n18998), .ZN(n19279) );
  AOI21_X1 U22107 ( .B1(n19000), .B2(n9715), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19002) );
  OAI22_X1 U22108 ( .A1(n19054), .A2(n19003), .B1(n19002), .B2(n19001), .ZN(
        n19004) );
  AOI21_X1 U22109 ( .B1(n19051), .B2(n19279), .A(n19004), .ZN(n19005) );
  NAND2_X1 U22110 ( .A1(n19268), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n19282) );
  OAI211_X1 U22111 ( .C1(n19040), .C2(n19284), .A(n19005), .B(n19282), .ZN(
        P3_U2825) );
  AOI21_X1 U22112 ( .B1(n19008), .B2(n19007), .A(n19006), .ZN(n19027) );
  OAI21_X1 U22113 ( .B1(n19011), .B2(n19010), .A(n19009), .ZN(n19012) );
  XNOR2_X1 U22114 ( .A(n19012), .B(n21879), .ZN(n19293) );
  OAI22_X1 U22115 ( .A1(n19040), .A2(n19293), .B1(n19156), .B2(n19862), .ZN(
        n19013) );
  AOI21_X1 U22116 ( .B1(n19730), .B2(n19014), .A(n19013), .ZN(n19021) );
  OR2_X1 U22117 ( .A1(n19016), .A2(n19015), .ZN(n19017) );
  AND2_X1 U22118 ( .A1(n19018), .A2(n19017), .ZN(n19292) );
  AOI22_X1 U22119 ( .A1(n19043), .A2(n19019), .B1(n19051), .B2(n19292), .ZN(
        n19020) );
  OAI211_X1 U22120 ( .C1(n19022), .C2(n19027), .A(n19021), .B(n19020), .ZN(
        P3_U2826) );
  OAI21_X1 U22121 ( .B1(n19025), .B2(n19024), .A(n19023), .ZN(n19301) );
  XOR2_X1 U22122 ( .A(n19026), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n19302) );
  AOI21_X1 U22123 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n9715), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19028) );
  OAI22_X1 U22124 ( .A1(n19054), .A2(n19029), .B1(n19028), .B2(n19027), .ZN(
        n19030) );
  AOI21_X1 U22125 ( .B1(n19051), .B2(n19302), .A(n19030), .ZN(n19031) );
  NAND2_X1 U22126 ( .A1(n19268), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n19303) );
  OAI211_X1 U22127 ( .C1(n19040), .C2(n19301), .A(n19031), .B(n19303), .ZN(
        P3_U2827) );
  OAI21_X1 U22128 ( .B1(n19034), .B2(n19033), .A(n19032), .ZN(n19320) );
  OAI21_X1 U22129 ( .B1(n19037), .B2(n19036), .A(n19035), .ZN(n19038) );
  INV_X1 U22130 ( .A(n19038), .ZN(n19322) );
  AND2_X1 U22131 ( .A1(n19268), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n19325) );
  AOI21_X1 U22132 ( .B1(n19051), .B2(n19322), .A(n19325), .ZN(n19039) );
  OAI21_X1 U22133 ( .B1(n19040), .B2(n19320), .A(n19039), .ZN(n19041) );
  AOI21_X1 U22134 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(n19044) );
  OAI221_X1 U22135 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19690), .C1(
        n19046), .C2(n9715), .A(n19044), .ZN(P3_U2828) );
  AOI22_X1 U22136 ( .A1(n19048), .A2(n19047), .B1(n19268), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n19053) );
  AOI22_X1 U22137 ( .A1(n19051), .A2(n19050), .B1(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19049), .ZN(n19052) );
  OAI211_X1 U22138 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19054), .A(
        n19053), .B(n19052), .ZN(P3_U2829) );
  OAI21_X1 U22139 ( .B1(n19055), .B2(n19060), .A(n19787), .ZN(n19056) );
  AOI21_X1 U22140 ( .B1(n19057), .B2(n19056), .A(n19070), .ZN(n19062) );
  INV_X1 U22141 ( .A(n19058), .ZN(n19059) );
  NOR3_X1 U22142 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n19060), .A3(
        n19059), .ZN(n19061) );
  AOI211_X1 U22143 ( .C1(n19063), .C2(n19786), .A(n19062), .B(n19061), .ZN(
        n19065) );
  OAI22_X1 U22144 ( .A1(n19065), .A2(n19336), .B1(n19249), .B2(n19064), .ZN(
        n19066) );
  AOI21_X1 U22145 ( .B1(n19193), .B2(n19067), .A(n19066), .ZN(n19069) );
  OAI211_X1 U22146 ( .C1(n19329), .C2(n19070), .A(n19069), .B(n19068), .ZN(
        P3_U2837) );
  OAI22_X1 U22147 ( .A1(n19072), .A2(n19200), .B1(n19071), .B2(n19321), .ZN(
        n19073) );
  OAI211_X1 U22148 ( .C1(n19075), .C2(n19314), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n19077), .ZN(n19076) );
  NAND2_X1 U22149 ( .A1(n19156), .A2(n19076), .ZN(n19086) );
  AOI211_X1 U22150 ( .C1(n19183), .C2(n19077), .A(n10061), .B(n19086), .ZN(
        n19081) );
  OAI22_X1 U22151 ( .A1(n19079), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n19078), .B2(n19249), .ZN(n19080) );
  OR3_X1 U22152 ( .A1(n19082), .A2(n19081), .A3(n19080), .ZN(P3_U2838) );
  AOI21_X1 U22153 ( .B1(n19083), .B2(n19329), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n19087) );
  AOI22_X1 U22154 ( .A1(n19268), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n19255), 
        .B2(n19084), .ZN(n19085) );
  OAI21_X1 U22155 ( .B1(n19087), .B2(n19086), .A(n19085), .ZN(P3_U2839) );
  AOI221_X1 U22156 ( .B1(n19106), .B2(n19089), .C1(n19088), .C2(n19089), .A(
        n19336), .ZN(n19101) );
  AOI22_X1 U22157 ( .A1(n19786), .A2(n19171), .B1(n19232), .B2(n19170), .ZN(
        n19109) );
  AOI21_X1 U22158 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n19142), .A(
        n19314), .ZN(n19090) );
  AOI221_X1 U22159 ( .B1(n19091), .B2(n19337), .C1(n19124), .C2(n19337), .A(
        n19090), .ZN(n19122) );
  NAND2_X1 U22160 ( .A1(n19321), .A2(n19200), .ZN(n19234) );
  AOI22_X1 U22161 ( .A1(n19337), .A2(n19093), .B1(n19092), .B2(n19234), .ZN(
        n19094) );
  NAND2_X1 U22162 ( .A1(n19122), .A2(n19094), .ZN(n19112) );
  INV_X1 U22163 ( .A(n19112), .ZN(n19099) );
  INV_X1 U22164 ( .A(n19095), .ZN(n19113) );
  INV_X1 U22165 ( .A(n19096), .ZN(n19199) );
  AOI22_X1 U22166 ( .A1(n19787), .A2(n19113), .B1(n19114), .B2(n19199), .ZN(
        n19098) );
  NAND4_X1 U22167 ( .A1(n19109), .A2(n19099), .A3(n19098), .A4(n19097), .ZN(
        n19100) );
  AOI22_X1 U22168 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n19290), .B1(
        n19101), .B2(n19100), .ZN(n19103) );
  OAI211_X1 U22169 ( .C1(n19104), .C2(n19249), .A(n19103), .B(n19102), .ZN(
        P3_U2840) );
  NOR3_X1 U22170 ( .A1(n19106), .A2(n19336), .A3(n19105), .ZN(n19131) );
  INV_X1 U22171 ( .A(n19107), .ZN(n19117) );
  NAND2_X1 U22172 ( .A1(n19108), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n19110) );
  NAND2_X1 U22173 ( .A1(n19323), .A2(n19109), .ZN(n19137) );
  AOI21_X1 U22174 ( .B1(n19121), .B2(n19113), .A(n19112), .ZN(n19115) );
  AOI211_X1 U22175 ( .C1(n19123), .C2(n19115), .A(n19268), .B(n19114), .ZN(
        n19116) );
  AOI21_X1 U22176 ( .B1(n19131), .B2(n19117), .A(n19116), .ZN(n19119) );
  OAI211_X1 U22177 ( .C1(n19120), .C2(n19249), .A(n19119), .B(n19118), .ZN(
        P3_U2841) );
  NAND2_X1 U22178 ( .A1(n19121), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19125) );
  AOI22_X1 U22179 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n19127), .B1(
        n19131), .B2(n19126), .ZN(n19129) );
  OAI211_X1 U22180 ( .C1(n19249), .C2(n19130), .A(n19129), .B(n19128), .ZN(
        P3_U2842) );
  AOI22_X1 U22181 ( .A1(n19255), .A2(n19132), .B1(n19131), .B2(n19136), .ZN(
        n19134) );
  OAI211_X1 U22182 ( .C1(n19136), .C2(n19135), .A(n19134), .B(n19133), .ZN(
        P3_U2843) );
  INV_X1 U22183 ( .A(n19137), .ZN(n19164) );
  NAND3_X1 U22184 ( .A1(n19138), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n19286), .ZN(n19139) );
  AOI22_X1 U22185 ( .A1(n19140), .A2(n19234), .B1(n19288), .B2(n19139), .ZN(
        n19141) );
  OAI211_X1 U22186 ( .C1(n19142), .C2(n19314), .A(n19164), .B(n19141), .ZN(
        n19155) );
  OAI221_X1 U22187 ( .B1(n19155), .B2(n19143), .C1(n19155), .C2(n19288), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n19151) );
  INV_X1 U22188 ( .A(n19144), .ZN(n19146) );
  NAND2_X1 U22189 ( .A1(n19145), .A2(n19263), .ZN(n19172) );
  NAND2_X1 U22190 ( .A1(n19146), .A2(n19172), .ZN(n19212) );
  NAND2_X1 U22191 ( .A1(n19323), .A2(n19212), .ZN(n19258) );
  NOR2_X1 U22192 ( .A1(n19147), .A2(n19258), .ZN(n19165) );
  AOI22_X1 U22193 ( .A1(n19149), .A2(n19255), .B1(n19148), .B2(n19165), .ZN(
        n19150) );
  OAI221_X1 U22194 ( .B1(n19268), .B2(n19151), .C1(n19156), .C2(n19885), .A(
        n19150), .ZN(P3_U2844) );
  AOI22_X1 U22195 ( .A1(n19153), .A2(n19255), .B1(n19165), .B2(n19152), .ZN(
        n19159) );
  INV_X1 U22196 ( .A(n19154), .ZN(n19158) );
  NAND3_X1 U22197 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n19156), .A3(
        n19155), .ZN(n19157) );
  NAND3_X1 U22198 ( .A1(n19159), .A2(n19158), .A3(n19157), .ZN(P3_U2845) );
  AOI21_X1 U22199 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n19237), .A(
        n19160), .ZN(n19162) );
  NAND2_X1 U22200 ( .A1(n19337), .A2(n19161), .ZN(n19222) );
  OAI21_X1 U22201 ( .B1(n19227), .B2(n19314), .A(n19222), .ZN(n19203) );
  AOI211_X1 U22202 ( .C1(n19163), .C2(n19199), .A(n19162), .B(n19203), .ZN(
        n19173) );
  AOI221_X1 U22203 ( .B1(n19183), .B2(n19164), .C1(n19173), .C2(n19164), .A(
        n19268), .ZN(n19166) );
  AOI22_X1 U22204 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n19166), .B1(
        n19165), .B2(n10542), .ZN(n19168) );
  OAI211_X1 U22205 ( .C1(n19169), .C2(n19249), .A(n19168), .B(n19167), .ZN(
        P3_U2846) );
  NAND2_X1 U22206 ( .A1(n19232), .A2(n19170), .ZN(n19178) );
  NAND2_X1 U22207 ( .A1(n19786), .A2(n19171), .ZN(n19176) );
  NOR2_X1 U22208 ( .A1(n19184), .A2(n19172), .ZN(n19186) );
  AOI21_X1 U22209 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n19186), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n19174) );
  OAI222_X1 U22210 ( .A1(n19178), .A2(n19177), .B1(n19176), .B2(n19175), .C1(
        n19174), .C2(n19173), .ZN(n19179) );
  AOI22_X1 U22211 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n19290), .B1(
        n19323), .B2(n19179), .ZN(n19181) );
  OAI211_X1 U22212 ( .C1(n19249), .C2(n19182), .A(n19181), .B(n19180), .ZN(
        P3_U2847) );
  INV_X1 U22213 ( .A(n19183), .ZN(n19185) );
  AOI21_X1 U22214 ( .B1(n19210), .B2(n19224), .A(n19237), .ZN(n19206) );
  AOI211_X1 U22215 ( .C1(n19185), .C2(n19184), .A(n19206), .B(n19203), .ZN(
        n19189) );
  INV_X1 U22216 ( .A(n19186), .ZN(n19188) );
  AOI221_X1 U22217 ( .B1(n19189), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n19188), .C2(n19187), .A(n19336), .ZN(n19190) );
  AOI211_X1 U22218 ( .C1(n19290), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n19191), .B(n19190), .ZN(n19196) );
  AOI22_X1 U22219 ( .A1(n19335), .A2(n19194), .B1(n19193), .B2(n19192), .ZN(
        n19195) );
  OAI211_X1 U22220 ( .C1(n19197), .C2(n19249), .A(n19196), .B(n19195), .ZN(
        P3_U2848) );
  AOI22_X1 U22221 ( .A1(n19268), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n19255), 
        .B2(n19198), .ZN(n19208) );
  NAND2_X1 U22222 ( .A1(n10312), .A2(n19199), .ZN(n19236) );
  OAI21_X1 U22223 ( .B1(n19201), .B2(n19200), .A(n19236), .ZN(n19202) );
  AOI211_X1 U22224 ( .C1(n19786), .C2(n19204), .A(n19203), .B(n19202), .ZN(
        n19216) );
  OAI211_X1 U22225 ( .C1(n19242), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n19323), .B(n19216), .ZN(n19205) );
  OAI211_X1 U22226 ( .C1(n19206), .C2(n19205), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n19156), .ZN(n19207) );
  OAI211_X1 U22227 ( .C1(n19258), .C2(n19209), .A(n19208), .B(n19207), .ZN(
        P3_U2849) );
  NAND2_X1 U22228 ( .A1(n19210), .A2(n19224), .ZN(n19211) );
  OAI21_X1 U22229 ( .B1(n17224), .B2(n19226), .A(n19211), .ZN(n19215) );
  AOI21_X1 U22230 ( .B1(n19213), .B2(n19212), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n19214) );
  AOI211_X1 U22231 ( .C1(n19216), .C2(n19215), .A(n19214), .B(n19336), .ZN(
        n19217) );
  AOI21_X1 U22232 ( .B1(n19255), .B2(n19218), .A(n19217), .ZN(n19220) );
  OAI211_X1 U22233 ( .C1(n19329), .C2(n17224), .A(n19220), .B(n19219), .ZN(
        P3_U2850) );
  AOI22_X1 U22234 ( .A1(n19268), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n19255), 
        .B2(n19221), .ZN(n19240) );
  NAND2_X1 U22235 ( .A1(n19323), .A2(n19222), .ZN(n19253) );
  NAND2_X1 U22236 ( .A1(n19786), .A2(n19223), .ZN(n19230) );
  INV_X1 U22237 ( .A(n19224), .ZN(n19225) );
  NAND2_X1 U22238 ( .A1(n19226), .A2(n19225), .ZN(n19229) );
  OR2_X1 U22239 ( .A1(n19227), .A2(n19314), .ZN(n19228) );
  NAND3_X1 U22240 ( .A1(n19230), .A2(n19229), .A3(n19228), .ZN(n19231) );
  AOI21_X1 U22241 ( .B1(n17105), .B2(n19232), .A(n19231), .ZN(n19251) );
  OAI21_X1 U22242 ( .B1(n19237), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n19251), .ZN(n19233) );
  AOI21_X1 U22243 ( .B1(n19235), .B2(n19234), .A(n19233), .ZN(n19245) );
  OAI211_X1 U22244 ( .C1(n19237), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n19245), .B(n19236), .ZN(n19238) );
  OAI211_X1 U22245 ( .C1(n19253), .C2(n19238), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n19156), .ZN(n19239) );
  OAI211_X1 U22246 ( .C1(n19241), .C2(n19258), .A(n19240), .B(n19239), .ZN(
        P3_U2851) );
  INV_X1 U22247 ( .A(n19242), .ZN(n19243) );
  OAI21_X1 U22248 ( .B1(n17259), .B2(n19253), .A(n19243), .ZN(n19244) );
  AOI21_X1 U22249 ( .B1(n19245), .B2(n19244), .A(n17080), .ZN(n19247) );
  NOR3_X1 U22250 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17259), .A3(
        n19258), .ZN(n19246) );
  AOI221_X1 U22251 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n19268), .C1(n19247), 
        .C2(n19156), .A(n19246), .ZN(n19248) );
  OAI21_X1 U22252 ( .B1(n19250), .B2(n19249), .A(n19248), .ZN(P3_U2852) );
  INV_X1 U22253 ( .A(n19251), .ZN(n19252) );
  OAI21_X1 U22254 ( .B1(n19253), .B2(n19252), .A(n19156), .ZN(n19257) );
  AOI22_X1 U22255 ( .A1(n19268), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n19255), 
        .B2(n19254), .ZN(n19256) );
  OAI221_X1 U22256 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n19258), .C1(
        n17259), .C2(n19257), .A(n19256), .ZN(P3_U2853) );
  AOI22_X1 U22257 ( .A1(n19259), .A2(n19331), .B1(n19268), .B2(
        P3_REIP_REG_7__SCAN_IN), .ZN(n19265) );
  OAI21_X1 U22258 ( .B1(n19261), .B2(n19329), .A(n19260), .ZN(n19262) );
  OAI221_X1 U22259 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n19263), .A(n19262), .ZN(
        n19264) );
  OAI211_X1 U22260 ( .C1(n19266), .C2(n19285), .A(n19265), .B(n19264), .ZN(
        P3_U2855) );
  NOR2_X1 U22261 ( .A1(n19290), .A2(n19267), .ZN(n19276) );
  NAND2_X1 U22262 ( .A1(n19268), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n19269) );
  OAI221_X1 U22263 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n19271), .C1(
        n19270), .C2(n19276), .A(n19269), .ZN(n19272) );
  AOI21_X1 U22264 ( .B1(n19273), .B2(n19331), .A(n19272), .ZN(n19274) );
  OAI21_X1 U22265 ( .B1(n19285), .B2(n19275), .A(n19274), .ZN(P3_U2856) );
  NAND3_X1 U22266 ( .A1(n19323), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n19308), .ZN(n19297) );
  NOR2_X1 U22267 ( .A1(n21879), .A2(n19297), .ZN(n19278) );
  INV_X1 U22268 ( .A(n19276), .ZN(n19277) );
  MUX2_X1 U22269 ( .A(n19278), .B(n19277), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n19281) );
  AND2_X1 U22270 ( .A1(n19331), .A2(n19279), .ZN(n19280) );
  NOR2_X1 U22271 ( .A1(n19281), .A2(n19280), .ZN(n19283) );
  OAI211_X1 U22272 ( .C1(n19285), .C2(n19284), .A(n19283), .B(n19282), .ZN(
        P3_U2857) );
  INV_X1 U22273 ( .A(n19286), .ZN(n19287) );
  AOI21_X1 U22274 ( .B1(n19289), .B2(n19288), .A(n19287), .ZN(n19311) );
  OAI211_X1 U22275 ( .C1(n19314), .C2(n19313), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n19311), .ZN(n19307) );
  AOI21_X1 U22276 ( .B1(n19291), .B2(n19307), .A(n19290), .ZN(n19300) );
  AOI22_X1 U22277 ( .A1(n19331), .A2(n19292), .B1(n19268), .B2(
        P3_REIP_REG_4__SCAN_IN), .ZN(n19296) );
  INV_X1 U22278 ( .A(n19293), .ZN(n19294) );
  NAND2_X1 U22279 ( .A1(n19335), .A2(n19294), .ZN(n19295) );
  OAI211_X1 U22280 ( .C1(n19297), .C2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n19296), .B(n19295), .ZN(n19298) );
  INV_X1 U22281 ( .A(n19298), .ZN(n19299) );
  OAI21_X1 U22282 ( .B1(n19300), .B2(n21879), .A(n19299), .ZN(P3_U2858) );
  INV_X1 U22283 ( .A(n19301), .ZN(n19306) );
  NAND2_X1 U22284 ( .A1(n19331), .A2(n19302), .ZN(n19304) );
  OAI211_X1 U22285 ( .C1(n19329), .C2(n21882), .A(n19304), .B(n19303), .ZN(
        n19305) );
  AOI21_X1 U22286 ( .B1(n19335), .B2(n19306), .A(n19305), .ZN(n19310) );
  OAI211_X1 U22287 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n19308), .A(
        n19323), .B(n19307), .ZN(n19309) );
  NAND2_X1 U22288 ( .A1(n19310), .A2(n19309), .ZN(P3_U2859) );
  NAND2_X1 U22289 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19312) );
  OAI21_X1 U22290 ( .B1(n19314), .B2(n19312), .A(n19311), .ZN(n19316) );
  NOR2_X1 U22291 ( .A1(n19314), .A2(n19313), .ZN(n19315) );
  AOI21_X1 U22292 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n19316), .A(
        n19315), .ZN(n19319) );
  NAND3_X1 U22293 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n19317), .A3(
        n19328), .ZN(n19318) );
  OAI211_X1 U22294 ( .C1(n19321), .C2(n19320), .A(n19319), .B(n19318), .ZN(
        n19324) );
  AOI22_X1 U22295 ( .A1(n19324), .A2(n19323), .B1(n19331), .B2(n19322), .ZN(
        n19327) );
  INV_X1 U22296 ( .A(n19325), .ZN(n19326) );
  OAI211_X1 U22297 ( .C1(n19329), .C2(n19328), .A(n19327), .B(n19326), .ZN(
        P3_U2860) );
  INV_X1 U22298 ( .A(n19330), .ZN(n19334) );
  INV_X1 U22299 ( .A(n19331), .ZN(n19332) );
  INV_X1 U22300 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19930) );
  OAI22_X1 U22301 ( .A1(n19332), .A2(n19334), .B1(n19930), .B2(n19156), .ZN(
        n19333) );
  AOI21_X1 U22302 ( .B1(n19335), .B2(n19334), .A(n19333), .ZN(n19340) );
  OAI211_X1 U22303 ( .C1(n19337), .C2(n19336), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n19156), .ZN(n19338) );
  NAND3_X1 U22304 ( .A1(n19340), .A2(n19339), .A3(n19338), .ZN(P3_U2862) );
  AOI21_X1 U22305 ( .B1(n19343), .B2(n19342), .A(n19341), .ZN(n19825) );
  OAI21_X1 U22306 ( .B1(n19825), .B2(n19428), .A(n19348), .ZN(n19344) );
  OAI221_X1 U22307 ( .B1(n19587), .B2(n19937), .C1(n19587), .C2(n19348), .A(
        n19344), .ZN(P3_U2863) );
  INV_X1 U22308 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19813) );
  NOR2_X1 U22309 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19813), .ZN(
        n19565) );
  NOR2_X1 U22310 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13797), .ZN(
        n19522) );
  NOR2_X1 U22311 ( .A1(n19565), .A2(n19522), .ZN(n19345) );
  OAI22_X1 U22312 ( .A1(n19347), .A2(n19813), .B1(n19346), .B2(n19345), .ZN(
        P3_U2866) );
  NOR2_X1 U22313 ( .A1(n19814), .A2(n19348), .ZN(P3_U2867) );
  NOR2_X1 U22314 ( .A1(n13797), .A2(n19813), .ZN(n19663) );
  NOR2_X1 U22315 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19587), .ZN(
        n19474) );
  NAND2_X1 U22316 ( .A1(n19663), .A2(n19474), .ZN(n19784) );
  NAND2_X1 U22317 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19730), .ZN(n19735) );
  NOR2_X1 U22318 ( .A1(n19813), .A2(n19497), .ZN(n19728) );
  NAND2_X1 U22319 ( .A1(n19587), .A2(n19728), .ZN(n19712) );
  INV_X1 U22320 ( .A(n19712), .ZN(n19719) );
  AND2_X1 U22321 ( .A1(n19730), .A2(BUF2_REG_16__SCAN_IN), .ZN(n19726) );
  NOR2_X2 U22322 ( .A1(n19635), .A2(n19349), .ZN(n19725) );
  NAND2_X1 U22323 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19800) );
  INV_X1 U22324 ( .A(n19663), .ZN(n19661) );
  NOR2_X2 U22325 ( .A1(n19800), .A2(n19661), .ZN(n19779) );
  NAND2_X1 U22326 ( .A1(n19806), .A2(n19587), .ZN(n19808) );
  NAND2_X1 U22327 ( .A1(n13797), .A2(n19813), .ZN(n19475) );
  NOR2_X2 U22328 ( .A1(n19808), .A2(n19475), .ZN(n19447) );
  NOR2_X1 U22329 ( .A1(n19779), .A2(n19447), .ZN(n19408) );
  NOR2_X1 U22330 ( .A1(n19688), .A2(n19408), .ZN(n19381) );
  AOI22_X1 U22331 ( .A1(n19719), .A2(n19726), .B1(n19725), .B2(n19381), .ZN(
        n19357) );
  AOI21_X1 U22332 ( .B1(n19784), .B2(n19712), .A(n19635), .ZN(n19693) );
  NOR2_X1 U22333 ( .A1(n19408), .A2(n19635), .ZN(n19351) );
  AOI22_X1 U22334 ( .A1(n19407), .A2(n19693), .B1(n19351), .B2(n19350), .ZN(
        n19384) );
  INV_X1 U22335 ( .A(n19352), .ZN(n19353) );
  NAND2_X1 U22336 ( .A1(n19354), .A2(n19353), .ZN(n19382) );
  NOR2_X1 U22337 ( .A1(n19355), .A2(n19382), .ZN(n19731) );
  AOI22_X1 U22338 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19731), .ZN(n19356) );
  OAI211_X1 U22339 ( .C1(n19784), .C2(n19735), .A(n19357), .B(n19356), .ZN(
        P3_U2868) );
  NAND2_X1 U22340 ( .A1(n19730), .A2(BUF2_REG_17__SCAN_IN), .ZN(n19670) );
  INV_X1 U22341 ( .A(n19784), .ZN(n19763) );
  AND2_X1 U22342 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19730), .ZN(n19738) );
  NOR2_X2 U22343 ( .A1(n19635), .A2(n19358), .ZN(n19736) );
  AOI22_X1 U22344 ( .A1(n19763), .A2(n19738), .B1(n19381), .B2(n19736), .ZN(
        n19360) );
  NOR2_X1 U22345 ( .A1(n19943), .A2(n19382), .ZN(n19667) );
  AOI22_X1 U22346 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19667), .ZN(n19359) );
  OAI211_X1 U22347 ( .C1(n19712), .C2(n19670), .A(n19360), .B(n19359), .ZN(
        P3_U2869) );
  NAND2_X1 U22348 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19730), .ZN(n19645) );
  AND2_X1 U22349 ( .A1(n19730), .A2(BUF2_REG_18__SCAN_IN), .ZN(n19744) );
  NOR2_X2 U22350 ( .A1(n19635), .A2(n19361), .ZN(n19742) );
  AOI22_X1 U22351 ( .A1(n19719), .A2(n19744), .B1(n19381), .B2(n19742), .ZN(
        n19363) );
  NOR2_X1 U22352 ( .A1(n13766), .A2(n19382), .ZN(n19642) );
  AOI22_X1 U22353 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19642), .ZN(n19362) );
  OAI211_X1 U22354 ( .C1(n19784), .C2(n19645), .A(n19363), .B(n19362), .ZN(
        P3_U2870) );
  NAND2_X1 U22355 ( .A1(n19730), .A2(BUF2_REG_19__SCAN_IN), .ZN(n19753) );
  AND2_X1 U22356 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19730), .ZN(n19749) );
  NOR2_X2 U22357 ( .A1(n19635), .A2(n19364), .ZN(n19748) );
  AOI22_X1 U22358 ( .A1(n19763), .A2(n19749), .B1(n19381), .B2(n19748), .ZN(
        n19367) );
  NOR2_X1 U22359 ( .A1(n19365), .A2(n19382), .ZN(n19750) );
  AOI22_X1 U22360 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19750), .ZN(n19366) );
  OAI211_X1 U22361 ( .C1(n19712), .C2(n19753), .A(n19367), .B(n19366), .ZN(
        P3_U2871) );
  NAND2_X1 U22362 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19730), .ZN(n19708) );
  AND2_X1 U22363 ( .A1(n19730), .A2(BUF2_REG_20__SCAN_IN), .ZN(n19756) );
  NOR2_X2 U22364 ( .A1(n19635), .A2(n19368), .ZN(n19754) );
  AOI22_X1 U22365 ( .A1(n19719), .A2(n19756), .B1(n19381), .B2(n19754), .ZN(
        n19371) );
  NOR2_X1 U22366 ( .A1(n19369), .A2(n19382), .ZN(n19705) );
  AOI22_X1 U22367 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19705), .ZN(n19370) );
  OAI211_X1 U22368 ( .C1(n19784), .C2(n19708), .A(n19371), .B(n19370), .ZN(
        P3_U2872) );
  NAND2_X1 U22369 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19730), .ZN(n19680) );
  AND2_X1 U22370 ( .A1(n19730), .A2(BUF2_REG_21__SCAN_IN), .ZN(n19762) );
  NOR2_X2 U22371 ( .A1(n19635), .A2(n19372), .ZN(n19760) );
  AOI22_X1 U22372 ( .A1(n19719), .A2(n19762), .B1(n19381), .B2(n19760), .ZN(
        n19375) );
  NOR2_X1 U22373 ( .A1(n19373), .A2(n19382), .ZN(n19677) );
  AOI22_X1 U22374 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19677), .ZN(n19374) );
  OAI211_X1 U22375 ( .C1(n19784), .C2(n19680), .A(n19375), .B(n19374), .ZN(
        P3_U2873) );
  NAND2_X1 U22376 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n19730), .ZN(n19773) );
  NOR2_X1 U22377 ( .A1(n14713), .A2(n19690), .ZN(n19769) );
  NOR2_X2 U22378 ( .A1(n19376), .A2(n19635), .ZN(n19768) );
  AOI22_X1 U22379 ( .A1(n19763), .A2(n19769), .B1(n19381), .B2(n19768), .ZN(
        n19379) );
  NOR2_X2 U22380 ( .A1(n19377), .A2(n19382), .ZN(n19770) );
  AOI22_X1 U22381 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19770), .ZN(n19378) );
  OAI211_X1 U22382 ( .C1(n19712), .C2(n19773), .A(n19379), .B(n19378), .ZN(
        P3_U2874) );
  NAND2_X1 U22383 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19730), .ZN(n19783) );
  NOR2_X1 U22384 ( .A1(n19690), .A2(n21701), .ZN(n19777) );
  NOR2_X2 U22385 ( .A1(n19380), .A2(n19635), .ZN(n19775) );
  AOI22_X1 U22386 ( .A1(n19763), .A2(n19777), .B1(n19381), .B2(n19775), .ZN(
        n19386) );
  NOR2_X2 U22387 ( .A1(n19383), .A2(n19382), .ZN(n19778) );
  AOI22_X1 U22388 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19384), .B1(
        n19447), .B2(n19778), .ZN(n19385) );
  OAI211_X1 U22389 ( .C1(n19712), .C2(n19783), .A(n19386), .B(n19385), .ZN(
        P3_U2875) );
  INV_X1 U22390 ( .A(n19475), .ZN(n19430) );
  NOR2_X1 U22391 ( .A1(n19428), .A2(n19635), .ZN(n19727) );
  AND2_X1 U22392 ( .A1(n19727), .A2(n19806), .ZN(n19662) );
  AOI22_X1 U22393 ( .A1(n19730), .A2(n19728), .B1(n19430), .B2(n19662), .ZN(
        n19404) );
  INV_X1 U22394 ( .A(n19404), .ZN(n19397) );
  INV_X1 U22395 ( .A(n19735), .ZN(n19689) );
  INV_X1 U22396 ( .A(n19688), .ZN(n19836) );
  NAND2_X1 U22397 ( .A1(n19806), .A2(n19836), .ZN(n19660) );
  NOR2_X1 U22398 ( .A1(n19475), .A2(n19660), .ZN(n19403) );
  AOI22_X1 U22399 ( .A1(n19689), .A2(n19719), .B1(n19725), .B2(n19403), .ZN(
        n19388) );
  INV_X1 U22400 ( .A(n19474), .ZN(n19567) );
  NOR2_X1 U22401 ( .A1(n19567), .A2(n19475), .ZN(n19459) );
  AOI22_X1 U22402 ( .A1(n19779), .A2(n19726), .B1(n19731), .B2(n19459), .ZN(
        n19387) );
  OAI211_X1 U22403 ( .C1(n18308), .C2(n19397), .A(n19388), .B(n19387), .ZN(
        P3_U2876) );
  INV_X1 U22404 ( .A(n19670), .ZN(n19737) );
  AOI22_X1 U22405 ( .A1(n19779), .A2(n19737), .B1(n19736), .B2(n19403), .ZN(
        n19390) );
  CLKBUF_X1 U22406 ( .A(n19459), .Z(n19462) );
  AOI22_X1 U22407 ( .A1(n19719), .A2(n19738), .B1(n19667), .B2(n19462), .ZN(
        n19389) );
  OAI211_X1 U22408 ( .C1(n18291), .C2(n19397), .A(n19390), .B(n19389), .ZN(
        P3_U2877) );
  INV_X1 U22409 ( .A(n19645), .ZN(n19743) );
  AOI22_X1 U22410 ( .A1(n19719), .A2(n19743), .B1(n19742), .B2(n19403), .ZN(
        n19392) );
  AOI22_X1 U22411 ( .A1(n19779), .A2(n19744), .B1(n19642), .B2(n19462), .ZN(
        n19391) );
  OAI211_X1 U22412 ( .C1(n13697), .C2(n19397), .A(n19392), .B(n19391), .ZN(
        P3_U2878) );
  INV_X1 U22413 ( .A(n19753), .ZN(n19701) );
  AOI22_X1 U22414 ( .A1(n19779), .A2(n19701), .B1(n19748), .B2(n19403), .ZN(
        n19394) );
  AOI22_X1 U22415 ( .A1(n19719), .A2(n19749), .B1(n19750), .B2(n19462), .ZN(
        n19393) );
  OAI211_X1 U22416 ( .C1(n18253), .C2(n19397), .A(n19394), .B(n19393), .ZN(
        P3_U2879) );
  INV_X1 U22417 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n19398) );
  INV_X1 U22418 ( .A(n19708), .ZN(n19755) );
  AOI22_X1 U22419 ( .A1(n19719), .A2(n19755), .B1(n19754), .B2(n19403), .ZN(
        n19396) );
  AOI22_X1 U22420 ( .A1(n19779), .A2(n19756), .B1(n19705), .B2(n19459), .ZN(
        n19395) );
  OAI211_X1 U22421 ( .C1(n19398), .C2(n19397), .A(n19396), .B(n19395), .ZN(
        P3_U2880) );
  AOI22_X1 U22422 ( .A1(n19779), .A2(n19762), .B1(n19760), .B2(n19403), .ZN(
        n19400) );
  AOI22_X1 U22423 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19404), .B1(
        n19677), .B2(n19459), .ZN(n19399) );
  OAI211_X1 U22424 ( .C1(n19712), .C2(n19680), .A(n19400), .B(n19399), .ZN(
        P3_U2881) );
  INV_X1 U22425 ( .A(n19769), .ZN(n19716) );
  INV_X1 U22426 ( .A(n19773), .ZN(n19713) );
  AOI22_X1 U22427 ( .A1(n19779), .A2(n19713), .B1(n19768), .B2(n19403), .ZN(
        n19402) );
  AOI22_X1 U22428 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19404), .B1(
        n19770), .B2(n19462), .ZN(n19401) );
  OAI211_X1 U22429 ( .C1(n19712), .C2(n19716), .A(n19402), .B(n19401), .ZN(
        P3_U2882) );
  INV_X1 U22430 ( .A(n19779), .ZN(n19767) );
  AOI22_X1 U22431 ( .A1(n19719), .A2(n19777), .B1(n19775), .B2(n19403), .ZN(
        n19406) );
  AOI22_X1 U22432 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19404), .B1(
        n19778), .B2(n19462), .ZN(n19405) );
  OAI211_X1 U22433 ( .C1(n19767), .C2(n19783), .A(n19406), .B(n19405), .ZN(
        P3_U2883) );
  NOR3_X1 U22434 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19806), .A3(
        n19475), .ZN(n19481) );
  INV_X1 U22435 ( .A(n19407), .ZN(n19588) );
  NOR2_X1 U22436 ( .A1(n19462), .A2(n19493), .ZN(n19451) );
  OAI21_X1 U22437 ( .B1(n19408), .B2(n19588), .A(n19451), .ZN(n19409) );
  OAI211_X1 U22438 ( .C1(n19493), .C2(n19923), .A(n19591), .B(n19409), .ZN(
        n19425) );
  NOR2_X1 U22439 ( .A1(n19688), .A2(n19451), .ZN(n19424) );
  AOI22_X1 U22440 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19425), .B1(
        n19725), .B2(n19424), .ZN(n19411) );
  AOI22_X1 U22441 ( .A1(n19447), .A2(n19726), .B1(n19731), .B2(n19493), .ZN(
        n19410) );
  OAI211_X1 U22442 ( .C1(n19735), .C2(n19767), .A(n19411), .B(n19410), .ZN(
        P3_U2884) );
  INV_X1 U22443 ( .A(n19447), .ZN(n19445) );
  AOI22_X1 U22444 ( .A1(n19779), .A2(n19738), .B1(n19736), .B2(n19424), .ZN(
        n19413) );
  AOI22_X1 U22445 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19425), .B1(
        n19667), .B2(n19493), .ZN(n19412) );
  OAI211_X1 U22446 ( .C1(n19445), .C2(n19670), .A(n19413), .B(n19412), .ZN(
        P3_U2885) );
  AOI22_X1 U22447 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19425), .B1(
        n19742), .B2(n19424), .ZN(n19415) );
  AOI22_X1 U22448 ( .A1(n19447), .A2(n19744), .B1(n19642), .B2(n19481), .ZN(
        n19414) );
  OAI211_X1 U22449 ( .C1(n19767), .C2(n19645), .A(n19415), .B(n19414), .ZN(
        P3_U2886) );
  AOI22_X1 U22450 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19425), .B1(
        n19748), .B2(n19424), .ZN(n19417) );
  AOI22_X1 U22451 ( .A1(n19779), .A2(n19749), .B1(n19750), .B2(n19481), .ZN(
        n19416) );
  OAI211_X1 U22452 ( .C1(n19445), .C2(n19753), .A(n19417), .B(n19416), .ZN(
        P3_U2887) );
  AOI22_X1 U22453 ( .A1(n19447), .A2(n19756), .B1(n19754), .B2(n19424), .ZN(
        n19419) );
  AOI22_X1 U22454 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19425), .B1(
        n19705), .B2(n19481), .ZN(n19418) );
  OAI211_X1 U22455 ( .C1(n19767), .C2(n19708), .A(n19419), .B(n19418), .ZN(
        P3_U2888) );
  AOI22_X1 U22456 ( .A1(n19447), .A2(n19762), .B1(n19760), .B2(n19424), .ZN(
        n19421) );
  AOI22_X1 U22457 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19425), .B1(
        n19677), .B2(n19493), .ZN(n19420) );
  OAI211_X1 U22458 ( .C1(n19767), .C2(n19680), .A(n19421), .B(n19420), .ZN(
        P3_U2889) );
  AOI22_X1 U22459 ( .A1(n19779), .A2(n19769), .B1(n19768), .B2(n19424), .ZN(
        n19423) );
  AOI22_X1 U22460 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19425), .B1(
        n19770), .B2(n19493), .ZN(n19422) );
  OAI211_X1 U22461 ( .C1(n19445), .C2(n19773), .A(n19423), .B(n19422), .ZN(
        P3_U2890) );
  AOI22_X1 U22462 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19425), .B1(
        n19775), .B2(n19424), .ZN(n19427) );
  AOI22_X1 U22463 ( .A1(n19779), .A2(n19777), .B1(n19778), .B2(n19493), .ZN(
        n19426) );
  OAI211_X1 U22464 ( .C1(n19445), .C2(n19783), .A(n19427), .B(n19426), .ZN(
        P3_U2891) );
  INV_X1 U22465 ( .A(n19731), .ZN(n19696) );
  NOR2_X2 U22466 ( .A1(n19800), .A2(n19475), .ZN(n19512) );
  INV_X1 U22467 ( .A(n19512), .ZN(n19519) );
  AOI22_X1 U22468 ( .A1(n19689), .A2(n19447), .B1(n19725), .B2(n19446), .ZN(
        n19432) );
  OR2_X1 U22469 ( .A1(n19806), .A2(n19428), .ZN(n19429) );
  AOI21_X1 U22470 ( .B1(n19588), .B2(n19429), .A(n19635), .ZN(n19521) );
  NAND2_X1 U22471 ( .A1(n19430), .A2(n19521), .ZN(n19448) );
  AOI22_X1 U22472 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19448), .B1(
        n19726), .B2(n19459), .ZN(n19431) );
  OAI211_X1 U22473 ( .C1(n19696), .C2(n19519), .A(n19432), .B(n19431), .ZN(
        P3_U2892) );
  AOI22_X1 U22474 ( .A1(n19737), .A2(n19459), .B1(n19736), .B2(n19446), .ZN(
        n19434) );
  AOI22_X1 U22475 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19448), .B1(
        n19447), .B2(n19738), .ZN(n19433) );
  OAI211_X1 U22476 ( .C1(n19741), .C2(n19519), .A(n19434), .B(n19433), .ZN(
        P3_U2893) );
  INV_X1 U22477 ( .A(n19642), .ZN(n19747) );
  AOI22_X1 U22478 ( .A1(n19447), .A2(n19743), .B1(n19742), .B2(n19446), .ZN(
        n19436) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19448), .B1(
        n19744), .B2(n19459), .ZN(n19435) );
  OAI211_X1 U22480 ( .C1(n19747), .C2(n19519), .A(n19436), .B(n19435), .ZN(
        P3_U2894) );
  INV_X1 U22481 ( .A(n19750), .ZN(n19704) );
  AOI22_X1 U22482 ( .A1(n19447), .A2(n19749), .B1(n19748), .B2(n19446), .ZN(
        n19438) );
  AOI22_X1 U22483 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19448), .B1(
        n19701), .B2(n19462), .ZN(n19437) );
  OAI211_X1 U22484 ( .C1(n19704), .C2(n19519), .A(n19438), .B(n19437), .ZN(
        P3_U2895) );
  INV_X1 U22485 ( .A(n19705), .ZN(n19759) );
  AOI22_X1 U22486 ( .A1(n19447), .A2(n19755), .B1(n19754), .B2(n19446), .ZN(
        n19440) );
  AOI22_X1 U22487 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19448), .B1(
        n19756), .B2(n19462), .ZN(n19439) );
  OAI211_X1 U22488 ( .C1(n19759), .C2(n19519), .A(n19440), .B(n19439), .ZN(
        P3_U2896) );
  AOI22_X1 U22489 ( .A1(n19762), .A2(n19459), .B1(n19760), .B2(n19446), .ZN(
        n19442) );
  AOI22_X1 U22490 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19448), .B1(
        n19677), .B2(n19512), .ZN(n19441) );
  OAI211_X1 U22491 ( .C1(n19445), .C2(n19680), .A(n19442), .B(n19441), .ZN(
        P3_U2897) );
  AOI22_X1 U22492 ( .A1(n19713), .A2(n19462), .B1(n19768), .B2(n19446), .ZN(
        n19444) );
  AOI22_X1 U22493 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19448), .B1(
        n19770), .B2(n19512), .ZN(n19443) );
  OAI211_X1 U22494 ( .C1(n19445), .C2(n19716), .A(n19444), .B(n19443), .ZN(
        P3_U2898) );
  INV_X1 U22495 ( .A(n19459), .ZN(n19473) );
  AOI22_X1 U22496 ( .A1(n19447), .A2(n19777), .B1(n19775), .B2(n19446), .ZN(
        n19450) );
  AOI22_X1 U22497 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19448), .B1(
        n19778), .B2(n19512), .ZN(n19449) );
  OAI211_X1 U22498 ( .C1(n19783), .C2(n19473), .A(n19450), .B(n19449), .ZN(
        P3_U2899) );
  INV_X1 U22499 ( .A(n19808), .ZN(n19634) );
  NAND2_X1 U22500 ( .A1(n19634), .A2(n19522), .ZN(n19537) );
  NOR2_X1 U22501 ( .A1(n19512), .A2(n19539), .ZN(n19498) );
  NOR2_X1 U22502 ( .A1(n19688), .A2(n19498), .ZN(n19469) );
  AOI22_X1 U22503 ( .A1(n19689), .A2(n19462), .B1(n19725), .B2(n19469), .ZN(
        n19454) );
  OAI21_X1 U22504 ( .B1(n19451), .B2(n19588), .A(n19498), .ZN(n19452) );
  OAI211_X1 U22505 ( .C1(n19539), .C2(n19923), .A(n19591), .B(n19452), .ZN(
        n19470) );
  AOI22_X1 U22506 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19470), .B1(
        n19726), .B2(n19493), .ZN(n19453) );
  OAI211_X1 U22507 ( .C1(n19696), .C2(n19537), .A(n19454), .B(n19453), .ZN(
        P3_U2900) );
  AOI22_X1 U22508 ( .A1(n19737), .A2(n19493), .B1(n19736), .B2(n19469), .ZN(
        n19456) );
  AOI22_X1 U22509 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19470), .B1(
        n19738), .B2(n19462), .ZN(n19455) );
  OAI211_X1 U22510 ( .C1(n19741), .C2(n19537), .A(n19456), .B(n19455), .ZN(
        P3_U2901) );
  AOI22_X1 U22511 ( .A1(n19743), .A2(n19459), .B1(n19742), .B2(n19469), .ZN(
        n19458) );
  AOI22_X1 U22512 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19470), .B1(
        n19744), .B2(n19493), .ZN(n19457) );
  OAI211_X1 U22513 ( .C1(n19747), .C2(n19537), .A(n19458), .B(n19457), .ZN(
        P3_U2902) );
  AOI22_X1 U22514 ( .A1(n19749), .A2(n19459), .B1(n19748), .B2(n19469), .ZN(
        n19461) );
  AOI22_X1 U22515 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19470), .B1(
        n19701), .B2(n19481), .ZN(n19460) );
  OAI211_X1 U22516 ( .C1(n19704), .C2(n19537), .A(n19461), .B(n19460), .ZN(
        P3_U2903) );
  AOI22_X1 U22517 ( .A1(n19755), .A2(n19462), .B1(n19754), .B2(n19469), .ZN(
        n19464) );
  AOI22_X1 U22518 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19470), .B1(
        n19756), .B2(n19481), .ZN(n19463) );
  OAI211_X1 U22519 ( .C1(n19759), .C2(n19537), .A(n19464), .B(n19463), .ZN(
        P3_U2904) );
  AOI22_X1 U22520 ( .A1(n19762), .A2(n19493), .B1(n19760), .B2(n19469), .ZN(
        n19466) );
  AOI22_X1 U22521 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19470), .B1(
        n19677), .B2(n19539), .ZN(n19465) );
  OAI211_X1 U22522 ( .C1(n19680), .C2(n19473), .A(n19466), .B(n19465), .ZN(
        P3_U2905) );
  AOI22_X1 U22523 ( .A1(n19713), .A2(n19493), .B1(n19768), .B2(n19469), .ZN(
        n19468) );
  AOI22_X1 U22524 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19470), .B1(
        n19770), .B2(n19539), .ZN(n19467) );
  OAI211_X1 U22525 ( .C1(n19716), .C2(n19473), .A(n19468), .B(n19467), .ZN(
        P3_U2906) );
  INV_X1 U22526 ( .A(n19777), .ZN(n19724) );
  INV_X1 U22527 ( .A(n19783), .ZN(n19718) );
  AOI22_X1 U22528 ( .A1(n19718), .A2(n19493), .B1(n19775), .B2(n19469), .ZN(
        n19472) );
  AOI22_X1 U22529 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19470), .B1(
        n19778), .B2(n19539), .ZN(n19471) );
  OAI211_X1 U22530 ( .C1(n19724), .C2(n19473), .A(n19472), .B(n19471), .ZN(
        P3_U2907) );
  NAND2_X1 U22531 ( .A1(n19522), .A2(n19474), .ZN(n19557) );
  INV_X1 U22532 ( .A(n19522), .ZN(n19520) );
  NOR2_X1 U22533 ( .A1(n19520), .A2(n19660), .ZN(n19492) );
  AOI22_X1 U22534 ( .A1(n19725), .A2(n19492), .B1(n19726), .B2(n19512), .ZN(
        n19478) );
  NOR2_X1 U22535 ( .A1(n19806), .A2(n19475), .ZN(n19476) );
  AOI22_X1 U22536 ( .A1(n19730), .A2(n19476), .B1(n19522), .B2(n19662), .ZN(
        n19494) );
  AOI22_X1 U22537 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19494), .B1(
        n19689), .B2(n19493), .ZN(n19477) );
  OAI211_X1 U22538 ( .C1(n19696), .C2(n19557), .A(n19478), .B(n19477), .ZN(
        P3_U2908) );
  AOI22_X1 U22539 ( .A1(n19738), .A2(n19493), .B1(n19736), .B2(n19492), .ZN(
        n19480) );
  AOI22_X1 U22540 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19494), .B1(
        n19737), .B2(n19512), .ZN(n19479) );
  OAI211_X1 U22541 ( .C1(n19741), .C2(n19557), .A(n19480), .B(n19479), .ZN(
        P3_U2909) );
  AOI22_X1 U22542 ( .A1(n19744), .A2(n19512), .B1(n19742), .B2(n19492), .ZN(
        n19483) );
  AOI22_X1 U22543 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19494), .B1(
        n19743), .B2(n19481), .ZN(n19482) );
  OAI211_X1 U22544 ( .C1(n19747), .C2(n19557), .A(n19483), .B(n19482), .ZN(
        P3_U2910) );
  AOI22_X1 U22545 ( .A1(n19701), .A2(n19512), .B1(n19748), .B2(n19492), .ZN(
        n19485) );
  AOI22_X1 U22546 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19494), .B1(
        n19749), .B2(n19493), .ZN(n19484) );
  OAI211_X1 U22547 ( .C1(n19704), .C2(n19557), .A(n19485), .B(n19484), .ZN(
        P3_U2911) );
  AOI22_X1 U22548 ( .A1(n19755), .A2(n19493), .B1(n19754), .B2(n19492), .ZN(
        n19487) );
  AOI22_X1 U22549 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19494), .B1(
        n19756), .B2(n19512), .ZN(n19486) );
  OAI211_X1 U22550 ( .C1(n19759), .C2(n19557), .A(n19487), .B(n19486), .ZN(
        P3_U2912) );
  INV_X1 U22551 ( .A(n19677), .ZN(n19766) );
  INV_X1 U22552 ( .A(n19680), .ZN(n19761) );
  AOI22_X1 U22553 ( .A1(n19761), .A2(n19493), .B1(n19760), .B2(n19492), .ZN(
        n19489) );
  AOI22_X1 U22554 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19494), .B1(
        n19762), .B2(n19512), .ZN(n19488) );
  OAI211_X1 U22555 ( .C1(n19766), .C2(n19557), .A(n19489), .B(n19488), .ZN(
        P3_U2913) );
  AOI22_X1 U22556 ( .A1(n19769), .A2(n19493), .B1(n19768), .B2(n19492), .ZN(
        n19491) );
  AOI22_X1 U22557 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19494), .B1(
        n19770), .B2(n19561), .ZN(n19490) );
  OAI211_X1 U22558 ( .C1(n19773), .C2(n19519), .A(n19491), .B(n19490), .ZN(
        P3_U2914) );
  AOI22_X1 U22559 ( .A1(n19777), .A2(n19493), .B1(n19775), .B2(n19492), .ZN(
        n19496) );
  AOI22_X1 U22560 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19494), .B1(
        n19778), .B2(n19561), .ZN(n19495) );
  OAI211_X1 U22561 ( .C1(n19783), .C2(n19519), .A(n19496), .B(n19495), .ZN(
        P3_U2915) );
  NOR2_X1 U22562 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19497), .ZN(
        n19566) );
  NAND2_X1 U22563 ( .A1(n19566), .A2(n19587), .ZN(n19582) );
  AOI21_X1 U22564 ( .B1(n19557), .B2(n19582), .A(n19688), .ZN(n19515) );
  AOI22_X1 U22565 ( .A1(n19725), .A2(n19515), .B1(n19726), .B2(n19539), .ZN(
        n19501) );
  INV_X1 U22566 ( .A(n19582), .ZN(n19583) );
  AOI221_X1 U22567 ( .B1(n19498), .B2(n19557), .C1(n19588), .C2(n19557), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19499) );
  OAI21_X1 U22568 ( .B1(n19583), .B2(n19499), .A(n19591), .ZN(n19516) );
  AOI22_X1 U22569 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19516), .B1(
        n19731), .B2(n19583), .ZN(n19500) );
  OAI211_X1 U22570 ( .C1(n19735), .C2(n19519), .A(n19501), .B(n19500), .ZN(
        P3_U2916) );
  AOI22_X1 U22571 ( .A1(n19737), .A2(n19539), .B1(n19736), .B2(n19515), .ZN(
        n19503) );
  AOI22_X1 U22572 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19516), .B1(
        n19738), .B2(n19512), .ZN(n19502) );
  OAI211_X1 U22573 ( .C1(n19741), .C2(n19582), .A(n19503), .B(n19502), .ZN(
        P3_U2917) );
  AOI22_X1 U22574 ( .A1(n19744), .A2(n19539), .B1(n19742), .B2(n19515), .ZN(
        n19505) );
  AOI22_X1 U22575 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19516), .B1(
        n19642), .B2(n19583), .ZN(n19504) );
  OAI211_X1 U22576 ( .C1(n19645), .C2(n19519), .A(n19505), .B(n19504), .ZN(
        P3_U2918) );
  AOI22_X1 U22577 ( .A1(n19701), .A2(n19539), .B1(n19748), .B2(n19515), .ZN(
        n19507) );
  AOI22_X1 U22578 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19516), .B1(
        n19749), .B2(n19512), .ZN(n19506) );
  OAI211_X1 U22579 ( .C1(n19704), .C2(n19582), .A(n19507), .B(n19506), .ZN(
        P3_U2919) );
  AOI22_X1 U22580 ( .A1(n19755), .A2(n19512), .B1(n19754), .B2(n19515), .ZN(
        n19509) );
  AOI22_X1 U22581 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19516), .B1(
        n19756), .B2(n19539), .ZN(n19508) );
  OAI211_X1 U22582 ( .C1(n19759), .C2(n19582), .A(n19509), .B(n19508), .ZN(
        P3_U2920) );
  AOI22_X1 U22583 ( .A1(n19762), .A2(n19539), .B1(n19760), .B2(n19515), .ZN(
        n19511) );
  AOI22_X1 U22584 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19516), .B1(
        n19677), .B2(n19583), .ZN(n19510) );
  OAI211_X1 U22585 ( .C1(n19680), .C2(n19519), .A(n19511), .B(n19510), .ZN(
        P3_U2921) );
  AOI22_X1 U22586 ( .A1(n19769), .A2(n19512), .B1(n19768), .B2(n19515), .ZN(
        n19514) );
  AOI22_X1 U22587 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19516), .B1(
        n19770), .B2(n19583), .ZN(n19513) );
  OAI211_X1 U22588 ( .C1(n19773), .C2(n19537), .A(n19514), .B(n19513), .ZN(
        P3_U2922) );
  AOI22_X1 U22589 ( .A1(n19718), .A2(n19539), .B1(n19775), .B2(n19515), .ZN(
        n19518) );
  AOI22_X1 U22590 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19516), .B1(
        n19778), .B2(n19583), .ZN(n19517) );
  OAI211_X1 U22591 ( .C1(n19724), .C2(n19519), .A(n19518), .B(n19517), .ZN(
        P3_U2923) );
  NOR2_X2 U22592 ( .A1(n19800), .A2(n19520), .ZN(n19609) );
  INV_X1 U22593 ( .A(n19609), .ZN(n19604) );
  AND2_X1 U22594 ( .A1(n19836), .A2(n19566), .ZN(n19538) );
  AOI22_X1 U22595 ( .A1(n19689), .A2(n19539), .B1(n19725), .B2(n19538), .ZN(
        n19524) );
  NAND2_X1 U22596 ( .A1(n19522), .A2(n19521), .ZN(n19540) );
  AOI22_X1 U22597 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19540), .B1(
        n19726), .B2(n19561), .ZN(n19523) );
  OAI211_X1 U22598 ( .C1(n19696), .C2(n19604), .A(n19524), .B(n19523), .ZN(
        P3_U2924) );
  AOI22_X1 U22599 ( .A1(n19738), .A2(n19539), .B1(n19736), .B2(n19538), .ZN(
        n19526) );
  AOI22_X1 U22600 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19540), .B1(
        n19737), .B2(n19561), .ZN(n19525) );
  OAI211_X1 U22601 ( .C1(n19741), .C2(n19604), .A(n19526), .B(n19525), .ZN(
        P3_U2925) );
  AOI22_X1 U22602 ( .A1(n19743), .A2(n19539), .B1(n19742), .B2(n19538), .ZN(
        n19528) );
  AOI22_X1 U22603 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19540), .B1(
        n19744), .B2(n19561), .ZN(n19527) );
  OAI211_X1 U22604 ( .C1(n19747), .C2(n19604), .A(n19528), .B(n19527), .ZN(
        P3_U2926) );
  AOI22_X1 U22605 ( .A1(n19701), .A2(n19561), .B1(n19748), .B2(n19538), .ZN(
        n19530) );
  AOI22_X1 U22606 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19540), .B1(
        n19749), .B2(n19539), .ZN(n19529) );
  OAI211_X1 U22607 ( .C1(n19704), .C2(n19604), .A(n19530), .B(n19529), .ZN(
        P3_U2927) );
  AOI22_X1 U22608 ( .A1(n19756), .A2(n19561), .B1(n19754), .B2(n19538), .ZN(
        n19532) );
  AOI22_X1 U22609 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19540), .B1(
        n19755), .B2(n19539), .ZN(n19531) );
  OAI211_X1 U22610 ( .C1(n19759), .C2(n19604), .A(n19532), .B(n19531), .ZN(
        P3_U2928) );
  AOI22_X1 U22611 ( .A1(n19762), .A2(n19561), .B1(n19760), .B2(n19538), .ZN(
        n19534) );
  AOI22_X1 U22612 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19540), .B1(
        n19761), .B2(n19539), .ZN(n19533) );
  OAI211_X1 U22613 ( .C1(n19766), .C2(n19604), .A(n19534), .B(n19533), .ZN(
        P3_U2929) );
  AOI22_X1 U22614 ( .A1(n19713), .A2(n19561), .B1(n19768), .B2(n19538), .ZN(
        n19536) );
  AOI22_X1 U22615 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19540), .B1(
        n19770), .B2(n19609), .ZN(n19535) );
  OAI211_X1 U22616 ( .C1(n19716), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P3_U2930) );
  AOI22_X1 U22617 ( .A1(n19777), .A2(n19539), .B1(n19775), .B2(n19538), .ZN(
        n19542) );
  AOI22_X1 U22618 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19540), .B1(
        n19778), .B2(n19609), .ZN(n19541) );
  OAI211_X1 U22619 ( .C1(n19783), .C2(n19557), .A(n19542), .B(n19541), .ZN(
        P3_U2931) );
  NAND2_X1 U22620 ( .A1(n19634), .A2(n19565), .ZN(n19633) );
  NOR2_X1 U22621 ( .A1(n19609), .A2(n19626), .ZN(n19589) );
  NOR2_X1 U22622 ( .A1(n19688), .A2(n19589), .ZN(n19560) );
  AOI22_X1 U22623 ( .A1(n19689), .A2(n19561), .B1(n19725), .B2(n19560), .ZN(
        n19546) );
  NOR2_X1 U22624 ( .A1(n19561), .A2(n19583), .ZN(n19543) );
  OAI21_X1 U22625 ( .B1(n19543), .B2(n19588), .A(n19589), .ZN(n19544) );
  OAI211_X1 U22626 ( .C1(n19626), .C2(n19923), .A(n19591), .B(n19544), .ZN(
        n19562) );
  AOI22_X1 U22627 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19562), .B1(
        n19726), .B2(n19583), .ZN(n19545) );
  OAI211_X1 U22628 ( .C1(n19696), .C2(n19633), .A(n19546), .B(n19545), .ZN(
        P3_U2932) );
  AOI22_X1 U22629 ( .A1(n19738), .A2(n19561), .B1(n19736), .B2(n19560), .ZN(
        n19548) );
  AOI22_X1 U22630 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19562), .B1(
        n19667), .B2(n19626), .ZN(n19547) );
  OAI211_X1 U22631 ( .C1(n19670), .C2(n19582), .A(n19548), .B(n19547), .ZN(
        P3_U2933) );
  AOI22_X1 U22632 ( .A1(n19744), .A2(n19583), .B1(n19742), .B2(n19560), .ZN(
        n19550) );
  AOI22_X1 U22633 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19562), .B1(
        n19642), .B2(n19626), .ZN(n19549) );
  OAI211_X1 U22634 ( .C1(n19645), .C2(n19557), .A(n19550), .B(n19549), .ZN(
        P3_U2934) );
  AOI22_X1 U22635 ( .A1(n19749), .A2(n19561), .B1(n19748), .B2(n19560), .ZN(
        n19552) );
  AOI22_X1 U22636 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19562), .B1(
        n19750), .B2(n19626), .ZN(n19551) );
  OAI211_X1 U22637 ( .C1(n19753), .C2(n19582), .A(n19552), .B(n19551), .ZN(
        P3_U2935) );
  AOI22_X1 U22638 ( .A1(n19755), .A2(n19561), .B1(n19754), .B2(n19560), .ZN(
        n19554) );
  AOI22_X1 U22639 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19562), .B1(
        n19756), .B2(n19583), .ZN(n19553) );
  OAI211_X1 U22640 ( .C1(n19759), .C2(n19633), .A(n19554), .B(n19553), .ZN(
        P3_U2936) );
  AOI22_X1 U22641 ( .A1(n19762), .A2(n19583), .B1(n19760), .B2(n19560), .ZN(
        n19556) );
  AOI22_X1 U22642 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19562), .B1(
        n19677), .B2(n19626), .ZN(n19555) );
  OAI211_X1 U22643 ( .C1(n19680), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P3_U2937) );
  AOI22_X1 U22644 ( .A1(n19769), .A2(n19561), .B1(n19768), .B2(n19560), .ZN(
        n19559) );
  AOI22_X1 U22645 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19562), .B1(
        n19770), .B2(n19626), .ZN(n19558) );
  OAI211_X1 U22646 ( .C1(n19773), .C2(n19582), .A(n19559), .B(n19558), .ZN(
        P3_U2938) );
  AOI22_X1 U22647 ( .A1(n19777), .A2(n19561), .B1(n19775), .B2(n19560), .ZN(
        n19564) );
  AOI22_X1 U22648 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19562), .B1(
        n19778), .B2(n19626), .ZN(n19563) );
  OAI211_X1 U22649 ( .C1(n19783), .C2(n19582), .A(n19564), .B(n19563), .ZN(
        P3_U2939) );
  INV_X1 U22650 ( .A(n19565), .ZN(n19613) );
  NOR2_X1 U22651 ( .A1(n19613), .A2(n19660), .ZN(n19612) );
  AOI22_X1 U22652 ( .A1(n19725), .A2(n19612), .B1(n19726), .B2(n19609), .ZN(
        n19569) );
  AOI22_X1 U22653 ( .A1(n19730), .A2(n19566), .B1(n19565), .B2(n19662), .ZN(
        n19584) );
  NOR2_X2 U22654 ( .A1(n19613), .A2(n19567), .ZN(n19656) );
  AOI22_X1 U22655 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19584), .B1(
        n19731), .B2(n19656), .ZN(n19568) );
  OAI211_X1 U22656 ( .C1(n19735), .C2(n19582), .A(n19569), .B(n19568), .ZN(
        P3_U2940) );
  INV_X1 U22657 ( .A(n19656), .ZN(n19654) );
  AOI22_X1 U22658 ( .A1(n19737), .A2(n19609), .B1(n19736), .B2(n19612), .ZN(
        n19571) );
  AOI22_X1 U22659 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19584), .B1(
        n19738), .B2(n19583), .ZN(n19570) );
  OAI211_X1 U22660 ( .C1(n19741), .C2(n19654), .A(n19571), .B(n19570), .ZN(
        P3_U2941) );
  AOI22_X1 U22661 ( .A1(n19744), .A2(n19609), .B1(n19742), .B2(n19612), .ZN(
        n19573) );
  AOI22_X1 U22662 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19584), .B1(
        n19642), .B2(n19656), .ZN(n19572) );
  OAI211_X1 U22663 ( .C1(n19645), .C2(n19582), .A(n19573), .B(n19572), .ZN(
        P3_U2942) );
  AOI22_X1 U22664 ( .A1(n19701), .A2(n19609), .B1(n19748), .B2(n19612), .ZN(
        n19575) );
  AOI22_X1 U22665 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19584), .B1(
        n19749), .B2(n19583), .ZN(n19574) );
  OAI211_X1 U22666 ( .C1(n19704), .C2(n19654), .A(n19575), .B(n19574), .ZN(
        P3_U2943) );
  AOI22_X1 U22667 ( .A1(n19755), .A2(n19583), .B1(n19754), .B2(n19612), .ZN(
        n19577) );
  AOI22_X1 U22668 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19584), .B1(
        n19756), .B2(n19609), .ZN(n19576) );
  OAI211_X1 U22669 ( .C1(n19759), .C2(n19654), .A(n19577), .B(n19576), .ZN(
        P3_U2944) );
  AOI22_X1 U22670 ( .A1(n19762), .A2(n19609), .B1(n19760), .B2(n19612), .ZN(
        n19579) );
  AOI22_X1 U22671 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19584), .B1(
        n19677), .B2(n19656), .ZN(n19578) );
  OAI211_X1 U22672 ( .C1(n19680), .C2(n19582), .A(n19579), .B(n19578), .ZN(
        P3_U2945) );
  AOI22_X1 U22673 ( .A1(n19713), .A2(n19609), .B1(n19768), .B2(n19612), .ZN(
        n19581) );
  AOI22_X1 U22674 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19584), .B1(
        n19770), .B2(n19656), .ZN(n19580) );
  OAI211_X1 U22675 ( .C1(n19716), .C2(n19582), .A(n19581), .B(n19580), .ZN(
        P3_U2946) );
  AOI22_X1 U22676 ( .A1(n19777), .A2(n19583), .B1(n19775), .B2(n19612), .ZN(
        n19586) );
  AOI22_X1 U22677 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19584), .B1(
        n19778), .B2(n19656), .ZN(n19585) );
  OAI211_X1 U22678 ( .C1(n19783), .C2(n19604), .A(n19586), .B(n19585), .ZN(
        P3_U2947) );
  NOR2_X1 U22679 ( .A1(n19806), .A2(n19613), .ZN(n19664) );
  NAND2_X1 U22680 ( .A1(n19587), .A2(n19664), .ZN(n19687) );
  INV_X1 U22681 ( .A(n19687), .ZN(n19681) );
  NOR2_X1 U22682 ( .A1(n19656), .A2(n19681), .ZN(n19636) );
  OAI21_X1 U22683 ( .B1(n19589), .B2(n19588), .A(n19636), .ZN(n19590) );
  OAI211_X1 U22684 ( .C1(n19681), .C2(n19923), .A(n19591), .B(n19590), .ZN(
        n19608) );
  NOR2_X1 U22685 ( .A1(n19688), .A2(n19636), .ZN(n19607) );
  AOI22_X1 U22686 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19608), .B1(
        n19725), .B2(n19607), .ZN(n19593) );
  AOI22_X1 U22687 ( .A1(n19731), .A2(n19681), .B1(n19726), .B2(n19626), .ZN(
        n19592) );
  OAI211_X1 U22688 ( .C1(n19735), .C2(n19604), .A(n19593), .B(n19592), .ZN(
        P3_U2948) );
  AOI22_X1 U22689 ( .A1(n19738), .A2(n19609), .B1(n19736), .B2(n19607), .ZN(
        n19595) );
  AOI22_X1 U22690 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19608), .B1(
        n19667), .B2(n19681), .ZN(n19594) );
  OAI211_X1 U22691 ( .C1(n19670), .C2(n19633), .A(n19595), .B(n19594), .ZN(
        P3_U2949) );
  AOI22_X1 U22692 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19608), .B1(
        n19742), .B2(n19607), .ZN(n19597) );
  AOI22_X1 U22693 ( .A1(n19642), .A2(n19681), .B1(n19744), .B2(n19626), .ZN(
        n19596) );
  OAI211_X1 U22694 ( .C1(n19645), .C2(n19604), .A(n19597), .B(n19596), .ZN(
        P3_U2950) );
  AOI22_X1 U22695 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19608), .B1(
        n19748), .B2(n19607), .ZN(n19599) );
  AOI22_X1 U22696 ( .A1(n19750), .A2(n19681), .B1(n19749), .B2(n19609), .ZN(
        n19598) );
  OAI211_X1 U22697 ( .C1(n19753), .C2(n19633), .A(n19599), .B(n19598), .ZN(
        P3_U2951) );
  AOI22_X1 U22698 ( .A1(n19755), .A2(n19609), .B1(n19754), .B2(n19607), .ZN(
        n19601) );
  AOI22_X1 U22699 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19608), .B1(
        n19756), .B2(n19626), .ZN(n19600) );
  OAI211_X1 U22700 ( .C1(n19759), .C2(n19687), .A(n19601), .B(n19600), .ZN(
        P3_U2952) );
  AOI22_X1 U22701 ( .A1(n19762), .A2(n19626), .B1(n19760), .B2(n19607), .ZN(
        n19603) );
  AOI22_X1 U22702 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19608), .B1(
        n19677), .B2(n19681), .ZN(n19602) );
  OAI211_X1 U22703 ( .C1(n19680), .C2(n19604), .A(n19603), .B(n19602), .ZN(
        P3_U2953) );
  AOI22_X1 U22704 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19608), .B1(
        n19768), .B2(n19607), .ZN(n19606) );
  AOI22_X1 U22705 ( .A1(n19770), .A2(n19681), .B1(n19769), .B2(n19609), .ZN(
        n19605) );
  OAI211_X1 U22706 ( .C1(n19773), .C2(n19633), .A(n19606), .B(n19605), .ZN(
        P3_U2954) );
  AOI22_X1 U22707 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19608), .B1(
        n19775), .B2(n19607), .ZN(n19611) );
  AOI22_X1 U22708 ( .A1(n19778), .A2(n19681), .B1(n19777), .B2(n19609), .ZN(
        n19610) );
  OAI211_X1 U22709 ( .C1(n19783), .C2(n19633), .A(n19611), .B(n19610), .ZN(
        P3_U2955) );
  AND2_X1 U22710 ( .A1(n19836), .A2(n19664), .ZN(n19629) );
  AOI22_X1 U22711 ( .A1(n19725), .A2(n19629), .B1(n19726), .B2(n19656), .ZN(
        n19615) );
  AOI22_X1 U22712 ( .A1(n19730), .A2(n19612), .B1(n19727), .B2(n19664), .ZN(
        n19630) );
  NOR2_X2 U22713 ( .A1(n19800), .A2(n19613), .ZN(n19709) );
  AOI22_X1 U22714 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19630), .B1(
        n19731), .B2(n19709), .ZN(n19614) );
  OAI211_X1 U22715 ( .C1(n19735), .C2(n19633), .A(n19615), .B(n19614), .ZN(
        P3_U2956) );
  INV_X1 U22716 ( .A(n19709), .ZN(n19723) );
  AOI22_X1 U22717 ( .A1(n19737), .A2(n19656), .B1(n19736), .B2(n19629), .ZN(
        n19617) );
  AOI22_X1 U22718 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19630), .B1(
        n19738), .B2(n19626), .ZN(n19616) );
  OAI211_X1 U22719 ( .C1(n19741), .C2(n19723), .A(n19617), .B(n19616), .ZN(
        P3_U2957) );
  AOI22_X1 U22720 ( .A1(n19744), .A2(n19656), .B1(n19742), .B2(n19629), .ZN(
        n19619) );
  AOI22_X1 U22721 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19630), .B1(
        n19642), .B2(n19709), .ZN(n19618) );
  OAI211_X1 U22722 ( .C1(n19645), .C2(n19633), .A(n19619), .B(n19618), .ZN(
        P3_U2958) );
  AOI22_X1 U22723 ( .A1(n19749), .A2(n19626), .B1(n19748), .B2(n19629), .ZN(
        n19621) );
  AOI22_X1 U22724 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19630), .B1(
        n19750), .B2(n19709), .ZN(n19620) );
  OAI211_X1 U22725 ( .C1(n19753), .C2(n19654), .A(n19621), .B(n19620), .ZN(
        P3_U2959) );
  AOI22_X1 U22726 ( .A1(n19756), .A2(n19656), .B1(n19754), .B2(n19629), .ZN(
        n19623) );
  AOI22_X1 U22727 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19630), .B1(
        n19705), .B2(n19709), .ZN(n19622) );
  OAI211_X1 U22728 ( .C1(n19708), .C2(n19633), .A(n19623), .B(n19622), .ZN(
        P3_U2960) );
  AOI22_X1 U22729 ( .A1(n19761), .A2(n19626), .B1(n19760), .B2(n19629), .ZN(
        n19625) );
  AOI22_X1 U22730 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19630), .B1(
        n19762), .B2(n19656), .ZN(n19624) );
  OAI211_X1 U22731 ( .C1(n19766), .C2(n19723), .A(n19625), .B(n19624), .ZN(
        P3_U2961) );
  AOI22_X1 U22732 ( .A1(n19769), .A2(n19626), .B1(n19768), .B2(n19629), .ZN(
        n19628) );
  AOI22_X1 U22733 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19630), .B1(
        n19770), .B2(n19709), .ZN(n19627) );
  OAI211_X1 U22734 ( .C1(n19773), .C2(n19654), .A(n19628), .B(n19627), .ZN(
        P3_U2962) );
  AOI22_X1 U22735 ( .A1(n19718), .A2(n19656), .B1(n19775), .B2(n19629), .ZN(
        n19632) );
  AOI22_X1 U22736 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19630), .B1(
        n19778), .B2(n19709), .ZN(n19631) );
  OAI211_X1 U22737 ( .C1(n19724), .C2(n19633), .A(n19632), .B(n19631), .ZN(
        P3_U2963) );
  NAND2_X1 U22738 ( .A1(n19634), .A2(n19663), .ZN(n19734) );
  INV_X1 U22739 ( .A(n19734), .ZN(n19776) );
  NOR2_X1 U22740 ( .A1(n19709), .A2(n19776), .ZN(n19691) );
  NOR2_X1 U22741 ( .A1(n19688), .A2(n19691), .ZN(n19655) );
  AOI22_X1 U22742 ( .A1(n19689), .A2(n19656), .B1(n19725), .B2(n19655), .ZN(
        n19639) );
  OAI22_X1 U22743 ( .A1(n19636), .A2(n19690), .B1(n19691), .B2(n19635), .ZN(
        n19637) );
  OAI21_X1 U22744 ( .B1(n19776), .B2(n19923), .A(n19637), .ZN(n19657) );
  AOI22_X1 U22745 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19657), .B1(
        n19726), .B2(n19681), .ZN(n19638) );
  OAI211_X1 U22746 ( .C1(n19696), .C2(n19734), .A(n19639), .B(n19638), .ZN(
        P3_U2964) );
  AOI22_X1 U22747 ( .A1(n19737), .A2(n19681), .B1(n19736), .B2(n19655), .ZN(
        n19641) );
  AOI22_X1 U22748 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19657), .B1(
        n19738), .B2(n19656), .ZN(n19640) );
  OAI211_X1 U22749 ( .C1(n19741), .C2(n19734), .A(n19641), .B(n19640), .ZN(
        P3_U2965) );
  AOI22_X1 U22750 ( .A1(n19744), .A2(n19681), .B1(n19742), .B2(n19655), .ZN(
        n19644) );
  AOI22_X1 U22751 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19657), .B1(
        n19642), .B2(n19776), .ZN(n19643) );
  OAI211_X1 U22752 ( .C1(n19645), .C2(n19654), .A(n19644), .B(n19643), .ZN(
        P3_U2966) );
  AOI22_X1 U22753 ( .A1(n19749), .A2(n19656), .B1(n19748), .B2(n19655), .ZN(
        n19647) );
  AOI22_X1 U22754 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19657), .B1(
        n19750), .B2(n19776), .ZN(n19646) );
  OAI211_X1 U22755 ( .C1(n19753), .C2(n19687), .A(n19647), .B(n19646), .ZN(
        P3_U2967) );
  AOI22_X1 U22756 ( .A1(n19755), .A2(n19656), .B1(n19754), .B2(n19655), .ZN(
        n19649) );
  AOI22_X1 U22757 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19657), .B1(
        n19756), .B2(n19681), .ZN(n19648) );
  OAI211_X1 U22758 ( .C1(n19759), .C2(n19734), .A(n19649), .B(n19648), .ZN(
        P3_U2968) );
  AOI22_X1 U22759 ( .A1(n19762), .A2(n19681), .B1(n19760), .B2(n19655), .ZN(
        n19651) );
  AOI22_X1 U22760 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19657), .B1(
        n19677), .B2(n19776), .ZN(n19650) );
  OAI211_X1 U22761 ( .C1(n19680), .C2(n19654), .A(n19651), .B(n19650), .ZN(
        P3_U2969) );
  AOI22_X1 U22762 ( .A1(n19713), .A2(n19681), .B1(n19768), .B2(n19655), .ZN(
        n19653) );
  AOI22_X1 U22763 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19657), .B1(
        n19770), .B2(n19776), .ZN(n19652) );
  OAI211_X1 U22764 ( .C1(n19716), .C2(n19654), .A(n19653), .B(n19652), .ZN(
        P3_U2970) );
  AOI22_X1 U22765 ( .A1(n19777), .A2(n19656), .B1(n19775), .B2(n19655), .ZN(
        n19659) );
  AOI22_X1 U22766 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19657), .B1(
        n19778), .B2(n19776), .ZN(n19658) );
  OAI211_X1 U22767 ( .C1(n19783), .C2(n19687), .A(n19659), .B(n19658), .ZN(
        P3_U2971) );
  NOR2_X1 U22768 ( .A1(n19661), .A2(n19660), .ZN(n19729) );
  AOI22_X1 U22769 ( .A1(n19689), .A2(n19681), .B1(n19725), .B2(n19729), .ZN(
        n19666) );
  AOI22_X1 U22770 ( .A1(n19730), .A2(n19664), .B1(n19663), .B2(n19662), .ZN(
        n19684) );
  AOI22_X1 U22771 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19684), .B1(
        n19726), .B2(n19709), .ZN(n19665) );
  OAI211_X1 U22772 ( .C1(n19784), .C2(n19696), .A(n19666), .B(n19665), .ZN(
        P3_U2972) );
  AOI22_X1 U22773 ( .A1(n19738), .A2(n19681), .B1(n19736), .B2(n19729), .ZN(
        n19669) );
  AOI22_X1 U22774 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19684), .B1(
        n19763), .B2(n19667), .ZN(n19668) );
  OAI211_X1 U22775 ( .C1(n19670), .C2(n19723), .A(n19669), .B(n19668), .ZN(
        P3_U2973) );
  AOI22_X1 U22776 ( .A1(n19743), .A2(n19681), .B1(n19742), .B2(n19729), .ZN(
        n19672) );
  AOI22_X1 U22777 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19684), .B1(
        n19744), .B2(n19709), .ZN(n19671) );
  OAI211_X1 U22778 ( .C1(n19784), .C2(n19747), .A(n19672), .B(n19671), .ZN(
        P3_U2974) );
  AOI22_X1 U22779 ( .A1(n19749), .A2(n19681), .B1(n19748), .B2(n19729), .ZN(
        n19674) );
  AOI22_X1 U22780 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19684), .B1(
        n19763), .B2(n19750), .ZN(n19673) );
  OAI211_X1 U22781 ( .C1(n19753), .C2(n19723), .A(n19674), .B(n19673), .ZN(
        P3_U2975) );
  AOI22_X1 U22782 ( .A1(n19755), .A2(n19681), .B1(n19754), .B2(n19729), .ZN(
        n19676) );
  AOI22_X1 U22783 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19684), .B1(
        n19756), .B2(n19709), .ZN(n19675) );
  OAI211_X1 U22784 ( .C1(n19784), .C2(n19759), .A(n19676), .B(n19675), .ZN(
        P3_U2976) );
  AOI22_X1 U22785 ( .A1(n19762), .A2(n19709), .B1(n19760), .B2(n19729), .ZN(
        n19679) );
  AOI22_X1 U22786 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19684), .B1(
        n19763), .B2(n19677), .ZN(n19678) );
  OAI211_X1 U22787 ( .C1(n19680), .C2(n19687), .A(n19679), .B(n19678), .ZN(
        P3_U2977) );
  AOI22_X1 U22788 ( .A1(n19769), .A2(n19681), .B1(n19768), .B2(n19729), .ZN(
        n19683) );
  AOI22_X1 U22789 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19684), .B1(
        n19763), .B2(n19770), .ZN(n19682) );
  OAI211_X1 U22790 ( .C1(n19773), .C2(n19723), .A(n19683), .B(n19682), .ZN(
        P3_U2978) );
  AOI22_X1 U22791 ( .A1(n19718), .A2(n19709), .B1(n19775), .B2(n19729), .ZN(
        n19686) );
  AOI22_X1 U22792 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19684), .B1(
        n19763), .B2(n19778), .ZN(n19685) );
  OAI211_X1 U22793 ( .C1(n19724), .C2(n19687), .A(n19686), .B(n19685), .ZN(
        P3_U2979) );
  AOI21_X1 U22794 ( .B1(n19784), .B2(n19712), .A(n19688), .ZN(n19717) );
  AOI22_X1 U22795 ( .A1(n19689), .A2(n19709), .B1(n19725), .B2(n19717), .ZN(
        n19695) );
  NOR2_X1 U22796 ( .A1(n19691), .A2(n19690), .ZN(n19692) );
  OAI22_X1 U22797 ( .A1(n19719), .A2(n19923), .B1(n19693), .B2(n19692), .ZN(
        n19720) );
  AOI22_X1 U22798 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19720), .B1(
        n19726), .B2(n19776), .ZN(n19694) );
  OAI211_X1 U22799 ( .C1(n19712), .C2(n19696), .A(n19695), .B(n19694), .ZN(
        P3_U2980) );
  AOI22_X1 U22800 ( .A1(n19737), .A2(n19776), .B1(n19736), .B2(n19717), .ZN(
        n19698) );
  AOI22_X1 U22801 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19720), .B1(
        n19738), .B2(n19709), .ZN(n19697) );
  OAI211_X1 U22802 ( .C1(n19712), .C2(n19741), .A(n19698), .B(n19697), .ZN(
        P3_U2981) );
  AOI22_X1 U22803 ( .A1(n19743), .A2(n19709), .B1(n19742), .B2(n19717), .ZN(
        n19700) );
  AOI22_X1 U22804 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19720), .B1(
        n19744), .B2(n19776), .ZN(n19699) );
  OAI211_X1 U22805 ( .C1(n19712), .C2(n19747), .A(n19700), .B(n19699), .ZN(
        P3_U2982) );
  AOI22_X1 U22806 ( .A1(n19701), .A2(n19776), .B1(n19748), .B2(n19717), .ZN(
        n19703) );
  AOI22_X1 U22807 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19720), .B1(
        n19749), .B2(n19709), .ZN(n19702) );
  OAI211_X1 U22808 ( .C1(n19712), .C2(n19704), .A(n19703), .B(n19702), .ZN(
        P3_U2983) );
  AOI22_X1 U22809 ( .A1(n19756), .A2(n19776), .B1(n19754), .B2(n19717), .ZN(
        n19707) );
  AOI22_X1 U22810 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n19705), .ZN(n19706) );
  OAI211_X1 U22811 ( .C1(n19708), .C2(n19723), .A(n19707), .B(n19706), .ZN(
        P3_U2984) );
  AOI22_X1 U22812 ( .A1(n19761), .A2(n19709), .B1(n19760), .B2(n19717), .ZN(
        n19711) );
  AOI22_X1 U22813 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19720), .B1(
        n19762), .B2(n19776), .ZN(n19710) );
  OAI211_X1 U22814 ( .C1(n19712), .C2(n19766), .A(n19711), .B(n19710), .ZN(
        P3_U2985) );
  AOI22_X1 U22815 ( .A1(n19713), .A2(n19776), .B1(n19768), .B2(n19717), .ZN(
        n19715) );
  AOI22_X1 U22816 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n19770), .ZN(n19714) );
  OAI211_X1 U22817 ( .C1(n19716), .C2(n19723), .A(n19715), .B(n19714), .ZN(
        P3_U2986) );
  AOI22_X1 U22818 ( .A1(n19718), .A2(n19776), .B1(n19775), .B2(n19717), .ZN(
        n19722) );
  AOI22_X1 U22819 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19720), .B1(
        n19719), .B2(n19778), .ZN(n19721) );
  OAI211_X1 U22820 ( .C1(n19724), .C2(n19723), .A(n19722), .B(n19721), .ZN(
        P3_U2987) );
  AND2_X1 U22821 ( .A1(n19836), .A2(n19728), .ZN(n19774) );
  AOI22_X1 U22822 ( .A1(n19763), .A2(n19726), .B1(n19725), .B2(n19774), .ZN(
        n19733) );
  AOI22_X1 U22823 ( .A1(n19730), .A2(n19729), .B1(n19728), .B2(n19727), .ZN(
        n19780) );
  AOI22_X1 U22824 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19780), .B1(
        n19779), .B2(n19731), .ZN(n19732) );
  OAI211_X1 U22825 ( .C1(n19735), .C2(n19734), .A(n19733), .B(n19732), .ZN(
        P3_U2988) );
  AOI22_X1 U22826 ( .A1(n19763), .A2(n19737), .B1(n19736), .B2(n19774), .ZN(
        n19740) );
  AOI22_X1 U22827 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19780), .B1(
        n19738), .B2(n19776), .ZN(n19739) );
  OAI211_X1 U22828 ( .C1(n19767), .C2(n19741), .A(n19740), .B(n19739), .ZN(
        P3_U2989) );
  AOI22_X1 U22829 ( .A1(n19743), .A2(n19776), .B1(n19742), .B2(n19774), .ZN(
        n19746) );
  AOI22_X1 U22830 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19780), .B1(
        n19763), .B2(n19744), .ZN(n19745) );
  OAI211_X1 U22831 ( .C1(n19767), .C2(n19747), .A(n19746), .B(n19745), .ZN(
        P3_U2990) );
  AOI22_X1 U22832 ( .A1(n19749), .A2(n19776), .B1(n19748), .B2(n19774), .ZN(
        n19752) );
  AOI22_X1 U22833 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19780), .B1(
        n19779), .B2(n19750), .ZN(n19751) );
  OAI211_X1 U22834 ( .C1(n19784), .C2(n19753), .A(n19752), .B(n19751), .ZN(
        P3_U2991) );
  AOI22_X1 U22835 ( .A1(n19755), .A2(n19776), .B1(n19754), .B2(n19774), .ZN(
        n19758) );
  AOI22_X1 U22836 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19780), .B1(
        n19763), .B2(n19756), .ZN(n19757) );
  OAI211_X1 U22837 ( .C1(n19767), .C2(n19759), .A(n19758), .B(n19757), .ZN(
        P3_U2992) );
  AOI22_X1 U22838 ( .A1(n19761), .A2(n19776), .B1(n19760), .B2(n19774), .ZN(
        n19765) );
  AOI22_X1 U22839 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19780), .B1(
        n19763), .B2(n19762), .ZN(n19764) );
  OAI211_X1 U22840 ( .C1(n19767), .C2(n19766), .A(n19765), .B(n19764), .ZN(
        P3_U2993) );
  AOI22_X1 U22841 ( .A1(n19769), .A2(n19776), .B1(n19768), .B2(n19774), .ZN(
        n19772) );
  AOI22_X1 U22842 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19780), .B1(
        n19779), .B2(n19770), .ZN(n19771) );
  OAI211_X1 U22843 ( .C1(n19784), .C2(n19773), .A(n19772), .B(n19771), .ZN(
        P3_U2994) );
  AOI22_X1 U22844 ( .A1(n19777), .A2(n19776), .B1(n19775), .B2(n19774), .ZN(
        n19782) );
  AOI22_X1 U22845 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19780), .B1(
        n19779), .B2(n19778), .ZN(n19781) );
  OAI211_X1 U22846 ( .C1(n19784), .C2(n19783), .A(n19782), .B(n19781), .ZN(
        P3_U2995) );
  NOR2_X1 U22847 ( .A1(n19787), .A2(n19786), .ZN(n19790) );
  OAI222_X1 U22848 ( .A1(n19791), .A2(n10238), .B1(n9870), .B2(n19790), .C1(
        n19789), .C2(n19788), .ZN(n19936) );
  OAI21_X1 U22849 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19792), .ZN(n19794) );
  OAI211_X1 U22850 ( .C1(n19798), .C2(n21661), .A(n19794), .B(n19793), .ZN(
        n19819) );
  OR2_X1 U22851 ( .A1(n19809), .A2(n19795), .ZN(n19796) );
  AOI22_X1 U22852 ( .A1(n19798), .A2(n19797), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19796), .ZN(n19817) );
  MUX2_X1 U22853 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n19799), .S(
        n19798), .Z(n19812) );
  INV_X1 U22854 ( .A(n19805), .ZN(n19803) );
  INV_X1 U22855 ( .A(n19800), .ZN(n19802) );
  AOI21_X1 U22856 ( .B1(n19803), .B2(n19802), .A(n19801), .ZN(n19804) );
  AOI21_X1 U22857 ( .B1(n19806), .B2(n19805), .A(n19804), .ZN(n19810) );
  NAND2_X1 U22858 ( .A1(n19812), .A2(n13797), .ZN(n19807) );
  OAI211_X1 U22859 ( .C1(n19810), .C2(n19809), .A(n19808), .B(n19807), .ZN(
        n19811) );
  OAI211_X1 U22860 ( .C1(n13797), .C2(n19812), .A(n19811), .B(n19814), .ZN(
        n19816) );
  AOI21_X1 U22861 ( .B1(n19814), .B2(n19813), .A(n19812), .ZN(n19815) );
  AOI222_X1 U22862 ( .A1(n19817), .A2(n19816), .B1(n19817), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19816), .C2(n19815), .ZN(
        n19818) );
  INV_X1 U22863 ( .A(n19842), .ZN(n19946) );
  AOI22_X1 U22864 ( .A1(n19821), .A2(n19946), .B1(n19844), .B2(n19940), .ZN(
        n19822) );
  INV_X1 U22865 ( .A(n19822), .ZN(n19827) );
  OAI211_X1 U22866 ( .C1(n19824), .C2(n19823), .A(n19938), .B(n19831), .ZN(
        n19922) );
  OAI21_X1 U22867 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19944), .A(n19922), 
        .ZN(n19833) );
  NOR2_X1 U22868 ( .A1(n19825), .A2(n19833), .ZN(n19826) );
  MUX2_X1 U22869 ( .A(n19827), .B(n19826), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19829) );
  OAI211_X1 U22870 ( .C1(n19831), .C2(n19830), .A(n19829), .B(n19828), .ZN(
        P3_U2996) );
  NAND2_X1 U22871 ( .A1(n19844), .A2(n19940), .ZN(n19838) );
  NAND4_X1 U22872 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n19844), .A4(n19832), .ZN(n19840) );
  INV_X1 U22873 ( .A(n19833), .ZN(n19834) );
  NAND3_X1 U22874 ( .A1(n19836), .A2(n19835), .A3(n19834), .ZN(n19837) );
  NAND4_X1 U22875 ( .A1(n19839), .A2(n19838), .A3(n19840), .A4(n19837), .ZN(
        P3_U2997) );
  AND4_X1 U22876 ( .A1(n19842), .A2(n19841), .A3(n19840), .A4(n19921), .ZN(
        P3_U2998) );
  INV_X1 U22877 ( .A(P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21739) );
  NOR2_X1 U22878 ( .A1(n21739), .A2(n19920), .ZN(P3_U2999) );
  AND2_X1 U22879 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19917), .ZN(
        P3_U3000) );
  AND2_X1 U22880 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19917), .ZN(
        P3_U3001) );
  AND2_X1 U22881 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19917), .ZN(
        P3_U3002) );
  AND2_X1 U22882 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19917), .ZN(
        P3_U3003) );
  AND2_X1 U22883 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19917), .ZN(
        P3_U3004) );
  AND2_X1 U22884 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19917), .ZN(
        P3_U3005) );
  AND2_X1 U22885 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19917), .ZN(
        P3_U3006) );
  AND2_X1 U22886 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19917), .ZN(
        P3_U3007) );
  AND2_X1 U22887 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19917), .ZN(
        P3_U3008) );
  AND2_X1 U22888 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19917), .ZN(
        P3_U3009) );
  AND2_X1 U22889 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19917), .ZN(
        P3_U3010) );
  AND2_X1 U22890 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19917), .ZN(
        P3_U3011) );
  AND2_X1 U22891 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19917), .ZN(
        P3_U3012) );
  INV_X1 U22892 ( .A(P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21844) );
  NOR2_X1 U22893 ( .A1(n21844), .A2(n19920), .ZN(P3_U3013) );
  AND2_X1 U22894 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19917), .ZN(
        P3_U3014) );
  AND2_X1 U22895 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19917), .ZN(
        P3_U3015) );
  AND2_X1 U22896 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19917), .ZN(
        P3_U3016) );
  AND2_X1 U22897 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19917), .ZN(
        P3_U3017) );
  AND2_X1 U22898 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19917), .ZN(
        P3_U3018) );
  AND2_X1 U22899 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19917), .ZN(
        P3_U3019) );
  AND2_X1 U22900 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19917), .ZN(
        P3_U3020) );
  AND2_X1 U22901 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19917), .ZN(P3_U3021) );
  AND2_X1 U22902 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19917), .ZN(P3_U3022) );
  AND2_X1 U22903 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19917), .ZN(P3_U3023) );
  INV_X1 U22904 ( .A(P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n21719) );
  NOR2_X1 U22905 ( .A1(n21719), .A2(n19920), .ZN(P3_U3024) );
  AND2_X1 U22906 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19917), .ZN(P3_U3025) );
  AND2_X1 U22907 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19917), .ZN(P3_U3026) );
  AND2_X1 U22908 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19917), .ZN(P3_U3027) );
  AND2_X1 U22909 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19917), .ZN(P3_U3028) );
  NOR2_X1 U22910 ( .A1(n19856), .A2(n21491), .ZN(n19851) );
  INV_X1 U22911 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19843) );
  AOI211_X1 U22912 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(HOLD), .A(n19851), .B(
        n19843), .ZN(n19847) );
  NAND2_X1 U22913 ( .A1(n19844), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19849) );
  AND2_X1 U22914 ( .A1(n19849), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n19855) );
  INV_X1 U22915 ( .A(NA), .ZN(n21485) );
  OAI21_X1 U22916 ( .B1(n21485), .B2(n19845), .A(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19854) );
  INV_X1 U22917 ( .A(n19854), .ZN(n19846) );
  OAI22_X1 U22918 ( .A1(n21589), .A2(n19847), .B1(n19855), .B2(n19846), .ZN(
        P3_U3029) );
  AOI22_X1 U22919 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .ZN(n19848) );
  OAI211_X1 U22920 ( .C1(n19851), .C2(n19848), .A(n19941), .B(n19849), .ZN(
        P3_U3030) );
  OAI22_X1 U22921 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19849), .ZN(n19850) );
  OAI22_X1 U22922 ( .A1(n19851), .A2(n19850), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19852) );
  OAI22_X1 U22923 ( .A1(n19855), .A2(n19854), .B1(n19853), .B2(n19852), .ZN(
        P3_U3031) );
  INV_X1 U22924 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19858) );
  NAND2_X1 U22925 ( .A1(n19856), .A2(n21589), .ZN(n19904) );
  CLKBUF_X1 U22926 ( .A(n19904), .Z(n21584) );
  OAI222_X1 U22927 ( .A1(n19924), .A2(n21587), .B1(n19857), .B2(n21589), .C1(
        n19858), .C2(n21584), .ZN(P3_U3032) );
  OAI222_X1 U22928 ( .A1(n21584), .A2(n19860), .B1(n19859), .B2(n21589), .C1(
        n19858), .C2(n21587), .ZN(P3_U3033) );
  OAI222_X1 U22929 ( .A1(n19904), .A2(n19862), .B1(n19861), .B2(n21589), .C1(
        n19860), .C2(n21587), .ZN(P3_U3034) );
  INV_X1 U22930 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19864) );
  OAI222_X1 U22931 ( .A1(n19904), .A2(n19864), .B1(n19863), .B2(n21589), .C1(
        n19862), .C2(n21587), .ZN(P3_U3035) );
  OAI222_X1 U22932 ( .A1(n19904), .A2(n19866), .B1(n19865), .B2(n21589), .C1(
        n19864), .C2(n21587), .ZN(P3_U3036) );
  OAI222_X1 U22933 ( .A1(n19904), .A2(n19868), .B1(n19867), .B2(n21589), .C1(
        n19866), .C2(n21587), .ZN(P3_U3037) );
  OAI222_X1 U22934 ( .A1(n19904), .A2(n19870), .B1(n19869), .B2(n21589), .C1(
        n19868), .C2(n21587), .ZN(P3_U3038) );
  OAI222_X1 U22935 ( .A1(n19904), .A2(n21816), .B1(n19871), .B2(n21589), .C1(
        n19870), .C2(n21587), .ZN(P3_U3039) );
  INV_X1 U22936 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U22937 ( .A1(n21584), .A2(n19873), .B1(n19872), .B2(n21589), .C1(
        n21816), .C2(n21587), .ZN(P3_U3040) );
  OAI222_X1 U22938 ( .A1(n21584), .A2(n19875), .B1(n19874), .B2(n21589), .C1(
        n19873), .C2(n21587), .ZN(P3_U3041) );
  INV_X1 U22939 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19878) );
  OAI222_X1 U22940 ( .A1(n21584), .A2(n19878), .B1(n19876), .B2(n21589), .C1(
        n19875), .C2(n21587), .ZN(P3_U3042) );
  OAI222_X1 U22941 ( .A1(n19878), .A2(n21587), .B1(n19877), .B2(n21589), .C1(
        n21778), .C2(n21584), .ZN(P3_U3043) );
  OAI222_X1 U22942 ( .A1(n21778), .A2(n21587), .B1(n19879), .B2(n21589), .C1(
        n19881), .C2(n21584), .ZN(P3_U3044) );
  OAI222_X1 U22943 ( .A1(n19881), .A2(n21587), .B1(n19880), .B2(n21589), .C1(
        n21819), .C2(n21584), .ZN(P3_U3045) );
  OAI222_X1 U22944 ( .A1(n21819), .A2(n21587), .B1(n19882), .B2(n21589), .C1(
        n19883), .C2(n21584), .ZN(P3_U3046) );
  OAI222_X1 U22945 ( .A1(n21584), .A2(n21717), .B1(n19884), .B2(n21589), .C1(
        n19883), .C2(n21587), .ZN(P3_U3047) );
  OAI222_X1 U22946 ( .A1(n21717), .A2(n21587), .B1(n21670), .B2(n21589), .C1(
        n19885), .C2(n21584), .ZN(P3_U3048) );
  OAI222_X1 U22947 ( .A1(n21584), .A2(n19887), .B1(n19886), .B2(n21589), .C1(
        n19885), .C2(n19909), .ZN(P3_U3049) );
  OAI222_X1 U22948 ( .A1(n21584), .A2(n19889), .B1(n19888), .B2(n21589), .C1(
        n19887), .C2(n19909), .ZN(P3_U3050) );
  OAI222_X1 U22949 ( .A1(n19889), .A2(n21587), .B1(n21850), .B2(n21589), .C1(
        n19890), .C2(n21584), .ZN(P3_U3051) );
  OAI222_X1 U22950 ( .A1(n21584), .A2(n19892), .B1(n19891), .B2(n21589), .C1(
        n19890), .C2(n19909), .ZN(P3_U3052) );
  INV_X1 U22951 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19895) );
  OAI222_X1 U22952 ( .A1(n19904), .A2(n19895), .B1(n19893), .B2(n21589), .C1(
        n19892), .C2(n19909), .ZN(P3_U3053) );
  OAI222_X1 U22953 ( .A1(n19895), .A2(n21587), .B1(n19894), .B2(n21589), .C1(
        n19896), .C2(n21584), .ZN(P3_U3054) );
  OAI222_X1 U22954 ( .A1(n21584), .A2(n19898), .B1(n19897), .B2(n21589), .C1(
        n19896), .C2(n19909), .ZN(P3_U3055) );
  INV_X1 U22955 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19900) );
  OAI222_X1 U22956 ( .A1(n19904), .A2(n19900), .B1(n19899), .B2(n21589), .C1(
        n19898), .C2(n21587), .ZN(P3_U3056) );
  OAI222_X1 U22957 ( .A1(n21584), .A2(n19902), .B1(n19901), .B2(n21589), .C1(
        n19900), .C2(n19909), .ZN(P3_U3057) );
  INV_X1 U22958 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n21586) );
  OAI222_X1 U22959 ( .A1(n19904), .A2(n21586), .B1(n19903), .B2(n21589), .C1(
        n19902), .C2(n21587), .ZN(P3_U3058) );
  OAI222_X1 U22960 ( .A1(n21584), .A2(n19908), .B1(n19905), .B2(n21589), .C1(
        n21585), .C2(n19909), .ZN(P3_U3060) );
  OAI222_X1 U22961 ( .A1(n19909), .A2(n19908), .B1(n19907), .B2(n21589), .C1(
        n19906), .C2(n21584), .ZN(P3_U3061) );
  INV_X1 U22962 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19910) );
  AOI22_X1 U22963 ( .A1(n21589), .A2(n19911), .B1(n19910), .B2(n19933), .ZN(
        P3_U3274) );
  INV_X1 U22964 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19926) );
  INV_X1 U22965 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19912) );
  AOI22_X1 U22966 ( .A1(n21589), .A2(n19926), .B1(n19912), .B2(n19933), .ZN(
        P3_U3275) );
  INV_X1 U22967 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19913) );
  AOI22_X1 U22968 ( .A1(n21589), .A2(n19914), .B1(n19913), .B2(n19933), .ZN(
        P3_U3276) );
  INV_X1 U22969 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19932) );
  INV_X1 U22970 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19915) );
  AOI22_X1 U22971 ( .A1(n21589), .A2(n19932), .B1(n19915), .B2(n19933), .ZN(
        P3_U3277) );
  INV_X1 U22972 ( .A(n19918), .ZN(n19916) );
  AOI21_X1 U22973 ( .B1(n19917), .B2(n21646), .A(n19916), .ZN(P3_U3280) );
  OAI21_X1 U22974 ( .B1(n19920), .B2(n19919), .A(n19918), .ZN(P3_U3281) );
  OAI221_X1 U22975 ( .B1(n19923), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19923), 
        .C2(n19922), .A(n19921), .ZN(P3_U3282) );
  AOI21_X1 U22976 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19925) );
  AOI22_X1 U22977 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19925), .B2(n19924), .ZN(n19927) );
  AOI22_X1 U22978 ( .A1(n19928), .A2(n19927), .B1(n19926), .B2(n19931), .ZN(
        P3_U3292) );
  NOR2_X1 U22979 ( .A1(n19931), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19929) );
  AOI22_X1 U22980 ( .A1(n19932), .A2(n19931), .B1(n19930), .B2(n19929), .ZN(
        P3_U3293) );
  INV_X1 U22981 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19934) );
  AOI22_X1 U22982 ( .A1(n21589), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19934), 
        .B2(n19933), .ZN(P3_U3294) );
  MUX2_X1 U22983 ( .A(P3_MORE_REG_SCAN_IN), .B(n19936), .S(n19935), .Z(
        P3_U3295) );
  OAI21_X1 U22984 ( .B1(n19938), .B2(n19937), .A(n19954), .ZN(n19939) );
  AOI21_X1 U22985 ( .B1(n19940), .B2(n19944), .A(n19939), .ZN(n19950) );
  AOI21_X1 U22986 ( .B1(n19943), .B2(n19942), .A(n19941), .ZN(n19945) );
  OAI211_X1 U22987 ( .C1(n19951), .C2(n19945), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19944), .ZN(n19947) );
  AOI21_X1 U22988 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19947), .A(n19946), 
        .ZN(n19949) );
  NAND2_X1 U22989 ( .A1(n19950), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19948) );
  OAI21_X1 U22990 ( .B1(n19950), .B2(n19949), .A(n19948), .ZN(P3_U3296) );
  MUX2_X1 U22991 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21589), .Z(P3_U3297) );
  INV_X1 U22992 ( .A(n19951), .ZN(n19953) );
  OAI21_X1 U22993 ( .B1(n19955), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19954), 
        .ZN(n19952) );
  OAI21_X1 U22994 ( .B1(n19954), .B2(n19953), .A(n19952), .ZN(P3_U3298) );
  NOR2_X1 U22995 ( .A1(n19955), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19957)
         );
  OAI21_X1 U22996 ( .B1(n19958), .B2(n19957), .A(n19956), .ZN(P3_U3299) );
  INV_X1 U22997 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19959) );
  NAND2_X1 U22998 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n21751), .ZN(n20681) );
  AOI22_X1 U22999 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20681), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20675), .ZN(n20745) );
  OAI21_X1 U23000 ( .B1(n20675), .B2(n19959), .A(n20674), .ZN(P2_U2815) );
  INV_X2 U23001 ( .A(n20818), .ZN(n20788) );
  NAND2_X1 U23002 ( .A1(n19961), .A2(n20818), .ZN(n20678) );
  AOI21_X1 U23003 ( .B1(n20675), .B2(n20678), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19960) );
  AOI21_X1 U23004 ( .B1(n20788), .B2(P2_CODEFETCH_REG_SCAN_IN), .A(n19960), 
        .ZN(P2_U2817) );
  INV_X1 U23005 ( .A(n19961), .ZN(n20683) );
  OAI21_X1 U23006 ( .B1(n20683), .B2(BS16), .A(n20745), .ZN(n20743) );
  OAI21_X1 U23007 ( .B1(n20745), .B2(n20395), .A(n20743), .ZN(P2_U2818) );
  NOR4_X1 U23008 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19971) );
  NOR4_X1 U23009 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19970) );
  NOR4_X1 U23010 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19962) );
  INV_X1 U23011 ( .A(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21801) );
  INV_X1 U23012 ( .A(P2_DATAWIDTH_REG_17__SCAN_IN), .ZN(n21668) );
  NAND3_X1 U23013 ( .A1(n19962), .A2(n21801), .A3(n21668), .ZN(n19968) );
  NOR4_X1 U23014 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19966) );
  NOR4_X1 U23015 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19965) );
  NOR4_X1 U23016 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19964) );
  NOR4_X1 U23017 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19963) );
  NAND4_X1 U23018 ( .A1(n19966), .A2(n19965), .A3(n19964), .A4(n19963), .ZN(
        n19967) );
  AOI211_X1 U23019 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19968), .B(n19967), .ZN(n19969) );
  NAND3_X1 U23020 ( .A1(n19971), .A2(n19970), .A3(n19969), .ZN(n19978) );
  NOR2_X1 U23021 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19978), .ZN(n19972) );
  INV_X1 U23022 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U23023 ( .A1(n19972), .A2(n19973), .B1(n19978), .B2(n20741), .ZN(
        P2_U2820) );
  OR3_X1 U23024 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19977) );
  INV_X1 U23025 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20739) );
  AOI22_X1 U23026 ( .A1(n19972), .A2(n19977), .B1(n19978), .B2(n20739), .ZN(
        P2_U2821) );
  INV_X1 U23027 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20744) );
  NAND2_X1 U23028 ( .A1(n19972), .A2(n20744), .ZN(n19976) );
  INV_X1 U23029 ( .A(n19978), .ZN(n19979) );
  OAI21_X1 U23030 ( .B1(n20692), .B2(n19973), .A(n19979), .ZN(n19974) );
  OAI21_X1 U23031 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19979), .A(n19974), 
        .ZN(n19975) );
  OAI221_X1 U23032 ( .B1(n19976), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19976), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19975), .ZN(P2_U2822) );
  INV_X1 U23033 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21707) );
  OAI221_X1 U23034 ( .B1(n19979), .B2(n21707), .C1(n19978), .C2(n19977), .A(
        n19976), .ZN(P2_U2823) );
  AOI22_X1 U23035 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19981), .B1(
        P2_EBX_REG_4__SCAN_IN), .B2(n19980), .ZN(n19999) );
  OAI22_X1 U23036 ( .A1(n20003), .A2(n19983), .B1(n19982), .B2(n12363), .ZN(
        n19984) );
  AOI211_X1 U23037 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19985), .A(n16754), .B(
        n19984), .ZN(n19998) );
  OAI22_X1 U23038 ( .A1(n20005), .A2(n19988), .B1(n19987), .B2(n19986), .ZN(
        n19989) );
  INV_X1 U23039 ( .A(n19989), .ZN(n19997) );
  NAND2_X1 U23040 ( .A1(n19990), .A2(n19991), .ZN(n19992) );
  MUX2_X1 U23041 ( .A(n19992), .B(n19991), .S(n10319), .Z(n19995) );
  NAND3_X1 U23042 ( .A1(n19995), .A2(n19994), .A3(n19993), .ZN(n19996) );
  NAND4_X1 U23043 ( .A1(n19999), .A2(n19998), .A3(n19997), .A4(n19996), .ZN(
        P2_U2851) );
  INV_X1 U23044 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20000) );
  OAI22_X1 U23045 ( .A1(n20003), .A2(n20002), .B1(n20001), .B2(n20000), .ZN(
        n20004) );
  INV_X1 U23046 ( .A(n20004), .ZN(n20009) );
  XNOR2_X1 U23047 ( .A(n20006), .B(n20005), .ZN(n20007) );
  NAND2_X1 U23048 ( .A1(n20007), .A2(n20020), .ZN(n20008) );
  OAI211_X1 U23049 ( .C1(n20124), .C2(n20024), .A(n20009), .B(n20008), .ZN(
        P2_U2915) );
  AOI22_X1 U23050 ( .A1(n20756), .A2(n20016), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n16191), .ZN(n20015) );
  OAI21_X1 U23051 ( .B1(n20012), .B2(n20011), .A(n20010), .ZN(n20013) );
  NAND2_X1 U23052 ( .A1(n20013), .A2(n20020), .ZN(n20014) );
  OAI211_X1 U23053 ( .C1(n20120), .C2(n20024), .A(n20015), .B(n20014), .ZN(
        P2_U2916) );
  AOI22_X1 U23054 ( .A1(n20016), .A2(n20772), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n16191), .ZN(n20023) );
  OAI21_X1 U23055 ( .B1(n20019), .B2(n20018), .A(n20017), .ZN(n20021) );
  NAND2_X1 U23056 ( .A1(n20021), .A2(n20020), .ZN(n20022) );
  OAI211_X1 U23057 ( .C1(n20025), .C2(n20024), .A(n20023), .B(n20022), .ZN(
        P2_U2918) );
  NAND2_X1 U23058 ( .A1(n20027), .A2(n20026), .ZN(n20029) );
  OAI21_X1 U23059 ( .B1(n20030), .B2(n20029), .A(n20028), .ZN(n20032) );
  INV_X1 U23060 ( .A(n20806), .ZN(n20031) );
  NOR2_X1 U23061 ( .A1(n20084), .A2(n21787), .ZN(P2_U2920) );
  INV_X1 U23062 ( .A(n20033), .ZN(n20034) );
  INV_X2 U23063 ( .A(n20084), .ZN(n20093) );
  AOI22_X1 U23064 ( .A1(n20799), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U23065 ( .B1(n20036), .B2(n20061), .A(n20035), .ZN(P2_U2921) );
  INV_X1 U23066 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n20038) );
  AOI22_X1 U23067 ( .A1(n20799), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U23068 ( .B1(n20038), .B2(n20061), .A(n20037), .ZN(P2_U2922) );
  AOI22_X1 U23069 ( .A1(n20799), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n20039) );
  OAI21_X1 U23070 ( .B1(n20040), .B2(n20061), .A(n20039), .ZN(P2_U2923) );
  INV_X1 U23071 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n21874) );
  AOI22_X1 U23072 ( .A1(n20799), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n20041) );
  OAI21_X1 U23073 ( .B1(n21874), .B2(n20061), .A(n20041), .ZN(P2_U2924) );
  AOI22_X1 U23074 ( .A1(n20799), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n20042) );
  OAI21_X1 U23075 ( .B1(n20043), .B2(n20061), .A(n20042), .ZN(P2_U2925) );
  INV_X1 U23076 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n21881) );
  AOI22_X1 U23077 ( .A1(n20799), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n20044) );
  OAI21_X1 U23078 ( .B1(n21881), .B2(n20061), .A(n20044), .ZN(P2_U2926) );
  INV_X1 U23079 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n20046) );
  AOI22_X1 U23080 ( .A1(n20799), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n20045) );
  OAI21_X1 U23081 ( .B1(n20046), .B2(n20061), .A(n20045), .ZN(P2_U2927) );
  INV_X1 U23082 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n20048) );
  AOI22_X1 U23083 ( .A1(n20799), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U23084 ( .B1(n20048), .B2(n20061), .A(n20047), .ZN(P2_U2928) );
  INV_X1 U23085 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U23086 ( .A1(n20799), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n20049) );
  OAI21_X1 U23087 ( .B1(n20050), .B2(n20061), .A(n20049), .ZN(P2_U2929) );
  INV_X1 U23088 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n21821) );
  AOI22_X1 U23089 ( .A1(n20799), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n20051) );
  OAI21_X1 U23090 ( .B1(n21821), .B2(n20061), .A(n20051), .ZN(P2_U2930) );
  INV_X1 U23091 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20053) );
  AOI22_X1 U23092 ( .A1(n20799), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n20052) );
  OAI21_X1 U23093 ( .B1(n20053), .B2(n20061), .A(n20052), .ZN(P2_U2931) );
  AOI22_X1 U23094 ( .A1(n20799), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U23095 ( .B1(n20055), .B2(n20061), .A(n20054), .ZN(P2_U2932) );
  INV_X1 U23096 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n20057) );
  AOI22_X1 U23097 ( .A1(n20799), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n20056) );
  OAI21_X1 U23098 ( .B1(n20057), .B2(n20061), .A(n20056), .ZN(P2_U2933) );
  INV_X1 U23099 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n20059) );
  AOI22_X1 U23100 ( .A1(n20799), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n20058) );
  OAI21_X1 U23101 ( .B1(n20059), .B2(n20061), .A(n20058), .ZN(P2_U2934) );
  AOI22_X1 U23102 ( .A1(n20799), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U23103 ( .B1(n20062), .B2(n20061), .A(n20060), .ZN(P2_U2935) );
  INV_X1 U23104 ( .A(n20082), .ZN(n20095) );
  AOI22_X1 U23105 ( .A1(n20799), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n20063) );
  OAI21_X1 U23106 ( .B1(n20064), .B2(n20095), .A(n20063), .ZN(P2_U2936) );
  AOI22_X1 U23107 ( .A1(n20799), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n20065) );
  OAI21_X1 U23108 ( .B1(n20066), .B2(n20095), .A(n20065), .ZN(P2_U2937) );
  AOI22_X1 U23109 ( .A1(n20086), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n20067) );
  OAI21_X1 U23110 ( .B1(n21804), .B2(n20095), .A(n20067), .ZN(P2_U2938) );
  AOI22_X1 U23111 ( .A1(n20086), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n20068) );
  OAI21_X1 U23112 ( .B1(n20069), .B2(n20095), .A(n20068), .ZN(P2_U2939) );
  AOI22_X1 U23113 ( .A1(n20086), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n20070) );
  OAI21_X1 U23114 ( .B1(n20071), .B2(n20095), .A(n20070), .ZN(P2_U2940) );
  AOI22_X1 U23115 ( .A1(n20086), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n20072) );
  OAI21_X1 U23116 ( .B1(n20073), .B2(n20095), .A(n20072), .ZN(P2_U2941) );
  AOI22_X1 U23117 ( .A1(n20086), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n20074) );
  OAI21_X1 U23118 ( .B1(n20075), .B2(n20095), .A(n20074), .ZN(P2_U2942) );
  AOI22_X1 U23119 ( .A1(n20086), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n20076) );
  OAI21_X1 U23120 ( .B1(n20077), .B2(n20095), .A(n20076), .ZN(P2_U2943) );
  AOI22_X1 U23121 ( .A1(n20086), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n20078) );
  OAI21_X1 U23122 ( .B1(n20079), .B2(n20095), .A(n20078), .ZN(P2_U2944) );
  AOI22_X1 U23123 ( .A1(n20086), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n20080) );
  OAI21_X1 U23124 ( .B1(n20081), .B2(n20095), .A(n20080), .ZN(P2_U2945) );
  AOI22_X1 U23125 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n20082), .B1(n20799), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n20083) );
  OAI21_X1 U23126 ( .B1(n20084), .B2(n21807), .A(n20083), .ZN(P2_U2946) );
  AOI22_X1 U23127 ( .A1(n20086), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n20085) );
  OAI21_X1 U23128 ( .B1(n20000), .B2(n20095), .A(n20085), .ZN(P2_U2947) );
  INV_X1 U23129 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n20088) );
  AOI22_X1 U23130 ( .A1(n20086), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n20087) );
  OAI21_X1 U23131 ( .B1(n20088), .B2(n20095), .A(n20087), .ZN(P2_U2948) );
  AOI22_X1 U23132 ( .A1(n20799), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n20089) );
  OAI21_X1 U23133 ( .B1(n20090), .B2(n20095), .A(n20089), .ZN(P2_U2949) );
  INV_X1 U23134 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n20092) );
  AOI22_X1 U23135 ( .A1(n20799), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n20091) );
  OAI21_X1 U23136 ( .B1(n20092), .B2(n20095), .A(n20091), .ZN(P2_U2950) );
  INV_X1 U23137 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n20096) );
  AOI22_X1 U23138 ( .A1(n20799), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n20093), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n20094) );
  OAI21_X1 U23139 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(P2_U2951) );
  NAND2_X1 U23140 ( .A1(n20758), .A2(n20766), .ZN(n20207) );
  NOR2_X1 U23141 ( .A1(n20247), .A2(n20207), .ZN(n20109) );
  AOI22_X1 U23142 ( .A1(n20621), .A2(n20668), .B1(n20613), .B2(n20109), .ZN(
        n20108) );
  AOI21_X1 U23143 ( .B1(n20625), .B2(n20173), .A(n20395), .ZN(n20097) );
  NOR2_X1 U23144 ( .A1(n20097), .A2(n20804), .ZN(n20102) );
  INV_X1 U23145 ( .A(n20098), .ZN(n20099) );
  NOR2_X1 U23146 ( .A1(n20663), .A2(n20109), .ZN(n20105) );
  NAND2_X1 U23147 ( .A1(n20102), .A2(n20105), .ZN(n20100) );
  INV_X1 U23148 ( .A(n20102), .ZN(n20106) );
  OAI21_X1 U23149 ( .B1(n20103), .B2(n20109), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20104) );
  AOI22_X1 U23150 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20144), .B1(
        n20614), .B2(n20143), .ZN(n20107) );
  OAI211_X1 U23151 ( .C1(n20626), .C2(n20173), .A(n20108), .B(n20107), .ZN(
        P2_U3048) );
  INV_X1 U23152 ( .A(n20109), .ZN(n20141) );
  OAI22_X1 U23153 ( .A1(n20632), .A2(n20625), .B1(n20572), .B2(n20141), .ZN(
        n20110) );
  INV_X1 U23154 ( .A(n20110), .ZN(n20112) );
  AOI22_X1 U23155 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20144), .B1(
        n20628), .B2(n20143), .ZN(n20111) );
  OAI211_X1 U23156 ( .C1(n20576), .C2(n20173), .A(n20112), .B(n20111), .ZN(
        P2_U3049) );
  AOI22_X1 U23157 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n20133), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n20134), .ZN(n20638) );
  NAND2_X1 U23158 ( .A1(n20136), .A2(n20113), .ZN(n20577) );
  OAI22_X1 U23159 ( .A1(n20638), .A2(n20625), .B1(n20577), .B2(n20141), .ZN(
        n20114) );
  INV_X1 U23160 ( .A(n20114), .ZN(n20117) );
  NOR2_X2 U23161 ( .A1(n20494), .A2(n20115), .ZN(n20634) );
  AOI22_X1 U23162 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20144), .B1(
        n20634), .B2(n20143), .ZN(n20116) );
  OAI211_X1 U23163 ( .C1(n20578), .C2(n20173), .A(n20117), .B(n20116), .ZN(
        P2_U3050) );
  AOI22_X2 U23164 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20133), .ZN(n20586) );
  AOI22_X1 U23165 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20133), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n20134), .ZN(n20644) );
  NAND2_X1 U23166 ( .A1(n20136), .A2(n20118), .ZN(n20582) );
  OAI22_X1 U23167 ( .A1(n20644), .A2(n20625), .B1(n20582), .B2(n20141), .ZN(
        n20119) );
  INV_X1 U23168 ( .A(n20119), .ZN(n20122) );
  NOR2_X2 U23169 ( .A1(n20494), .A2(n20120), .ZN(n20640) );
  AOI22_X1 U23170 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20144), .B1(
        n20640), .B2(n20143), .ZN(n20121) );
  OAI211_X1 U23171 ( .C1(n20586), .C2(n20173), .A(n20122), .B(n20121), .ZN(
        P2_U3051) );
  AOI22_X1 U23172 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n20133), .ZN(n20588) );
  AOI22_X1 U23173 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n20133), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n20134), .ZN(n20650) );
  OAI22_X1 U23174 ( .A1(n20650), .A2(n20625), .B1(n20587), .B2(n20141), .ZN(
        n20123) );
  INV_X1 U23175 ( .A(n20123), .ZN(n20126) );
  NOR2_X2 U23176 ( .A1(n20494), .A2(n20124), .ZN(n20646) );
  AOI22_X1 U23177 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20144), .B1(
        n20646), .B2(n20143), .ZN(n20125) );
  OAI211_X1 U23178 ( .C1(n20588), .C2(n20173), .A(n20126), .B(n20125), .ZN(
        P2_U3052) );
  AOI22_X2 U23179 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n20133), .ZN(n20596) );
  AOI22_X1 U23180 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n20133), .ZN(n20656) );
  NAND2_X1 U23181 ( .A1(n20136), .A2(n20127), .ZN(n20592) );
  OAI22_X1 U23182 ( .A1(n20656), .A2(n20625), .B1(n20592), .B2(n20141), .ZN(
        n20128) );
  INV_X1 U23183 ( .A(n20128), .ZN(n20132) );
  INV_X1 U23184 ( .A(n20129), .ZN(n20130) );
  NOR2_X2 U23185 ( .A1(n20494), .A2(n20130), .ZN(n20652) );
  AOI22_X1 U23186 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20144), .B1(
        n20652), .B2(n20143), .ZN(n20131) );
  OAI211_X1 U23187 ( .C1(n20596), .C2(n20173), .A(n20132), .B(n20131), .ZN(
        P2_U3053) );
  AOI22_X1 U23188 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n20133), .ZN(n20601) );
  AOI22_X1 U23189 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20134), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20133), .ZN(n20662) );
  NAND2_X1 U23190 ( .A1(n20136), .A2(n20135), .ZN(n20597) );
  OAI22_X1 U23191 ( .A1(n9921), .A2(n20625), .B1(n20597), .B2(n20141), .ZN(
        n20137) );
  INV_X1 U23192 ( .A(n20137), .ZN(n20140) );
  NOR2_X2 U23193 ( .A1(n20494), .A2(n20138), .ZN(n20658) );
  AOI22_X1 U23194 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20144), .B1(
        n20658), .B2(n20143), .ZN(n20139) );
  OAI211_X1 U23195 ( .C1(n20601), .C2(n20173), .A(n20140), .B(n20139), .ZN(
        P2_U3054) );
  OAI22_X1 U23196 ( .A1(n20673), .A2(n20625), .B1(n20141), .B2(n20602), .ZN(
        n20142) );
  INV_X1 U23197 ( .A(n20142), .ZN(n20146) );
  AOI22_X1 U23198 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20144), .B1(
        n20665), .B2(n20143), .ZN(n20145) );
  OAI211_X1 U23199 ( .C1(n20610), .C2(n20173), .A(n20146), .B(n20145), .ZN(
        P2_U3055) );
  NOR3_X2 U23200 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20786), .A3(
        n20207), .ZN(n20168) );
  OR2_X1 U23201 ( .A1(n20168), .A2(n20489), .ZN(n20147) );
  OR2_X1 U23202 ( .A1(n20207), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20150) );
  OAI21_X1 U23203 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20150), .A(n20489), 
        .ZN(n20149) );
  AOI22_X1 U23204 ( .A1(n20169), .A2(n20614), .B1(n20613), .B2(n20168), .ZN(
        n20155) );
  NAND2_X1 U23205 ( .A1(n20751), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20753) );
  OAI21_X1 U23206 ( .B1(n20753), .B2(n20396), .A(n20150), .ZN(n20153) );
  OR2_X1 U23207 ( .A1(n20168), .A2(n20800), .ZN(n20151) );
  NAND4_X1 U23208 ( .A1(n20153), .A2(n20619), .A3(n20152), .A4(n20151), .ZN(
        n20170) );
  AOI22_X1 U23209 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20558), .ZN(n20154) );
  OAI211_X1 U23210 ( .C1(n20571), .C2(n20173), .A(n20155), .B(n20154), .ZN(
        P2_U3056) );
  AOI22_X1 U23211 ( .A1(n20169), .A2(n20628), .B1(n20627), .B2(n20168), .ZN(
        n20157) );
  AOI22_X1 U23212 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20629), .ZN(n20156) );
  OAI211_X1 U23213 ( .C1(n20632), .C2(n20173), .A(n20157), .B(n20156), .ZN(
        P2_U3057) );
  AOI22_X1 U23214 ( .A1(n20169), .A2(n20634), .B1(n20633), .B2(n20168), .ZN(
        n20159) );
  INV_X1 U23215 ( .A(n20578), .ZN(n20635) );
  AOI22_X1 U23216 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20635), .ZN(n20158) );
  OAI211_X1 U23217 ( .C1(n20638), .C2(n20173), .A(n20159), .B(n20158), .ZN(
        P2_U3058) );
  AOI22_X1 U23218 ( .A1(n20169), .A2(n20640), .B1(n20639), .B2(n20168), .ZN(
        n20161) );
  INV_X1 U23219 ( .A(n20586), .ZN(n20641) );
  AOI22_X1 U23220 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20641), .ZN(n20160) );
  OAI211_X1 U23221 ( .C1(n20644), .C2(n20173), .A(n20161), .B(n20160), .ZN(
        P2_U3059) );
  AOI22_X1 U23222 ( .A1(n20169), .A2(n20646), .B1(n20645), .B2(n20168), .ZN(
        n20163) );
  INV_X1 U23223 ( .A(n20588), .ZN(n20647) );
  AOI22_X1 U23224 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20647), .ZN(n20162) );
  OAI211_X1 U23225 ( .C1(n20650), .C2(n20173), .A(n20163), .B(n20162), .ZN(
        P2_U3060) );
  AOI22_X1 U23226 ( .A1(n20169), .A2(n20652), .B1(n20651), .B2(n20168), .ZN(
        n20165) );
  INV_X1 U23227 ( .A(n20596), .ZN(n20653) );
  AOI22_X1 U23228 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20653), .ZN(n20164) );
  OAI211_X1 U23229 ( .C1(n20656), .C2(n20173), .A(n20165), .B(n20164), .ZN(
        P2_U3061) );
  AOI22_X1 U23230 ( .A1(n20169), .A2(n20658), .B1(n20657), .B2(n20168), .ZN(
        n20167) );
  INV_X1 U23231 ( .A(n20601), .ZN(n20659) );
  AOI22_X1 U23232 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20659), .ZN(n20166) );
  OAI211_X1 U23233 ( .C1(n9921), .C2(n20173), .A(n20167), .B(n20166), .ZN(
        P2_U3062) );
  AOI22_X1 U23234 ( .A1(n20169), .A2(n20665), .B1(n20664), .B2(n20168), .ZN(
        n20172) );
  INV_X1 U23235 ( .A(n20610), .ZN(n20667) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20170), .B1(
        n20201), .B2(n20667), .ZN(n20171) );
  OAI211_X1 U23237 ( .C1(n20673), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        P2_U3063) );
  NOR3_X2 U23238 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20776), .A3(
        n20207), .ZN(n20199) );
  OAI21_X1 U23239 ( .B1(n20174), .B2(n20199), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20176) );
  INV_X1 U23240 ( .A(n20207), .ZN(n20206) );
  NAND2_X1 U23241 ( .A1(n20175), .A2(n20206), .ZN(n20180) );
  NAND2_X1 U23242 ( .A1(n20176), .A2(n20180), .ZN(n20200) );
  AOI22_X1 U23243 ( .A1(n20200), .A2(n20614), .B1(n20613), .B2(n20199), .ZN(
        n20186) );
  INV_X1 U23244 ( .A(n20199), .ZN(n20177) );
  OAI21_X1 U23245 ( .B1(n20178), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20177), 
        .ZN(n20183) );
  OAI21_X1 U23246 ( .B1(n20179), .B2(n20201), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20181) );
  NAND2_X1 U23247 ( .A1(n20181), .A2(n20180), .ZN(n20182) );
  MUX2_X1 U23248 ( .A(n20183), .B(n20182), .S(n20749), .Z(n20184) );
  NAND2_X1 U23249 ( .A1(n20184), .A2(n20619), .ZN(n20202) );
  AOI22_X1 U23250 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20621), .ZN(n20185) );
  OAI211_X1 U23251 ( .C1(n20626), .C2(n20243), .A(n20186), .B(n20185), .ZN(
        P2_U3064) );
  AOI22_X1 U23252 ( .A1(n20200), .A2(n20628), .B1(n20627), .B2(n20199), .ZN(
        n20188) );
  AOI22_X1 U23253 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20499), .ZN(n20187) );
  OAI211_X1 U23254 ( .C1(n20576), .C2(n20243), .A(n20188), .B(n20187), .ZN(
        P2_U3065) );
  AOI22_X1 U23255 ( .A1(n20200), .A2(n20634), .B1(n20633), .B2(n20199), .ZN(
        n20190) );
  INV_X1 U23256 ( .A(n20638), .ZN(n20502) );
  AOI22_X1 U23257 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20502), .ZN(n20189) );
  OAI211_X1 U23258 ( .C1(n20578), .C2(n20243), .A(n20190), .B(n20189), .ZN(
        P2_U3066) );
  AOI22_X1 U23259 ( .A1(n20200), .A2(n20640), .B1(n20639), .B2(n20199), .ZN(
        n20192) );
  INV_X1 U23260 ( .A(n20644), .ZN(n20505) );
  AOI22_X1 U23261 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20505), .ZN(n20191) );
  OAI211_X1 U23262 ( .C1(n20586), .C2(n20243), .A(n20192), .B(n20191), .ZN(
        P2_U3067) );
  AOI22_X1 U23263 ( .A1(n20200), .A2(n20646), .B1(n20645), .B2(n20199), .ZN(
        n20194) );
  INV_X1 U23264 ( .A(n20650), .ZN(n20508) );
  AOI22_X1 U23265 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20508), .ZN(n20193) );
  OAI211_X1 U23266 ( .C1(n20588), .C2(n20243), .A(n20194), .B(n20193), .ZN(
        P2_U3068) );
  AOI22_X1 U23267 ( .A1(n20200), .A2(n20652), .B1(n20651), .B2(n20199), .ZN(
        n20196) );
  INV_X1 U23268 ( .A(n20656), .ZN(n20511) );
  AOI22_X1 U23269 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20511), .ZN(n20195) );
  OAI211_X1 U23270 ( .C1(n20596), .C2(n20243), .A(n20196), .B(n20195), .ZN(
        P2_U3069) );
  AOI22_X1 U23271 ( .A1(n20200), .A2(n20658), .B1(n20657), .B2(n20199), .ZN(
        n20198) );
  INV_X1 U23272 ( .A(n20662), .ZN(n20514) );
  AOI22_X1 U23273 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20514), .ZN(n20197) );
  OAI211_X1 U23274 ( .C1(n20601), .C2(n20243), .A(n20198), .B(n20197), .ZN(
        P2_U3070) );
  AOI22_X1 U23275 ( .A1(n20200), .A2(n20665), .B1(n20664), .B2(n20199), .ZN(
        n20204) );
  INV_X1 U23276 ( .A(n20673), .ZN(n20519) );
  AOI22_X1 U23277 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20202), .B1(
        n20201), .B2(n20519), .ZN(n20203) );
  OAI211_X1 U23278 ( .C1(n20610), .C2(n20243), .A(n20204), .B(n20203), .ZN(
        P2_U3071) );
  NAND2_X1 U23279 ( .A1(n20457), .A2(n20206), .ZN(n20236) );
  INV_X1 U23280 ( .A(n20236), .ZN(n20211) );
  AOI22_X1 U23281 ( .A1(n20558), .A2(n20270), .B1(n20613), .B2(n20211), .ZN(
        n20217) );
  OAI21_X1 U23282 ( .B1(n20453), .B2(n20753), .A(n20749), .ZN(n20215) );
  NOR2_X1 U23283 ( .A1(n20776), .A2(n20207), .ZN(n20210) );
  OAI21_X1 U23284 ( .B1(n20212), .B2(n20489), .A(n20800), .ZN(n20208) );
  AOI21_X1 U23285 ( .B1(n20208), .B2(n20236), .A(n20494), .ZN(n20209) );
  INV_X1 U23286 ( .A(n20210), .ZN(n20214) );
  OAI21_X1 U23287 ( .B1(n20212), .B2(n20211), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20213) );
  AOI22_X1 U23288 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20240), .B1(
        n20614), .B2(n20239), .ZN(n20216) );
  OAI211_X1 U23289 ( .C1(n20571), .C2(n20243), .A(n20217), .B(n20216), .ZN(
        P2_U3072) );
  OAI22_X1 U23290 ( .A1(n20576), .A2(n20237), .B1(n20236), .B2(n20572), .ZN(
        n20218) );
  INV_X1 U23291 ( .A(n20218), .ZN(n20220) );
  AOI22_X1 U23292 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20240), .B1(
        n20628), .B2(n20239), .ZN(n20219) );
  OAI211_X1 U23293 ( .C1(n20632), .C2(n20243), .A(n20220), .B(n20219), .ZN(
        P2_U3073) );
  OAI22_X1 U23294 ( .A1(n20578), .A2(n20237), .B1(n20236), .B2(n20577), .ZN(
        n20221) );
  INV_X1 U23295 ( .A(n20221), .ZN(n20223) );
  AOI22_X1 U23296 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20240), .B1(
        n20634), .B2(n20239), .ZN(n20222) );
  OAI211_X1 U23297 ( .C1(n20638), .C2(n20243), .A(n20223), .B(n20222), .ZN(
        P2_U3074) );
  OAI22_X1 U23298 ( .A1(n20586), .A2(n20237), .B1(n20236), .B2(n20582), .ZN(
        n20224) );
  INV_X1 U23299 ( .A(n20224), .ZN(n20226) );
  AOI22_X1 U23300 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20240), .B1(
        n20640), .B2(n20239), .ZN(n20225) );
  OAI211_X1 U23301 ( .C1(n20644), .C2(n20243), .A(n20226), .B(n20225), .ZN(
        P2_U3075) );
  OAI22_X1 U23302 ( .A1(n20650), .A2(n20243), .B1(n20236), .B2(n20587), .ZN(
        n20227) );
  INV_X1 U23303 ( .A(n20227), .ZN(n20229) );
  AOI22_X1 U23304 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20240), .B1(
        n20646), .B2(n20239), .ZN(n20228) );
  OAI211_X1 U23305 ( .C1(n20588), .C2(n20237), .A(n20229), .B(n20228), .ZN(
        P2_U3076) );
  OAI22_X1 U23306 ( .A1(n20656), .A2(n20243), .B1(n20236), .B2(n20592), .ZN(
        n20230) );
  INV_X1 U23307 ( .A(n20230), .ZN(n20232) );
  AOI22_X1 U23308 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20240), .B1(
        n20652), .B2(n20239), .ZN(n20231) );
  OAI211_X1 U23309 ( .C1(n20596), .C2(n20237), .A(n20232), .B(n20231), .ZN(
        P2_U3077) );
  OAI22_X1 U23310 ( .A1(n20601), .A2(n20237), .B1(n20236), .B2(n20597), .ZN(
        n20233) );
  INV_X1 U23311 ( .A(n20233), .ZN(n20235) );
  AOI22_X1 U23312 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20240), .B1(
        n20658), .B2(n20239), .ZN(n20234) );
  OAI211_X1 U23313 ( .C1(n9921), .C2(n20243), .A(n20235), .B(n20234), .ZN(
        P2_U3078) );
  OAI22_X1 U23314 ( .A1(n20610), .A2(n20237), .B1(n20236), .B2(n20602), .ZN(
        n20238) );
  INV_X1 U23315 ( .A(n20238), .ZN(n20242) );
  AOI22_X1 U23316 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20240), .B1(
        n20665), .B2(n20239), .ZN(n20241) );
  OAI211_X1 U23317 ( .C1(n20673), .C2(n20243), .A(n20242), .B(n20241), .ZN(
        P2_U3079) );
  NOR2_X1 U23318 ( .A1(n20246), .A2(n20245), .ZN(n20492) );
  NAND2_X1 U23319 ( .A1(n20492), .A2(n20758), .ZN(n20252) );
  NOR2_X1 U23320 ( .A1(n20274), .A2(n20247), .ZN(n20268) );
  OAI21_X1 U23321 ( .B1(n20249), .B2(n20268), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20248) );
  OAI21_X1 U23322 ( .B1(n20252), .B2(n20804), .A(n20248), .ZN(n20269) );
  AOI22_X1 U23323 ( .A1(n20269), .A2(n20614), .B1(n20613), .B2(n20268), .ZN(
        n20255) );
  OAI21_X1 U23324 ( .B1(n20270), .B2(n20275), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20251) );
  AOI211_X1 U23325 ( .C1(n20249), .C2(n20800), .A(n20749), .B(n20268), .ZN(
        n20250) );
  AOI211_X1 U23326 ( .C1(n20252), .C2(n20251), .A(n20494), .B(n20250), .ZN(
        n20253) );
  AOI22_X1 U23327 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20621), .ZN(n20254) );
  OAI211_X1 U23328 ( .C1(n20626), .C2(n20306), .A(n20255), .B(n20254), .ZN(
        P2_U3080) );
  AOI22_X1 U23329 ( .A1(n20269), .A2(n20628), .B1(n20627), .B2(n20268), .ZN(
        n20257) );
  AOI22_X1 U23330 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20499), .ZN(n20256) );
  OAI211_X1 U23331 ( .C1(n20576), .C2(n20306), .A(n20257), .B(n20256), .ZN(
        P2_U3081) );
  AOI22_X1 U23332 ( .A1(n20269), .A2(n20634), .B1(n20633), .B2(n20268), .ZN(
        n20259) );
  AOI22_X1 U23333 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20502), .ZN(n20258) );
  OAI211_X1 U23334 ( .C1(n20578), .C2(n20306), .A(n20259), .B(n20258), .ZN(
        P2_U3082) );
  AOI22_X1 U23335 ( .A1(n20269), .A2(n20640), .B1(n20639), .B2(n20268), .ZN(
        n20261) );
  AOI22_X1 U23336 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20505), .ZN(n20260) );
  OAI211_X1 U23337 ( .C1(n20586), .C2(n20306), .A(n20261), .B(n20260), .ZN(
        P2_U3083) );
  AOI22_X1 U23338 ( .A1(n20269), .A2(n20646), .B1(n20645), .B2(n20268), .ZN(
        n20263) );
  AOI22_X1 U23339 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20508), .ZN(n20262) );
  OAI211_X1 U23340 ( .C1(n20588), .C2(n20306), .A(n20263), .B(n20262), .ZN(
        P2_U3084) );
  AOI22_X1 U23341 ( .A1(n20269), .A2(n20652), .B1(n20651), .B2(n20268), .ZN(
        n20265) );
  AOI22_X1 U23342 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20511), .ZN(n20264) );
  OAI211_X1 U23343 ( .C1(n20596), .C2(n20306), .A(n20265), .B(n20264), .ZN(
        P2_U3085) );
  AOI22_X1 U23344 ( .A1(n20269), .A2(n20658), .B1(n20657), .B2(n20268), .ZN(
        n20267) );
  AOI22_X1 U23345 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20514), .ZN(n20266) );
  OAI211_X1 U23346 ( .C1(n20601), .C2(n20306), .A(n20267), .B(n20266), .ZN(
        P2_U3086) );
  AOI22_X1 U23347 ( .A1(n20269), .A2(n20665), .B1(n20664), .B2(n20268), .ZN(
        n20273) );
  AOI22_X1 U23348 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20271), .B1(
        n20270), .B2(n20519), .ZN(n20272) );
  OAI211_X1 U23349 ( .C1(n20610), .C2(n20306), .A(n20273), .B(n20272), .ZN(
        P2_U3087) );
  NOR3_X1 U23350 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20786), .A3(
        n20274), .ZN(n20280) );
  AOI22_X1 U23351 ( .A1(n20621), .A2(n20275), .B1(n20613), .B2(n20280), .ZN(
        n20285) );
  OAI21_X1 U23352 ( .B1(n20753), .B2(n20535), .A(n20749), .ZN(n20283) );
  NAND2_X1 U23353 ( .A1(n20776), .A2(n20276), .ZN(n20282) );
  INV_X1 U23354 ( .A(n20282), .ZN(n20279) );
  INV_X1 U23355 ( .A(n20280), .ZN(n20305) );
  AOI21_X1 U23356 ( .B1(n20277), .B2(n20305), .A(n20494), .ZN(n20278) );
  AOI22_X1 U23357 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20309), .B1(
        n20614), .B2(n20308), .ZN(n20284) );
  OAI211_X1 U23358 ( .C1(n20626), .C2(n20298), .A(n20285), .B(n20284), .ZN(
        P2_U3088) );
  OAI22_X1 U23359 ( .A1(n20632), .A2(n20306), .B1(n20305), .B2(n20572), .ZN(
        n20286) );
  INV_X1 U23360 ( .A(n20286), .ZN(n20288) );
  AOI22_X1 U23361 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20309), .B1(
        n20628), .B2(n20308), .ZN(n20287) );
  OAI211_X1 U23362 ( .C1(n20576), .C2(n20298), .A(n20288), .B(n20287), .ZN(
        P2_U3089) );
  OAI22_X1 U23363 ( .A1(n20578), .A2(n20298), .B1(n20305), .B2(n20577), .ZN(
        n20289) );
  INV_X1 U23364 ( .A(n20289), .ZN(n20291) );
  AOI22_X1 U23365 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20309), .B1(
        n20634), .B2(n20308), .ZN(n20290) );
  OAI211_X1 U23366 ( .C1(n20638), .C2(n20306), .A(n20291), .B(n20290), .ZN(
        P2_U3090) );
  OAI22_X1 U23367 ( .A1(n20644), .A2(n20306), .B1(n20305), .B2(n20582), .ZN(
        n20292) );
  INV_X1 U23368 ( .A(n20292), .ZN(n20294) );
  AOI22_X1 U23369 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20309), .B1(
        n20640), .B2(n20308), .ZN(n20293) );
  OAI211_X1 U23370 ( .C1(n20586), .C2(n20298), .A(n20294), .B(n20293), .ZN(
        P2_U3091) );
  OAI22_X1 U23371 ( .A1(n20650), .A2(n20306), .B1(n20587), .B2(n20305), .ZN(
        n20295) );
  INV_X1 U23372 ( .A(n20295), .ZN(n20297) );
  AOI22_X1 U23373 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20309), .B1(
        n20646), .B2(n20308), .ZN(n20296) );
  OAI211_X1 U23374 ( .C1(n20588), .C2(n20298), .A(n20297), .B(n20296), .ZN(
        P2_U3092) );
  OAI22_X1 U23375 ( .A1(n20596), .A2(n20298), .B1(n20592), .B2(n20305), .ZN(
        n20299) );
  INV_X1 U23376 ( .A(n20299), .ZN(n20301) );
  AOI22_X1 U23377 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20309), .B1(
        n20652), .B2(n20308), .ZN(n20300) );
  OAI211_X1 U23378 ( .C1(n20656), .C2(n20306), .A(n20301), .B(n20300), .ZN(
        P2_U3093) );
  OAI22_X1 U23379 ( .A1(n9921), .A2(n20306), .B1(n20305), .B2(n20597), .ZN(
        n20302) );
  INV_X1 U23380 ( .A(n20302), .ZN(n20304) );
  AOI22_X1 U23381 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20309), .B1(
        n20658), .B2(n20308), .ZN(n20303) );
  OAI211_X1 U23382 ( .C1(n20601), .C2(n20298), .A(n20304), .B(n20303), .ZN(
        P2_U3094) );
  OAI22_X1 U23383 ( .A1(n20673), .A2(n20306), .B1(n20305), .B2(n20602), .ZN(
        n20307) );
  INV_X1 U23384 ( .A(n20307), .ZN(n20311) );
  AOI22_X1 U23385 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20309), .B1(
        n20665), .B2(n20308), .ZN(n20310) );
  OAI211_X1 U23386 ( .C1(n20610), .C2(n20298), .A(n20311), .B(n20310), .ZN(
        P2_U3095) );
  INV_X1 U23387 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n20315) );
  AOI22_X1 U23388 ( .A1(n20328), .A2(n20628), .B1(n20327), .B2(n20627), .ZN(
        n20314) );
  AOI22_X1 U23389 ( .A1(n20312), .A2(n20499), .B1(n20362), .B2(n20629), .ZN(
        n20313) );
  OAI211_X1 U23390 ( .C1(n20316), .C2(n20315), .A(n20314), .B(n20313), .ZN(
        P2_U3097) );
  AOI22_X1 U23391 ( .A1(n20328), .A2(n20634), .B1(n20327), .B2(n20633), .ZN(
        n20318) );
  AOI22_X1 U23392 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20635), .ZN(n20317) );
  OAI211_X1 U23393 ( .C1(n20638), .C2(n20298), .A(n20318), .B(n20317), .ZN(
        P2_U3098) );
  AOI22_X1 U23394 ( .A1(n20328), .A2(n20640), .B1(n20327), .B2(n20639), .ZN(
        n20320) );
  AOI22_X1 U23395 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20641), .ZN(n20319) );
  OAI211_X1 U23396 ( .C1(n20644), .C2(n20298), .A(n20320), .B(n20319), .ZN(
        P2_U3099) );
  AOI22_X1 U23397 ( .A1(n20328), .A2(n20646), .B1(n20327), .B2(n20645), .ZN(
        n20322) );
  AOI22_X1 U23398 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20647), .ZN(n20321) );
  OAI211_X1 U23399 ( .C1(n20650), .C2(n20298), .A(n20322), .B(n20321), .ZN(
        P2_U3100) );
  AOI22_X1 U23400 ( .A1(n20328), .A2(n20652), .B1(n20327), .B2(n20651), .ZN(
        n20324) );
  AOI22_X1 U23401 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20653), .ZN(n20323) );
  OAI211_X1 U23402 ( .C1(n20656), .C2(n20298), .A(n20324), .B(n20323), .ZN(
        P2_U3101) );
  AOI22_X1 U23403 ( .A1(n20328), .A2(n20658), .B1(n20327), .B2(n20657), .ZN(
        n20326) );
  AOI22_X1 U23404 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20659), .ZN(n20325) );
  OAI211_X1 U23405 ( .C1(n9921), .C2(n20298), .A(n20326), .B(n20325), .ZN(
        P2_U3102) );
  AOI22_X1 U23406 ( .A1(n20328), .A2(n20665), .B1(n20327), .B2(n20664), .ZN(
        n20331) );
  AOI22_X1 U23407 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20329), .B1(
        n20362), .B2(n20667), .ZN(n20330) );
  OAI211_X1 U23408 ( .C1(n20673), .C2(n20298), .A(n20331), .B(n20330), .ZN(
        P2_U3103) );
  INV_X1 U23409 ( .A(n20753), .ZN(n20333) );
  INV_X1 U23410 ( .A(n20752), .ZN(n20332) );
  NAND2_X1 U23411 ( .A1(n20333), .A2(n20332), .ZN(n20335) );
  AOI211_X1 U23412 ( .C1(n20336), .C2(n20800), .A(n20749), .B(n20360), .ZN(
        n20334) );
  INV_X1 U23413 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n20341) );
  OAI21_X1 U23414 ( .B1(n20336), .B2(n20360), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20337) );
  OAI21_X1 U23415 ( .B1(n20338), .B2(n20804), .A(n20337), .ZN(n20361) );
  AOI22_X1 U23416 ( .A1(n20361), .A2(n20614), .B1(n20360), .B2(n20613), .ZN(
        n20340) );
  AOI22_X1 U23417 ( .A1(n20362), .A2(n20621), .B1(n20388), .B2(n20558), .ZN(
        n20339) );
  OAI211_X1 U23418 ( .C1(n20365), .C2(n20341), .A(n20340), .B(n20339), .ZN(
        P2_U3104) );
  INV_X1 U23419 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20344) );
  AOI22_X1 U23420 ( .A1(n20361), .A2(n20628), .B1(n20360), .B2(n20627), .ZN(
        n20343) );
  AOI22_X1 U23421 ( .A1(n20362), .A2(n20499), .B1(n20388), .B2(n20629), .ZN(
        n20342) );
  OAI211_X1 U23422 ( .C1(n20365), .C2(n20344), .A(n20343), .B(n20342), .ZN(
        P2_U3105) );
  INV_X1 U23423 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20347) );
  AOI22_X1 U23424 ( .A1(n20361), .A2(n20634), .B1(n20360), .B2(n20633), .ZN(
        n20346) );
  AOI22_X1 U23425 ( .A1(n20362), .A2(n20502), .B1(n20388), .B2(n20635), .ZN(
        n20345) );
  OAI211_X1 U23426 ( .C1(n20365), .C2(n20347), .A(n20346), .B(n20345), .ZN(
        P2_U3106) );
  INV_X1 U23427 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n20350) );
  AOI22_X1 U23428 ( .A1(n20361), .A2(n20640), .B1(n20360), .B2(n20639), .ZN(
        n20349) );
  AOI22_X1 U23429 ( .A1(n20362), .A2(n20505), .B1(n20388), .B2(n20641), .ZN(
        n20348) );
  OAI211_X1 U23430 ( .C1(n20365), .C2(n20350), .A(n20349), .B(n20348), .ZN(
        P2_U3107) );
  INV_X1 U23431 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n20353) );
  AOI22_X1 U23432 ( .A1(n20361), .A2(n20646), .B1(n20360), .B2(n20645), .ZN(
        n20352) );
  AOI22_X1 U23433 ( .A1(n20362), .A2(n20508), .B1(n20388), .B2(n20647), .ZN(
        n20351) );
  OAI211_X1 U23434 ( .C1(n20365), .C2(n20353), .A(n20352), .B(n20351), .ZN(
        P2_U3108) );
  INV_X1 U23435 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n20356) );
  AOI22_X1 U23436 ( .A1(n20361), .A2(n20652), .B1(n20360), .B2(n20651), .ZN(
        n20355) );
  AOI22_X1 U23437 ( .A1(n20362), .A2(n20511), .B1(n20388), .B2(n20653), .ZN(
        n20354) );
  OAI211_X1 U23438 ( .C1(n20365), .C2(n20356), .A(n20355), .B(n20354), .ZN(
        P2_U3109) );
  INV_X1 U23439 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n20359) );
  AOI22_X1 U23440 ( .A1(n20361), .A2(n20658), .B1(n20360), .B2(n20657), .ZN(
        n20358) );
  AOI22_X1 U23441 ( .A1(n20362), .A2(n20514), .B1(n20388), .B2(n20659), .ZN(
        n20357) );
  OAI211_X1 U23442 ( .C1(n20365), .C2(n20359), .A(n20358), .B(n20357), .ZN(
        P2_U3110) );
  AOI22_X1 U23443 ( .A1(n20361), .A2(n20665), .B1(n20360), .B2(n20664), .ZN(
        n20364) );
  AOI22_X1 U23444 ( .A1(n20362), .A2(n20519), .B1(n20388), .B2(n20667), .ZN(
        n20363) );
  OAI211_X1 U23445 ( .C1(n20365), .C2(n11642), .A(n20364), .B(n20363), .ZN(
        P2_U3111) );
  INV_X1 U23446 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20369) );
  OAI22_X1 U23447 ( .A1(n20576), .A2(n20426), .B1(n20386), .B2(n20572), .ZN(
        n20366) );
  INV_X1 U23448 ( .A(n20366), .ZN(n20368) );
  AOI22_X1 U23449 ( .A1(n20628), .A2(n20389), .B1(n20388), .B2(n20499), .ZN(
        n20367) );
  OAI211_X1 U23450 ( .C1(n20393), .C2(n20369), .A(n20368), .B(n20367), .ZN(
        P2_U3113) );
  INV_X1 U23451 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20373) );
  OAI22_X1 U23452 ( .A1(n20578), .A2(n20426), .B1(n20386), .B2(n20577), .ZN(
        n20370) );
  INV_X1 U23453 ( .A(n20370), .ZN(n20372) );
  AOI22_X1 U23454 ( .A1(n20634), .A2(n20389), .B1(n20388), .B2(n20502), .ZN(
        n20371) );
  OAI211_X1 U23455 ( .C1(n20393), .C2(n20373), .A(n20372), .B(n20371), .ZN(
        P2_U3114) );
  INV_X1 U23456 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20377) );
  OAI22_X1 U23457 ( .A1(n20586), .A2(n20426), .B1(n20386), .B2(n20582), .ZN(
        n20374) );
  INV_X1 U23458 ( .A(n20374), .ZN(n20376) );
  AOI22_X1 U23459 ( .A1(n20640), .A2(n20389), .B1(n20388), .B2(n20505), .ZN(
        n20375) );
  OAI211_X1 U23460 ( .C1(n20393), .C2(n20377), .A(n20376), .B(n20375), .ZN(
        P2_U3115) );
  OAI22_X1 U23461 ( .A1(n20588), .A2(n20426), .B1(n20386), .B2(n20587), .ZN(
        n20378) );
  INV_X1 U23462 ( .A(n20378), .ZN(n20380) );
  AOI22_X1 U23463 ( .A1(n20646), .A2(n20389), .B1(n20388), .B2(n20508), .ZN(
        n20379) );
  OAI211_X1 U23464 ( .C1(n20393), .C2(n20381), .A(n20380), .B(n20379), .ZN(
        P2_U3116) );
  INV_X1 U23465 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20385) );
  OAI22_X1 U23466 ( .A1(n20596), .A2(n20426), .B1(n20386), .B2(n20592), .ZN(
        n20382) );
  INV_X1 U23467 ( .A(n20382), .ZN(n20384) );
  AOI22_X1 U23468 ( .A1(n20652), .A2(n20389), .B1(n20388), .B2(n20511), .ZN(
        n20383) );
  OAI211_X1 U23469 ( .C1(n20393), .C2(n20385), .A(n20384), .B(n20383), .ZN(
        P2_U3117) );
  INV_X1 U23470 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n20392) );
  OAI22_X1 U23471 ( .A1(n20601), .A2(n20426), .B1(n20386), .B2(n20597), .ZN(
        n20387) );
  INV_X1 U23472 ( .A(n20387), .ZN(n20391) );
  AOI22_X1 U23473 ( .A1(n20658), .A2(n20389), .B1(n20388), .B2(n20514), .ZN(
        n20390) );
  OAI211_X1 U23474 ( .C1(n20393), .C2(n20392), .A(n20391), .B(n20390), .ZN(
        P2_U3118) );
  INV_X1 U23475 ( .A(n20425), .ZN(n20400) );
  AOI22_X1 U23476 ( .A1(n20621), .A2(n20394), .B1(n20613), .B2(n20400), .ZN(
        n20406) );
  OR2_X1 U23477 ( .A1(n20751), .A2(n20395), .ZN(n20616) );
  OAI21_X1 U23478 ( .B1(n20616), .B2(n20396), .A(n20749), .ZN(n20404) );
  INV_X1 U23479 ( .A(n20401), .ZN(n20397) );
  OAI211_X1 U23480 ( .C1(n20397), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20425), 
        .B(n20804), .ZN(n20398) );
  OAI211_X1 U23481 ( .C1(n20404), .C2(n20399), .A(n20619), .B(n20398), .ZN(
        n20429) );
  INV_X1 U23482 ( .A(n20399), .ZN(n20403) );
  OAI21_X1 U23483 ( .B1(n20401), .B2(n20400), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20402) );
  AOI22_X1 U23484 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20429), .B1(
        n20614), .B2(n20428), .ZN(n20405) );
  OAI211_X1 U23485 ( .C1(n20626), .C2(n20432), .A(n20406), .B(n20405), .ZN(
        P2_U3120) );
  OAI22_X1 U23486 ( .A1(n20632), .A2(n20426), .B1(n20572), .B2(n20425), .ZN(
        n20407) );
  INV_X1 U23487 ( .A(n20407), .ZN(n20409) );
  AOI22_X1 U23488 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20429), .B1(
        n20628), .B2(n20428), .ZN(n20408) );
  OAI211_X1 U23489 ( .C1(n20576), .C2(n20432), .A(n20409), .B(n20408), .ZN(
        P2_U3121) );
  OAI22_X1 U23490 ( .A1(n20578), .A2(n20432), .B1(n20425), .B2(n20577), .ZN(
        n20410) );
  INV_X1 U23491 ( .A(n20410), .ZN(n20412) );
  AOI22_X1 U23492 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20429), .B1(
        n20634), .B2(n20428), .ZN(n20411) );
  OAI211_X1 U23493 ( .C1(n20638), .C2(n20426), .A(n20412), .B(n20411), .ZN(
        P2_U3122) );
  OAI22_X1 U23494 ( .A1(n20586), .A2(n20432), .B1(n20582), .B2(n20425), .ZN(
        n20413) );
  INV_X1 U23495 ( .A(n20413), .ZN(n20415) );
  AOI22_X1 U23496 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20429), .B1(
        n20640), .B2(n20428), .ZN(n20414) );
  OAI211_X1 U23497 ( .C1(n20644), .C2(n20426), .A(n20415), .B(n20414), .ZN(
        P2_U3123) );
  OAI22_X1 U23498 ( .A1(n20588), .A2(n20432), .B1(n20587), .B2(n20425), .ZN(
        n20416) );
  INV_X1 U23499 ( .A(n20416), .ZN(n20418) );
  AOI22_X1 U23500 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20429), .B1(
        n20646), .B2(n20428), .ZN(n20417) );
  OAI211_X1 U23501 ( .C1(n20650), .C2(n20426), .A(n20418), .B(n20417), .ZN(
        P2_U3124) );
  OAI22_X1 U23502 ( .A1(n20596), .A2(n20432), .B1(n20592), .B2(n20425), .ZN(
        n20419) );
  INV_X1 U23503 ( .A(n20419), .ZN(n20421) );
  AOI22_X1 U23504 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20429), .B1(
        n20652), .B2(n20428), .ZN(n20420) );
  OAI211_X1 U23505 ( .C1(n20656), .C2(n20426), .A(n20421), .B(n20420), .ZN(
        P2_U3125) );
  OAI22_X1 U23506 ( .A1(n20662), .A2(n20426), .B1(n20597), .B2(n20425), .ZN(
        n20422) );
  INV_X1 U23507 ( .A(n20422), .ZN(n20424) );
  AOI22_X1 U23508 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20429), .B1(
        n20658), .B2(n20428), .ZN(n20423) );
  OAI211_X1 U23509 ( .C1(n20601), .C2(n20432), .A(n20424), .B(n20423), .ZN(
        P2_U3126) );
  OAI22_X1 U23510 ( .A1(n20673), .A2(n20426), .B1(n20602), .B2(n20425), .ZN(
        n20427) );
  INV_X1 U23511 ( .A(n20427), .ZN(n20431) );
  AOI22_X1 U23512 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20429), .B1(
        n20665), .B2(n20428), .ZN(n20430) );
  OAI211_X1 U23513 ( .C1(n20610), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P2_U3127) );
  INV_X1 U23514 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n21657) );
  AOI22_X1 U23515 ( .A1(n20448), .A2(n20614), .B1(n20613), .B2(n20447), .ZN(
        n20434) );
  AOI22_X1 U23516 ( .A1(n20449), .A2(n20621), .B1(n20475), .B2(n20558), .ZN(
        n20433) );
  OAI211_X1 U23517 ( .C1(n20438), .C2(n21657), .A(n20434), .B(n20433), .ZN(
        P2_U3128) );
  INV_X1 U23518 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20437) );
  AOI22_X1 U23519 ( .A1(n20448), .A2(n20634), .B1(n20633), .B2(n20447), .ZN(
        n20436) );
  AOI22_X1 U23520 ( .A1(n20449), .A2(n20502), .B1(n20475), .B2(n20635), .ZN(
        n20435) );
  OAI211_X1 U23521 ( .C1(n20438), .C2(n20437), .A(n20436), .B(n20435), .ZN(
        P2_U3130) );
  AOI22_X1 U23522 ( .A1(n20448), .A2(n20640), .B1(n20639), .B2(n20447), .ZN(
        n20440) );
  AOI22_X1 U23523 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20505), .ZN(n20439) );
  OAI211_X1 U23524 ( .C1(n20586), .C2(n20485), .A(n20440), .B(n20439), .ZN(
        P2_U3131) );
  AOI22_X1 U23525 ( .A1(n20448), .A2(n20646), .B1(n20645), .B2(n20447), .ZN(
        n20442) );
  AOI22_X1 U23526 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20508), .ZN(n20441) );
  OAI211_X1 U23527 ( .C1(n20485), .C2(n20588), .A(n20442), .B(n20441), .ZN(
        P2_U3132) );
  AOI22_X1 U23528 ( .A1(n20448), .A2(n20652), .B1(n20651), .B2(n20447), .ZN(
        n20444) );
  AOI22_X1 U23529 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20511), .ZN(n20443) );
  OAI211_X1 U23530 ( .C1(n20596), .C2(n20485), .A(n20444), .B(n20443), .ZN(
        P2_U3133) );
  AOI22_X1 U23531 ( .A1(n20448), .A2(n20658), .B1(n20657), .B2(n20447), .ZN(
        n20446) );
  AOI22_X1 U23532 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20514), .ZN(n20445) );
  OAI211_X1 U23533 ( .C1(n20485), .C2(n20601), .A(n20446), .B(n20445), .ZN(
        P2_U3134) );
  AOI22_X1 U23534 ( .A1(n20448), .A2(n20665), .B1(n20664), .B2(n20447), .ZN(
        n20452) );
  AOI22_X1 U23535 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20450), .B1(
        n20449), .B2(n20519), .ZN(n20451) );
  OAI211_X1 U23536 ( .C1(n20485), .C2(n20610), .A(n20452), .B(n20451), .ZN(
        P2_U3135) );
  OR2_X1 U23537 ( .A1(n20454), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20459) );
  INV_X1 U23538 ( .A(n20455), .ZN(n20456) );
  NAND2_X1 U23539 ( .A1(n20457), .A2(n20456), .ZN(n20460) );
  NAND2_X1 U23540 ( .A1(n20460), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20458) );
  INV_X1 U23541 ( .A(n20460), .ZN(n20480) );
  AOI22_X1 U23542 ( .A1(n20481), .A2(n20614), .B1(n20613), .B2(n20480), .ZN(
        n20466) );
  INV_X1 U23543 ( .A(n20616), .ZN(n20530) );
  OAI21_X1 U23544 ( .B1(n20480), .B2(n20800), .A(n20619), .ZN(n20461) );
  NOR2_X1 U23545 ( .A1(n20462), .A2(n20461), .ZN(n20463) );
  OAI221_X1 U23546 ( .B1(n20464), .B2(n20746), .C1(n20464), .C2(n20530), .A(
        n20463), .ZN(n20482) );
  AOI22_X1 U23547 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20482), .B1(
        n20475), .B2(n20621), .ZN(n20465) );
  OAI211_X1 U23548 ( .C1(n20626), .C2(n20490), .A(n20466), .B(n20465), .ZN(
        P2_U3136) );
  AOI22_X1 U23549 ( .A1(n20481), .A2(n20628), .B1(n20627), .B2(n20480), .ZN(
        n20468) );
  AOI22_X1 U23550 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20482), .B1(
        n20475), .B2(n20499), .ZN(n20467) );
  OAI211_X1 U23551 ( .C1(n20490), .C2(n20576), .A(n20468), .B(n20467), .ZN(
        P2_U3137) );
  AOI22_X1 U23552 ( .A1(n20481), .A2(n20634), .B1(n20633), .B2(n20480), .ZN(
        n20470) );
  AOI22_X1 U23553 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20482), .B1(
        n20475), .B2(n20502), .ZN(n20469) );
  OAI211_X1 U23554 ( .C1(n20490), .C2(n20578), .A(n20470), .B(n20469), .ZN(
        P2_U3138) );
  AOI22_X1 U23555 ( .A1(n20481), .A2(n20640), .B1(n20639), .B2(n20480), .ZN(
        n20472) );
  AOI22_X1 U23556 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20482), .B1(
        n20475), .B2(n20505), .ZN(n20471) );
  OAI211_X1 U23557 ( .C1(n20586), .C2(n20490), .A(n20472), .B(n20471), .ZN(
        P2_U3139) );
  AOI22_X1 U23558 ( .A1(n20481), .A2(n20646), .B1(n20645), .B2(n20480), .ZN(
        n20474) );
  AOI22_X1 U23559 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20482), .B1(
        n20520), .B2(n20647), .ZN(n20473) );
  OAI211_X1 U23560 ( .C1(n20485), .C2(n20650), .A(n20474), .B(n20473), .ZN(
        P2_U3140) );
  AOI22_X1 U23561 ( .A1(n20481), .A2(n20652), .B1(n20651), .B2(n20480), .ZN(
        n20477) );
  AOI22_X1 U23562 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20482), .B1(
        n20475), .B2(n20511), .ZN(n20476) );
  OAI211_X1 U23563 ( .C1(n20596), .C2(n20490), .A(n20477), .B(n20476), .ZN(
        P2_U3141) );
  AOI22_X1 U23564 ( .A1(n20481), .A2(n20658), .B1(n20657), .B2(n20480), .ZN(
        n20479) );
  AOI22_X1 U23565 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20482), .B1(
        n20520), .B2(n20659), .ZN(n20478) );
  OAI211_X1 U23566 ( .C1(n9921), .C2(n20485), .A(n20479), .B(n20478), .ZN(
        P2_U3142) );
  AOI22_X1 U23567 ( .A1(n20481), .A2(n20665), .B1(n20664), .B2(n20480), .ZN(
        n20484) );
  AOI22_X1 U23568 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20482), .B1(
        n20520), .B2(n20667), .ZN(n20483) );
  OAI211_X1 U23569 ( .C1(n20673), .C2(n20485), .A(n20484), .B(n20483), .ZN(
        P2_U3143) );
  NAND3_X1 U23570 ( .A1(n20776), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20531) );
  NOR2_X1 U23571 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20531), .ZN(
        n20517) );
  INV_X1 U23572 ( .A(n20486), .ZN(n20488) );
  INV_X1 U23573 ( .A(n20492), .ZN(n20487) );
  OAI22_X1 U23574 ( .A1(n20495), .A2(n20489), .B1(n20488), .B2(n20487), .ZN(
        n20518) );
  AOI22_X1 U23575 ( .A1(n20518), .A2(n20614), .B1(n20613), .B2(n20517), .ZN(
        n20498) );
  AOI21_X1 U23576 ( .B1(n20555), .B2(n20490), .A(n20395), .ZN(n20491) );
  AOI21_X1 U23577 ( .B1(n20492), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n20491), .ZN(n20493) );
  AOI211_X1 U23578 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20495), .A(n20494), 
        .B(n20493), .ZN(n20496) );
  AOI22_X1 U23579 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20621), .ZN(n20497) );
  OAI211_X1 U23580 ( .C1(n20626), .C2(n20555), .A(n20498), .B(n20497), .ZN(
        P2_U3144) );
  AOI22_X1 U23581 ( .A1(n20518), .A2(n20628), .B1(n20627), .B2(n20517), .ZN(
        n20501) );
  AOI22_X1 U23582 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20499), .ZN(n20500) );
  OAI211_X1 U23583 ( .C1(n20576), .C2(n20555), .A(n20501), .B(n20500), .ZN(
        P2_U3145) );
  AOI22_X1 U23584 ( .A1(n20518), .A2(n20634), .B1(n20633), .B2(n20517), .ZN(
        n20504) );
  AOI22_X1 U23585 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20502), .ZN(n20503) );
  OAI211_X1 U23586 ( .C1(n20578), .C2(n20555), .A(n20504), .B(n20503), .ZN(
        P2_U3146) );
  AOI22_X1 U23587 ( .A1(n20518), .A2(n20640), .B1(n20639), .B2(n20517), .ZN(
        n20507) );
  AOI22_X1 U23588 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20505), .ZN(n20506) );
  OAI211_X1 U23589 ( .C1(n20586), .C2(n20555), .A(n20507), .B(n20506), .ZN(
        P2_U3147) );
  AOI22_X1 U23590 ( .A1(n20518), .A2(n20646), .B1(n20645), .B2(n20517), .ZN(
        n20510) );
  AOI22_X1 U23591 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20508), .ZN(n20509) );
  OAI211_X1 U23592 ( .C1(n20588), .C2(n20555), .A(n20510), .B(n20509), .ZN(
        P2_U3148) );
  AOI22_X1 U23593 ( .A1(n20518), .A2(n20652), .B1(n20651), .B2(n20517), .ZN(
        n20513) );
  AOI22_X1 U23594 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20511), .ZN(n20512) );
  OAI211_X1 U23595 ( .C1(n20596), .C2(n20555), .A(n20513), .B(n20512), .ZN(
        P2_U3149) );
  AOI22_X1 U23596 ( .A1(n20518), .A2(n20658), .B1(n20657), .B2(n20517), .ZN(
        n20516) );
  AOI22_X1 U23597 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20514), .ZN(n20515) );
  OAI211_X1 U23598 ( .C1(n20601), .C2(n20555), .A(n20516), .B(n20515), .ZN(
        P2_U3150) );
  AOI22_X1 U23599 ( .A1(n20518), .A2(n20665), .B1(n20664), .B2(n20517), .ZN(
        n20523) );
  AOI22_X1 U23600 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20521), .B1(
        n20520), .B2(n20519), .ZN(n20522) );
  OAI211_X1 U23601 ( .C1(n20610), .C2(n20555), .A(n20523), .B(n20522), .ZN(
        P2_U3151) );
  OR2_X1 U23602 ( .A1(n20531), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20528) );
  INV_X1 U23603 ( .A(n20524), .ZN(n20526) );
  NOR2_X1 U23604 ( .A1(n20786), .A2(n20531), .ZN(n20562) );
  INV_X1 U23605 ( .A(n20562), .ZN(n20525) );
  NAND3_X1 U23606 ( .A1(n20526), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20525), 
        .ZN(n20533) );
  INV_X1 U23607 ( .A(n20533), .ZN(n20527) );
  AOI22_X1 U23608 ( .A1(n20551), .A2(n20614), .B1(n20613), .B2(n20562), .ZN(
        n20538) );
  INV_X1 U23609 ( .A(n20535), .ZN(n20529) );
  NAND2_X1 U23610 ( .A1(n20530), .A2(n20529), .ZN(n20532) );
  AOI21_X1 U23611 ( .B1(n20532), .B2(n20531), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n20534) );
  AOI22_X1 U23612 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20558), .ZN(n20537) );
  OAI211_X1 U23613 ( .C1(n20571), .C2(n20555), .A(n20538), .B(n20537), .ZN(
        P2_U3152) );
  AOI22_X1 U23614 ( .A1(n20551), .A2(n20628), .B1(n20627), .B2(n20562), .ZN(
        n20540) );
  AOI22_X1 U23615 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20629), .ZN(n20539) );
  OAI211_X1 U23616 ( .C1(n20632), .C2(n20555), .A(n20540), .B(n20539), .ZN(
        P2_U3153) );
  AOI22_X1 U23617 ( .A1(n20551), .A2(n20634), .B1(n20633), .B2(n20562), .ZN(
        n20542) );
  AOI22_X1 U23618 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20635), .ZN(n20541) );
  OAI211_X1 U23619 ( .C1(n20638), .C2(n20555), .A(n20542), .B(n20541), .ZN(
        P2_U3154) );
  AOI22_X1 U23620 ( .A1(n20551), .A2(n20640), .B1(n20639), .B2(n20562), .ZN(
        n20544) );
  AOI22_X1 U23621 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20641), .ZN(n20543) );
  OAI211_X1 U23622 ( .C1(n20644), .C2(n20555), .A(n20544), .B(n20543), .ZN(
        P2_U3155) );
  AOI22_X1 U23623 ( .A1(n20551), .A2(n20646), .B1(n20645), .B2(n20562), .ZN(
        n20546) );
  AOI22_X1 U23624 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20647), .ZN(n20545) );
  OAI211_X1 U23625 ( .C1(n20650), .C2(n20555), .A(n20546), .B(n20545), .ZN(
        P2_U3156) );
  AOI22_X1 U23626 ( .A1(n20551), .A2(n20652), .B1(n20651), .B2(n20562), .ZN(
        n20548) );
  AOI22_X1 U23627 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20653), .ZN(n20547) );
  OAI211_X1 U23628 ( .C1(n20656), .C2(n20555), .A(n20548), .B(n20547), .ZN(
        P2_U3157) );
  AOI22_X1 U23629 ( .A1(n20551), .A2(n20658), .B1(n20657), .B2(n20562), .ZN(
        n20550) );
  AOI22_X1 U23630 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20659), .ZN(n20549) );
  OAI211_X1 U23631 ( .C1(n9921), .C2(n20555), .A(n20550), .B(n20549), .ZN(
        P2_U3158) );
  AOI22_X1 U23632 ( .A1(n20551), .A2(n20665), .B1(n20664), .B2(n20562), .ZN(
        n20554) );
  AOI22_X1 U23633 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20552), .B1(
        n20559), .B2(n20667), .ZN(n20553) );
  OAI211_X1 U23634 ( .C1(n20673), .C2(n20555), .A(n20554), .B(n20553), .ZN(
        P2_U3159) );
  NAND2_X1 U23635 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20557), .ZN(
        n20615) );
  NOR2_X1 U23636 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20615), .ZN(
        n20565) );
  AOI22_X1 U23637 ( .A1(n20558), .A2(n20622), .B1(n20613), .B2(n20565), .ZN(
        n20570) );
  NOR3_X1 U23638 ( .A1(n20622), .A2(n20559), .A3(n20804), .ZN(n20561) );
  INV_X1 U23639 ( .A(n20748), .ZN(n20560) );
  NOR2_X1 U23640 ( .A1(n20561), .A2(n20560), .ZN(n20568) );
  NOR2_X1 U23641 ( .A1(n20565), .A2(n20562), .ZN(n20567) );
  INV_X1 U23642 ( .A(n20567), .ZN(n20564) );
  INV_X1 U23643 ( .A(n20565), .ZN(n20603) );
  OAI211_X1 U23644 ( .C1(n20568), .C2(n20564), .A(n20619), .B(n20563), .ZN(
        n20607) );
  OAI21_X1 U23645 ( .B1(n9801), .B2(n20565), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20566) );
  AOI22_X1 U23646 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20607), .B1(
        n20614), .B2(n20606), .ZN(n20569) );
  OAI211_X1 U23647 ( .C1(n20571), .C2(n20604), .A(n20570), .B(n20569), .ZN(
        P2_U3160) );
  OAI22_X1 U23648 ( .A1(n20632), .A2(n20604), .B1(n20572), .B2(n20603), .ZN(
        n20573) );
  INV_X1 U23649 ( .A(n20573), .ZN(n20575) );
  AOI22_X1 U23650 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20607), .B1(
        n20628), .B2(n20606), .ZN(n20574) );
  OAI211_X1 U23651 ( .C1(n20576), .C2(n20672), .A(n20575), .B(n20574), .ZN(
        P2_U3161) );
  OAI22_X1 U23652 ( .A1(n20578), .A2(n20672), .B1(n20577), .B2(n20603), .ZN(
        n20579) );
  INV_X1 U23653 ( .A(n20579), .ZN(n20581) );
  AOI22_X1 U23654 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20607), .B1(
        n20634), .B2(n20606), .ZN(n20580) );
  OAI211_X1 U23655 ( .C1(n20638), .C2(n20604), .A(n20581), .B(n20580), .ZN(
        P2_U3162) );
  OAI22_X1 U23656 ( .A1(n20644), .A2(n20604), .B1(n20582), .B2(n20603), .ZN(
        n20583) );
  INV_X1 U23657 ( .A(n20583), .ZN(n20585) );
  AOI22_X1 U23658 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20607), .B1(
        n20640), .B2(n20606), .ZN(n20584) );
  OAI211_X1 U23659 ( .C1(n20586), .C2(n20672), .A(n20585), .B(n20584), .ZN(
        P2_U3163) );
  OAI22_X1 U23660 ( .A1(n20588), .A2(n20672), .B1(n20587), .B2(n20603), .ZN(
        n20589) );
  INV_X1 U23661 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23662 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20607), .B1(
        n20646), .B2(n20606), .ZN(n20590) );
  OAI211_X1 U23663 ( .C1(n20650), .C2(n20604), .A(n20591), .B(n20590), .ZN(
        P2_U3164) );
  OAI22_X1 U23664 ( .A1(n20656), .A2(n20604), .B1(n20592), .B2(n20603), .ZN(
        n20593) );
  INV_X1 U23665 ( .A(n20593), .ZN(n20595) );
  AOI22_X1 U23666 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20607), .B1(
        n20652), .B2(n20606), .ZN(n20594) );
  OAI211_X1 U23667 ( .C1(n20596), .C2(n20672), .A(n20595), .B(n20594), .ZN(
        P2_U3165) );
  OAI22_X1 U23668 ( .A1(n9921), .A2(n20604), .B1(n20597), .B2(n20603), .ZN(
        n20598) );
  INV_X1 U23669 ( .A(n20598), .ZN(n20600) );
  AOI22_X1 U23670 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20607), .B1(
        n20658), .B2(n20606), .ZN(n20599) );
  OAI211_X1 U23671 ( .C1(n20601), .C2(n20672), .A(n20600), .B(n20599), .ZN(
        P2_U3166) );
  OAI22_X1 U23672 ( .A1(n20673), .A2(n20604), .B1(n20603), .B2(n20602), .ZN(
        n20605) );
  INV_X1 U23673 ( .A(n20605), .ZN(n20609) );
  AOI22_X1 U23674 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20607), .B1(
        n20665), .B2(n20606), .ZN(n20608) );
  OAI211_X1 U23675 ( .C1(n20610), .C2(n20672), .A(n20609), .B(n20608), .ZN(
        P2_U3167) );
  OR2_X1 U23676 ( .A1(n20663), .A2(n20489), .ZN(n20611) );
  OAI21_X1 U23677 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20615), .A(n20489), 
        .ZN(n20612) );
  AND2_X1 U23678 ( .A1(n20618), .A2(n20612), .ZN(n20666) );
  AOI22_X1 U23679 ( .A1(n20666), .A2(n20614), .B1(n20613), .B2(n20663), .ZN(
        n20624) );
  OAI21_X1 U23680 ( .B1(n20616), .B2(n20752), .A(n20615), .ZN(n20620) );
  OR2_X1 U23681 ( .A1(n20663), .A2(n20800), .ZN(n20617) );
  NAND4_X1 U23682 ( .A1(n20620), .A2(n20619), .A3(n20618), .A4(n20617), .ZN(
        n20669) );
  AOI22_X1 U23683 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20669), .B1(
        n20622), .B2(n20621), .ZN(n20623) );
  OAI211_X1 U23684 ( .C1(n20626), .C2(n20625), .A(n20624), .B(n20623), .ZN(
        P2_U3168) );
  AOI22_X1 U23685 ( .A1(n20666), .A2(n20628), .B1(n20627), .B2(n20663), .ZN(
        n20631) );
  AOI22_X1 U23686 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20629), .ZN(n20630) );
  OAI211_X1 U23687 ( .C1(n20632), .C2(n20672), .A(n20631), .B(n20630), .ZN(
        P2_U3169) );
  AOI22_X1 U23688 ( .A1(n20666), .A2(n20634), .B1(n20633), .B2(n20663), .ZN(
        n20637) );
  AOI22_X1 U23689 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20635), .ZN(n20636) );
  OAI211_X1 U23690 ( .C1(n20638), .C2(n20672), .A(n20637), .B(n20636), .ZN(
        P2_U3170) );
  AOI22_X1 U23691 ( .A1(n20666), .A2(n20640), .B1(n20639), .B2(n20663), .ZN(
        n20643) );
  AOI22_X1 U23692 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20641), .ZN(n20642) );
  OAI211_X1 U23693 ( .C1(n20644), .C2(n20672), .A(n20643), .B(n20642), .ZN(
        P2_U3171) );
  AOI22_X1 U23694 ( .A1(n20666), .A2(n20646), .B1(n20645), .B2(n20663), .ZN(
        n20649) );
  AOI22_X1 U23695 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20647), .ZN(n20648) );
  OAI211_X1 U23696 ( .C1(n20650), .C2(n20672), .A(n20649), .B(n20648), .ZN(
        P2_U3172) );
  AOI22_X1 U23697 ( .A1(n20666), .A2(n20652), .B1(n20651), .B2(n20663), .ZN(
        n20655) );
  AOI22_X1 U23698 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20653), .ZN(n20654) );
  OAI211_X1 U23699 ( .C1(n20656), .C2(n20672), .A(n20655), .B(n20654), .ZN(
        P2_U3173) );
  AOI22_X1 U23700 ( .A1(n20666), .A2(n20658), .B1(n20657), .B2(n20663), .ZN(
        n20661) );
  AOI22_X1 U23701 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20659), .ZN(n20660) );
  OAI211_X1 U23702 ( .C1(n9921), .C2(n20672), .A(n20661), .B(n20660), .ZN(
        P2_U3174) );
  AOI22_X1 U23703 ( .A1(n20666), .A2(n20665), .B1(n20664), .B2(n20663), .ZN(
        n20671) );
  AOI22_X1 U23704 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20669), .B1(
        n20668), .B2(n20667), .ZN(n20670) );
  OAI211_X1 U23705 ( .C1(n20673), .C2(n20672), .A(n20671), .B(n20670), .ZN(
        P2_U3175) );
  AND2_X1 U23706 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20674), .ZN(
        P2_U3179) );
  AND2_X1 U23707 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20674), .ZN(
        P2_U3180) );
  AND2_X1 U23708 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20674), .ZN(
        P2_U3181) );
  AND2_X1 U23709 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20674), .ZN(
        P2_U3182) );
  AND2_X1 U23710 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20674), .ZN(
        P2_U3183) );
  AND2_X1 U23711 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20674), .ZN(
        P2_U3184) );
  AND2_X1 U23712 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20674), .ZN(
        P2_U3185) );
  AND2_X1 U23713 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20674), .ZN(
        P2_U3186) );
  AND2_X1 U23714 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20674), .ZN(
        P2_U3187) );
  AND2_X1 U23715 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20674), .ZN(
        P2_U3188) );
  AND2_X1 U23716 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20674), .ZN(
        P2_U3189) );
  AND2_X1 U23717 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20674), .ZN(
        P2_U3190) );
  AND2_X1 U23718 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20674), .ZN(
        P2_U3191) );
  AND2_X1 U23719 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20674), .ZN(
        P2_U3192) );
  NOR2_X1 U23720 ( .A1(n21668), .A2(n20745), .ZN(P2_U3193) );
  AND2_X1 U23721 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20674), .ZN(
        P2_U3194) );
  AND2_X1 U23722 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20674), .ZN(
        P2_U3195) );
  AND2_X1 U23723 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20674), .ZN(
        P2_U3196) );
  AND2_X1 U23724 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20674), .ZN(
        P2_U3197) );
  AND2_X1 U23725 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20674), .ZN(
        P2_U3198) );
  AND2_X1 U23726 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20674), .ZN(
        P2_U3199) );
  AND2_X1 U23727 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20674), .ZN(
        P2_U3200) );
  NOR2_X1 U23728 ( .A1(n21801), .A2(n20745), .ZN(P2_U3201) );
  AND2_X1 U23729 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20674), .ZN(P2_U3202) );
  AND2_X1 U23730 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20674), .ZN(P2_U3203) );
  AND2_X1 U23731 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20674), .ZN(P2_U3204) );
  AND2_X1 U23732 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20674), .ZN(P2_U3205) );
  AND2_X1 U23733 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20674), .ZN(P2_U3206) );
  AND2_X1 U23734 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20674), .ZN(P2_U3207) );
  AND2_X1 U23735 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20674), .ZN(P2_U3208) );
  INV_X1 U23736 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20816) );
  NOR2_X1 U23737 ( .A1(n20812), .A2(n20684), .ZN(n20682) );
  OR3_X1 U23738 ( .A1(n20816), .A2(n20675), .A3(n20682), .ZN(n20676) );
  NOR3_X1 U23739 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21485), .ZN(n20689) );
  AOI21_X1 U23740 ( .B1(n21751), .B2(n20676), .A(n20689), .ZN(n20677) );
  OAI221_X1 U23741 ( .B1(n20678), .B2(P2_REQUESTPENDING_REG_SCAN_IN), .C1(
        n20678), .C2(n21491), .A(n20677), .ZN(P2_U3209) );
  AOI21_X1 U23742 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21491), .A(n21751), 
        .ZN(n20685) );
  NOR3_X1 U23743 ( .A1(n20685), .A2(n20816), .A3(n20675), .ZN(n20679) );
  NOR2_X1 U23744 ( .A1(n20679), .A2(n20682), .ZN(n20680) );
  OAI211_X1 U23745 ( .C1(n21491), .C2(n20681), .A(n20680), .B(n20806), .ZN(
        P2_U3210) );
  AOI22_X1 U23746 ( .A1(n20683), .A2(n20816), .B1(n20682), .B2(n21485), .ZN(
        n20691) );
  OAI21_X1 U23747 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20690) );
  NOR2_X1 U23748 ( .A1(n21751), .A2(n20684), .ZN(n20687) );
  AOI21_X1 U23749 ( .B1(n20687), .B2(n20686), .A(n20685), .ZN(n20688) );
  OAI22_X1 U23750 ( .A1(n20691), .A2(n20690), .B1(n20689), .B2(n20688), .ZN(
        P2_U3211) );
  OAI222_X1 U23751 ( .A1(n20733), .A2(n20694), .B1(n20693), .B2(n20788), .C1(
        n20692), .C2(n20734), .ZN(P2_U3212) );
  OAI222_X1 U23752 ( .A1(n20733), .A2(n11505), .B1(n20695), .B2(n20788), .C1(
        n20694), .C2(n20734), .ZN(P2_U3213) );
  OAI222_X1 U23753 ( .A1(n20733), .A2(n16465), .B1(n20696), .B2(n20788), .C1(
        n11505), .C2(n20734), .ZN(P2_U3214) );
  OAI222_X1 U23754 ( .A1(n20733), .A2(n15925), .B1(n20697), .B2(n20788), .C1(
        n16465), .C2(n20734), .ZN(P2_U3215) );
  OAI222_X1 U23755 ( .A1(n20733), .A2(n20698), .B1(n21790), .B2(n20788), .C1(
        n15925), .C2(n20734), .ZN(P2_U3216) );
  OAI222_X1 U23756 ( .A1(n20733), .A2(n20700), .B1(n20699), .B2(n20788), .C1(
        n20698), .C2(n20734), .ZN(P2_U3217) );
  OAI222_X1 U23757 ( .A1(n20733), .A2(n20702), .B1(n20701), .B2(n20788), .C1(
        n20700), .C2(n20734), .ZN(P2_U3218) );
  OAI222_X1 U23758 ( .A1(n20733), .A2(n15879), .B1(n20703), .B2(n20788), .C1(
        n20702), .C2(n20734), .ZN(P2_U3219) );
  OAI222_X1 U23759 ( .A1(n20733), .A2(n20705), .B1(n20704), .B2(n20788), .C1(
        n15879), .C2(n20734), .ZN(P2_U3220) );
  OAI222_X1 U23760 ( .A1(n20733), .A2(n21738), .B1(n20706), .B2(n20788), .C1(
        n20705), .C2(n20734), .ZN(P2_U3221) );
  OAI222_X1 U23761 ( .A1(n20733), .A2(n20708), .B1(n20707), .B2(n20788), .C1(
        n21738), .C2(n20734), .ZN(P2_U3222) );
  OAI222_X1 U23762 ( .A1(n20733), .A2(n11973), .B1(n20709), .B2(n20788), .C1(
        n20708), .C2(n20734), .ZN(P2_U3223) );
  OAI222_X1 U23763 ( .A1(n20733), .A2(n15833), .B1(n20710), .B2(n20788), .C1(
        n11973), .C2(n20734), .ZN(P2_U3224) );
  OAI222_X1 U23764 ( .A1(n20733), .A2(n20712), .B1(n20711), .B2(n20788), .C1(
        n15833), .C2(n20734), .ZN(P2_U3225) );
  OAI222_X1 U23765 ( .A1(n20733), .A2(n15798), .B1(n20713), .B2(n20788), .C1(
        n20712), .C2(n20734), .ZN(P2_U3226) );
  OAI222_X1 U23766 ( .A1(n20733), .A2(n20715), .B1(n20714), .B2(n20788), .C1(
        n15798), .C2(n20734), .ZN(P2_U3227) );
  OAI222_X1 U23767 ( .A1(n20733), .A2(n12228), .B1(n20716), .B2(n20788), .C1(
        n20715), .C2(n20734), .ZN(P2_U3228) );
  OAI222_X1 U23768 ( .A1(n20733), .A2(n20718), .B1(n20717), .B2(n20788), .C1(
        n12228), .C2(n20734), .ZN(P2_U3229) );
  OAI222_X1 U23769 ( .A1(n20733), .A2(n11996), .B1(n20719), .B2(n20788), .C1(
        n20718), .C2(n20734), .ZN(P2_U3230) );
  OAI222_X1 U23770 ( .A1(n20733), .A2(n21847), .B1(n20720), .B2(n20788), .C1(
        n11996), .C2(n20734), .ZN(P2_U3231) );
  OAI222_X1 U23771 ( .A1(n20733), .A2(n12238), .B1(n20721), .B2(n20788), .C1(
        n21847), .C2(n20734), .ZN(P2_U3232) );
  OAI222_X1 U23772 ( .A1(n20733), .A2(n21725), .B1(n20722), .B2(n20788), .C1(
        n12238), .C2(n20734), .ZN(P2_U3233) );
  OAI222_X1 U23773 ( .A1(n20733), .A2(n21822), .B1(n20723), .B2(n20788), .C1(
        n21725), .C2(n20734), .ZN(P2_U3234) );
  OAI222_X1 U23774 ( .A1(n20733), .A2(n20725), .B1(n20724), .B2(n20788), .C1(
        n21822), .C2(n20734), .ZN(P2_U3235) );
  OAI222_X1 U23775 ( .A1(n20733), .A2(n20726), .B1(n21817), .B2(n20788), .C1(
        n20725), .C2(n20734), .ZN(P2_U3236) );
  OAI222_X1 U23776 ( .A1(n20733), .A2(n20729), .B1(n20727), .B2(n20788), .C1(
        n20726), .C2(n20734), .ZN(P2_U3237) );
  OAI222_X1 U23777 ( .A1(n20734), .A2(n20729), .B1(n20728), .B2(n20788), .C1(
        n12369), .C2(n20733), .ZN(P2_U3238) );
  OAI222_X1 U23778 ( .A1(n20733), .A2(n20731), .B1(n20730), .B2(n20788), .C1(
        n12369), .C2(n20734), .ZN(P2_U3239) );
  OAI222_X1 U23779 ( .A1(n20733), .A2(n16218), .B1(n20732), .B2(n20788), .C1(
        n20731), .C2(n20734), .ZN(P2_U3240) );
  OAI222_X1 U23780 ( .A1(n20733), .A2(n12381), .B1(n20735), .B2(n20788), .C1(
        n16218), .C2(n20734), .ZN(P2_U3241) );
  INV_X1 U23781 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20736) );
  AOI22_X1 U23782 ( .A1(n20788), .A2(n21707), .B1(n20736), .B2(n20818), .ZN(
        P2_U3585) );
  INV_X1 U23783 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21673) );
  INV_X1 U23784 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n20737) );
  AOI22_X1 U23785 ( .A1(n20788), .A2(n21673), .B1(n20737), .B2(n20818), .ZN(
        P2_U3586) );
  INV_X1 U23786 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20738) );
  AOI22_X1 U23787 ( .A1(n20788), .A2(n20739), .B1(n20738), .B2(n20818), .ZN(
        P2_U3587) );
  INV_X1 U23788 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20740) );
  AOI22_X1 U23789 ( .A1(n20788), .A2(n20741), .B1(n20740), .B2(n20818), .ZN(
        P2_U3588) );
  OAI21_X1 U23790 ( .B1(n20745), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20743), 
        .ZN(n20742) );
  INV_X1 U23791 ( .A(n20742), .ZN(P2_U3591) );
  OAI21_X1 U23792 ( .B1(n20745), .B2(n20744), .A(n20743), .ZN(P2_U3592) );
  NAND2_X1 U23793 ( .A1(n20746), .A2(n20767), .ZN(n20764) );
  NAND2_X1 U23794 ( .A1(n20748), .A2(n20747), .ZN(n20768) );
  AOI21_X1 U23795 ( .B1(n20750), .B2(n20749), .A(n20768), .ZN(n20759) );
  AOI21_X1 U23796 ( .B1(n20764), .B2(n20759), .A(n20751), .ZN(n20755) );
  NOR3_X1 U23797 ( .A1(n20753), .A2(n20804), .A3(n20752), .ZN(n20754) );
  AOI211_X1 U23798 ( .C1(n20756), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n20755), 
        .B(n20754), .ZN(n20757) );
  INV_X1 U23799 ( .A(n20784), .ZN(n20785) );
  AOI22_X1 U23800 ( .A1(n20784), .A2(n20758), .B1(n20757), .B2(n20785), .ZN(
        P2_U3602) );
  INV_X1 U23801 ( .A(n20759), .ZN(n20761) );
  AOI22_X1 U23802 ( .A1(n20762), .A2(n20761), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20760), .ZN(n20763) );
  AND2_X1 U23803 ( .A1(n20764), .A2(n20763), .ZN(n20765) );
  AOI22_X1 U23804 ( .A1(n20784), .A2(n20766), .B1(n20765), .B2(n20785), .ZN(
        P2_U3603) );
  INV_X1 U23805 ( .A(n20767), .ZN(n20771) );
  INV_X1 U23806 ( .A(n20768), .ZN(n20770) );
  MUX2_X1 U23807 ( .A(n20771), .B(n20770), .S(n20769), .Z(n20774) );
  NAND2_X1 U23808 ( .A1(n20772), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20773) );
  AND2_X1 U23809 ( .A1(n20774), .A2(n20773), .ZN(n20775) );
  AOI22_X1 U23810 ( .A1(n20784), .A2(n20776), .B1(n20775), .B2(n20785), .ZN(
        P2_U3604) );
  INV_X1 U23811 ( .A(n20777), .ZN(n20780) );
  OAI22_X1 U23812 ( .A1(n20781), .A2(n20780), .B1(n20779), .B2(n20778), .ZN(
        n20782) );
  AOI21_X1 U23813 ( .B1(n20786), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20782), 
        .ZN(n20783) );
  OAI22_X1 U23814 ( .A1(n20786), .A2(n20785), .B1(n20784), .B2(n20783), .ZN(
        P2_U3605) );
  INV_X1 U23815 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20787) );
  AOI22_X1 U23816 ( .A1(n20788), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20787), 
        .B2(n20818), .ZN(P2_U3608) );
  INV_X1 U23817 ( .A(n20789), .ZN(n20792) );
  OAI22_X1 U23818 ( .A1(n20793), .A2(n20792), .B1(n20791), .B2(n20790), .ZN(
        n20794) );
  INV_X1 U23819 ( .A(n20794), .ZN(n20795) );
  NAND2_X1 U23820 ( .A1(n20796), .A2(n20795), .ZN(n20798) );
  MUX2_X1 U23821 ( .A(P2_MORE_REG_SCAN_IN), .B(n20798), .S(n20797), .Z(
        P2_U3609) );
  NAND2_X1 U23822 ( .A1(n20799), .A2(n20812), .ZN(n20803) );
  NAND2_X1 U23823 ( .A1(n20801), .A2(n20800), .ZN(n20802) );
  NAND4_X1 U23824 ( .A1(n20805), .A2(n20804), .A3(n20803), .A4(n20802), .ZN(
        n20817) );
  AOI21_X1 U23825 ( .B1(n20807), .B2(n20395), .A(n20806), .ZN(n20809) );
  NOR3_X1 U23826 ( .A1(n20810), .A2(n20809), .A3(n20808), .ZN(n20814) );
  AOI21_X1 U23827 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20812), .A(n20811), 
        .ZN(n20813) );
  OAI21_X1 U23828 ( .B1(n20814), .B2(n20813), .A(n20817), .ZN(n20815) );
  OAI21_X1 U23829 ( .B1(n20817), .B2(n20816), .A(n20815), .ZN(P2_U3610) );
  INV_X1 U23830 ( .A(P2_M_IO_N_REG_SCAN_IN), .ZN(n20819) );
  AOI22_X1 U23831 ( .A1(n20788), .A2(n20820), .B1(n20819), .B2(n20818), .ZN(
        P2_U3611) );
  AOI21_X1 U23832 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21494), .A(n21486), 
        .ZN(n21489) );
  INV_X1 U23833 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20821) );
  INV_X2 U23834 ( .A(n21570), .ZN(n21583) );
  AOI21_X1 U23835 ( .B1(n21489), .B2(n20821), .A(n21583), .ZN(P1_U2802) );
  OAI21_X1 U23836 ( .B1(n20823), .B2(n20822), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20824) );
  OAI21_X1 U23837 ( .B1(n20826), .B2(n20825), .A(n20824), .ZN(P1_U2803) );
  NOR2_X1 U23838 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20828) );
  OAI21_X1 U23839 ( .B1(n20828), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21570), .ZN(
        n20827) );
  OAI21_X1 U23840 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21570), .A(n20827), 
        .ZN(P1_U2804) );
  NOR2_X1 U23841 ( .A1(n21489), .A2(n21583), .ZN(n21560) );
  OAI21_X1 U23842 ( .B1(BS16), .B2(n20828), .A(n21560), .ZN(n21558) );
  OAI21_X1 U23843 ( .B1(n21560), .B2(n21173), .A(n21558), .ZN(P1_U2805) );
  OAI21_X1 U23844 ( .B1(n20831), .B2(n20830), .A(n20829), .ZN(P1_U2806) );
  NOR4_X1 U23845 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20835) );
  NOR4_X1 U23846 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20834) );
  NOR4_X1 U23847 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20833) );
  NOR4_X1 U23848 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20832) );
  NAND4_X1 U23849 ( .A1(n20835), .A2(n20834), .A3(n20833), .A4(n20832), .ZN(
        n20841) );
  NOR4_X1 U23850 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20839) );
  AOI211_X1 U23851 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20838) );
  NOR4_X1 U23852 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20837) );
  NOR4_X1 U23853 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20836) );
  NAND4_X1 U23854 ( .A1(n20839), .A2(n20838), .A3(n20837), .A4(n20836), .ZN(
        n20840) );
  NOR2_X1 U23855 ( .A1(n20841), .A2(n20840), .ZN(n21569) );
  INV_X1 U23856 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21555) );
  NOR3_X1 U23857 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20843) );
  OAI21_X1 U23858 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20843), .A(n21569), .ZN(
        n20842) );
  OAI21_X1 U23859 ( .B1(n21569), .B2(n21555), .A(n20842), .ZN(P1_U2807) );
  INV_X1 U23860 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21552) );
  NOR2_X1 U23861 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21563) );
  OAI21_X1 U23862 ( .B1(n20843), .B2(n21563), .A(n21569), .ZN(n20844) );
  OAI21_X1 U23863 ( .B1(n21569), .B2(n21552), .A(n20844), .ZN(P1_U2808) );
  AOI22_X1 U23864 ( .A1(n20909), .A2(n20846), .B1(n20845), .B2(n21509), .ZN(
        n20855) );
  INV_X1 U23865 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20929) );
  OAI22_X1 U23866 ( .A1(n20883), .A2(n20929), .B1(n20882), .B2(n20847), .ZN(
        n20848) );
  AOI211_X1 U23867 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20849), .A(n17539), .B(
        n20848), .ZN(n20854) );
  OAI22_X1 U23868 ( .A1(n20926), .A2(n20851), .B1(n20850), .B2(n20897), .ZN(
        n20852) );
  INV_X1 U23869 ( .A(n20852), .ZN(n20853) );
  NAND3_X1 U23870 ( .A1(n20855), .A2(n20854), .A3(n20853), .ZN(P1_U2831) );
  AOI21_X1 U23871 ( .B1(n20858), .B2(n20857), .A(n20856), .ZN(n20886) );
  INV_X1 U23872 ( .A(n20886), .ZN(n20902) );
  AOI21_X1 U23873 ( .B1(n20860), .B2(n20859), .A(n20902), .ZN(n20881) );
  NAND2_X1 U23874 ( .A1(n20907), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n20861) );
  OAI211_X1 U23875 ( .C1(n20882), .C2(n20862), .A(n20861), .B(n20904), .ZN(
        n20865) );
  NOR2_X1 U23876 ( .A1(n20897), .A2(n20863), .ZN(n20864) );
  AOI211_X1 U23877 ( .C1(n20866), .C2(n20909), .A(n20865), .B(n20864), .ZN(
        n20870) );
  AOI22_X1 U23878 ( .A1(n20879), .A2(n20868), .B1(n20867), .B2(n21506), .ZN(
        n20869) );
  OAI211_X1 U23879 ( .C1(n20881), .C2(n21506), .A(n20870), .B(n20869), .ZN(
        P1_U2833) );
  INV_X1 U23880 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21792) );
  AOI22_X1 U23881 ( .A1(n20909), .A2(n20871), .B1(n20907), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20872) );
  OAI21_X1 U23882 ( .B1(n20897), .B2(n20873), .A(n20872), .ZN(n20877) );
  INV_X1 U23883 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21503) );
  NOR3_X1 U23884 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n21503), .A3(n20887), .ZN(
        n20874) );
  AOI211_X1 U23885 ( .C1(n20912), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17539), .B(n20874), .ZN(n20875) );
  INV_X1 U23886 ( .A(n20875), .ZN(n20876) );
  AOI211_X1 U23887 ( .C1(n20879), .C2(n20878), .A(n20877), .B(n20876), .ZN(
        n20880) );
  OAI21_X1 U23888 ( .B1(n20881), .B2(n21792), .A(n20880), .ZN(P1_U2834) );
  INV_X1 U23889 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20935) );
  OAI22_X1 U23890 ( .A1(n20883), .A2(n20935), .B1(n20882), .B2(n21775), .ZN(
        n20884) );
  AOI211_X1 U23891 ( .C1(n20909), .C2(n20930), .A(n17539), .B(n20884), .ZN(
        n20885) );
  OAI221_X1 U23892 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20887), .C1(n21503), 
        .C2(n20886), .A(n20885), .ZN(n20888) );
  AOI21_X1 U23893 ( .B1(n20933), .B2(n20889), .A(n20888), .ZN(n20890) );
  OAI21_X1 U23894 ( .B1(n20891), .B2(n20897), .A(n20890), .ZN(P1_U2835) );
  AOI22_X1 U23895 ( .A1(n20907), .A2(P1_EBX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20912), .ZN(n20906) );
  INV_X1 U23896 ( .A(n20892), .ZN(n20896) );
  OAI22_X1 U23897 ( .A1(n20896), .A2(n20895), .B1(n20894), .B2(n20893), .ZN(
        n20901) );
  OAI22_X1 U23898 ( .A1(n20899), .A2(n20917), .B1(n20898), .B2(n20897), .ZN(
        n20900) );
  AOI211_X1 U23899 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n20902), .A(n20901), .B(
        n20900), .ZN(n20905) );
  NAND4_X1 U23900 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .A3(n20911), .A4(n21500), .ZN(n20903) );
  NAND4_X1 U23901 ( .A1(n20906), .A2(n20905), .A3(n20904), .A4(n20903), .ZN(
        P1_U2836) );
  AOI22_X1 U23902 ( .A1(n20909), .A2(n20908), .B1(n20907), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20922) );
  NAND2_X1 U23903 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20910) );
  OAI211_X1 U23904 ( .C1(P1_REIP_REG_3__SCAN_IN), .C2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20911), .B(n20910), .ZN(n20915) );
  AOI22_X1 U23905 ( .A1(n21167), .A2(n20913), .B1(n20912), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20914) );
  OAI211_X1 U23906 ( .C1(n20917), .C2(n20916), .A(n20915), .B(n20914), .ZN(
        n20918) );
  AOI21_X1 U23907 ( .B1(n20920), .B2(n20919), .A(n20918), .ZN(n20921) );
  OAI211_X1 U23908 ( .C1(n20923), .C2(n14137), .A(n20922), .B(n20921), .ZN(
        P1_U2837) );
  OAI22_X1 U23909 ( .A1(n20926), .A2(n15079), .B1(n20925), .B2(n20924), .ZN(
        n20927) );
  INV_X1 U23910 ( .A(n20927), .ZN(n20928) );
  OAI21_X1 U23911 ( .B1(n20936), .B2(n20929), .A(n20928), .ZN(P1_U2863) );
  AOI22_X1 U23912 ( .A1(n20933), .A2(n20932), .B1(n20931), .B2(n20930), .ZN(
        n20934) );
  OAI21_X1 U23913 ( .B1(n20936), .B2(n20935), .A(n20934), .ZN(P1_U2867) );
  AOI22_X1 U23914 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20940), .B1(n20966), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20937) );
  OAI21_X1 U23915 ( .B1(n20939), .B2(n20938), .A(n20937), .ZN(P1_U2921) );
  INV_X1 U23916 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U23917 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20941) );
  OAI21_X1 U23918 ( .B1(n20942), .B2(n20969), .A(n20941), .ZN(P1_U2922) );
  INV_X1 U23919 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20944) );
  AOI22_X1 U23920 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20943) );
  OAI21_X1 U23921 ( .B1(n20944), .B2(n20969), .A(n20943), .ZN(P1_U2923) );
  AOI22_X1 U23922 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20945) );
  OAI21_X1 U23923 ( .B1(n21643), .B2(n20969), .A(n20945), .ZN(P1_U2924) );
  INV_X1 U23924 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20947) );
  AOI22_X1 U23925 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20946) );
  OAI21_X1 U23926 ( .B1(n20947), .B2(n20969), .A(n20946), .ZN(P1_U2925) );
  INV_X1 U23927 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20949) );
  AOI22_X1 U23928 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20948) );
  OAI21_X1 U23929 ( .B1(n20949), .B2(n20969), .A(n20948), .ZN(P1_U2926) );
  INV_X1 U23930 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U23931 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20950) );
  OAI21_X1 U23932 ( .B1(n20951), .B2(n20969), .A(n20950), .ZN(P1_U2927) );
  AOI22_X1 U23933 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20952) );
  OAI21_X1 U23934 ( .B1(n20953), .B2(n20969), .A(n20952), .ZN(P1_U2928) );
  AOI22_X1 U23935 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20954) );
  OAI21_X1 U23936 ( .B1(n12881), .B2(n20969), .A(n20954), .ZN(P1_U2929) );
  AOI22_X1 U23937 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20955) );
  OAI21_X1 U23938 ( .B1(n12876), .B2(n20969), .A(n20955), .ZN(P1_U2930) );
  AOI22_X1 U23939 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20956) );
  OAI21_X1 U23940 ( .B1(n20957), .B2(n20969), .A(n20956), .ZN(P1_U2931) );
  AOI22_X1 U23941 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20958) );
  OAI21_X1 U23942 ( .B1(n20959), .B2(n20969), .A(n20958), .ZN(P1_U2932) );
  AOI22_X1 U23943 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20960) );
  OAI21_X1 U23944 ( .B1(n20961), .B2(n20969), .A(n20960), .ZN(P1_U2933) );
  AOI22_X1 U23945 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20962) );
  OAI21_X1 U23946 ( .B1(n20963), .B2(n20969), .A(n20962), .ZN(P1_U2934) );
  AOI22_X1 U23947 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20964) );
  OAI21_X1 U23948 ( .B1(n20965), .B2(n20969), .A(n20964), .ZN(P1_U2935) );
  AOI22_X1 U23949 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20967), .B1(n20966), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20968) );
  OAI21_X1 U23950 ( .B1(n20970), .B2(n20969), .A(n20968), .ZN(P1_U2936) );
  AOI22_X1 U23951 ( .A1(n20993), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20988), .ZN(n20972) );
  NAND2_X1 U23952 ( .A1(n20980), .A2(n20971), .ZN(n20982) );
  NAND2_X1 U23953 ( .A1(n20972), .A2(n20982), .ZN(P1_U2946) );
  AOI22_X1 U23954 ( .A1(n20993), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20988), .ZN(n20974) );
  NAND2_X1 U23955 ( .A1(n20980), .A2(n20973), .ZN(n20986) );
  NAND2_X1 U23956 ( .A1(n20974), .A2(n20986), .ZN(P1_U2948) );
  AOI22_X1 U23957 ( .A1(n20993), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20988), .ZN(n20976) );
  NAND2_X1 U23958 ( .A1(n20980), .A2(n20975), .ZN(n20989) );
  NAND2_X1 U23959 ( .A1(n20976), .A2(n20989), .ZN(P1_U2949) );
  AOI22_X1 U23960 ( .A1(n20993), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20988), .ZN(n20978) );
  NAND2_X1 U23961 ( .A1(n20980), .A2(n20977), .ZN(n20991) );
  NAND2_X1 U23962 ( .A1(n20978), .A2(n20991), .ZN(P1_U2950) );
  AOI22_X1 U23963 ( .A1(n20993), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20988), .ZN(n20981) );
  NAND2_X1 U23964 ( .A1(n20980), .A2(n20979), .ZN(n20994) );
  NAND2_X1 U23965 ( .A1(n20981), .A2(n20994), .ZN(P1_U2951) );
  AOI22_X1 U23966 ( .A1(n20993), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20988), .ZN(n20983) );
  NAND2_X1 U23967 ( .A1(n20983), .A2(n20982), .ZN(P1_U2961) );
  AOI22_X1 U23968 ( .A1(n20993), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20988), .ZN(n20985) );
  NAND2_X1 U23969 ( .A1(n20985), .A2(n20984), .ZN(P1_U2962) );
  AOI22_X1 U23970 ( .A1(n20993), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20988), .ZN(n20987) );
  NAND2_X1 U23971 ( .A1(n20987), .A2(n20986), .ZN(P1_U2963) );
  AOI22_X1 U23972 ( .A1(n20993), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20988), .ZN(n20990) );
  NAND2_X1 U23973 ( .A1(n20990), .A2(n20989), .ZN(P1_U2964) );
  AOI22_X1 U23974 ( .A1(n20993), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20988), .ZN(n20992) );
  NAND2_X1 U23975 ( .A1(n20992), .A2(n20991), .ZN(P1_U2965) );
  AOI22_X1 U23976 ( .A1(n20993), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20988), .ZN(n20995) );
  NAND2_X1 U23977 ( .A1(n20995), .A2(n20994), .ZN(P1_U2966) );
  INV_X1 U23978 ( .A(n20996), .ZN(n20997) );
  AOI22_X1 U23979 ( .A1(n21000), .A2(n20999), .B1(n20998), .B2(n20997), .ZN(
        n21006) );
  OAI22_X1 U23980 ( .A1(n21003), .A2(n21002), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21001), .ZN(n21004) );
  NAND3_X1 U23981 ( .A1(n21006), .A2(n21005), .A3(n21004), .ZN(P1_U3031) );
  NOR2_X1 U23982 ( .A1(n21008), .A2(n21007), .ZN(P1_U3032) );
  INV_X1 U23983 ( .A(n21257), .ZN(n21081) );
  OR2_X1 U23984 ( .A1(n21294), .A2(n21085), .ZN(n21010) );
  INV_X1 U23985 ( .A(n21010), .ZN(n21032) );
  AOI22_X1 U23986 ( .A1(n21446), .A2(n21378), .B1(n21412), .B2(n21032), .ZN(
        n21016) );
  OAI21_X1 U23987 ( .B1(n21061), .B2(n21446), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21009) );
  NAND2_X1 U23988 ( .A1(n21009), .A2(n21420), .ZN(n21014) );
  NOR2_X1 U23989 ( .A1(n21079), .A2(n21369), .ZN(n21012) );
  OR2_X1 U23990 ( .A1(n21169), .A2(n21168), .ZN(n21112) );
  AOI22_X1 U23991 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21112), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n21010), .ZN(n21011) );
  INV_X1 U23992 ( .A(n21012), .ZN(n21013) );
  AOI22_X1 U23993 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n21034), .B1(
        n21411), .B2(n21033), .ZN(n21015) );
  OAI211_X1 U23994 ( .C1(n21381), .C2(n21058), .A(n21016), .B(n21015), .ZN(
        P1_U3033) );
  AOI22_X1 U23995 ( .A1(n21446), .A2(n21382), .B1(n21426), .B2(n21032), .ZN(
        n21018) );
  AOI22_X1 U23996 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n21034), .B1(
        n21425), .B2(n21033), .ZN(n21017) );
  OAI211_X1 U23997 ( .C1(n21385), .C2(n21058), .A(n21018), .B(n21017), .ZN(
        P1_U3034) );
  AOI22_X1 U23998 ( .A1(n21446), .A2(n21433), .B1(n21432), .B2(n21032), .ZN(
        n21021) );
  AOI22_X1 U23999 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n21034), .B1(
        n21431), .B2(n21033), .ZN(n21020) );
  OAI211_X1 U24000 ( .C1(n21436), .C2(n21058), .A(n21021), .B(n21020), .ZN(
        P1_U3035) );
  AOI22_X1 U24001 ( .A1(n21446), .A2(n21388), .B1(n21438), .B2(n21032), .ZN(
        n21024) );
  AOI22_X1 U24002 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n21034), .B1(
        n21437), .B2(n21033), .ZN(n21023) );
  OAI211_X1 U24003 ( .C1(n21391), .C2(n21058), .A(n21024), .B(n21023), .ZN(
        P1_U3036) );
  AOI22_X1 U24004 ( .A1(n21446), .A2(n21392), .B1(n21444), .B2(n21032), .ZN(
        n21026) );
  AOI22_X1 U24005 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n21034), .B1(
        n21443), .B2(n21033), .ZN(n21025) );
  OAI211_X1 U24006 ( .C1(n21395), .C2(n21058), .A(n21026), .B(n21025), .ZN(
        P1_U3037) );
  AOI22_X1 U24007 ( .A1(n21446), .A2(n21453), .B1(n21452), .B2(n21032), .ZN(
        n21028) );
  AOI22_X1 U24008 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n21034), .B1(
        n21451), .B2(n21033), .ZN(n21027) );
  OAI211_X1 U24009 ( .C1(n21456), .C2(n21058), .A(n21028), .B(n21027), .ZN(
        P1_U3038) );
  AOI22_X1 U24010 ( .A1(n21446), .A2(n21459), .B1(n21458), .B2(n21032), .ZN(
        n21031) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n21034), .B1(
        n21457), .B2(n21033), .ZN(n21030) );
  OAI211_X1 U24012 ( .C1(n21462), .C2(n21058), .A(n21031), .B(n21030), .ZN(
        P1_U3039) );
  AOI22_X1 U24013 ( .A1(n21446), .A2(n21467), .B1(n21466), .B2(n21032), .ZN(
        n21036) );
  AOI22_X1 U24014 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21034), .B1(
        n21464), .B2(n21033), .ZN(n21035) );
  OAI211_X1 U24015 ( .C1(n21473), .C2(n21058), .A(n21036), .B(n21035), .ZN(
        P1_U3040) );
  NOR2_X1 U24016 ( .A1(n21085), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21042) );
  INV_X1 U24017 ( .A(n21042), .ZN(n21039) );
  NOR2_X1 U24018 ( .A1(n21329), .A2(n21039), .ZN(n21060) );
  INV_X1 U24019 ( .A(n21037), .ZN(n21331) );
  AOI21_X1 U24020 ( .B1(n21038), .B2(n21331), .A(n21060), .ZN(n21040) );
  OAI22_X1 U24021 ( .A1(n21040), .A2(n21418), .B1(n21039), .B2(n21578), .ZN(
        n21059) );
  AOI22_X1 U24022 ( .A1(n21412), .A2(n21060), .B1(n21411), .B2(n21059), .ZN(
        n21044) );
  OAI21_X1 U24023 ( .B1(n21082), .B2(n21201), .A(n21040), .ZN(n21041) );
  OAI221_X1 U24024 ( .B1(n21420), .B2(n21042), .C1(n21418), .C2(n21041), .A(
        n21416), .ZN(n21062) );
  AOI22_X1 U24025 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21378), .ZN(n21043) );
  OAI211_X1 U24026 ( .C1(n21381), .C2(n21074), .A(n21044), .B(n21043), .ZN(
        P1_U3041) );
  AOI22_X1 U24027 ( .A1(n21426), .A2(n21060), .B1(n21425), .B2(n21059), .ZN(
        n21046) );
  AOI22_X1 U24028 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21382), .ZN(n21045) );
  OAI211_X1 U24029 ( .C1(n21385), .C2(n21074), .A(n21046), .B(n21045), .ZN(
        P1_U3042) );
  AOI22_X1 U24030 ( .A1(n21432), .A2(n21060), .B1(n21431), .B2(n21059), .ZN(
        n21048) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21433), .ZN(n21047) );
  OAI211_X1 U24032 ( .C1(n21436), .C2(n21074), .A(n21048), .B(n21047), .ZN(
        P1_U3043) );
  AOI22_X1 U24033 ( .A1(n21438), .A2(n21060), .B1(n21437), .B2(n21059), .ZN(
        n21050) );
  INV_X1 U24034 ( .A(n21391), .ZN(n21439) );
  AOI22_X1 U24035 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n21062), .B1(
        n21055), .B2(n21439), .ZN(n21049) );
  OAI211_X1 U24036 ( .C1(n21442), .C2(n21058), .A(n21050), .B(n21049), .ZN(
        P1_U3044) );
  AOI22_X1 U24037 ( .A1(n21444), .A2(n21060), .B1(n21443), .B2(n21059), .ZN(
        n21052) );
  AOI22_X1 U24038 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21392), .ZN(n21051) );
  OAI211_X1 U24039 ( .C1(n21395), .C2(n21074), .A(n21052), .B(n21051), .ZN(
        P1_U3045) );
  AOI22_X1 U24040 ( .A1(n21452), .A2(n21060), .B1(n21451), .B2(n21059), .ZN(
        n21054) );
  AOI22_X1 U24041 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21453), .ZN(n21053) );
  OAI211_X1 U24042 ( .C1(n21456), .C2(n21074), .A(n21054), .B(n21053), .ZN(
        P1_U3046) );
  AOI22_X1 U24043 ( .A1(n21458), .A2(n21060), .B1(n21457), .B2(n21059), .ZN(
        n21057) );
  INV_X1 U24044 ( .A(n21462), .ZN(n21356) );
  AOI22_X1 U24045 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n21062), .B1(
        n21055), .B2(n21356), .ZN(n21056) );
  OAI211_X1 U24046 ( .C1(n21359), .C2(n21058), .A(n21057), .B(n21056), .ZN(
        P1_U3047) );
  AOI22_X1 U24047 ( .A1(n21466), .A2(n21060), .B1(n21464), .B2(n21059), .ZN(
        n21064) );
  AOI22_X1 U24048 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n21062), .B1(
        n21061), .B2(n21467), .ZN(n21063) );
  OAI211_X1 U24049 ( .C1(n21473), .C2(n21074), .A(n21064), .B(n21063), .ZN(
        P1_U3048) );
  INV_X1 U24050 ( .A(n21436), .ZN(n21344) );
  AOI22_X1 U24051 ( .A1(n21104), .A2(n21344), .B1(n21432), .B2(n21069), .ZN(
        n21066) );
  AOI22_X1 U24052 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21071), .B1(
        n21431), .B2(n21070), .ZN(n21065) );
  OAI211_X1 U24053 ( .C1(n21347), .C2(n21074), .A(n21066), .B(n21065), .ZN(
        P1_U3051) );
  AOI22_X1 U24054 ( .A1(n21104), .A2(n21439), .B1(n21438), .B2(n21069), .ZN(
        n21068) );
  AOI22_X1 U24055 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21071), .B1(
        n21437), .B2(n21070), .ZN(n21067) );
  OAI211_X1 U24056 ( .C1(n21442), .C2(n21074), .A(n21068), .B(n21067), .ZN(
        P1_U3052) );
  AOI22_X1 U24057 ( .A1(n21104), .A2(n21356), .B1(n21458), .B2(n21069), .ZN(
        n21073) );
  AOI22_X1 U24058 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21071), .B1(
        n21457), .B2(n21070), .ZN(n21072) );
  OAI211_X1 U24059 ( .C1(n21359), .C2(n21074), .A(n21073), .B(n21072), .ZN(
        P1_U3055) );
  NOR2_X1 U24060 ( .A1(n21409), .A2(n21085), .ZN(n21080) );
  AOI21_X1 U24061 ( .B1(n21076), .B2(n21075), .A(n21418), .ZN(n21084) );
  INV_X1 U24062 ( .A(n21085), .ZN(n21077) );
  NAND2_X1 U24063 ( .A1(n21078), .A2(n21077), .ZN(n21083) );
  OAI21_X1 U24064 ( .B1(n21079), .B2(n21260), .A(n21083), .ZN(n21087) );
  INV_X1 U24065 ( .A(n21083), .ZN(n21103) );
  AOI22_X1 U24066 ( .A1(n21132), .A2(n21421), .B1(n21412), .B2(n21103), .ZN(
        n21090) );
  INV_X1 U24067 ( .A(n21084), .ZN(n21088) );
  OAI21_X1 U24068 ( .B1(n21409), .B2(n21085), .A(n21418), .ZN(n21086) );
  AOI22_X1 U24069 ( .A1(n21105), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n21104), .B2(n21378), .ZN(n21089) );
  OAI211_X1 U24070 ( .C1(n21108), .C2(n21303), .A(n21090), .B(n21089), .ZN(
        P1_U3057) );
  AOI22_X1 U24071 ( .A1(n21132), .A2(n21427), .B1(n21426), .B2(n21103), .ZN(
        n21092) );
  AOI22_X1 U24072 ( .A1(n21105), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n21104), .B2(n21382), .ZN(n21091) );
  OAI211_X1 U24073 ( .C1(n21108), .C2(n21306), .A(n21092), .B(n21091), .ZN(
        P1_U3058) );
  AOI22_X1 U24074 ( .A1(n21104), .A2(n21433), .B1(n21103), .B2(n21432), .ZN(
        n21094) );
  AOI22_X1 U24075 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n21105), .B1(
        n21132), .B2(n21344), .ZN(n21093) );
  OAI211_X1 U24076 ( .C1(n21108), .C2(n21309), .A(n21094), .B(n21093), .ZN(
        P1_U3059) );
  AOI22_X1 U24077 ( .A1(n21104), .A2(n21388), .B1(n21103), .B2(n21438), .ZN(
        n21096) );
  AOI22_X1 U24078 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n21105), .B1(
        n21132), .B2(n21439), .ZN(n21095) );
  OAI211_X1 U24079 ( .C1(n21108), .C2(n21312), .A(n21096), .B(n21095), .ZN(
        P1_U3060) );
  AOI22_X1 U24080 ( .A1(n21104), .A2(n21392), .B1(n21103), .B2(n21444), .ZN(
        n21098) );
  AOI22_X1 U24081 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n21105), .B1(
        n21132), .B2(n21445), .ZN(n21097) );
  OAI211_X1 U24082 ( .C1(n21108), .C2(n21315), .A(n21098), .B(n21097), .ZN(
        P1_U3061) );
  AOI22_X1 U24083 ( .A1(n21132), .A2(n21352), .B1(n21452), .B2(n21103), .ZN(
        n21100) );
  AOI22_X1 U24084 ( .A1(n21105), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n21104), .B2(n21453), .ZN(n21099) );
  OAI211_X1 U24085 ( .C1(n21108), .C2(n21318), .A(n21100), .B(n21099), .ZN(
        P1_U3062) );
  AOI22_X1 U24086 ( .A1(n21104), .A2(n21459), .B1(n21103), .B2(n21458), .ZN(
        n21102) );
  AOI22_X1 U24087 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n21105), .B1(
        n21132), .B2(n21356), .ZN(n21101) );
  OAI211_X1 U24088 ( .C1(n21108), .C2(n21321), .A(n21102), .B(n21101), .ZN(
        P1_U3063) );
  AOI22_X1 U24089 ( .A1(n21132), .A2(n21362), .B1(n21466), .B2(n21103), .ZN(
        n21107) );
  AOI22_X1 U24090 ( .A1(n21105), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n21104), .B2(n21467), .ZN(n21106) );
  OAI211_X1 U24091 ( .C1(n21108), .C2(n21327), .A(n21107), .B(n21106), .ZN(
        P1_U3064) );
  INV_X1 U24092 ( .A(n21293), .ZN(n21372) );
  NAND3_X1 U24093 ( .A1(n21137), .A2(n21420), .A3(n14378), .ZN(n21111) );
  OAI21_X1 U24094 ( .B1(n21112), .B2(n21372), .A(n21111), .ZN(n21131) );
  AOI22_X1 U24095 ( .A1(n21412), .A2(n9906), .B1(n21411), .B2(n21131), .ZN(
        n21118) );
  AOI21_X1 U24096 ( .B1(n21113), .B2(n21164), .A(n21173), .ZN(n21114) );
  AOI21_X1 U24097 ( .B1(n21137), .B2(n14378), .A(n21114), .ZN(n21115) );
  NOR2_X1 U24098 ( .A1(n21115), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21116) );
  AOI22_X1 U24099 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21378), .ZN(n21117) );
  OAI211_X1 U24100 ( .C1(n21381), .C2(n21164), .A(n21118), .B(n21117), .ZN(
        P1_U3065) );
  AOI22_X1 U24101 ( .A1(n21426), .A2(n9906), .B1(n21425), .B2(n21131), .ZN(
        n21120) );
  AOI22_X1 U24102 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21382), .ZN(n21119) );
  OAI211_X1 U24103 ( .C1(n21385), .C2(n21164), .A(n21120), .B(n21119), .ZN(
        P1_U3066) );
  AOI22_X1 U24104 ( .A1(n21432), .A2(n9906), .B1(n21431), .B2(n21131), .ZN(
        n21122) );
  AOI22_X1 U24105 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21433), .ZN(n21121) );
  OAI211_X1 U24106 ( .C1(n21436), .C2(n21164), .A(n21122), .B(n21121), .ZN(
        P1_U3067) );
  AOI22_X1 U24107 ( .A1(n21438), .A2(n9906), .B1(n21437), .B2(n21131), .ZN(
        n21124) );
  AOI22_X1 U24108 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21388), .ZN(n21123) );
  OAI211_X1 U24109 ( .C1(n21391), .C2(n21164), .A(n21124), .B(n21123), .ZN(
        P1_U3068) );
  AOI22_X1 U24110 ( .A1(n21444), .A2(n9906), .B1(n21443), .B2(n21131), .ZN(
        n21126) );
  AOI22_X1 U24111 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21392), .ZN(n21125) );
  OAI211_X1 U24112 ( .C1(n21395), .C2(n21164), .A(n21126), .B(n21125), .ZN(
        P1_U3069) );
  AOI22_X1 U24113 ( .A1(n21452), .A2(n9906), .B1(n21451), .B2(n21131), .ZN(
        n21128) );
  AOI22_X1 U24114 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21453), .ZN(n21127) );
  OAI211_X1 U24115 ( .C1(n21456), .C2(n21164), .A(n21128), .B(n21127), .ZN(
        P1_U3070) );
  AOI22_X1 U24116 ( .A1(n21458), .A2(n9906), .B1(n21457), .B2(n21131), .ZN(
        n21130) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21459), .ZN(n21129) );
  OAI211_X1 U24118 ( .C1(n21462), .C2(n21164), .A(n21130), .B(n21129), .ZN(
        P1_U3071) );
  AOI22_X1 U24119 ( .A1(n21466), .A2(n9906), .B1(n21464), .B2(n21131), .ZN(
        n21135) );
  AOI22_X1 U24120 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n21133), .B1(
        n21132), .B2(n21467), .ZN(n21134) );
  OAI211_X1 U24121 ( .C1(n21473), .C2(n21164), .A(n21135), .B(n21134), .ZN(
        P1_U3072) );
  NOR2_X1 U24122 ( .A1(n21136), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21143) );
  INV_X1 U24123 ( .A(n21143), .ZN(n21138) );
  NOR2_X1 U24124 ( .A1(n21329), .A2(n21138), .ZN(n21159) );
  AOI21_X1 U24125 ( .B1(n21137), .B2(n21331), .A(n21159), .ZN(n21140) );
  OAI22_X1 U24126 ( .A1(n21140), .A2(n21418), .B1(n21138), .B2(n21578), .ZN(
        n21158) );
  AOI22_X1 U24127 ( .A1(n21412), .A2(n21159), .B1(n21411), .B2(n21158), .ZN(
        n21145) );
  INV_X1 U24128 ( .A(n21139), .ZN(n21141) );
  OAI21_X1 U24129 ( .B1(n21141), .B2(n21201), .A(n21140), .ZN(n21142) );
  OAI221_X1 U24130 ( .B1(n21420), .B2(n21143), .C1(n21418), .C2(n21142), .A(
        n21416), .ZN(n21161) );
  AOI22_X1 U24131 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21421), .ZN(n21144) );
  OAI211_X1 U24132 ( .C1(n21424), .C2(n21164), .A(n21145), .B(n21144), .ZN(
        P1_U3073) );
  AOI22_X1 U24133 ( .A1(n21426), .A2(n21159), .B1(n21425), .B2(n21158), .ZN(
        n21147) );
  AOI22_X1 U24134 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21427), .ZN(n21146) );
  OAI211_X1 U24135 ( .C1(n21430), .C2(n21164), .A(n21147), .B(n21146), .ZN(
        P1_U3074) );
  AOI22_X1 U24136 ( .A1(n21432), .A2(n21159), .B1(n21431), .B2(n21158), .ZN(
        n21149) );
  AOI22_X1 U24137 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21344), .ZN(n21148) );
  OAI211_X1 U24138 ( .C1(n21347), .C2(n21164), .A(n21149), .B(n21148), .ZN(
        P1_U3075) );
  AOI22_X1 U24139 ( .A1(n21438), .A2(n21159), .B1(n21437), .B2(n21158), .ZN(
        n21151) );
  AOI22_X1 U24140 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21439), .ZN(n21150) );
  OAI211_X1 U24141 ( .C1(n21442), .C2(n21164), .A(n21151), .B(n21150), .ZN(
        P1_U3076) );
  AOI22_X1 U24142 ( .A1(n21444), .A2(n21159), .B1(n21443), .B2(n21158), .ZN(
        n21153) );
  AOI22_X1 U24143 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21445), .ZN(n21152) );
  OAI211_X1 U24144 ( .C1(n21450), .C2(n21164), .A(n21153), .B(n21152), .ZN(
        P1_U3077) );
  AOI22_X1 U24145 ( .A1(n21452), .A2(n21159), .B1(n21451), .B2(n21158), .ZN(
        n21155) );
  AOI22_X1 U24146 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21352), .ZN(n21154) );
  OAI211_X1 U24147 ( .C1(n21355), .C2(n21164), .A(n21155), .B(n21154), .ZN(
        P1_U3078) );
  AOI22_X1 U24148 ( .A1(n21458), .A2(n21159), .B1(n21457), .B2(n21158), .ZN(
        n21157) );
  AOI22_X1 U24149 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21356), .ZN(n21156) );
  OAI211_X1 U24150 ( .C1(n21359), .C2(n21164), .A(n21157), .B(n21156), .ZN(
        P1_U3079) );
  AOI22_X1 U24151 ( .A1(n21466), .A2(n21159), .B1(n21464), .B2(n21158), .ZN(
        n21163) );
  AOI22_X1 U24152 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21161), .B1(
        n21160), .B2(n21362), .ZN(n21162) );
  OAI211_X1 U24153 ( .C1(n21367), .C2(n21164), .A(n21163), .B(n21162), .ZN(
        P1_U3080) );
  NAND2_X1 U24154 ( .A1(n21166), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21259) );
  OR2_X1 U24155 ( .A1(n21294), .A2(n21259), .ZN(n21174) );
  INV_X1 U24156 ( .A(n21174), .ZN(n21194) );
  NAND2_X1 U24157 ( .A1(n21167), .A2(n21291), .ZN(n21227) );
  OAI21_X1 U24158 ( .B1(n21227), .B2(n21369), .A(n21174), .ZN(n21176) );
  INV_X1 U24159 ( .A(n21176), .ZN(n21172) );
  INV_X1 U24160 ( .A(n21168), .ZN(n21170) );
  NOR2_X1 U24161 ( .A1(n21170), .A2(n21169), .ZN(n21292) );
  INV_X1 U24162 ( .A(n21292), .ZN(n21296) );
  OAI22_X1 U24163 ( .A1(n21172), .A2(n21418), .B1(n21171), .B2(n21296), .ZN(
        n21193) );
  AOI22_X1 U24164 ( .A1(n21412), .A2(n21194), .B1(n21411), .B2(n21193), .ZN(
        n21180) );
  AOI21_X1 U24165 ( .B1(n21223), .B2(n21178), .A(n21173), .ZN(n21177) );
  NAND2_X1 U24166 ( .A1(n21174), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21175) );
  AOI22_X1 U24167 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n21195), .B2(n21378), .ZN(n21179) );
  OAI211_X1 U24168 ( .C1(n21381), .C2(n21223), .A(n21180), .B(n21179), .ZN(
        P1_U3097) );
  AOI22_X1 U24169 ( .A1(n21426), .A2(n21194), .B1(n21425), .B2(n21193), .ZN(
        n21182) );
  AOI22_X1 U24170 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n21195), .B2(n21382), .ZN(n21181) );
  OAI211_X1 U24171 ( .C1(n21385), .C2(n21223), .A(n21182), .B(n21181), .ZN(
        P1_U3098) );
  AOI22_X1 U24172 ( .A1(n21432), .A2(n21194), .B1(n21431), .B2(n21193), .ZN(
        n21184) );
  AOI22_X1 U24173 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n21195), .B2(n21433), .ZN(n21183) );
  OAI211_X1 U24174 ( .C1(n21436), .C2(n21223), .A(n21184), .B(n21183), .ZN(
        P1_U3099) );
  AOI22_X1 U24175 ( .A1(n21438), .A2(n21194), .B1(n21437), .B2(n21193), .ZN(
        n21186) );
  AOI22_X1 U24176 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n21195), .B2(n21388), .ZN(n21185) );
  OAI211_X1 U24177 ( .C1(n21391), .C2(n21223), .A(n21186), .B(n21185), .ZN(
        P1_U3100) );
  AOI22_X1 U24178 ( .A1(n21444), .A2(n21194), .B1(n21443), .B2(n21193), .ZN(
        n21188) );
  AOI22_X1 U24179 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n21195), .B2(n21392), .ZN(n21187) );
  OAI211_X1 U24180 ( .C1(n21395), .C2(n21223), .A(n21188), .B(n21187), .ZN(
        P1_U3101) );
  AOI22_X1 U24181 ( .A1(n21452), .A2(n21194), .B1(n21451), .B2(n21193), .ZN(
        n21190) );
  AOI22_X1 U24182 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n21195), .B2(n21453), .ZN(n21189) );
  OAI211_X1 U24183 ( .C1(n21456), .C2(n21223), .A(n21190), .B(n21189), .ZN(
        P1_U3102) );
  AOI22_X1 U24184 ( .A1(n21458), .A2(n21194), .B1(n21457), .B2(n21193), .ZN(
        n21192) );
  AOI22_X1 U24185 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n21195), .B2(n21459), .ZN(n21191) );
  OAI211_X1 U24186 ( .C1(n21462), .C2(n21223), .A(n21192), .B(n21191), .ZN(
        P1_U3103) );
  AOI22_X1 U24187 ( .A1(n21466), .A2(n21194), .B1(n21464), .B2(n21193), .ZN(
        n21198) );
  AOI22_X1 U24188 ( .A1(n21196), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n21195), .B2(n21467), .ZN(n21197) );
  OAI211_X1 U24189 ( .C1(n21473), .C2(n21223), .A(n21198), .B(n21197), .ZN(
        P1_U3104) );
  NOR2_X1 U24190 ( .A1(n21259), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21203) );
  INV_X1 U24191 ( .A(n21203), .ZN(n21199) );
  NOR2_X1 U24192 ( .A1(n21329), .A2(n21199), .ZN(n21219) );
  INV_X1 U24193 ( .A(n21227), .ZN(n21261) );
  AOI21_X1 U24194 ( .B1(n21261), .B2(n21331), .A(n21219), .ZN(n21200) );
  OAI22_X1 U24195 ( .A1(n21200), .A2(n21418), .B1(n21199), .B2(n21578), .ZN(
        n21218) );
  AOI22_X1 U24196 ( .A1(n21412), .A2(n21219), .B1(n21411), .B2(n21218), .ZN(
        n21205) );
  OAI21_X1 U24197 ( .B1(n21264), .B2(n21201), .A(n21200), .ZN(n21202) );
  OAI221_X1 U24198 ( .B1(n21420), .B2(n21203), .C1(n21418), .C2(n21202), .A(
        n21416), .ZN(n21220) );
  AOI22_X1 U24199 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21421), .ZN(n21204) );
  OAI211_X1 U24200 ( .C1(n21424), .C2(n21223), .A(n21205), .B(n21204), .ZN(
        P1_U3105) );
  AOI22_X1 U24201 ( .A1(n21426), .A2(n21219), .B1(n21425), .B2(n21218), .ZN(
        n21207) );
  AOI22_X1 U24202 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21427), .ZN(n21206) );
  OAI211_X1 U24203 ( .C1(n21430), .C2(n21223), .A(n21207), .B(n21206), .ZN(
        P1_U3106) );
  AOI22_X1 U24204 ( .A1(n21432), .A2(n21219), .B1(n21431), .B2(n21218), .ZN(
        n21209) );
  AOI22_X1 U24205 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21344), .ZN(n21208) );
  OAI211_X1 U24206 ( .C1(n21347), .C2(n21223), .A(n21209), .B(n21208), .ZN(
        P1_U3107) );
  AOI22_X1 U24207 ( .A1(n21438), .A2(n21219), .B1(n21437), .B2(n21218), .ZN(
        n21211) );
  AOI22_X1 U24208 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21439), .ZN(n21210) );
  OAI211_X1 U24209 ( .C1(n21442), .C2(n21223), .A(n21211), .B(n21210), .ZN(
        P1_U3108) );
  AOI22_X1 U24210 ( .A1(n21444), .A2(n21219), .B1(n21443), .B2(n21218), .ZN(
        n21213) );
  AOI22_X1 U24211 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21445), .ZN(n21212) );
  OAI211_X1 U24212 ( .C1(n21450), .C2(n21223), .A(n21213), .B(n21212), .ZN(
        P1_U3109) );
  AOI22_X1 U24213 ( .A1(n21452), .A2(n21219), .B1(n21451), .B2(n21218), .ZN(
        n21215) );
  AOI22_X1 U24214 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21352), .ZN(n21214) );
  OAI211_X1 U24215 ( .C1(n21355), .C2(n21223), .A(n21215), .B(n21214), .ZN(
        P1_U3110) );
  AOI22_X1 U24216 ( .A1(n21458), .A2(n21219), .B1(n21457), .B2(n21218), .ZN(
        n21217) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21356), .ZN(n21216) );
  OAI211_X1 U24218 ( .C1(n21359), .C2(n21223), .A(n21217), .B(n21216), .ZN(
        P1_U3111) );
  AOI22_X1 U24219 ( .A1(n21466), .A2(n21219), .B1(n21464), .B2(n21218), .ZN(
        n21222) );
  AOI22_X1 U24220 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21220), .B1(
        n21252), .B2(n21362), .ZN(n21221) );
  OAI211_X1 U24221 ( .C1(n21367), .C2(n21223), .A(n21222), .B(n21221), .ZN(
        P1_U3112) );
  INV_X1 U24222 ( .A(n21252), .ZN(n21224) );
  NAND2_X1 U24223 ( .A1(n21224), .A2(n21420), .ZN(n21226) );
  OAI21_X1 U24224 ( .B1(n21226), .B2(n21283), .A(n21288), .ZN(n21232) );
  NOR2_X1 U24225 ( .A1(n21227), .A2(n14378), .ZN(n21229) );
  NOR2_X1 U24226 ( .A1(n21233), .A2(n21234), .ZN(n21370) );
  NOR2_X1 U24227 ( .A1(n21409), .A2(n21259), .ZN(n21266) );
  INV_X1 U24228 ( .A(n21266), .ZN(n21262) );
  NOR2_X1 U24229 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21262), .ZN(
        n21251) );
  AOI22_X1 U24230 ( .A1(n21283), .A2(n21421), .B1(n21412), .B2(n21251), .ZN(
        n21238) );
  INV_X1 U24231 ( .A(n21229), .ZN(n21231) );
  INV_X1 U24232 ( .A(n21251), .ZN(n21230) );
  AOI22_X1 U24233 ( .A1(n21232), .A2(n21231), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21230), .ZN(n21235) );
  OAI21_X1 U24234 ( .B1(n21234), .B2(n21233), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21375) );
  NAND3_X1 U24235 ( .A1(n21236), .A2(n21235), .A3(n21375), .ZN(n21253) );
  AOI22_X1 U24236 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21378), .ZN(n21237) );
  OAI211_X1 U24237 ( .C1(n21256), .C2(n21303), .A(n21238), .B(n21237), .ZN(
        P1_U3113) );
  AOI22_X1 U24238 ( .A1(n21283), .A2(n21427), .B1(n21426), .B2(n21251), .ZN(
        n21240) );
  AOI22_X1 U24239 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21382), .ZN(n21239) );
  OAI211_X1 U24240 ( .C1(n21256), .C2(n21306), .A(n21240), .B(n21239), .ZN(
        P1_U3114) );
  AOI22_X1 U24241 ( .A1(n21283), .A2(n21344), .B1(n21432), .B2(n21251), .ZN(
        n21242) );
  AOI22_X1 U24242 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21433), .ZN(n21241) );
  OAI211_X1 U24243 ( .C1(n21256), .C2(n21309), .A(n21242), .B(n21241), .ZN(
        P1_U3115) );
  AOI22_X1 U24244 ( .A1(n21283), .A2(n21439), .B1(n21438), .B2(n21251), .ZN(
        n21244) );
  AOI22_X1 U24245 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21388), .ZN(n21243) );
  OAI211_X1 U24246 ( .C1(n21256), .C2(n21312), .A(n21244), .B(n21243), .ZN(
        P1_U3116) );
  AOI22_X1 U24247 ( .A1(n21283), .A2(n21445), .B1(n21444), .B2(n21251), .ZN(
        n21246) );
  AOI22_X1 U24248 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21392), .ZN(n21245) );
  OAI211_X1 U24249 ( .C1(n21256), .C2(n21315), .A(n21246), .B(n21245), .ZN(
        P1_U3117) );
  AOI22_X1 U24250 ( .A1(n21283), .A2(n21352), .B1(n21452), .B2(n21251), .ZN(
        n21248) );
  AOI22_X1 U24251 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21453), .ZN(n21247) );
  OAI211_X1 U24252 ( .C1(n21256), .C2(n21318), .A(n21248), .B(n21247), .ZN(
        P1_U3118) );
  AOI22_X1 U24253 ( .A1(n21252), .A2(n21459), .B1(n21251), .B2(n21458), .ZN(
        n21250) );
  AOI22_X1 U24254 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21253), .B1(
        n21283), .B2(n21356), .ZN(n21249) );
  OAI211_X1 U24255 ( .C1(n21256), .C2(n21321), .A(n21250), .B(n21249), .ZN(
        P1_U3119) );
  AOI22_X1 U24256 ( .A1(n21283), .A2(n21362), .B1(n21466), .B2(n21251), .ZN(
        n21255) );
  AOI22_X1 U24257 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21253), .B1(
        n21252), .B2(n21467), .ZN(n21254) );
  OAI211_X1 U24258 ( .C1(n21256), .C2(n21327), .A(n21255), .B(n21254), .ZN(
        P1_U3120) );
  NOR2_X1 U24259 ( .A1(n21405), .A2(n21259), .ZN(n21282) );
  INV_X1 U24260 ( .A(n21260), .ZN(n21406) );
  AOI21_X1 U24261 ( .B1(n21261), .B2(n21406), .A(n21282), .ZN(n21263) );
  OAI22_X1 U24262 ( .A1(n21263), .A2(n21418), .B1(n21262), .B2(n21578), .ZN(
        n21281) );
  AOI22_X1 U24263 ( .A1(n21412), .A2(n21282), .B1(n21411), .B2(n21281), .ZN(
        n21268) );
  OAI21_X1 U24264 ( .B1(n21264), .B2(n21414), .A(n21263), .ZN(n21265) );
  OAI221_X1 U24265 ( .B1(n21420), .B2(n21266), .C1(n21418), .C2(n21265), .A(
        n21416), .ZN(n21284) );
  AOI22_X1 U24266 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21378), .ZN(n21267) );
  OAI211_X1 U24267 ( .C1(n21381), .C2(n21300), .A(n21268), .B(n21267), .ZN(
        P1_U3121) );
  AOI22_X1 U24268 ( .A1(n21426), .A2(n21282), .B1(n21425), .B2(n21281), .ZN(
        n21270) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21382), .ZN(n21269) );
  OAI211_X1 U24270 ( .C1(n21385), .C2(n21300), .A(n21270), .B(n21269), .ZN(
        P1_U3122) );
  AOI22_X1 U24271 ( .A1(n21432), .A2(n21282), .B1(n21431), .B2(n21281), .ZN(
        n21272) );
  AOI22_X1 U24272 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21433), .ZN(n21271) );
  OAI211_X1 U24273 ( .C1(n21436), .C2(n21300), .A(n21272), .B(n21271), .ZN(
        P1_U3123) );
  AOI22_X1 U24274 ( .A1(n21438), .A2(n21282), .B1(n21437), .B2(n21281), .ZN(
        n21274) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21388), .ZN(n21273) );
  OAI211_X1 U24276 ( .C1(n21391), .C2(n21300), .A(n21274), .B(n21273), .ZN(
        P1_U3124) );
  AOI22_X1 U24277 ( .A1(n21444), .A2(n21282), .B1(n21443), .B2(n21281), .ZN(
        n21276) );
  AOI22_X1 U24278 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21392), .ZN(n21275) );
  OAI211_X1 U24279 ( .C1(n21395), .C2(n21300), .A(n21276), .B(n21275), .ZN(
        P1_U3125) );
  AOI22_X1 U24280 ( .A1(n21452), .A2(n21282), .B1(n21451), .B2(n21281), .ZN(
        n21278) );
  AOI22_X1 U24281 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21453), .ZN(n21277) );
  OAI211_X1 U24282 ( .C1(n21456), .C2(n21300), .A(n21278), .B(n21277), .ZN(
        P1_U3126) );
  AOI22_X1 U24283 ( .A1(n21458), .A2(n21282), .B1(n21457), .B2(n21281), .ZN(
        n21280) );
  AOI22_X1 U24284 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21459), .ZN(n21279) );
  OAI211_X1 U24285 ( .C1(n21462), .C2(n21300), .A(n21280), .B(n21279), .ZN(
        P1_U3127) );
  AOI22_X1 U24286 ( .A1(n21466), .A2(n21282), .B1(n21464), .B2(n21281), .ZN(
        n21286) );
  AOI22_X1 U24287 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21284), .B1(
        n21283), .B2(n21467), .ZN(n21285) );
  OAI211_X1 U24288 ( .C1(n21473), .C2(n21300), .A(n21286), .B(n21285), .ZN(
        P1_U3128) );
  OR2_X1 U24289 ( .A1(n21415), .A2(n14113), .ZN(n21335) );
  NAND3_X1 U24290 ( .A1(n21300), .A2(n21420), .A3(n21366), .ZN(n21289) );
  NAND2_X1 U24291 ( .A1(n21289), .A2(n21288), .ZN(n21298) );
  NOR2_X1 U24292 ( .A1(n21330), .A2(n21369), .ZN(n21295) );
  NAND2_X1 U24293 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21408) );
  AOI22_X1 U24294 ( .A1(n21322), .A2(n21421), .B1(n21412), .B2(n9907), .ZN(
        n21302) );
  INV_X1 U24295 ( .A(n21295), .ZN(n21297) );
  AOI22_X1 U24296 ( .A1(n21298), .A2(n21297), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21296), .ZN(n21299) );
  AOI22_X1 U24297 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21378), .ZN(n21301) );
  OAI211_X1 U24298 ( .C1(n21328), .C2(n21303), .A(n21302), .B(n21301), .ZN(
        P1_U3129) );
  AOI22_X1 U24299 ( .A1(n21322), .A2(n21427), .B1(n21426), .B2(n9907), .ZN(
        n21305) );
  AOI22_X1 U24300 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21382), .ZN(n21304) );
  OAI211_X1 U24301 ( .C1(n21328), .C2(n21306), .A(n21305), .B(n21304), .ZN(
        P1_U3130) );
  AOI22_X1 U24302 ( .A1(n21322), .A2(n21344), .B1(n21432), .B2(n9907), .ZN(
        n21308) );
  AOI22_X1 U24303 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21433), .ZN(n21307) );
  OAI211_X1 U24304 ( .C1(n21328), .C2(n21309), .A(n21308), .B(n21307), .ZN(
        P1_U3131) );
  AOI22_X1 U24305 ( .A1(n21322), .A2(n21439), .B1(n21438), .B2(n9907), .ZN(
        n21311) );
  AOI22_X1 U24306 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21388), .ZN(n21310) );
  OAI211_X1 U24307 ( .C1(n21328), .C2(n21312), .A(n21311), .B(n21310), .ZN(
        P1_U3132) );
  AOI22_X1 U24308 ( .A1(n21322), .A2(n21445), .B1(n21444), .B2(n9907), .ZN(
        n21314) );
  AOI22_X1 U24309 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21392), .ZN(n21313) );
  OAI211_X1 U24310 ( .C1(n21328), .C2(n21315), .A(n21314), .B(n21313), .ZN(
        P1_U3133) );
  AOI22_X1 U24311 ( .A1(n21322), .A2(n21352), .B1(n21452), .B2(n9907), .ZN(
        n21317) );
  AOI22_X1 U24312 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21453), .ZN(n21316) );
  OAI211_X1 U24313 ( .C1(n21328), .C2(n21318), .A(n21317), .B(n21316), .ZN(
        P1_U3134) );
  AOI22_X1 U24314 ( .A1(n21322), .A2(n21356), .B1(n21458), .B2(n9907), .ZN(
        n21320) );
  AOI22_X1 U24315 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21459), .ZN(n21319) );
  OAI211_X1 U24316 ( .C1(n21328), .C2(n21321), .A(n21320), .B(n21319), .ZN(
        P1_U3135) );
  AOI22_X1 U24317 ( .A1(n21322), .A2(n21362), .B1(n21466), .B2(n9907), .ZN(
        n21326) );
  AOI22_X1 U24318 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21324), .B1(
        n21323), .B2(n21467), .ZN(n21325) );
  OAI211_X1 U24319 ( .C1(n21328), .C2(n21327), .A(n21326), .B(n21325), .ZN(
        P1_U3136) );
  NOR3_X2 U24320 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21329), .A3(
        n21408), .ZN(n21361) );
  AOI21_X1 U24321 ( .B1(n21407), .B2(n21331), .A(n21361), .ZN(n21333) );
  NOR2_X1 U24322 ( .A1(n21408), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n21337) );
  INV_X1 U24323 ( .A(n21337), .ZN(n21332) );
  OAI22_X1 U24324 ( .A1(n21333), .A2(n21418), .B1(n21332), .B2(n21578), .ZN(
        n21360) );
  AOI22_X1 U24325 ( .A1(n21412), .A2(n21361), .B1(n21411), .B2(n21360), .ZN(
        n21341) );
  INV_X1 U24326 ( .A(n21334), .ZN(n21336) );
  NOR2_X1 U24327 ( .A1(n21336), .A2(n21335), .ZN(n21338) );
  AOI22_X1 U24328 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21421), .ZN(n21340) );
  OAI211_X1 U24329 ( .C1(n21424), .C2(n21366), .A(n21341), .B(n21340), .ZN(
        P1_U3137) );
  AOI22_X1 U24330 ( .A1(n21426), .A2(n21361), .B1(n21425), .B2(n21360), .ZN(
        n21343) );
  AOI22_X1 U24331 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21427), .ZN(n21342) );
  OAI211_X1 U24332 ( .C1(n21430), .C2(n21366), .A(n21343), .B(n21342), .ZN(
        P1_U3138) );
  AOI22_X1 U24333 ( .A1(n21432), .A2(n21361), .B1(n21431), .B2(n21360), .ZN(
        n21346) );
  AOI22_X1 U24334 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21344), .ZN(n21345) );
  OAI211_X1 U24335 ( .C1(n21347), .C2(n21366), .A(n21346), .B(n21345), .ZN(
        P1_U3139) );
  AOI22_X1 U24336 ( .A1(n21438), .A2(n21361), .B1(n21437), .B2(n21360), .ZN(
        n21349) );
  AOI22_X1 U24337 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21439), .ZN(n21348) );
  OAI211_X1 U24338 ( .C1(n21442), .C2(n21366), .A(n21349), .B(n21348), .ZN(
        P1_U3140) );
  AOI22_X1 U24339 ( .A1(n21444), .A2(n21361), .B1(n21443), .B2(n21360), .ZN(
        n21351) );
  AOI22_X1 U24340 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21445), .ZN(n21350) );
  OAI211_X1 U24341 ( .C1(n21450), .C2(n21366), .A(n21351), .B(n21350), .ZN(
        P1_U3141) );
  AOI22_X1 U24342 ( .A1(n21452), .A2(n21361), .B1(n21451), .B2(n21360), .ZN(
        n21354) );
  AOI22_X1 U24343 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21352), .ZN(n21353) );
  OAI211_X1 U24344 ( .C1(n21355), .C2(n21366), .A(n21354), .B(n21353), .ZN(
        P1_U3142) );
  AOI22_X1 U24345 ( .A1(n21458), .A2(n21361), .B1(n21457), .B2(n21360), .ZN(
        n21358) );
  AOI22_X1 U24346 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21356), .ZN(n21357) );
  OAI211_X1 U24347 ( .C1(n21359), .C2(n21366), .A(n21358), .B(n21357), .ZN(
        P1_U3143) );
  AOI22_X1 U24348 ( .A1(n21466), .A2(n21361), .B1(n21464), .B2(n21360), .ZN(
        n21365) );
  AOI22_X1 U24349 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21363), .B1(
        n10743), .B2(n21362), .ZN(n21364) );
  OAI211_X1 U24350 ( .C1(n21367), .C2(n21366), .A(n21365), .B(n21364), .ZN(
        P1_U3144) );
  NOR3_X2 U24351 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21409), .A3(
        n21408), .ZN(n21401) );
  NAND2_X1 U24352 ( .A1(n21407), .A2(n21369), .ZN(n21373) );
  INV_X1 U24353 ( .A(n21370), .ZN(n21371) );
  OAI22_X1 U24354 ( .A1(n21373), .A2(n21418), .B1(n21372), .B2(n21371), .ZN(
        n21400) );
  AOI22_X1 U24355 ( .A1(n21412), .A2(n21401), .B1(n21411), .B2(n21400), .ZN(
        n21380) );
  OAI21_X1 U24356 ( .B1(n21468), .B2(n10743), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21374) );
  AOI21_X1 U24357 ( .B1(n21374), .B2(n21373), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21377) );
  AOI22_X1 U24358 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21378), .ZN(n21379) );
  OAI211_X1 U24359 ( .C1(n21381), .C2(n21449), .A(n21380), .B(n21379), .ZN(
        P1_U3145) );
  AOI22_X1 U24360 ( .A1(n21426), .A2(n21401), .B1(n21425), .B2(n21400), .ZN(
        n21384) );
  AOI22_X1 U24361 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21382), .ZN(n21383) );
  OAI211_X1 U24362 ( .C1(n21385), .C2(n21449), .A(n21384), .B(n21383), .ZN(
        P1_U3146) );
  AOI22_X1 U24363 ( .A1(n21432), .A2(n21401), .B1(n21431), .B2(n21400), .ZN(
        n21387) );
  AOI22_X1 U24364 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21433), .ZN(n21386) );
  OAI211_X1 U24365 ( .C1(n21436), .C2(n21449), .A(n21387), .B(n21386), .ZN(
        P1_U3147) );
  AOI22_X1 U24366 ( .A1(n21438), .A2(n21401), .B1(n21437), .B2(n21400), .ZN(
        n21390) );
  AOI22_X1 U24367 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21388), .ZN(n21389) );
  OAI211_X1 U24368 ( .C1(n21391), .C2(n21449), .A(n21390), .B(n21389), .ZN(
        P1_U3148) );
  AOI22_X1 U24369 ( .A1(n21444), .A2(n21401), .B1(n21443), .B2(n21400), .ZN(
        n21394) );
  AOI22_X1 U24370 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21392), .ZN(n21393) );
  OAI211_X1 U24371 ( .C1(n21395), .C2(n21449), .A(n21394), .B(n21393), .ZN(
        P1_U3149) );
  AOI22_X1 U24372 ( .A1(n21452), .A2(n21401), .B1(n21451), .B2(n21400), .ZN(
        n21397) );
  AOI22_X1 U24373 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21453), .ZN(n21396) );
  OAI211_X1 U24374 ( .C1(n21456), .C2(n21449), .A(n21397), .B(n21396), .ZN(
        P1_U3150) );
  AOI22_X1 U24375 ( .A1(n21458), .A2(n21401), .B1(n21457), .B2(n21400), .ZN(
        n21399) );
  AOI22_X1 U24376 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21459), .ZN(n21398) );
  OAI211_X1 U24377 ( .C1(n21462), .C2(n21449), .A(n21399), .B(n21398), .ZN(
        P1_U3151) );
  AOI22_X1 U24378 ( .A1(n21466), .A2(n21401), .B1(n21464), .B2(n21400), .ZN(
        n21404) );
  AOI22_X1 U24379 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21402), .B1(
        n10743), .B2(n21467), .ZN(n21403) );
  OAI211_X1 U24380 ( .C1(n21473), .C2(n21449), .A(n21404), .B(n21403), .ZN(
        P1_U3152) );
  NOR2_X1 U24381 ( .A1(n21405), .A2(n21408), .ZN(n21465) );
  AOI21_X1 U24382 ( .B1(n21407), .B2(n21406), .A(n21465), .ZN(n21413) );
  NOR2_X1 U24383 ( .A1(n21409), .A2(n21408), .ZN(n21419) );
  INV_X1 U24384 ( .A(n21419), .ZN(n21410) );
  OAI22_X1 U24385 ( .A1(n21413), .A2(n21418), .B1(n21410), .B2(n21578), .ZN(
        n21463) );
  AOI22_X1 U24386 ( .A1(n21412), .A2(n21465), .B1(n21411), .B2(n21463), .ZN(
        n21423) );
  OAI21_X1 U24387 ( .B1(n21415), .B2(n21414), .A(n21413), .ZN(n21417) );
  OAI221_X1 U24388 ( .B1(n21420), .B2(n21419), .C1(n21418), .C2(n21417), .A(
        n21416), .ZN(n21469) );
  AOI22_X1 U24389 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21469), .B1(
        n21446), .B2(n21421), .ZN(n21422) );
  OAI211_X1 U24390 ( .C1(n21424), .C2(n21449), .A(n21423), .B(n21422), .ZN(
        P1_U3153) );
  AOI22_X1 U24391 ( .A1(n21426), .A2(n21465), .B1(n21425), .B2(n21463), .ZN(
        n21429) );
  AOI22_X1 U24392 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21469), .B1(
        n21446), .B2(n21427), .ZN(n21428) );
  OAI211_X1 U24393 ( .C1(n21430), .C2(n21449), .A(n21429), .B(n21428), .ZN(
        P1_U3154) );
  AOI22_X1 U24394 ( .A1(n21432), .A2(n21465), .B1(n21431), .B2(n21463), .ZN(
        n21435) );
  AOI22_X1 U24395 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21469), .B1(
        n21468), .B2(n21433), .ZN(n21434) );
  OAI211_X1 U24396 ( .C1(n21436), .C2(n21472), .A(n21435), .B(n21434), .ZN(
        P1_U3155) );
  AOI22_X1 U24397 ( .A1(n21438), .A2(n21465), .B1(n21437), .B2(n21463), .ZN(
        n21441) );
  AOI22_X1 U24398 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21469), .B1(
        n21446), .B2(n21439), .ZN(n21440) );
  OAI211_X1 U24399 ( .C1(n21442), .C2(n21449), .A(n21441), .B(n21440), .ZN(
        P1_U3156) );
  AOI22_X1 U24400 ( .A1(n21444), .A2(n21465), .B1(n21443), .B2(n21463), .ZN(
        n21448) );
  AOI22_X1 U24401 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21469), .B1(
        n21446), .B2(n21445), .ZN(n21447) );
  OAI211_X1 U24402 ( .C1(n21450), .C2(n21449), .A(n21448), .B(n21447), .ZN(
        P1_U3157) );
  AOI22_X1 U24403 ( .A1(n21452), .A2(n21465), .B1(n21451), .B2(n21463), .ZN(
        n21455) );
  AOI22_X1 U24404 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21469), .B1(
        n21468), .B2(n21453), .ZN(n21454) );
  OAI211_X1 U24405 ( .C1(n21456), .C2(n21472), .A(n21455), .B(n21454), .ZN(
        P1_U3158) );
  AOI22_X1 U24406 ( .A1(n21458), .A2(n21465), .B1(n21457), .B2(n21463), .ZN(
        n21461) );
  AOI22_X1 U24407 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21469), .B1(
        n21468), .B2(n21459), .ZN(n21460) );
  OAI211_X1 U24408 ( .C1(n21462), .C2(n21472), .A(n21461), .B(n21460), .ZN(
        P1_U3159) );
  AOI22_X1 U24409 ( .A1(n21466), .A2(n21465), .B1(n21464), .B2(n21463), .ZN(
        n21471) );
  AOI22_X1 U24410 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21469), .B1(
        n21468), .B2(n21467), .ZN(n21470) );
  OAI211_X1 U24411 ( .C1(n21473), .C2(n21472), .A(n21471), .B(n21470), .ZN(
        P1_U3160) );
  AOI21_X1 U24412 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20825), .A(n21474), 
        .ZN(n21476) );
  NAND2_X1 U24413 ( .A1(n21476), .A2(n21475), .ZN(P1_U3163) );
  AND2_X1 U24414 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21477), .ZN(
        P1_U3164) );
  AND2_X1 U24415 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21477), .ZN(
        P1_U3165) );
  AND2_X1 U24416 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21477), .ZN(
        P1_U3166) );
  AND2_X1 U24417 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21477), .ZN(
        P1_U3167) );
  AND2_X1 U24418 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21477), .ZN(
        P1_U3168) );
  AND2_X1 U24419 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21477), .ZN(
        P1_U3169) );
  AND2_X1 U24420 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21477), .ZN(
        P1_U3170) );
  AND2_X1 U24421 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21477), .ZN(
        P1_U3171) );
  AND2_X1 U24422 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21477), .ZN(
        P1_U3172) );
  AND2_X1 U24423 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21477), .ZN(
        P1_U3173) );
  AND2_X1 U24424 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21477), .ZN(
        P1_U3174) );
  AND2_X1 U24425 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21477), .ZN(
        P1_U3175) );
  AND2_X1 U24426 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21477), .ZN(
        P1_U3176) );
  AND2_X1 U24427 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21477), .ZN(
        P1_U3177) );
  AND2_X1 U24428 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21477), .ZN(
        P1_U3178) );
  AND2_X1 U24429 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21477), .ZN(
        P1_U3179) );
  AND2_X1 U24430 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21477), .ZN(
        P1_U3180) );
  AND2_X1 U24431 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21477), .ZN(
        P1_U3181) );
  AND2_X1 U24432 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21477), .ZN(
        P1_U3182) );
  AND2_X1 U24433 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21477), .ZN(
        P1_U3183) );
  AND2_X1 U24434 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21477), .ZN(
        P1_U3184) );
  AND2_X1 U24435 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21477), .ZN(
        P1_U3185) );
  AND2_X1 U24436 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21477), .ZN(P1_U3186) );
  AND2_X1 U24437 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21477), .ZN(P1_U3187) );
  AND2_X1 U24438 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21477), .ZN(P1_U3188) );
  AND2_X1 U24439 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21477), .ZN(P1_U3189) );
  AND2_X1 U24440 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21477), .ZN(P1_U3190) );
  AND2_X1 U24441 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21477), .ZN(P1_U3191) );
  AND2_X1 U24442 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21477), .ZN(P1_U3192) );
  AND2_X1 U24443 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21477), .ZN(P1_U3193) );
  AOI21_X1 U24444 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21478), .A(n21486), 
        .ZN(n21493) );
  NOR2_X1 U24445 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21480) );
  NAND2_X1 U24446 ( .A1(n21486), .A2(NA), .ZN(n21479) );
  OAI211_X1 U24447 ( .C1(n21491), .C2(n21480), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .B(n21479), .ZN(n21481) );
  INV_X1 U24448 ( .A(n21481), .ZN(n21482) );
  OAI22_X1 U24449 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21493), .B1(n21583), 
        .B2(n21482), .ZN(P1_U3194) );
  INV_X1 U24450 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21487) );
  NOR3_X1 U24451 ( .A1(NA), .A2(n21487), .A3(n21486), .ZN(n21484) );
  OAI22_X1 U24452 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21485), .B1(
        P1_STATE_REG_2__SCAN_IN), .B2(n21484), .ZN(n21492) );
  NOR3_X1 U24453 ( .A1(NA), .A2(n21486), .A3(n21574), .ZN(n21488) );
  OAI22_X1 U24454 ( .A1(n21489), .A2(n21488), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n21487), .ZN(n21490) );
  OAI22_X1 U24455 ( .A1(n21493), .A2(n21492), .B1(n21491), .B2(n21490), .ZN(
        P1_U3196) );
  NAND2_X1 U24456 ( .A1(n21583), .A2(n21494), .ZN(n21539) );
  INV_X1 U24457 ( .A(n21539), .ZN(n21530) );
  INV_X1 U24458 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n21496) );
  INV_X2 U24459 ( .A(n21533), .ZN(n21551) );
  OAI222_X1 U24460 ( .A1(n21547), .A2(n21498), .B1(n21496), .B2(n21583), .C1(
        n21495), .C2(n21551), .ZN(P1_U3197) );
  INV_X1 U24461 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n21497) );
  OAI222_X1 U24462 ( .A1(n21551), .A2(n21498), .B1(n21497), .B2(n21583), .C1(
        n14137), .C2(n21539), .ZN(P1_U3198) );
  OAI222_X1 U24463 ( .A1(n21551), .A2(n14137), .B1(n21499), .B2(n21583), .C1(
        n21500), .C2(n21539), .ZN(P1_U3199) );
  INV_X1 U24464 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21501) );
  OAI222_X1 U24465 ( .A1(n21539), .A2(n21503), .B1(n21501), .B2(n21583), .C1(
        n21500), .C2(n21551), .ZN(P1_U3200) );
  INV_X1 U24466 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21502) );
  OAI222_X1 U24467 ( .A1(n21551), .A2(n21503), .B1(n21502), .B2(n21583), .C1(
        n21792), .C2(n21539), .ZN(P1_U3201) );
  INV_X1 U24468 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21504) );
  OAI222_X1 U24469 ( .A1(n21551), .A2(n21792), .B1(n21504), .B2(n21583), .C1(
        n21506), .C2(n21539), .ZN(P1_U3202) );
  INV_X1 U24470 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21505) );
  OAI222_X1 U24471 ( .A1(n21551), .A2(n21506), .B1(n21505), .B2(n21583), .C1(
        n21507), .C2(n21539), .ZN(P1_U3203) );
  INV_X1 U24472 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21802) );
  OAI222_X1 U24473 ( .A1(n21539), .A2(n21509), .B1(n21802), .B2(n21583), .C1(
        n21507), .C2(n21551), .ZN(P1_U3204) );
  INV_X1 U24474 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n21508) );
  OAI222_X1 U24475 ( .A1(n21551), .A2(n21509), .B1(n21508), .B2(n21583), .C1(
        n21511), .C2(n21539), .ZN(P1_U3205) );
  INV_X1 U24476 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n21510) );
  OAI222_X1 U24477 ( .A1(n21551), .A2(n21511), .B1(n21510), .B2(n21583), .C1(
        n21513), .C2(n21539), .ZN(P1_U3206) );
  AOI22_X1 U24478 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21530), .ZN(n21512) );
  OAI21_X1 U24479 ( .B1(n21513), .B2(n21551), .A(n21512), .ZN(P1_U3207) );
  AOI22_X1 U24480 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n21533), .ZN(n21514) );
  OAI21_X1 U24481 ( .B1(n21516), .B2(n21547), .A(n21514), .ZN(P1_U3208) );
  INV_X1 U24482 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n21515) );
  OAI222_X1 U24483 ( .A1(n21551), .A2(n21516), .B1(n21515), .B2(n21583), .C1(
        n21518), .C2(n21539), .ZN(P1_U3209) );
  INV_X1 U24484 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n21517) );
  OAI222_X1 U24485 ( .A1(n21551), .A2(n21518), .B1(n21517), .B2(n21583), .C1(
        n21520), .C2(n21547), .ZN(P1_U3210) );
  INV_X1 U24486 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n21519) );
  INV_X1 U24487 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21522) );
  OAI222_X1 U24488 ( .A1(n21551), .A2(n21520), .B1(n21519), .B2(n21583), .C1(
        n21522), .C2(n21539), .ZN(P1_U3211) );
  INV_X1 U24489 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n21521) );
  OAI222_X1 U24490 ( .A1(n21551), .A2(n21522), .B1(n21521), .B2(n21583), .C1(
        n21523), .C2(n21547), .ZN(P1_U3212) );
  INV_X1 U24491 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n21524) );
  OAI222_X1 U24492 ( .A1(n21539), .A2(n21526), .B1(n21524), .B2(n21583), .C1(
        n21523), .C2(n21551), .ZN(P1_U3213) );
  INV_X1 U24493 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n21525) );
  OAI222_X1 U24494 ( .A1(n21551), .A2(n21526), .B1(n21525), .B2(n21583), .C1(
        n21771), .C2(n21547), .ZN(P1_U3214) );
  AOI22_X1 U24495 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21530), .ZN(n21527) );
  OAI21_X1 U24496 ( .B1(n21771), .B2(n21551), .A(n21527), .ZN(P1_U3215) );
  AOI22_X1 U24497 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n21533), .ZN(n21528) );
  OAI21_X1 U24498 ( .B1(n14858), .B2(n21547), .A(n21528), .ZN(P1_U3216) );
  INV_X1 U24499 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21529) );
  OAI222_X1 U24500 ( .A1(n21551), .A2(n14858), .B1(n21529), .B2(n21583), .C1(
        n21532), .C2(n21547), .ZN(P1_U3217) );
  AOI22_X1 U24501 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21530), .ZN(n21531) );
  OAI21_X1 U24502 ( .B1(n21532), .B2(n21551), .A(n21531), .ZN(P1_U3218) );
  AOI22_X1 U24503 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21570), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21533), .ZN(n21534) );
  OAI21_X1 U24504 ( .B1(n21536), .B2(n21547), .A(n21534), .ZN(P1_U3219) );
  INV_X1 U24505 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21535) );
  OAI222_X1 U24506 ( .A1(n21551), .A2(n21536), .B1(n21535), .B2(n21583), .C1(
        n21537), .C2(n21547), .ZN(P1_U3220) );
  INV_X1 U24507 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21538) );
  OAI222_X1 U24508 ( .A1(n21539), .A2(n21541), .B1(n21538), .B2(n21583), .C1(
        n21537), .C2(n21551), .ZN(P1_U3221) );
  INV_X1 U24509 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21540) );
  OAI222_X1 U24510 ( .A1(n21551), .A2(n21541), .B1(n21540), .B2(n21583), .C1(
        n21542), .C2(n21547), .ZN(P1_U3222) );
  INV_X1 U24511 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21848) );
  INV_X1 U24512 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21543) );
  OAI222_X1 U24513 ( .A1(n21547), .A2(n21848), .B1(n21543), .B2(n21583), .C1(
        n21542), .C2(n21551), .ZN(P1_U3223) );
  INV_X1 U24514 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21544) );
  OAI222_X1 U24515 ( .A1(n21551), .A2(n21848), .B1(n21544), .B2(n21583), .C1(
        n21546), .C2(n21547), .ZN(P1_U3224) );
  INV_X1 U24516 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n21545) );
  OAI222_X1 U24517 ( .A1(n21551), .A2(n21546), .B1(n21545), .B2(n21583), .C1(
        n21550), .C2(n21547), .ZN(P1_U3225) );
  INV_X1 U24518 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n21549) );
  OAI222_X1 U24519 ( .A1(n21551), .A2(n21550), .B1(n21549), .B2(n21583), .C1(
        n21548), .C2(n21547), .ZN(P1_U3226) );
  INV_X1 U24520 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21682) );
  AOI22_X1 U24521 ( .A1(n21583), .A2(n21552), .B1(n21682), .B2(n21570), .ZN(
        P1_U3458) );
  INV_X1 U24522 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21564) );
  INV_X1 U24523 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21553) );
  AOI22_X1 U24524 ( .A1(n21583), .A2(n21564), .B1(n21553), .B2(n21570), .ZN(
        P1_U3459) );
  INV_X1 U24525 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21554) );
  AOI22_X1 U24526 ( .A1(n21583), .A2(n21555), .B1(n21554), .B2(n21570), .ZN(
        P1_U3460) );
  INV_X1 U24527 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21567) );
  INV_X1 U24528 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21556) );
  AOI22_X1 U24529 ( .A1(n21583), .A2(n21567), .B1(n21556), .B2(n21570), .ZN(
        P1_U3461) );
  OAI21_X1 U24530 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n21560), .A(n21558), 
        .ZN(n21557) );
  INV_X1 U24531 ( .A(n21557), .ZN(P1_U3464) );
  INV_X1 U24532 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21559) );
  OAI21_X1 U24533 ( .B1(n21560), .B2(n21559), .A(n21558), .ZN(P1_U3465) );
  INV_X1 U24534 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21562) );
  NOR3_X1 U24535 ( .A1(n21562), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n21561) );
  AOI221_X1 U24536 ( .B1(n21563), .B2(n21562), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n21561), .ZN(n21565) );
  INV_X1 U24537 ( .A(n21569), .ZN(n21566) );
  AOI22_X1 U24538 ( .A1(n21569), .A2(n21565), .B1(n21564), .B2(n21566), .ZN(
        P1_U3481) );
  NOR2_X1 U24539 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21568) );
  AOI22_X1 U24540 ( .A1(n21569), .A2(n21568), .B1(n21567), .B2(n21566), .ZN(
        P1_U3482) );
  AOI22_X1 U24541 ( .A1(n21583), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21571), 
        .B2(n21570), .ZN(P1_U3483) );
  AOI211_X1 U24542 ( .C1(n20967), .C2(n21574), .A(n21573), .B(n21572), .ZN(
        n21582) );
  INV_X1 U24543 ( .A(n21575), .ZN(n21577) );
  NAND3_X1 U24544 ( .A1(n21577), .A2(n21576), .A3(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21579) );
  AOI22_X1 U24545 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21579), .B1(n21578), 
        .B2(n13446), .ZN(n21581) );
  NAND2_X1 U24546 ( .A1(n21582), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n21580) );
  OAI21_X1 U24547 ( .B1(n21582), .B2(n21581), .A(n21580), .ZN(P1_U3485) );
  MUX2_X1 U24548 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21583), .Z(P1_U3486) );
  OAI222_X1 U24549 ( .A1(n21589), .A2(n21588), .B1(n21587), .B2(n21586), .C1(
        n21585), .C2(n21584), .ZN(n21899) );
  INV_X1 U24550 ( .A(keyinput17), .ZN(n21897) );
  NOR4_X1 U24551 ( .A1(P3_DATAO_REG_30__SCAN_IN), .A2(n16103), .A3(n16095), 
        .A4(n21867), .ZN(n21600) );
  INV_X1 U24552 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n21861) );
  NOR4_X1 U24553 ( .A1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        BUF1_REG_26__SCAN_IN), .A3(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(
        n21861), .ZN(n21599) );
  NAND4_X1 U24554 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P1_DATAO_REG_12__SCAN_IN), .A4(P3_ADDRESS_REG_19__SCAN_IN), .ZN(
        n21594) );
  INV_X1 U24555 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n21591) );
  NOR4_X1 U24556 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n21874), .A3(n21873), .A4(
        n21882), .ZN(n21590) );
  NAND4_X1 U24557 ( .A1(n21591), .A2(n15295), .A3(n21590), .A4(
        P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n21593) );
  NAND4_X1 U24558 ( .A1(n21835), .A2(P2_EBX_REG_29__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .A4(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n21592) );
  NOR4_X1 U24559 ( .A1(n21594), .A2(n21593), .A3(n21592), .A4(
        P3_UWORD_REG_7__SCAN_IN), .ZN(n21598) );
  NOR3_X1 U24560 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(P3_DATAO_REG_27__SCAN_IN), .A3(n14128), .ZN(n21595) );
  AND4_X1 U24561 ( .A1(n21596), .A2(n21595), .A3(n21847), .A4(n21848), .ZN(
        n21597) );
  AND4_X1 U24562 ( .A1(n21600), .A2(n21599), .A3(n21598), .A4(n21597), .ZN(
        n21635) );
  INV_X1 U24563 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21789) );
  NOR4_X1 U24564 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(BS16), .A3(
        n21768), .A4(n21771), .ZN(n21601) );
  NAND3_X1 U24565 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n21601), .A3(n21778), 
        .ZN(n21610) );
  NAND4_X1 U24566 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_DATAO_REG_23__SCAN_IN), .A4(n21816), .ZN(n21602) );
  NOR3_X1 U24567 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(
        P3_D_C_N_REG_SCAN_IN), .A3(n21602), .ZN(n21608) );
  NAND4_X1 U24568 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(n21792), .A4(n21784), .ZN(n21606) );
  NAND4_X1 U24569 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_4__7__SCAN_IN), .A3(BUF1_REG_15__SCAN_IN), .A4(
        P2_DATAO_REG_31__SCAN_IN), .ZN(n21605) );
  NAND4_X1 U24570 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .A3(P2_REIP_REG_4__SCAN_IN), .A4(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n21604) );
  NAND4_X1 U24571 ( .A1(P1_EBX_REG_15__SCAN_IN), .A2(P1_ADDRESS_REG_7__SCAN_IN), .A3(P3_REIP_REG_15__SCAN_IN), .A4(P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n21603)
         );
  NOR4_X1 U24572 ( .A1(n21606), .A2(n21605), .A3(n21604), .A4(n21603), .ZN(
        n21607) );
  NAND4_X1 U24573 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n21608), .A3(n21607), 
        .A4(n21821), .ZN(n21609) );
  NOR4_X1 U24574 ( .A1(P2_ADDRESS_REG_4__SCAN_IN), .A2(n21789), .A3(n21610), 
        .A4(n21609), .ZN(n21634) );
  NOR4_X1 U24575 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(
        BUF2_REG_22__SCAN_IN), .A3(P1_UWORD_REG_11__SCAN_IN), .A4(n21646), 
        .ZN(n21611) );
  NAND3_X1 U24576 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(
        P1_REIP_REG_0__SCAN_IN), .A3(n21611), .ZN(n21621) );
  NAND4_X1 U24577 ( .A1(P1_EAX_REG_12__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A3(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A4(n21641), .ZN(n21612) );
  NOR3_X1 U24578 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(n21638), .A3(n21612), 
        .ZN(n21619) );
  NAND4_X1 U24579 ( .A1(P2_BYTEENABLE_REG_2__SCAN_IN), .A2(n21671), .A3(n21674), .A4(n21670), .ZN(n21617) );
  NAND4_X1 U24580 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A4(n21668), .ZN(n21616) );
  NAND4_X1 U24581 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(
        P3_EAX_REG_15__SCAN_IN), .A3(P3_DATAO_REG_22__SCAN_IN), .A4(
        P1_BE_N_REG_3__SCAN_IN), .ZN(n21615) );
  INV_X1 U24582 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n21613) );
  NAND4_X1 U24583 ( .A1(n21613), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_11__4__SCAN_IN), .A4(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n21614) );
  NOR4_X1 U24584 ( .A1(n21617), .A2(n21616), .A3(n21615), .A4(n21614), .ZN(
        n21618) );
  NAND4_X1 U24585 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_EAX_REG_13__SCAN_IN), .A3(n21619), .A4(n21618), .ZN(n21620) );
  NOR4_X1 U24586 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(
        P3_LWORD_REG_2__SCAN_IN), .A3(n21621), .A4(n21620), .ZN(n21633) );
  NOR4_X1 U24587 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(
        P2_BYTEENABLE_REG_3__SCAN_IN), .A3(n21704), .A4(n21706), .ZN(n21622)
         );
  NAND3_X1 U24588 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_DATAO_REG_5__SCAN_IN), .A3(n21622), .ZN(n21631) );
  NOR4_X1 U24589 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), 
        .A4(n21720), .ZN(n21629) );
  NOR4_X1 U24590 ( .A1(P2_REIP_REG_20__SCAN_IN), .A2(DATAI_20_), .A3(n21701), 
        .A4(n21717), .ZN(n21628) );
  NAND4_X1 U24591 ( .A1(READY21_REG_SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .A3(n21738), .A4(n21733), .ZN(n21626) );
  NAND4_X1 U24592 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(
        P3_DATAO_REG_15__SCAN_IN), .A3(n21725), .A4(n21726), .ZN(n21625) );
  NAND4_X1 U24593 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .A3(P3_INSTQUEUE_REG_8__3__SCAN_IN), 
        .A4(n21751), .ZN(n21624) );
  INV_X1 U24594 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n21742) );
  INV_X1 U24595 ( .A(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n21754) );
  NAND4_X1 U24596 ( .A1(n21742), .A2(n21754), .A3(n21756), .A4(n21753), .ZN(
        n21623) );
  NOR4_X1 U24597 ( .A1(n21626), .A2(n21625), .A3(n21624), .A4(n21623), .ZN(
        n21627) );
  NAND3_X1 U24598 ( .A1(n21629), .A2(n21628), .A3(n21627), .ZN(n21630) );
  NOR4_X1 U24599 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_3__5__SCAN_IN), .A3(n21631), .A4(n21630), .ZN(n21632)
         );
  NAND4_X1 U24600 ( .A1(n21635), .A2(n21634), .A3(n21633), .A4(n21632), .ZN(
        n21896) );
  INV_X1 U24601 ( .A(P3_DATAO_REG_9__SCAN_IN), .ZN(n21637) );
  AOI22_X1 U24602 ( .A1(n21638), .A2(keyinput114), .B1(keyinput102), .B2(
        n21637), .ZN(n21636) );
  OAI221_X1 U24603 ( .B1(n21638), .B2(keyinput114), .C1(n21637), .C2(
        keyinput102), .A(n21636), .ZN(n21651) );
  INV_X1 U24604 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n21640) );
  AOI22_X1 U24605 ( .A1(n21641), .A2(keyinput30), .B1(keyinput117), .B2(n21640), .ZN(n21639) );
  OAI221_X1 U24606 ( .B1(n21641), .B2(keyinput30), .C1(n21640), .C2(
        keyinput117), .A(n21639), .ZN(n21650) );
  AOI22_X1 U24607 ( .A1(n21644), .A2(keyinput35), .B1(keyinput0), .B2(n21643), 
        .ZN(n21642) );
  OAI221_X1 U24608 ( .B1(n21644), .B2(keyinput35), .C1(n21643), .C2(keyinput0), 
        .A(n21642), .ZN(n21649) );
  INV_X1 U24609 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n21647) );
  AOI22_X1 U24610 ( .A1(n21647), .A2(keyinput92), .B1(keyinput54), .B2(n21646), 
        .ZN(n21645) );
  OAI221_X1 U24611 ( .B1(n21647), .B2(keyinput92), .C1(n21646), .C2(keyinput54), .A(n21645), .ZN(n21648) );
  NOR4_X1 U24612 ( .A1(n21651), .A2(n21650), .A3(n21649), .A4(n21648), .ZN(
        n21699) );
  INV_X1 U24613 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n21653) );
  AOI22_X1 U24614 ( .A1(n21654), .A2(keyinput87), .B1(n21653), .B2(keyinput16), 
        .ZN(n21652) );
  OAI221_X1 U24615 ( .B1(n21654), .B2(keyinput87), .C1(n21653), .C2(keyinput16), .A(n21652), .ZN(n21666) );
  INV_X1 U24616 ( .A(P3_LWORD_REG_2__SCAN_IN), .ZN(n21656) );
  AOI22_X1 U24617 ( .A1(n21657), .A2(keyinput45), .B1(keyinput100), .B2(n21656), .ZN(n21655) );
  OAI221_X1 U24618 ( .B1(n21657), .B2(keyinput45), .C1(n21656), .C2(
        keyinput100), .A(n21655), .ZN(n21665) );
  INV_X1 U24619 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n21659) );
  AOI22_X1 U24620 ( .A1(n21659), .A2(keyinput108), .B1(n18343), .B2(keyinput26), .ZN(n21658) );
  OAI221_X1 U24621 ( .B1(n21659), .B2(keyinput108), .C1(n18343), .C2(
        keyinput26), .A(n21658), .ZN(n21664) );
  INV_X1 U24622 ( .A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n21662) );
  AOI22_X1 U24623 ( .A1(n21662), .A2(keyinput122), .B1(keyinput78), .B2(n21661), .ZN(n21660) );
  OAI221_X1 U24624 ( .B1(n21662), .B2(keyinput122), .C1(n21661), .C2(
        keyinput78), .A(n21660), .ZN(n21663) );
  NOR4_X1 U24625 ( .A1(n21666), .A2(n21665), .A3(n21664), .A4(n21663), .ZN(
        n21698) );
  AOI22_X1 U24626 ( .A1(n18286), .A2(keyinput55), .B1(keyinput61), .B2(n21668), 
        .ZN(n21667) );
  OAI221_X1 U24627 ( .B1(n18286), .B2(keyinput55), .C1(n21668), .C2(keyinput61), .A(n21667), .ZN(n21680) );
  AOI22_X1 U24628 ( .A1(n21671), .A2(keyinput75), .B1(keyinput119), .B2(n21670), .ZN(n21669) );
  OAI221_X1 U24629 ( .B1(n21671), .B2(keyinput75), .C1(n21670), .C2(
        keyinput119), .A(n21669), .ZN(n21679) );
  AOI22_X1 U24630 ( .A1(n21674), .A2(keyinput2), .B1(keyinput47), .B2(n21673), 
        .ZN(n21672) );
  OAI221_X1 U24631 ( .B1(n21674), .B2(keyinput2), .C1(n21673), .C2(keyinput47), 
        .A(n21672), .ZN(n21678) );
  AOI22_X1 U24632 ( .A1(n18228), .A2(keyinput21), .B1(keyinput53), .B2(n21676), 
        .ZN(n21675) );
  OAI221_X1 U24633 ( .B1(n18228), .B2(keyinput21), .C1(n21676), .C2(keyinput53), .A(n21675), .ZN(n21677) );
  NOR4_X1 U24634 ( .A1(n21680), .A2(n21679), .A3(n21678), .A4(n21677), .ZN(
        n21697) );
  INV_X1 U24635 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n21683) );
  AOI22_X1 U24636 ( .A1(n21683), .A2(keyinput113), .B1(keyinput79), .B2(n21682), .ZN(n21681) );
  OAI221_X1 U24637 ( .B1(n21683), .B2(keyinput113), .C1(n21682), .C2(
        keyinput79), .A(n21681), .ZN(n21695) );
  INV_X1 U24638 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n21686) );
  AOI22_X1 U24639 ( .A1(n21686), .A2(keyinput23), .B1(keyinput65), .B2(n21685), 
        .ZN(n21684) );
  OAI221_X1 U24640 ( .B1(n21686), .B2(keyinput23), .C1(n21685), .C2(keyinput65), .A(n21684), .ZN(n21694) );
  INV_X1 U24641 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n21688) );
  AOI22_X1 U24642 ( .A1(n21689), .A2(keyinput98), .B1(keyinput49), .B2(n21688), 
        .ZN(n21687) );
  OAI221_X1 U24643 ( .B1(n21689), .B2(keyinput98), .C1(n21688), .C2(keyinput49), .A(n21687), .ZN(n21693) );
  XNOR2_X1 U24644 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B(keyinput94), .ZN(
        n21691) );
  XNOR2_X1 U24645 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B(keyinput68), 
        .ZN(n21690) );
  NAND2_X1 U24646 ( .A1(n21691), .A2(n21690), .ZN(n21692) );
  NOR4_X1 U24647 ( .A1(n21695), .A2(n21694), .A3(n21693), .A4(n21692), .ZN(
        n21696) );
  NAND4_X1 U24648 ( .A1(n21699), .A2(n21698), .A3(n21697), .A4(n21696), .ZN(
        n21894) );
  AOI22_X1 U24649 ( .A1(n21701), .A2(keyinput27), .B1(n11996), .B2(keyinput24), 
        .ZN(n21700) );
  OAI221_X1 U24650 ( .B1(n21701), .B2(keyinput27), .C1(n11996), .C2(keyinput24), .A(n21700), .ZN(n21714) );
  INV_X1 U24651 ( .A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n21703) );
  AOI22_X1 U24652 ( .A1(n21704), .A2(keyinput62), .B1(keyinput22), .B2(n21703), 
        .ZN(n21702) );
  OAI221_X1 U24653 ( .B1(n21704), .B2(keyinput62), .C1(n21703), .C2(keyinput22), .A(n21702), .ZN(n21713) );
  AOI22_X1 U24654 ( .A1(n21707), .A2(keyinput110), .B1(n21706), .B2(
        keyinput121), .ZN(n21705) );
  OAI221_X1 U24655 ( .B1(n21707), .B2(keyinput110), .C1(n21706), .C2(
        keyinput121), .A(n21705), .ZN(n21712) );
  INV_X1 U24656 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n21708) );
  XOR2_X1 U24657 ( .A(n21708), .B(keyinput81), .Z(n21710) );
  XNOR2_X1 U24658 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B(keyinput44), .ZN(
        n21709) );
  NAND2_X1 U24659 ( .A1(n21710), .A2(n21709), .ZN(n21711) );
  NOR4_X1 U24660 ( .A1(n21714), .A2(n21713), .A3(n21712), .A4(n21711), .ZN(
        n21766) );
  INV_X1 U24661 ( .A(DATAI_20_), .ZN(n21716) );
  AOI22_X1 U24662 ( .A1(n21717), .A2(keyinput69), .B1(n21716), .B2(keyinput39), 
        .ZN(n21715) );
  OAI221_X1 U24663 ( .B1(n21717), .B2(keyinput69), .C1(n21716), .C2(keyinput39), .A(n21715), .ZN(n21730) );
  AOI22_X1 U24664 ( .A1(n21720), .A2(keyinput59), .B1(keyinput120), .B2(n21719), .ZN(n21718) );
  OAI221_X1 U24665 ( .B1(n21720), .B2(keyinput59), .C1(n21719), .C2(
        keyinput120), .A(n21718), .ZN(n21729) );
  INV_X1 U24666 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n21723) );
  AOI22_X1 U24667 ( .A1(n21723), .A2(keyinput104), .B1(keyinput1), .B2(n21722), 
        .ZN(n21721) );
  OAI221_X1 U24668 ( .B1(n21723), .B2(keyinput104), .C1(n21722), .C2(keyinput1), .A(n21721), .ZN(n21728) );
  AOI22_X1 U24669 ( .A1(n21726), .A2(keyinput57), .B1(n21725), .B2(keyinput6), 
        .ZN(n21724) );
  OAI221_X1 U24670 ( .B1(n21726), .B2(keyinput57), .C1(n21725), .C2(keyinput6), 
        .A(n21724), .ZN(n21727) );
  NOR4_X1 U24671 ( .A1(n21730), .A2(n21729), .A3(n21728), .A4(n21727), .ZN(
        n21765) );
  INV_X1 U24672 ( .A(READY21_REG_SCAN_IN), .ZN(n21732) );
  AOI22_X1 U24673 ( .A1(n21733), .A2(keyinput5), .B1(n21732), .B2(keyinput118), 
        .ZN(n21731) );
  OAI221_X1 U24674 ( .B1(n21733), .B2(keyinput5), .C1(n21732), .C2(keyinput118), .A(n21731), .ZN(n21736) );
  INV_X1 U24675 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n21734) );
  XNOR2_X1 U24676 ( .A(n21734), .B(keyinput127), .ZN(n21735) );
  NOR2_X1 U24677 ( .A1(n21736), .A2(n21735), .ZN(n21748) );
  AOI22_X1 U24678 ( .A1(n21739), .A2(keyinput105), .B1(n21738), .B2(keyinput90), .ZN(n21737) );
  OAI221_X1 U24679 ( .B1(n21739), .B2(keyinput105), .C1(n21738), .C2(
        keyinput90), .A(n21737), .ZN(n21740) );
  INV_X1 U24680 ( .A(n21740), .ZN(n21747) );
  AOI22_X1 U24681 ( .A1(n21743), .A2(keyinput25), .B1(n21742), .B2(keyinput10), 
        .ZN(n21741) );
  OAI221_X1 U24682 ( .B1(n21743), .B2(keyinput25), .C1(n21742), .C2(keyinput10), .A(n21741), .ZN(n21744) );
  INV_X1 U24683 ( .A(n21744), .ZN(n21746) );
  XNOR2_X1 U24684 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B(keyinput9), .ZN(
        n21745) );
  AND4_X1 U24685 ( .A1(n21748), .A2(n21747), .A3(n21746), .A4(n21745), .ZN(
        n21764) );
  INV_X1 U24686 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n21750) );
  AOI22_X1 U24687 ( .A1(n21751), .A2(keyinput88), .B1(keyinput51), .B2(n21750), 
        .ZN(n21749) );
  OAI221_X1 U24688 ( .B1(n21751), .B2(keyinput88), .C1(n21750), .C2(keyinput51), .A(n21749), .ZN(n21762) );
  AOI22_X1 U24689 ( .A1(n21754), .A2(keyinput38), .B1(keyinput31), .B2(n21753), 
        .ZN(n21752) );
  OAI221_X1 U24690 ( .B1(n21754), .B2(keyinput38), .C1(n21753), .C2(keyinput31), .A(n21752), .ZN(n21761) );
  AOI22_X1 U24691 ( .A1(n21756), .A2(keyinput46), .B1(n18378), .B2(keyinput33), 
        .ZN(n21755) );
  OAI221_X1 U24692 ( .B1(n21756), .B2(keyinput46), .C1(n18378), .C2(keyinput33), .A(n21755), .ZN(n21760) );
  XOR2_X1 U24693 ( .A(n16242), .B(keyinput52), .Z(n21758) );
  XNOR2_X1 U24694 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B(keyinput126), .ZN(
        n21757) );
  NAND2_X1 U24695 ( .A1(n21758), .A2(n21757), .ZN(n21759) );
  NOR4_X1 U24696 ( .A1(n21762), .A2(n21761), .A3(n21760), .A4(n21759), .ZN(
        n21763) );
  NAND4_X1 U24697 ( .A1(n21766), .A2(n21765), .A3(n21764), .A4(n21763), .ZN(
        n21893) );
  INV_X1 U24698 ( .A(BS16), .ZN(n21769) );
  AOI22_X1 U24699 ( .A1(n21769), .A2(keyinput67), .B1(n21768), .B2(keyinput101), .ZN(n21767) );
  OAI221_X1 U24700 ( .B1(n21769), .B2(keyinput67), .C1(n21768), .C2(
        keyinput101), .A(n21767), .ZN(n21782) );
  INV_X1 U24701 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21772) );
  AOI22_X1 U24702 ( .A1(n21772), .A2(keyinput73), .B1(keyinput28), .B2(n21771), 
        .ZN(n21770) );
  OAI221_X1 U24703 ( .B1(n21772), .B2(keyinput73), .C1(n21771), .C2(keyinput28), .A(n21770), .ZN(n21781) );
  AOI22_X1 U24704 ( .A1(n21775), .A2(keyinput15), .B1(keyinput14), .B2(n21774), 
        .ZN(n21773) );
  OAI221_X1 U24705 ( .B1(n21775), .B2(keyinput15), .C1(n21774), .C2(keyinput14), .A(n21773), .ZN(n21780) );
  INV_X1 U24706 ( .A(P1_LWORD_REG_1__SCAN_IN), .ZN(n21777) );
  AOI22_X1 U24707 ( .A1(n21778), .A2(keyinput103), .B1(keyinput70), .B2(n21777), .ZN(n21776) );
  OAI221_X1 U24708 ( .B1(n21778), .B2(keyinput103), .C1(n21777), .C2(
        keyinput70), .A(n21776), .ZN(n21779) );
  NOR4_X1 U24709 ( .A1(n21782), .A2(n21781), .A3(n21780), .A4(n21779), .ZN(
        n21830) );
  AOI22_X1 U24710 ( .A1(n21785), .A2(keyinput36), .B1(keyinput42), .B2(n21784), 
        .ZN(n21783) );
  OAI221_X1 U24711 ( .B1(n21785), .B2(keyinput36), .C1(n21784), .C2(keyinput42), .A(n21783), .ZN(n21797) );
  AOI22_X1 U24712 ( .A1(n21787), .A2(keyinput99), .B1(n13448), .B2(keyinput83), 
        .ZN(n21786) );
  OAI221_X1 U24713 ( .B1(n21787), .B2(keyinput99), .C1(n13448), .C2(keyinput83), .A(n21786), .ZN(n21796) );
  AOI22_X1 U24714 ( .A1(n21790), .A2(keyinput74), .B1(n21789), .B2(keyinput32), 
        .ZN(n21788) );
  OAI221_X1 U24715 ( .B1(n21790), .B2(keyinput74), .C1(n21789), .C2(keyinput32), .A(n21788), .ZN(n21795) );
  AOI22_X1 U24716 ( .A1(n21793), .A2(keyinput125), .B1(n21792), .B2(keyinput18), .ZN(n21791) );
  OAI221_X1 U24717 ( .B1(n21793), .B2(keyinput125), .C1(n21792), .C2(
        keyinput18), .A(n21791), .ZN(n21794) );
  NOR4_X1 U24718 ( .A1(n21797), .A2(n21796), .A3(n21795), .A4(n21794), .ZN(
        n21829) );
  INV_X1 U24719 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n21799) );
  AOI22_X1 U24720 ( .A1(n21799), .A2(keyinput34), .B1(keyinput97), .B2(n16465), 
        .ZN(n21798) );
  OAI221_X1 U24721 ( .B1(n21799), .B2(keyinput34), .C1(n16465), .C2(keyinput97), .A(n21798), .ZN(n21811) );
  AOI22_X1 U24722 ( .A1(n21802), .A2(keyinput4), .B1(keyinput7), .B2(n21801), 
        .ZN(n21800) );
  OAI221_X1 U24723 ( .B1(n21802), .B2(keyinput4), .C1(n21801), .C2(keyinput7), 
        .A(n21800), .ZN(n21810) );
  AOI22_X1 U24724 ( .A1(n21805), .A2(keyinput96), .B1(keyinput20), .B2(n21804), 
        .ZN(n21803) );
  OAI221_X1 U24725 ( .B1(n21805), .B2(keyinput96), .C1(n21804), .C2(keyinput20), .A(n21803), .ZN(n21809) );
  AOI22_X1 U24726 ( .A1(n21807), .A2(keyinput64), .B1(n11610), .B2(keyinput84), 
        .ZN(n21806) );
  OAI221_X1 U24727 ( .B1(n21807), .B2(keyinput64), .C1(n11610), .C2(keyinput84), .A(n21806), .ZN(n21808) );
  NOR4_X1 U24728 ( .A1(n21811), .A2(n21810), .A3(n21809), .A4(n21808), .ZN(
        n21828) );
  INV_X1 U24729 ( .A(P3_D_C_N_REG_SCAN_IN), .ZN(n21814) );
  AOI22_X1 U24730 ( .A1(n21814), .A2(keyinput3), .B1(n21813), .B2(keyinput72), 
        .ZN(n21812) );
  OAI221_X1 U24731 ( .B1(n21814), .B2(keyinput3), .C1(n21813), .C2(keyinput72), 
        .A(n21812), .ZN(n21826) );
  AOI22_X1 U24732 ( .A1(n21817), .A2(keyinput37), .B1(keyinput63), .B2(n21816), 
        .ZN(n21815) );
  OAI221_X1 U24733 ( .B1(n21817), .B2(keyinput37), .C1(n21816), .C2(keyinput63), .A(n21815), .ZN(n21825) );
  AOI22_X1 U24734 ( .A1(n15074), .A2(keyinput124), .B1(keyinput111), .B2(
        n21819), .ZN(n21818) );
  OAI221_X1 U24735 ( .B1(n15074), .B2(keyinput124), .C1(n21819), .C2(
        keyinput111), .A(n21818), .ZN(n21824) );
  AOI22_X1 U24736 ( .A1(n21822), .A2(keyinput11), .B1(keyinput93), .B2(n21821), 
        .ZN(n21820) );
  OAI221_X1 U24737 ( .B1(n21822), .B2(keyinput11), .C1(n21821), .C2(keyinput93), .A(n21820), .ZN(n21823) );
  NOR4_X1 U24738 ( .A1(n21826), .A2(n21825), .A3(n21824), .A4(n21823), .ZN(
        n21827) );
  NAND4_X1 U24739 ( .A1(n21830), .A2(n21829), .A3(n21828), .A4(n21827), .ZN(
        n21892) );
  AOI22_X1 U24740 ( .A1(n21833), .A2(keyinput85), .B1(n21832), .B2(keyinput115), .ZN(n21831) );
  OAI221_X1 U24741 ( .B1(n21833), .B2(keyinput85), .C1(n21832), .C2(
        keyinput115), .A(n21831), .ZN(n21842) );
  AOI22_X1 U24742 ( .A1(n21835), .A2(keyinput86), .B1(keyinput82), .B2(n15295), 
        .ZN(n21834) );
  OAI221_X1 U24743 ( .B1(n21835), .B2(keyinput86), .C1(n15295), .C2(keyinput82), .A(n21834), .ZN(n21841) );
  XNOR2_X1 U24744 ( .A(P2_EBX_REG_29__SCAN_IN), .B(keyinput91), .ZN(n21839) );
  XNOR2_X1 U24745 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B(keyinput48), .ZN(
        n21838) );
  XNOR2_X1 U24746 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput76), .ZN(
        n21837) );
  XNOR2_X1 U24747 ( .A(keyinput50), .B(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n21836) );
  NAND4_X1 U24748 ( .A1(n21839), .A2(n21838), .A3(n21837), .A4(n21836), .ZN(
        n21840) );
  NOR3_X1 U24749 ( .A1(n21842), .A2(n21841), .A3(n21840), .ZN(n21890) );
  NAND2_X1 U24750 ( .A1(n21844), .A2(keyinput19), .ZN(n21843) );
  OAI221_X1 U24751 ( .B1(n21845), .B2(keyinput17), .C1(n21844), .C2(keyinput19), .A(n21843), .ZN(n21857) );
  AOI22_X1 U24752 ( .A1(n21848), .A2(keyinput12), .B1(n21847), .B2(keyinput8), 
        .ZN(n21846) );
  OAI221_X1 U24753 ( .B1(n21848), .B2(keyinput12), .C1(n21847), .C2(keyinput8), 
        .A(n21846), .ZN(n21856) );
  AOI22_X1 U24754 ( .A1(n21851), .A2(keyinput107), .B1(keyinput106), .B2(
        n21850), .ZN(n21849) );
  OAI221_X1 U24755 ( .B1(n21851), .B2(keyinput107), .C1(n21850), .C2(
        keyinput106), .A(n21849), .ZN(n21855) );
  AOI22_X1 U24756 ( .A1(n21853), .A2(keyinput40), .B1(n14128), .B2(keyinput123), .ZN(n21852) );
  OAI221_X1 U24757 ( .B1(n21853), .B2(keyinput40), .C1(n14128), .C2(
        keyinput123), .A(n21852), .ZN(n21854) );
  NOR4_X1 U24758 ( .A1(n21857), .A2(n21856), .A3(n21855), .A4(n21854), .ZN(
        n21889) );
  AOI22_X1 U24759 ( .A1(n16103), .A2(keyinput41), .B1(n16095), .B2(keyinput109), .ZN(n21858) );
  OAI221_X1 U24760 ( .B1(n16103), .B2(keyinput41), .C1(n16095), .C2(
        keyinput109), .A(n21858), .ZN(n21871) );
  AOI22_X1 U24761 ( .A1(n21861), .A2(keyinput60), .B1(n21860), .B2(keyinput71), 
        .ZN(n21859) );
  OAI221_X1 U24762 ( .B1(n21861), .B2(keyinput60), .C1(n21860), .C2(keyinput71), .A(n21859), .ZN(n21870) );
  INV_X1 U24763 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n21864) );
  INV_X1 U24764 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n21863) );
  AOI22_X1 U24765 ( .A1(n21864), .A2(keyinput95), .B1(keyinput56), .B2(n21863), 
        .ZN(n21862) );
  OAI221_X1 U24766 ( .B1(n21864), .B2(keyinput95), .C1(n21863), .C2(keyinput56), .A(n21862), .ZN(n21869) );
  AOI22_X1 U24767 ( .A1(n21867), .A2(keyinput66), .B1(keyinput58), .B2(n21866), 
        .ZN(n21865) );
  OAI221_X1 U24768 ( .B1(n21867), .B2(keyinput66), .C1(n21866), .C2(keyinput58), .A(n21865), .ZN(n21868) );
  NOR4_X1 U24769 ( .A1(n21871), .A2(n21870), .A3(n21869), .A4(n21868), .ZN(
        n21888) );
  AOI22_X1 U24770 ( .A1(n21874), .A2(keyinput112), .B1(keyinput89), .B2(n21873), .ZN(n21872) );
  OAI221_X1 U24771 ( .B1(n21874), .B2(keyinput112), .C1(n21873), .C2(
        keyinput89), .A(n21872), .ZN(n21886) );
  INV_X1 U24772 ( .A(P3_UWORD_REG_7__SCAN_IN), .ZN(n21877) );
  AOI22_X1 U24773 ( .A1(n21877), .A2(keyinput13), .B1(n21876), .B2(keyinput80), 
        .ZN(n21875) );
  OAI221_X1 U24774 ( .B1(n21877), .B2(keyinput13), .C1(n21876), .C2(keyinput80), .A(n21875), .ZN(n21885) );
  AOI22_X1 U24775 ( .A1(n16118), .A2(keyinput43), .B1(keyinput29), .B2(n21879), 
        .ZN(n21878) );
  OAI221_X1 U24776 ( .B1(n16118), .B2(keyinput43), .C1(n21879), .C2(keyinput29), .A(n21878), .ZN(n21884) );
  AOI22_X1 U24777 ( .A1(n21882), .A2(keyinput116), .B1(n21881), .B2(keyinput77), .ZN(n21880) );
  OAI221_X1 U24778 ( .B1(n21882), .B2(keyinput116), .C1(n21881), .C2(
        keyinput77), .A(n21880), .ZN(n21883) );
  NOR4_X1 U24779 ( .A1(n21886), .A2(n21885), .A3(n21884), .A4(n21883), .ZN(
        n21887) );
  NAND4_X1 U24780 ( .A1(n21890), .A2(n21889), .A3(n21888), .A4(n21887), .ZN(
        n21891) );
  NOR4_X1 U24781 ( .A1(n21894), .A2(n21893), .A3(n21892), .A4(n21891), .ZN(
        n21895) );
  OAI221_X1 U24782 ( .B1(n21897), .B2(DATAI_8_), .C1(n21897), .C2(n21896), .A(
        n21895), .ZN(n21898) );
  XNOR2_X1 U24783 ( .A(n21899), .B(n21898), .ZN(P3_U3059) );
  AND4_X2 U14012 ( .A1(n10857), .A2(n10856), .A3(n10855), .A4(n10854), .ZN(
        n10867) );
  AND2_X1 U13123 ( .A1(n10281), .A2(n10280), .ZN(n10871) );
  BUF_X1 U11304 ( .A(n9727), .Z(n20127) );
  INV_X1 U11173 ( .A(n18455), .ZN(n18424) );
  INV_X1 U11167 ( .A(n18502), .ZN(n19377) );
  AND2_X2 U14649 ( .A1(n9731), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11567) );
  NOR2_X1 U11191 ( .A1(n11195), .A2(n10217), .ZN(n11323) );
  AND2_X1 U11212 ( .A1(n10871), .A2(n11152), .ZN(n13356) );
  CLKBUF_X1 U11214 ( .A(n10877), .Z(n15586) );
  CLKBUF_X1 U11247 ( .A(n10865), .Z(n14290) );
  NAND2_X1 U11264 ( .A1(n10284), .A2(n10272), .ZN(n11457) );
  CLKBUF_X1 U11265 ( .A(n13893), .Z(n16817) );
  CLKBUF_X1 U11270 ( .A(n19045), .Z(n9714) );
  CLKBUF_X1 U11318 ( .A(n18734), .Z(n18755) );
  CLKBUF_X2 U11467 ( .A(n11522), .Z(n13869) );
  CLKBUF_X1 U11606 ( .A(n19045), .Z(n9715) );
  CLKBUF_X1 U11607 ( .A(n17694), .Z(n17693) );
  CLKBUF_X1 U11608 ( .A(n13452), .Z(n13523) );
endmodule

