

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4876, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022;

  NAND2_X1 U2372 ( .A1(n4417), .A2(n3988), .ZN(n4411) );
  INV_X1 U2374 ( .A(n2654), .ZN(n2282) );
  CLKBUF_X2 U2375 ( .A(n2547), .Z(n2131) );
  INV_X2 U2376 ( .A(n2134), .ZN(n3973) );
  NAND2_X1 U2377 ( .A1(n2640), .A2(n4277), .ZN(n2686) );
  AND2_X1 U2378 ( .A1(n2686), .A2(n2687), .ZN(n3976) );
  OAI21_X1 U2379 ( .B1(n2135), .B2(n4873), .A(n2744), .ZN(n3404) );
  INV_X1 U2380 ( .A(n3976), .ZN(n3986) );
  BUF_X1 U2381 ( .A(n2769), .Z(n3014) );
  NAND2_X1 U2382 ( .A1(n4682), .A2(n2159), .ZN(n4580) );
  OAI21_X1 U2383 ( .B1(n4138), .B2(n4140), .A(n4139), .ZN(n4018) );
  OAI21_X1 U2384 ( .B1(n2135), .B2(n2354), .A(n2694), .ZN(n3242) );
  AND2_X1 U2385 ( .A1(n2215), .A2(n2213), .ZN(n4933) );
  NAND2_X1 U2386 ( .A1(n4558), .A2(n2234), .ZN(n4504) );
  XNOR2_X1 U2387 ( .A(n2428), .B(IR_REG_22__SCAN_IN), .ZN(n4345) );
  NAND2_X1 U2388 ( .A1(n4933), .A2(n2537), .ZN(n3950) );
  AND4_X1 U2389 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n2130)
         );
  NAND2_X1 U2390 ( .A1(n2445), .A2(n2444), .ZN(n4209) );
  AND2_X2 U2391 ( .A1(n2296), .A2(n2297), .ZN(n2424) );
  OAI21_X2 U2392 ( .B1(n3602), .B2(n3120), .A(n4299), .ZN(n3391) );
  INV_X1 U2393 ( .A(n3392), .ZN(n3441) );
  NOR2_X2 U2394 ( .A1(n4897), .A2(n4898), .ZN(n4896) );
  NOR2_X2 U2395 ( .A1(n3350), .A2(n3349), .ZN(n3348) );
  NAND2_X1 U2396 ( .A1(n3972), .A2(n3971), .ZN(n3985) );
  NAND2_X1 U2397 ( .A1(n3112), .A2(n4278), .ZN(n3243) );
  NAND2_X1 U2398 ( .A1(n3119), .A2(n4299), .ZN(n4249) );
  NAND2_X2 U2399 ( .A1(n3441), .A2(n3603), .ZN(n4299) );
  AND4_X1 U2400 ( .A1(n2820), .A2(n2819), .A3(n2818), .A4(n2817), .ZN(n4062)
         );
  NAND4_X1 U2401 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2712), .ZN(n3551)
         );
  AND4_X1 U2402 ( .A1(n2773), .A2(n2772), .A3(n2771), .A4(n2770), .ZN(n3392)
         );
  AND4_X1 U2403 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n3478)
         );
  NAND2_X1 U2404 ( .A1(n2732), .A2(REG0_REG_2__SCAN_IN), .ZN(n2712) );
  INV_X1 U2405 ( .A(n2699), .ZN(n2641) );
  NAND2_X1 U2406 ( .A1(n2239), .A2(n2240), .ZN(n2535) );
  NAND2_X1 U2407 ( .A1(n3517), .A2(n2778), .ZN(n3439) );
  XNOR2_X1 U2408 ( .A(n2514), .B(n2564), .ZN(n3651) );
  NAND2_X1 U2409 ( .A1(n3069), .A2(n2409), .ZN(n3071) );
  AOI21_X1 U2410 ( .B1(n3345), .B2(n3344), .A(n2397), .ZN(n2562) );
  NAND2_X1 U2412 ( .A1(n3036), .A2(n3035), .ZN(n3113) );
  NAND4_X1 U2413 ( .A1(n2756), .A2(n2755), .A3(n2754), .A4(n2753), .ZN(n4356)
         );
  AND2_X2 U2414 ( .A1(n3218), .A2(n2632), .ZN(n4998) );
  NAND2_X1 U2415 ( .A1(n2642), .A2(n2641), .ZN(n3990) );
  NOR2_X1 U2416 ( .A1(n3233), .A2(n3235), .ZN(n3234) );
  INV_X1 U2417 ( .A(n3035), .ZN(n3305) );
  AND2_X1 U2418 ( .A1(n2674), .A2(n2675), .ZN(n3218) );
  AOI21_X1 U2419 ( .B1(n4882), .B2(REG2_REG_4__SCAN_IN), .A(n2554), .ZN(n3233)
         );
  INV_X2 U2420 ( .A(n2281), .ZN(n2769) );
  XNOR2_X1 U2421 ( .A(n2463), .B(n3213), .ZN(n3210) );
  NAND2_X1 U2422 ( .A1(n4369), .A2(n2458), .ZN(n2463) );
  OAI21_X1 U2423 ( .B1(n2532), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2541) );
  INV_X2 U2424 ( .A(IR_REG_31__SCAN_IN), .ZN(n2517) );
  XNOR2_X1 U2425 ( .A(n4408), .B(n4407), .ZN(n4017) );
  AOI21_X1 U2426 ( .B1(n2147), .B2(n3955), .A(n3954), .ZN(n3956) );
  OAI21_X1 U2427 ( .B1(n4432), .B2(n3100), .A(n3099), .ZN(n4416) );
  AND2_X1 U2428 ( .A1(n3160), .A2(n3159), .ZN(n4012) );
  OR2_X1 U2429 ( .A1(n4932), .A2(n2214), .ZN(n2213) );
  NAND2_X1 U2430 ( .A1(n4921), .A2(n2536), .ZN(n2215) );
  XNOR2_X1 U2431 ( .A(n2535), .B(n4978), .ZN(n4921) );
  NAND2_X1 U2432 ( .A1(n4922), .A2(n2573), .ZN(n4937) );
  NAND2_X1 U2433 ( .A1(n2347), .A2(n2348), .ZN(n2571) );
  OAI21_X1 U2434 ( .B1(n4548), .B2(n3137), .A(n4203), .ZN(n4492) );
  NAND3_X1 U2435 ( .A1(n2212), .A2(n2211), .A3(n2177), .ZN(n2210) );
  NAND2_X1 U2436 ( .A1(n2515), .A2(n2512), .ZN(n2211) );
  NAND2_X1 U2437 ( .A1(n2379), .A2(n2154), .ZN(n3517) );
  NAND2_X1 U2438 ( .A1(n3651), .A2(n2513), .ZN(n2212) );
  NAND2_X1 U2439 ( .A1(n3381), .A2(REG1_REG_10__SCAN_IN), .ZN(n3380) );
  OAI21_X1 U2440 ( .B1(n3280), .B2(n3493), .A(n2561), .ZN(n3345) );
  AOI21_X1 U2441 ( .B1(n2314), .B2(n2315), .A(n2161), .ZN(n2313) );
  INV_X2 U2442 ( .A(n4955), .ZN(n2132) );
  AND3_X1 U2443 ( .A1(n2325), .A2(n2172), .A3(n2328), .ZN(n2559) );
  NAND2_X1 U2444 ( .A1(n2237), .A2(n2477), .ZN(n2483) );
  AND2_X1 U2445 ( .A1(n4274), .A2(n4309), .ZN(n4240) );
  INV_X4 U2446 ( .A(n2730), .ZN(n2823) );
  NAND2_X1 U2447 ( .A1(n3113), .A2(n4275), .ZN(n3110) );
  INV_X1 U2448 ( .A(n2133), .ZN(n2140) );
  INV_X1 U2449 ( .A(n2133), .ZN(n2141) );
  INV_X1 U2450 ( .A(n3367), .ZN(n3475) );
  AND2_X1 U2451 ( .A1(n3115), .A2(n4281), .ZN(n4238) );
  NAND2_X1 U2452 ( .A1(n2251), .A2(n3305), .ZN(n4275) );
  AND3_X1 U2453 ( .A1(n2722), .A2(n2322), .A3(n2725), .ZN(n3367) );
  NAND2_X1 U2454 ( .A1(n2693), .A2(n2692), .ZN(n2698) );
  INV_X1 U2455 ( .A(n3989), .ZN(n2726) );
  NAND2_X1 U2456 ( .A1(n2203), .A2(n2204), .ZN(n2474) );
  INV_X2 U2457 ( .A(n4358), .ZN(U4043) );
  INV_X1 U2458 ( .A(n3365), .ZN(n3374) );
  INV_X1 U2459 ( .A(n2686), .ZN(n2642) );
  INV_X1 U2460 ( .A(n3550), .ZN(n3047) );
  INV_X1 U2461 ( .A(n3609), .ZN(n3603) );
  AND2_X1 U2462 ( .A1(n2553), .A2(n4884), .ZN(n2554) );
  XNOR2_X1 U2463 ( .A(n2553), .B(n2552), .ZN(n4882) );
  NAND2_X1 U2464 ( .A1(n2551), .A2(n2550), .ZN(n2553) );
  CLKBUF_X3 U2465 ( .A(n2875), .Z(n2136) );
  BUF_X2 U2466 ( .A(n2875), .Z(n2137) );
  AND2_X1 U2467 ( .A1(n2602), .A2(n2427), .ZN(n2699) );
  NAND2_X1 U2468 ( .A1(n2324), .A2(n2548), .ZN(n2549) );
  AOI21_X1 U2469 ( .B1(n2443), .B2(n2442), .A(n2441), .ZN(n2444) );
  XNOR2_X1 U2470 ( .A(n2426), .B(n2583), .ZN(n4861) );
  NAND2_X1 U2471 ( .A1(n3962), .A2(IR_REG_31__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U2472 ( .A1(n2195), .A2(n2451), .ZN(n3230) );
  NOR2_X1 U2473 ( .A1(n2507), .A2(n2415), .ZN(n2296) );
  OR2_X1 U2474 ( .A1(n2454), .A2(n2517), .ZN(n2455) );
  NOR2_X1 U2475 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2422)
         );
  INV_X1 U2476 ( .A(IR_REG_27__SCAN_IN), .ZN(n2585) );
  NOR2_X1 U2477 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2421)
         );
  NOR2_X1 U2478 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2420)
         );
  INV_X1 U2479 ( .A(IR_REG_3__SCAN_IN), .ZN(n2460) );
  INV_X1 U2480 ( .A(IR_REG_15__SCAN_IN), .ZN(n2525) );
  INV_X1 U2482 ( .A(IR_REG_16__SCAN_IN), .ZN(n2529) );
  INV_X1 U2483 ( .A(IR_REG_14__SCAN_IN), .ZN(n2518) );
  NOR2_X1 U2484 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2414)
         );
  NOR2_X1 U2485 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2413)
         );
  NOR2_X1 U2486 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2412)
         );
  NOR2_X2 U2487 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2485)
         );
  XNOR2_X1 U2488 ( .A(n2569), .B(n4980), .ZN(n4897) );
  BUF_X4 U2489 ( .A(n3990), .Z(n2133) );
  NAND2_X2 U2490 ( .A1(n3064), .A2(n3063), .ZN(n3397) );
  AOI21_X2 U2491 ( .B1(n4614), .B2(n3086), .A(n2399), .ZN(n4595) );
  NAND2_X2 U2492 ( .A1(n4642), .A2(n3085), .ZN(n4614) );
  INV_X1 U2493 ( .A(n2655), .ZN(n4858) );
  BUF_X4 U2494 ( .A(n4209), .Z(n2135) );
  NAND2_X2 U2495 ( .A1(n4858), .A2(n2282), .ZN(n2281) );
  AND2_X2 U2496 ( .A1(n4858), .A2(n2654), .ZN(n2875) );
  NAND2_X1 U2497 ( .A1(n2445), .A2(n2444), .ZN(n2138) );
  INV_X1 U2498 ( .A(n2680), .ZN(n2139) );
  NAND2_X1 U2499 ( .A1(n2655), .A2(n2654), .ZN(n2680) );
  AND2_X1 U2500 ( .A1(n2364), .A2(n4055), .ZN(n2363) );
  NAND2_X1 U2501 ( .A1(n4162), .A2(n2365), .ZN(n2364) );
  AND2_X1 U2502 ( .A1(n3094), .A2(n2292), .ZN(n2291) );
  NAND2_X1 U2503 ( .A1(n3093), .A2(n3092), .ZN(n3094) );
  NAND2_X1 U2504 ( .A1(n2293), .A2(n3091), .ZN(n2292) );
  AND2_X1 U2505 ( .A1(n4345), .A2(n4277), .ZN(n3156) );
  INV_X1 U2506 ( .A(IR_REG_18__SCAN_IN), .ZN(n2417) );
  NOR2_X1 U2507 ( .A1(n3281), .A2(n2209), .ZN(n3350) );
  AND2_X1 U2508 ( .A1(n2484), .A2(n2558), .ZN(n2209) );
  OAI21_X1 U2509 ( .B1(n3933), .B2(n2351), .A(n2350), .ZN(n2569) );
  NAND2_X1 U2510 ( .A1(n3945), .A2(n2568), .ZN(n2350) );
  NOR2_X1 U2511 ( .A1(n3945), .A2(n2568), .ZN(n2351) );
  NAND2_X1 U2512 ( .A1(n2600), .A2(n2185), .ZN(n2991) );
  AND2_X1 U2513 ( .A1(n4517), .A2(n4537), .ZN(n3088) );
  NAND2_X1 U2514 ( .A1(n2143), .A2(n3145), .ZN(n2261) );
  INV_X1 U2515 ( .A(n4409), .ZN(n4397) );
  NAND2_X1 U2516 ( .A1(n2272), .A2(n2271), .ZN(n4398) );
  NAND2_X1 U2517 ( .A1(n2647), .A2(n2264), .ZN(n2652) );
  NOR2_X1 U2518 ( .A1(n2648), .A2(n2517), .ZN(n2264) );
  NAND2_X1 U2519 ( .A1(n2429), .A2(n2432), .ZN(n2435) );
  AND2_X1 U2520 ( .A1(n2590), .A2(n2589), .ZN(n3199) );
  AND2_X1 U2521 ( .A1(n3199), .A2(n4360), .ZN(n4940) );
  INV_X1 U2522 ( .A(n3117), .ZN(n2258) );
  AOI21_X1 U2523 ( .B1(n4395), .B2(n2277), .A(n4394), .ZN(n2276) );
  INV_X1 U2524 ( .A(n4206), .ZN(n2277) );
  OR2_X1 U2525 ( .A1(n3436), .A2(n3437), .ZN(n2373) );
  NOR2_X1 U2526 ( .A1(n2949), .A2(n2391), .ZN(n2390) );
  INV_X1 U2527 ( .A(n2898), .ZN(n2391) );
  INV_X1 U2528 ( .A(IR_REG_20__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U2529 ( .A1(n2353), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  NAND2_X1 U2530 ( .A1(n4879), .A2(REG1_REG_4__SCAN_IN), .ZN(n2208) );
  NOR2_X1 U2531 ( .A1(n3234), .A2(n2406), .ZN(n2556) );
  AOI21_X1 U2532 ( .B1(n2570), .B2(n2349), .A(n2187), .ZN(n2348) );
  OAI21_X1 U2533 ( .B1(n2306), .B2(n2305), .A(n2179), .ZN(n2304) );
  NAND2_X1 U2534 ( .A1(n4406), .A2(n3988), .ZN(n4395) );
  NAND2_X1 U2535 ( .A1(n4479), .A2(n4458), .ZN(n3097) );
  INV_X1 U2536 ( .A(n2991), .ZN(n2601) );
  OR2_X1 U2537 ( .A1(n4555), .A2(n4537), .ZN(n4493) );
  AND2_X1 U2538 ( .A1(n3156), .A2(n2635), .ZN(n3161) );
  AOI21_X1 U2539 ( .B1(n2269), .B2(n2267), .A(n2164), .ZN(n2266) );
  INV_X1 U2540 ( .A(n2269), .ZN(n2268) );
  INV_X1 U2541 ( .A(n4240), .ZN(n2319) );
  AND2_X1 U2542 ( .A1(n3070), .A2(n2166), .ZN(n2318) );
  NAND2_X1 U2543 ( .A1(n4354), .A2(n3539), .ZN(n2320) );
  OAI21_X1 U2544 ( .B1(n2142), .B2(n2258), .A(n4297), .ZN(n2257) );
  INV_X1 U2545 ( .A(n2258), .ZN(n2254) );
  NOR2_X1 U2546 ( .A1(n4861), .A2(n2395), .ZN(n2427) );
  AND2_X1 U2547 ( .A1(n3121), .A2(n3603), .ZN(n2233) );
  NAND2_X1 U2548 ( .A1(n2419), .A2(IR_REG_31__SCAN_IN), .ZN(n2604) );
  INV_X1 U2549 ( .A(IR_REG_23__SCAN_IN), .ZN(n2603) );
  INV_X1 U2550 ( .A(IR_REG_6__SCAN_IN), .ZN(n2476) );
  NAND2_X1 U2551 ( .A1(n2761), .A2(n2760), .ZN(n2379) );
  OR2_X1 U2552 ( .A1(n2933), .A2(n4133), .ZN(n2916) );
  OR2_X1 U2553 ( .A1(n2633), .A2(n4672), .ZN(n3029) );
  AND2_X1 U2554 ( .A1(n2368), .A2(n4162), .ZN(n2367) );
  INV_X1 U2555 ( .A(n4055), .ZN(n2368) );
  NAND2_X1 U2556 ( .A1(n2359), .A2(n2358), .ZN(n2357) );
  INV_X1 U2557 ( .A(n2363), .ZN(n2358) );
  INV_X1 U2558 ( .A(n2360), .ZN(n2359) );
  INV_X1 U2559 ( .A(n4162), .ZN(n2366) );
  AOI21_X1 U2560 ( .B1(n2367), .B2(n2365), .A(n2361), .ZN(n2360) );
  INV_X1 U2561 ( .A(n4056), .ZN(n2361) );
  NOR2_X1 U2562 ( .A1(n2396), .A2(n2895), .ZN(n2896) );
  INV_X1 U2563 ( .A(n2742), .ZN(n2378) );
  INV_X1 U2564 ( .A(n4874), .ZN(n3213) );
  NAND2_X1 U2565 ( .A1(n2208), .A2(n2149), .ZN(n2207) );
  INV_X1 U2566 ( .A(IR_REG_4__SCAN_IN), .ZN(n2410) );
  XNOR2_X1 U2567 ( .A(n2556), .B(n4872), .ZN(n3203) );
  NAND2_X1 U2568 ( .A1(n3203), .A2(n2330), .ZN(n2328) );
  NOR2_X1 U2569 ( .A1(n3264), .A2(n2331), .ZN(n2330) );
  NAND2_X1 U2570 ( .A1(n2327), .A2(n2326), .ZN(n2325) );
  INV_X1 U2571 ( .A(n3264), .ZN(n2326) );
  INV_X1 U2572 ( .A(n2332), .ZN(n2327) );
  NAND2_X1 U2573 ( .A1(n2236), .A2(n2157), .ZN(n2237) );
  NAND2_X1 U2574 ( .A1(n3379), .A2(REG2_REG_10__SCAN_IN), .ZN(n2339) );
  INV_X1 U2575 ( .A(n3413), .ZN(n2336) );
  AOI21_X1 U2576 ( .B1(n2523), .B2(n2241), .A(n2186), .ZN(n2240) );
  INV_X1 U2577 ( .A(n4909), .ZN(n2241) );
  NAND2_X1 U2578 ( .A1(n4924), .A2(n4923), .ZN(n4922) );
  NOR2_X1 U2579 ( .A1(n2304), .A2(n2302), .ZN(n2301) );
  INV_X1 U2580 ( .A(n3097), .ZN(n2302) );
  INV_X1 U2581 ( .A(n2304), .ZN(n2300) );
  AND2_X1 U2582 ( .A1(n2312), .A2(n2307), .ZN(n2306) );
  NAND2_X1 U2583 ( .A1(n4268), .A2(n4423), .ZN(n2312) );
  NAND2_X1 U2584 ( .A1(n2309), .A2(n2308), .ZN(n2307) );
  INV_X1 U2585 ( .A(n3101), .ZN(n2309) );
  NOR2_X1 U2586 ( .A1(n3101), .A2(n2311), .ZN(n2310) );
  INV_X1 U2587 ( .A(n3099), .ZN(n2311) );
  INV_X1 U2588 ( .A(n4406), .ZN(n4426) );
  INV_X1 U2589 ( .A(n4433), .ZN(n4454) );
  NAND2_X1 U2590 ( .A1(n4351), .A2(n3090), .ZN(n3091) );
  AND2_X1 U2591 ( .A1(n2176), .A2(n4524), .ZN(n2235) );
  NAND2_X1 U2592 ( .A1(n4513), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U2593 ( .A1(n2599), .A2(n2220), .ZN(n2931) );
  NAND2_X1 U2594 ( .A1(n2599), .A2(REG3_REG_17__SCAN_IN), .ZN(n2899) );
  OAI21_X1 U2595 ( .B1(n4656), .B2(n4270), .A(n4316), .ZN(n4624) );
  NAND2_X1 U2596 ( .A1(n4624), .A2(n4645), .ZN(n4623) );
  OR2_X1 U2597 ( .A1(n2874), .A2(n2860), .ZN(n2862) );
  INV_X1 U2598 ( .A(n4672), .ZN(n4700) );
  INV_X1 U2599 ( .A(n4654), .ZN(n4697) );
  CLKBUF_X1 U2600 ( .A(n3046), .Z(n3482) );
  INV_X1 U2601 ( .A(IR_REG_19__SCAN_IN), .ZN(n3791) );
  AND2_X1 U2602 ( .A1(n4283), .A2(n4280), .ZN(n4245) );
  OR2_X1 U2603 ( .A1(n4973), .A2(n2699), .ZN(n3162) );
  AND2_X1 U2604 ( .A1(n2723), .A2(n2724), .ZN(n2322) );
  AND2_X1 U2605 ( .A1(n3218), .A2(n4863), .ZN(n4672) );
  INV_X1 U2606 ( .A(n4405), .ZN(n3988) );
  NOR2_X2 U2607 ( .A1(n4504), .A2(n4115), .ZN(n4482) );
  AND2_X1 U2608 ( .A1(n4707), .A2(n4706), .ZN(n4682) );
  NOR2_X2 U2609 ( .A1(n3632), .A2(n4059), .ZN(n4707) );
  NAND3_X1 U2610 ( .A1(n2602), .A2(n2610), .A3(n2609), .ZN(n3188) );
  NAND2_X1 U2611 ( .A1(n2424), .A2(n2146), .ZN(n2647) );
  INV_X1 U2612 ( .A(IR_REG_17__SCAN_IN), .ZN(n2416) );
  INV_X1 U2613 ( .A(IR_REG_11__SCAN_IN), .ZN(n3669) );
  NOR2_X1 U2614 ( .A1(n2469), .A2(IR_REG_5__SCAN_IN), .ZN(n2509) );
  NOR2_X1 U2615 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2454)
         );
  AND4_X1 U2616 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(n3516)
         );
  INV_X1 U2617 ( .A(n4498), .ZN(n4072) );
  INV_X1 U2618 ( .A(n2384), .ZN(n2383) );
  OAI22_X1 U2619 ( .A1(n2998), .A2(n2385), .B1(n3002), .B2(n3003), .ZN(n2384)
         );
  INV_X1 U2620 ( .A(n4479), .ZN(n4117) );
  AND2_X1 U2621 ( .A1(n2991), .A2(n2990), .ZN(n4486) );
  AND2_X1 U2622 ( .A1(n2912), .A2(n2911), .ZN(n4517) );
  INV_X1 U2623 ( .A(n4165), .ZN(n4194) );
  XNOR2_X1 U2624 ( .A(n2474), .B(n4872), .ZN(n3202) );
  NAND2_X1 U2625 ( .A1(n2197), .A2(n2196), .ZN(n3381) );
  XNOR2_X1 U2626 ( .A(n2562), .B(n4869), .ZN(n3379) );
  OR2_X1 U2627 ( .A1(n2565), .A2(n2564), .ZN(n2566) );
  NAND2_X1 U2628 ( .A1(n2341), .A2(n2340), .ZN(n2579) );
  NAND2_X1 U2629 ( .A1(n2246), .A2(n2249), .ZN(n2245) );
  NAND2_X1 U2630 ( .A1(n2543), .A2(n2250), .ZN(n2249) );
  INV_X1 U2631 ( .A(n3949), .ZN(n2250) );
  NAND2_X1 U2632 ( .A1(n2259), .A2(n2261), .ZN(n2283) );
  AOI21_X1 U2633 ( .B1(n4721), .B2(n4787), .A(n2217), .ZN(n2259) );
  NAND2_X1 U2634 ( .A1(n4403), .A2(n2260), .ZN(n2217) );
  INV_X1 U2635 ( .A(n4906), .ZN(n2349) );
  INV_X1 U2636 ( .A(n4291), .ZN(n2267) );
  XNOR2_X1 U2637 ( .A(IR_REG_27__SCAN_IN), .B(IR_REG_28__SCAN_IN), .ZN(n2439)
         );
  NOR2_X1 U2638 ( .A1(n2751), .A2(n2216), .ZN(n2749) );
  NAND2_X1 U2639 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_5__SCAN_IN), .ZN(
        n2216) );
  AND2_X1 U2640 ( .A1(n3100), .A2(n3099), .ZN(n2308) );
  NAND2_X1 U2641 ( .A1(n4420), .A2(n4206), .ZN(n4396) );
  NOR2_X1 U2642 ( .A1(n4442), .A2(n3157), .ZN(n3158) );
  NOR2_X1 U2643 ( .A1(n2219), .A2(n4156), .ZN(n2218) );
  INV_X1 U2644 ( .A(n2957), .ZN(n2600) );
  OR2_X1 U2645 ( .A1(n4351), .A2(n4524), .ZN(n4494) );
  AND2_X1 U2646 ( .A1(n2405), .A2(n4201), .ZN(n2280) );
  NOR2_X1 U2647 ( .A1(n3951), .A2(n2221), .ZN(n2220) );
  INV_X1 U2648 ( .A(n2884), .ZN(n2599) );
  NOR2_X1 U2649 ( .A1(n2226), .A2(n2225), .ZN(n2224) );
  INV_X1 U2650 ( .A(n2815), .ZN(n2597) );
  INV_X1 U2651 ( .A(n4308), .ZN(n2270) );
  NAND2_X1 U2652 ( .A1(n3047), .A2(n3367), .ZN(n2321) );
  INV_X1 U2653 ( .A(n3244), .ZN(n4278) );
  AND2_X1 U2654 ( .A1(n2276), .A2(n3143), .ZN(n2273) );
  OAI21_X1 U2655 ( .B1(n3142), .B2(n2275), .A(n2276), .ZN(n2271) );
  NAND2_X1 U2656 ( .A1(n4395), .A2(n4422), .ZN(n2275) );
  NOR2_X1 U2657 ( .A1(n3171), .A2(n4673), .ZN(n2229) );
  INV_X1 U2658 ( .A(n3373), .ZN(n3168) );
  OR2_X1 U2659 ( .A1(n3188), .A2(n2621), .ZN(n3164) );
  INV_X1 U2660 ( .A(IR_REG_28__SCAN_IN), .ZN(n2582) );
  NOR2_X1 U2661 ( .A1(IR_REG_29__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2649)
         );
  INV_X1 U2662 ( .A(n4112), .ZN(n2385) );
  AND2_X1 U2663 ( .A1(n2985), .A2(n2180), .ZN(n2381) );
  NAND2_X1 U2664 ( .A1(n3436), .A2(n3437), .ZN(n2371) );
  OR2_X1 U2665 ( .A1(n2786), .A2(n2596), .ZN(n2797) );
  NAND2_X1 U2666 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2596) );
  NAND2_X1 U2667 ( .A1(n2749), .A2(REG3_REG_7__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U2668 ( .A1(n2597), .A2(n2224), .ZN(n2840) );
  AOI21_X1 U2669 ( .B1(n2390), .B2(n2388), .A(n2162), .ZN(n2387) );
  INV_X1 U2670 ( .A(n2390), .ZN(n2389) );
  INV_X1 U2671 ( .A(n2896), .ZN(n2388) );
  OR2_X1 U2672 ( .A1(n2916), .A2(n4049), .ZN(n2957) );
  OR2_X1 U2673 ( .A1(n2797), .A2(n3382), .ZN(n2815) );
  NAND2_X1 U2674 ( .A1(n2597), .A2(REG3_REG_11__SCAN_IN), .ZN(n2828) );
  OAI22_X1 U2675 ( .A1(n3036), .A2(n3990), .B1(n3305), .B2(n3989), .ZN(n2688)
         );
  OAI22_X1 U2676 ( .A1(n2730), .A2(n3036), .B1(n3305), .B2(n2133), .ZN(n2705)
         );
  INV_X1 U2677 ( .A(n4598), .ZN(n4179) );
  INV_X1 U2678 ( .A(REG3_REG_18__SCAN_IN), .ZN(n3951) );
  INV_X1 U2679 ( .A(n3406), .ZN(n3616) );
  NAND2_X1 U2680 ( .A1(n2629), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  AND2_X1 U2681 ( .A1(n3153), .A2(n3152), .ZN(n4207) );
  AND4_X1 U2682 ( .A1(n2879), .A2(n2878), .A3(n2877), .A4(n2876), .ZN(n3076)
         );
  NAND2_X1 U2683 ( .A1(n3231), .A2(n2144), .ZN(n2204) );
  NAND2_X1 U2684 ( .A1(n2205), .A2(n2208), .ZN(n2203) );
  AND2_X1 U2685 ( .A1(n2149), .A2(n2144), .ZN(n2205) );
  AND2_X1 U2686 ( .A1(n3283), .A2(REG1_REG_8__SCAN_IN), .ZN(n3281) );
  OR2_X1 U2687 ( .A1(n2487), .A2(n2486), .ZN(n2489) );
  NAND2_X1 U2688 ( .A1(n2200), .A2(n2398), .ZN(n2199) );
  NAND2_X1 U2689 ( .A1(n2202), .A2(n4869), .ZN(n2201) );
  INV_X1 U2690 ( .A(n2398), .ZN(n2202) );
  INV_X1 U2691 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U2692 ( .A1(n2334), .A2(n2333), .ZN(n2565) );
  NAND2_X1 U2693 ( .A1(n3413), .A2(n2174), .ZN(n2333) );
  NAND2_X1 U2694 ( .A1(n2339), .A2(n2335), .ZN(n2334) );
  AND2_X1 U2695 ( .A1(n2338), .A2(n2174), .ZN(n2335) );
  INV_X1 U2696 ( .A(n2210), .ZN(n2522) );
  INV_X1 U2697 ( .A(n4935), .ZN(n2214) );
  NOR2_X1 U2698 ( .A1(n2577), .A2(n2343), .ZN(n2342) );
  INV_X1 U2699 ( .A(n4938), .ZN(n2343) );
  NAND2_X1 U2700 ( .A1(n2345), .A2(n2346), .ZN(n2340) );
  OAI21_X1 U2701 ( .B1(n2248), .B2(n2543), .A(n2247), .ZN(n2246) );
  AND2_X1 U2702 ( .A1(n2539), .A2(n3949), .ZN(n2248) );
  NAND2_X1 U2703 ( .A1(n2543), .A2(n2539), .ZN(n2247) );
  NOR2_X1 U2704 ( .A1(n2664), .A2(n4071), .ZN(n2228) );
  NAND2_X1 U2705 ( .A1(n2278), .A2(n2279), .ZN(n4420) );
  NOR2_X1 U2706 ( .A1(n3142), .A2(n2274), .ZN(n2278) );
  INV_X1 U2707 ( .A(n4422), .ZN(n2274) );
  INV_X1 U2708 ( .A(n4445), .ZN(n4439) );
  AOI21_X1 U2709 ( .B1(n2291), .B2(n2294), .A(n2152), .ZN(n2290) );
  INV_X1 U2710 ( .A(n3091), .ZN(n2294) );
  NAND2_X1 U2711 ( .A1(n2600), .A2(REG3_REG_22__SCAN_IN), .ZN(n2972) );
  NAND2_X1 U2712 ( .A1(n2600), .A2(n2218), .ZN(n2989) );
  AND2_X1 U2713 ( .A1(n4228), .A2(n4493), .ZN(n4531) );
  NAND2_X1 U2714 ( .A1(n4623), .A2(n4201), .ZN(n4607) );
  OR2_X1 U2715 ( .A1(n2862), .A2(n4088), .ZN(n2884) );
  INV_X1 U2716 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4088) );
  OAI21_X1 U2717 ( .B1(n4634), .B2(n3081), .A(n3080), .ZN(n3084) );
  AND2_X1 U2718 ( .A1(n4201), .A2(n4317), .ZN(n4645) );
  AND3_X1 U2719 ( .A1(n2888), .A2(n2887), .A3(n2886), .ZN(n4622) );
  INV_X1 U2720 ( .A(n4629), .ZN(n4653) );
  NAND2_X1 U2721 ( .A1(n3127), .A2(n4272), .ZN(n4656) );
  NAND2_X1 U2722 ( .A1(n2597), .A2(n2223), .ZN(n2872) );
  AND2_X1 U2723 ( .A1(n2224), .A2(REG3_REG_13__SCAN_IN), .ZN(n2223) );
  NAND2_X1 U2724 ( .A1(n2598), .A2(REG3_REG_14__SCAN_IN), .ZN(n2874) );
  INV_X1 U2725 ( .A(n2872), .ZN(n2598) );
  INV_X1 U2726 ( .A(n2318), .ZN(n2314) );
  NAND2_X1 U2727 ( .A1(n2265), .A2(n2269), .ZN(n3571) );
  NAND2_X1 U2728 ( .A1(n3457), .A2(n4291), .ZN(n2265) );
  NAND2_X1 U2729 ( .A1(n2317), .A2(n2320), .ZN(n3574) );
  NAND2_X1 U2730 ( .A1(n3071), .A2(n2318), .ZN(n2317) );
  NAND3_X1 U2731 ( .A1(n3397), .A2(n2408), .A3(n2287), .ZN(n2286) );
  INV_X1 U2732 ( .A(n2173), .ZN(n2252) );
  NAND2_X1 U2733 ( .A1(n2254), .A2(n2173), .ZN(n2253) );
  INV_X1 U2734 ( .A(n2257), .ZN(n2256) );
  NAND2_X1 U2735 ( .A1(n2255), .A2(n3117), .ZN(n3502) );
  NAND2_X1 U2736 ( .A1(n3548), .A2(n2142), .ZN(n2255) );
  NAND2_X1 U2737 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2751) );
  AND2_X1 U2738 ( .A1(n2235), .A2(n3092), .ZN(n2234) );
  INV_X1 U2739 ( .A(n4533), .ZN(n4537) );
  AND2_X1 U2740 ( .A1(n4558), .A2(n4553), .ZN(n4560) );
  AND2_X1 U2741 ( .A1(n4682), .A2(n2150), .ZN(n2401) );
  NAND2_X1 U2742 ( .A1(n2233), .A2(n3595), .ZN(n2232) );
  NAND2_X1 U2743 ( .A1(n3170), .A2(n3603), .ZN(n3611) );
  INV_X1 U2744 ( .A(n3610), .ZN(n3170) );
  NAND2_X1 U2745 ( .A1(n3241), .A2(n3374), .ZN(n3373) );
  INV_X1 U2746 ( .A(n4995), .ZN(n4987) );
  AND2_X1 U2747 ( .A1(n4946), .A2(n2674), .ZN(n4995) );
  AND2_X1 U2748 ( .A1(n2130), .A2(n2583), .ZN(n2386) );
  NAND2_X1 U2749 ( .A1(n2446), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  XNOR2_X1 U2750 ( .A(n2607), .B(n2606), .ZN(n2624) );
  INV_X1 U2751 ( .A(IR_REG_24__SCAN_IN), .ZN(n2606) );
  NAND2_X1 U2752 ( .A1(n2605), .A2(IR_REG_31__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U2753 ( .A1(n2379), .A2(n3335), .ZN(n3519) );
  AND2_X1 U2754 ( .A1(n3019), .A2(n3018), .ZN(n4461) );
  AND4_X1 U2755 ( .A1(n2845), .A2(n2844), .A3(n2843), .A4(n2842), .ZN(n4677)
         );
  INV_X1 U2756 ( .A(n4355), .ZN(n3444) );
  INV_X1 U2757 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4049) );
  NAND2_X1 U2758 ( .A1(n2369), .A2(n4162), .ZN(n4054) );
  NAND2_X1 U2759 ( .A1(n3325), .A2(n2742), .ZN(n3319) );
  AND2_X1 U2760 ( .A1(n2905), .A2(n2904), .ZN(n4610) );
  NAND2_X1 U2761 ( .A1(n4026), .A2(n2998), .ZN(n4110) );
  NAND2_X1 U2762 ( .A1(n4026), .A2(n3002), .ZN(n2382) );
  NAND2_X1 U2763 ( .A1(n3326), .A2(n2738), .ZN(n3325) );
  NAND2_X1 U2764 ( .A1(n3439), .A2(n3437), .ZN(n2375) );
  NAND2_X1 U2765 ( .A1(n2370), .A2(n3436), .ZN(n2374) );
  OR2_X1 U2766 ( .A1(n3439), .A2(n3437), .ZN(n2370) );
  INV_X1 U2767 ( .A(n3242), .ZN(n3968) );
  INV_X1 U2768 ( .A(n4191), .ZN(n4180) );
  AND2_X1 U2769 ( .A1(n3031), .A2(n3030), .ZN(n4102) );
  INV_X1 U2770 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4133) );
  AOI21_X1 U2771 ( .B1(n2360), .B2(n2362), .A(n2165), .ZN(n2355) );
  INV_X1 U2772 ( .A(n2367), .ZN(n2362) );
  NAND2_X1 U2773 ( .A1(n2897), .A2(n2896), .ZN(n2392) );
  INV_X1 U2774 ( .A(n4169), .ZN(n4192) );
  AND2_X1 U2775 ( .A1(n3031), .A2(n2673), .ZN(n4165) );
  AOI21_X1 U2776 ( .B1(n2378), .B2(n3318), .A(n2158), .ZN(n2377) );
  NAND2_X1 U2777 ( .A1(n3108), .A2(n3107), .ZN(n4406) );
  OR2_X1 U2778 ( .A1(n4011), .A2(n2281), .ZN(n3108) );
  INV_X1 U2779 ( .A(n4461), .ZN(n4350) );
  NAND2_X1 U2780 ( .A1(n2660), .A2(n2659), .ZN(n4479) );
  OR2_X1 U2781 ( .A1(n4465), .A2(n2281), .ZN(n2660) );
  NAND2_X1 U2782 ( .A1(n2996), .A2(n2995), .ZN(n4498) );
  INV_X1 U2783 ( .A(n4517), .ZN(n4555) );
  NAND2_X1 U2784 ( .A1(n2921), .A2(n2920), .ZN(n4576) );
  OR2_X1 U2785 ( .A1(n4132), .A2(n2281), .ZN(n2921) );
  NAND2_X1 U2786 ( .A1(n2938), .A2(n2937), .ZN(n4352) );
  INV_X1 U2787 ( .A(n4610), .ZN(n4035) );
  OAI211_X1 U2788 ( .C1(n4650), .C2(n2281), .A(n2866), .B(n2865), .ZN(n4674)
         );
  INV_X1 U2789 ( .A(n3076), .ZN(n4698) );
  INV_X1 U2790 ( .A(n4677), .ZN(n4058) );
  INV_X1 U2791 ( .A(n4062), .ZN(n4353) );
  INV_X1 U2792 ( .A(n3516), .ZN(n3606) );
  NAND2_X1 U2793 ( .A1(n2137), .A2(REG2_REG_6__SCAN_IN), .ZN(n2754) );
  OR2_X1 U2794 ( .A1(n4973), .A2(n2641), .ZN(n4358) );
  NAND2_X1 U2795 ( .A1(n2450), .A2(n2145), .ZN(n2193) );
  INV_X1 U2796 ( .A(n3231), .ZN(n2206) );
  INV_X1 U2797 ( .A(n2207), .ZN(n3232) );
  AND2_X1 U2798 ( .A1(n2236), .A2(n2238), .ZN(n3260) );
  AND2_X1 U2799 ( .A1(n2329), .A2(n2332), .ZN(n3265) );
  NAND2_X1 U2800 ( .A1(n3203), .A2(REG2_REG_6__SCAN_IN), .ZN(n2329) );
  XNOR2_X1 U2801 ( .A(n2483), .B(n2558), .ZN(n3283) );
  NAND2_X1 U2802 ( .A1(n2560), .A2(n2558), .ZN(n2561) );
  NAND2_X1 U2803 ( .A1(n3380), .A2(n2493), .ZN(n3421) );
  INV_X1 U2804 ( .A(n2337), .ZN(n3414) );
  NAND2_X1 U2805 ( .A1(n2339), .A2(n2338), .ZN(n2337) );
  NAND2_X1 U2806 ( .A1(n2212), .A2(n2211), .ZN(n3938) );
  NOR2_X1 U2807 ( .A1(n4894), .A2(n4895), .ZN(n4893) );
  XNOR2_X1 U2808 ( .A(n2210), .B(n4901), .ZN(n4894) );
  NOR2_X1 U2809 ( .A1(n4896), .A2(n2570), .ZN(n4907) );
  NOR2_X1 U2810 ( .A1(n4893), .A2(n2523), .ZN(n4910) );
  AND2_X1 U2811 ( .A1(n3199), .A2(n3154), .ZN(n4914) );
  INV_X1 U2812 ( .A(n4914), .ZN(n4945) );
  NAND2_X1 U2813 ( .A1(n4936), .A2(n2576), .ZN(n3946) );
  XNOR2_X1 U2814 ( .A(n4410), .B(n4409), .ZN(n4721) );
  NAND2_X1 U2815 ( .A1(n2300), .A2(n2163), .ZN(n2299) );
  NAND2_X1 U2816 ( .A1(n2303), .A2(n2306), .ZN(n4408) );
  NAND2_X1 U2817 ( .A1(n4432), .A2(n2310), .ZN(n2303) );
  NAND2_X1 U2818 ( .A1(n4511), .A2(n3091), .ZN(n4491) );
  AND2_X1 U2819 ( .A1(n4521), .A2(n4520), .ZN(n4744) );
  OAI21_X1 U2820 ( .B1(n3427), .B2(n3426), .A(n4649), .ZN(n4652) );
  NAND2_X1 U2821 ( .A1(n2629), .A2(n2542), .ZN(n4341) );
  NAND2_X1 U2822 ( .A1(n3548), .A2(n4283), .ZN(n3468) );
  OR2_X1 U2823 ( .A1(n3162), .A2(n3163), .ZN(n4649) );
  INV_X1 U2824 ( .A(n4668), .ZN(n4711) );
  AND2_X1 U2825 ( .A1(n4600), .A2(n4998), .ZN(n4668) );
  INV_X1 U2826 ( .A(n4649), .ZN(n4950) );
  XOR2_X1 U2827 ( .A(n4377), .B(n4382), .Z(n4798) );
  NAND2_X1 U2828 ( .A1(n3188), .A2(n3302), .ZN(n4972) );
  AND2_X1 U2829 ( .A1(n2297), .A2(n2648), .ZN(n2295) );
  INV_X1 U2830 ( .A(IR_REG_30__SCAN_IN), .ZN(n3959) );
  INV_X1 U2831 ( .A(n2624), .ZN(n3193) );
  NAND2_X1 U2832 ( .A1(n2638), .A2(STATE_REG_SCAN_IN), .ZN(n4973) );
  NAND2_X1 U2833 ( .A1(n2432), .A2(IR_REG_31__SCAN_IN), .ZN(n2433) );
  AND2_X1 U2834 ( .A1(n2528), .A2(n2527), .ZN(n4913) );
  INV_X1 U2835 ( .A(n2506), .ZN(n2511) );
  XNOR2_X1 U2836 ( .A(n2501), .B(IR_REG_12__SCAN_IN), .ZN(n4867) );
  XNOR2_X1 U2837 ( .A(n2479), .B(IR_REG_7__SCAN_IN), .ZN(n4871) );
  XNOR2_X1 U2838 ( .A(n2473), .B(IR_REG_6__SCAN_IN), .ZN(n4872) );
  AND2_X1 U2839 ( .A1(n2466), .A2(n2462), .ZN(n4874) );
  NAND2_X1 U2840 ( .A1(n4942), .A2(n2245), .ZN(n2243) );
  NAND2_X1 U2841 ( .A1(n2263), .A2(n2175), .ZN(U3547) );
  NAND2_X1 U2842 ( .A1(n2283), .A2(n5022), .ZN(n2263) );
  INV_X1 U2843 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2262) );
  OR2_X1 U2844 ( .A1(n4010), .A2(n4794), .ZN(n3172) );
  NAND2_X1 U2845 ( .A1(n2282), .A2(STATE_REG_SCAN_IN), .ZN(n3183) );
  AND2_X1 U2846 ( .A1(n3116), .A2(n4283), .ZN(n2142) );
  XOR2_X1 U2847 ( .A(n4398), .B(n4397), .Z(n2143) );
  NAND2_X1 U2848 ( .A1(n4873), .A2(REG1_REG_5__SCAN_IN), .ZN(n2144) );
  AND2_X1 U2849 ( .A1(n2449), .A2(REG1_REG_1__SCAN_IN), .ZN(n2145) );
  AND2_X1 U2850 ( .A1(n2130), .A2(n2151), .ZN(n2146) );
  INV_X1 U2851 ( .A(n2316), .ZN(n2315) );
  NAND2_X1 U2852 ( .A1(n2319), .A2(n2320), .ZN(n2316) );
  INV_X4 U2853 ( .A(n2680), .ZN(n2732) );
  NAND2_X1 U2854 ( .A1(n4393), .A2(n4395), .ZN(n4407) );
  INV_X1 U2855 ( .A(n4407), .ZN(n2305) );
  INV_X1 U2856 ( .A(n4104), .ZN(n2230) );
  INV_X1 U2857 ( .A(n4942), .ZN(n4908) );
  AND2_X1 U2858 ( .A1(n3199), .A2(n4359), .ZN(n4942) );
  INV_X1 U2859 ( .A(n2137), .ZN(n3150) );
  NAND2_X1 U2860 ( .A1(n2392), .A2(n2898), .ZN(n4033) );
  OR2_X1 U2861 ( .A1(n3950), .A2(n3949), .ZN(n2147) );
  OR2_X1 U2862 ( .A1(n3032), .A2(n4199), .ZN(n2148) );
  NAND2_X1 U2863 ( .A1(n2468), .A2(n4884), .ZN(n2149) );
  AND2_X1 U2864 ( .A1(n2229), .A2(n4104), .ZN(n2150) );
  INV_X1 U2865 ( .A(n4161), .ZN(n2365) );
  AND4_X1 U2866 ( .A1(n2584), .A2(n2585), .A3(n2582), .A4(n2583), .ZN(n2151)
         );
  AND2_X1 U2867 ( .A1(n4519), .A2(n4502), .ZN(n2152) );
  AND2_X1 U2868 ( .A1(n3516), .A2(n3121), .ZN(n2153) );
  NAND2_X1 U2869 ( .A1(n4623), .A2(n2280), .ZN(n4548) );
  NAND2_X1 U2870 ( .A1(n2382), .A2(n3004), .ZN(n4109) );
  AND2_X1 U2871 ( .A1(n3335), .A2(n2775), .ZN(n2154) );
  NOR2_X1 U2872 ( .A1(n4907), .A2(n4906), .ZN(n2155) );
  NOR2_X1 U2873 ( .A1(n4910), .A2(n4909), .ZN(n2156) );
  AND2_X1 U2874 ( .A1(n2238), .A2(n2393), .ZN(n2157) );
  INV_X1 U2875 ( .A(n4354), .ZN(n4170) );
  AND2_X1 U2876 ( .A1(n2748), .A2(n2747), .ZN(n2158) );
  AND2_X1 U2877 ( .A1(n2150), .A2(n4179), .ZN(n2159) );
  AND2_X1 U2878 ( .A1(n2796), .A2(n2371), .ZN(n2160) );
  AND2_X1 U2879 ( .A1(n4062), .A2(n3573), .ZN(n2161) );
  NOR2_X1 U2880 ( .A1(n2956), .A2(n2955), .ZN(n2162) );
  NAND2_X1 U2881 ( .A1(n4407), .A2(n2310), .ZN(n2163) );
  NAND2_X1 U2882 ( .A1(n4305), .A2(n4274), .ZN(n2164) );
  AND2_X1 U2883 ( .A1(n2363), .A2(n2366), .ZN(n2165) );
  OR2_X1 U2884 ( .A1(n4354), .A2(n3539), .ZN(n2166) );
  INV_X1 U2885 ( .A(n3121), .ZN(n3440) );
  AND2_X1 U2886 ( .A1(n4936), .A2(n2344), .ZN(n2167) );
  INV_X1 U2887 ( .A(n4329), .ZN(n3142) );
  AND2_X1 U2888 ( .A1(n2683), .A2(n2682), .ZN(n2168) );
  AND2_X1 U2889 ( .A1(n3318), .A2(n2738), .ZN(n2169) );
  AND2_X1 U2890 ( .A1(n2595), .A2(n2594), .ZN(n2170) );
  OR2_X1 U2891 ( .A1(n2451), .A2(n2194), .ZN(n2171) );
  INV_X1 U2892 ( .A(IR_REG_25__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U2893 ( .A1(n4871), .A2(REG2_REG_7__SCAN_IN), .ZN(n2172) );
  INV_X1 U2894 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2194) );
  NAND2_X1 U2895 ( .A1(n4682), .A2(n4683), .ZN(n4628) );
  XNOR2_X1 U2896 ( .A(n2491), .B(IR_REG_10__SCAN_IN), .ZN(n4869) );
  INV_X1 U2897 ( .A(n4512), .ZN(n2293) );
  NAND2_X1 U2898 ( .A1(n2567), .A2(n2566), .ZN(n3933) );
  NAND2_X1 U2899 ( .A1(n4357), .A2(n3404), .ZN(n2173) );
  NAND2_X1 U2900 ( .A1(n2511), .A2(n2510), .ZN(n3945) );
  NAND2_X1 U2901 ( .A1(n2424), .A2(n2386), .ZN(n2446) );
  NAND2_X1 U2902 ( .A1(n2372), .A2(n2160), .ZN(n3592) );
  XNOR2_X1 U2903 ( .A(n2631), .B(n2630), .ZN(n2640) );
  NAND2_X1 U2904 ( .A1(n4868), .A2(REG2_REG_11__SCAN_IN), .ZN(n2174) );
  NAND2_X1 U2905 ( .A1(n2356), .A2(n2355), .ZN(n4138) );
  NAND2_X1 U2906 ( .A1(n3071), .A2(n3070), .ZN(n3535) );
  XNOR2_X1 U2907 ( .A(n2565), .B(n4867), .ZN(n3650) );
  NAND2_X1 U2908 ( .A1(n2376), .A2(n2377), .ZN(n3334) );
  OR2_X1 U2909 ( .A1(n5022), .A2(n2262), .ZN(n2175) );
  NAND2_X1 U2910 ( .A1(n4558), .A2(n2235), .ZN(n4501) );
  AND2_X1 U2911 ( .A1(n4553), .A2(n4537), .ZN(n2176) );
  NAND2_X1 U2912 ( .A1(n2374), .A2(n2375), .ZN(n3591) );
  INV_X1 U2913 ( .A(n2424), .ZN(n2586) );
  OR2_X1 U2914 ( .A1(n3945), .A2(n4783), .ZN(n2177) );
  INV_X1 U2915 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2225) );
  NAND2_X1 U2916 ( .A1(n4682), .A2(n2229), .ZN(n2231) );
  INV_X1 U2917 ( .A(IR_REG_0__SCAN_IN), .ZN(n2354) );
  AND2_X1 U2918 ( .A1(n2317), .A2(n2315), .ZN(n2178) );
  NAND2_X1 U2919 ( .A1(n4406), .A2(n4405), .ZN(n2179) );
  OR2_X1 U2920 ( .A1(n4112), .A2(n3004), .ZN(n2180) );
  AND2_X1 U2921 ( .A1(n2882), .A2(n2881), .ZN(n2181) );
  AND2_X1 U2922 ( .A1(n4558), .A2(n2176), .ZN(n4523) );
  AND2_X1 U2923 ( .A1(n2220), .A2(REG3_REG_19__SCAN_IN), .ZN(n2182) );
  AND2_X1 U2924 ( .A1(n2500), .A2(n2498), .ZN(n4868) );
  AND2_X1 U2925 ( .A1(n2337), .A2(n2336), .ZN(n2183) );
  NOR2_X1 U2926 ( .A1(n3610), .A2(n2232), .ZN(n3461) );
  NOR2_X1 U2927 ( .A1(n3035), .A2(n3242), .ZN(n3241) );
  NOR2_X1 U2928 ( .A1(n3481), .A2(n3482), .ZN(n3403) );
  NAND2_X1 U2929 ( .A1(n2288), .A2(n3067), .ZN(n3390) );
  OR2_X1 U2930 ( .A1(n2543), .A2(n2540), .ZN(n2184) );
  NAND2_X1 U2931 ( .A1(n2328), .A2(n2325), .ZN(n3263) );
  AND2_X1 U2932 ( .A1(n2218), .A2(REG3_REG_24__SCAN_IN), .ZN(n2185) );
  INV_X1 U2933 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2221) );
  INV_X1 U2934 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2222) );
  INV_X1 U2935 ( .A(n2577), .ZN(n2346) );
  AND2_X1 U2936 ( .A1(n4865), .A2(REG2_REG_18__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U2937 ( .A1(n2246), .A2(n2184), .ZN(n2244) );
  AND2_X1 U2938 ( .A1(n4913), .A2(REG1_REG_15__SCAN_IN), .ZN(n2186) );
  AND2_X1 U2939 ( .A1(n4913), .A2(REG2_REG_15__SCAN_IN), .ZN(n2187) );
  INV_X1 U2940 ( .A(n2345), .ZN(n2344) );
  OR2_X1 U2941 ( .A1(n3947), .A2(n2575), .ZN(n2345) );
  AND2_X1 U2942 ( .A1(n3170), .A2(n2233), .ZN(n2188) );
  AND2_X1 U2943 ( .A1(n4942), .A2(n2244), .ZN(n2189) );
  AND2_X1 U2944 ( .A1(n2545), .A2(n2546), .ZN(n2190) );
  AND2_X1 U2945 ( .A1(n2207), .A2(n2206), .ZN(n2191) );
  INV_X1 U2946 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U2947 ( .A1(n3223), .A2(n3222), .ZN(n2453) );
  NAND3_X1 U2948 ( .A1(n2171), .A2(n2192), .A3(n2193), .ZN(n3223) );
  NAND3_X1 U2949 ( .A1(n2451), .A2(n2195), .A3(n2194), .ZN(n2192) );
  NAND2_X1 U2950 ( .A1(n2450), .A2(n2449), .ZN(n2195) );
  NAND2_X1 U2951 ( .A1(n3348), .A2(n2200), .ZN(n2196) );
  INV_X1 U2952 ( .A(n2198), .ZN(n2197) );
  OAI21_X1 U2953 ( .B1(n3348), .B2(n2201), .A(n2199), .ZN(n2198) );
  NOR2_X1 U2954 ( .A1(n3348), .A2(n2398), .ZN(n2492) );
  INV_X1 U2955 ( .A(n4869), .ZN(n2200) );
  INV_X1 U2956 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2219) );
  NAND2_X1 U2957 ( .A1(n2599), .A2(n2182), .ZN(n2933) );
  INV_X1 U2958 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2959 ( .A1(n2601), .A2(n2228), .ZN(n3103) );
  NAND2_X1 U2960 ( .A1(n3103), .A2(n3832), .ZN(n2227) );
  NAND2_X1 U2961 ( .A1(n2601), .A2(REG3_REG_25__SCAN_IN), .ZN(n2665) );
  NAND2_X1 U2962 ( .A1(n4392), .A2(n2227), .ZN(n4011) );
  INV_X1 U2963 ( .A(n2231), .ZN(n4615) );
  NOR2_X2 U2964 ( .A1(n4411), .A2(n4412), .ZN(n4384) );
  NOR2_X4 U2965 ( .A1(n4444), .A2(n4423), .ZN(n4417) );
  NAND2_X1 U2966 ( .A1(n3202), .A2(REG1_REG_6__SCAN_IN), .ZN(n2236) );
  NAND2_X1 U2967 ( .A1(n2475), .A2(n4872), .ZN(n2238) );
  NAND2_X1 U2968 ( .A1(n4893), .A2(n2241), .ZN(n2239) );
  INV_X1 U2969 ( .A(n2535), .ZN(n2531) );
  NAND2_X1 U2970 ( .A1(n3950), .A2(n2189), .ZN(n2242) );
  OAI211_X1 U2971 ( .C1(n3950), .C2(n2243), .A(n2242), .B(n2170), .ZN(U3259)
         );
  NAND2_X1 U2972 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2448)
         );
  AND3_X2 U2973 ( .A1(n2684), .A2(n2168), .A3(n2681), .ZN(n3036) );
  NAND2_X1 U2974 ( .A1(n2251), .A2(n3035), .ZN(n3037) );
  INV_X2 U2975 ( .A(n3036), .ZN(n2251) );
  OAI22_X1 U2976 ( .A1(n3548), .A2(n2253), .B1(n2256), .B2(n2252), .ZN(n3398)
         );
  NAND2_X1 U2977 ( .A1(n3398), .A2(n4301), .ZN(n3118) );
  NAND2_X1 U2978 ( .A1(n2261), .A2(n4403), .ZN(n4720) );
  NAND2_X1 U2979 ( .A1(n4719), .A2(n4998), .ZN(n2260) );
  OAI21_X1 U2980 ( .B1(n3457), .B2(n2268), .A(n2266), .ZN(n3627) );
  OAI21_X1 U2981 ( .B1(n3457), .B2(n4303), .A(n4291), .ZN(n3531) );
  AOI21_X1 U2982 ( .B1(n4303), .B2(n4291), .A(n2270), .ZN(n2269) );
  NAND2_X1 U2983 ( .A1(n4433), .A2(n2273), .ZN(n2272) );
  NAND2_X1 U2984 ( .A1(n4433), .A2(n3143), .ZN(n2279) );
  AND2_X1 U2985 ( .A1(n2279), .A2(n4329), .ZN(n4421) );
  AND2_X4 U2986 ( .A1(n2282), .A2(n2655), .ZN(n3270) );
  NAND2_X1 U2987 ( .A1(n2651), .A2(n2652), .ZN(n2654) );
  MUX2_X1 U2988 ( .A(REG0_REG_29__SCAN_IN), .B(n2283), .S(n5013), .Z(U3515) );
  NAND2_X1 U2989 ( .A1(n3397), .A2(n2408), .ZN(n2288) );
  NAND2_X1 U2990 ( .A1(n2286), .A2(n2284), .ZN(n3456) );
  INV_X1 U2991 ( .A(n2285), .ZN(n2284) );
  OAI21_X1 U2992 ( .B1(n3067), .B2(n2153), .A(n3068), .ZN(n2285) );
  INV_X1 U2993 ( .A(n2153), .ZN(n2287) );
  NAND2_X1 U2994 ( .A1(n2289), .A2(n2290), .ZN(n4470) );
  NAND2_X1 U2995 ( .A1(n4513), .A2(n2291), .ZN(n2289) );
  INV_X1 U2996 ( .A(n2469), .ZN(n2297) );
  NAND3_X1 U2997 ( .A1(n2146), .A2(n2296), .A3(n2295), .ZN(n3962) );
  NAND2_X1 U2998 ( .A1(n3098), .A2(n2301), .ZN(n2298) );
  NAND2_X1 U2999 ( .A1(n3098), .A2(n3097), .ZN(n4432) );
  NAND2_X1 U3000 ( .A1(n2298), .A2(n2299), .ZN(n4410) );
  OAI21_X1 U3001 ( .B1(n3071), .B2(n2316), .A(n2313), .ZN(n3631) );
  AND2_X1 U3002 ( .A1(n3546), .A2(n2321), .ZN(n3469) );
  NAND2_X1 U3003 ( .A1(n4366), .A2(n4367), .ZN(n2324) );
  XNOR2_X1 U3004 ( .A(n2547), .B(n3449), .ZN(n4367) );
  XNOR2_X2 U3005 ( .A(n2455), .B(IR_REG_2__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U3006 ( .A1(n2323), .A2(n2546), .ZN(n4366) );
  INV_X1 U3007 ( .A(n2545), .ZN(n2323) );
  NAND2_X1 U3008 ( .A1(n2557), .A2(n4872), .ZN(n2332) );
  NAND2_X1 U3009 ( .A1(n2563), .A2(n4869), .ZN(n2338) );
  NAND2_X1 U3010 ( .A1(n4937), .A2(n2342), .ZN(n2341) );
  NAND2_X1 U3011 ( .A1(n4937), .A2(n4938), .ZN(n4936) );
  NAND2_X1 U3012 ( .A1(n4896), .A2(n2349), .ZN(n2347) );
  XNOR2_X1 U3013 ( .A(n2571), .B(n4978), .ZN(n4924) );
  INV_X1 U3014 ( .A(IR_REG_1__SCAN_IN), .ZN(n2353) );
  INV_X1 U3015 ( .A(IR_REG_2__SCAN_IN), .ZN(n2352) );
  NAND3_X1 U3016 ( .A1(n2354), .A2(n2353), .A3(n2352), .ZN(n2459) );
  NAND2_X1 U3017 ( .A1(n4163), .A2(n2357), .ZN(n2356) );
  NAND2_X1 U3018 ( .A1(n4163), .A2(n4161), .ZN(n2369) );
  NAND2_X1 U3019 ( .A1(n3439), .A2(n2373), .ZN(n2372) );
  NAND2_X1 U3020 ( .A1(n3326), .A2(n2169), .ZN(n2376) );
  NAND2_X1 U3021 ( .A1(n4024), .A2(n2985), .ZN(n4026) );
  NAND2_X1 U3022 ( .A1(n2380), .A2(n2383), .ZN(n4069) );
  NAND2_X1 U3023 ( .A1(n4024), .A2(n2381), .ZN(n2380) );
  NAND2_X1 U3024 ( .A1(n2424), .A2(n2130), .ZN(n2425) );
  OAI21_X1 U3025 ( .B1(n2897), .B2(n2389), .A(n2387), .ZN(n4151) );
  OR2_X2 U3026 ( .A1(n4443), .A2(n4439), .ZN(n4444) );
  NAND2_X1 U3027 ( .A1(n4482), .A2(n4462), .ZN(n4443) );
  NAND2_X1 U3028 ( .A1(n4452), .A2(n3096), .ZN(n3098) );
  INV_X1 U3029 ( .A(n2571), .ZN(n2572) );
  NAND2_X1 U3030 ( .A1(n3168), .A2(n3047), .ZN(n3481) );
  XNOR2_X1 U3031 ( .A(n2437), .B(IR_REG_26__SCAN_IN), .ZN(n2602) );
  INV_X1 U3032 ( .A(n2559), .ZN(n2560) );
  XNOR2_X1 U3033 ( .A(n2559), .B(n3284), .ZN(n3280) );
  AND2_X1 U3034 ( .A1(n3242), .A2(n2698), .ZN(n3251) );
  AND2_X1 U3035 ( .A1(n2135), .A2(DATAI_27_), .ZN(n4423) );
  OAI21_X1 U3036 ( .B1(n2135), .B2(n2552), .A(n2733), .ZN(n3046) );
  NAND2_X1 U3037 ( .A1(n2135), .A2(DATAI_4_), .ZN(n2733) );
  OAI21_X1 U3038 ( .B1(n2135), .B2(n2710), .A(n2709), .ZN(n3365) );
  NAND2_X1 U3039 ( .A1(n2135), .A2(DATAI_2_), .ZN(n2709) );
  NAND2_X1 U3040 ( .A1(n2135), .A2(DATAI_0_), .ZN(n2694) );
  OAI21_X1 U3041 ( .B1(n2138), .B2(n3230), .A(n2685), .ZN(n3035) );
  OAI21_X1 U3042 ( .B1(n2131), .B2(n2456), .A(n2457), .ZN(n4371) );
  NAND2_X1 U3043 ( .A1(n2645), .A2(n3301), .ZN(n4196) );
  OR2_X1 U3044 ( .A1(n3175), .A2(n3425), .ZN(n5019) );
  OR2_X1 U3045 ( .A1(n3262), .A2(n5020), .ZN(n2393) );
  AND2_X1 U3046 ( .A1(n4660), .A2(n4659), .ZN(n2394) );
  XOR2_X1 U3047 ( .A(n2603), .B(IR_REG_24__SCAN_IN), .Z(n2395) );
  NOR3_X1 U3048 ( .A1(n2883), .A2(n4079), .A3(n4080), .ZN(n2396) );
  AND2_X1 U3049 ( .A1(n4870), .A2(REG2_REG_9__SCAN_IN), .ZN(n2397) );
  AND2_X1 U3050 ( .A1(n4870), .A2(REG1_REG_9__SCAN_IN), .ZN(n2398) );
  AND2_X1 U3051 ( .A1(n4590), .A2(n2230), .ZN(n2399) );
  AND2_X1 U3052 ( .A1(n2460), .A2(n2410), .ZN(n2400) );
  INV_X1 U3053 ( .A(n4238), .ZN(n3038) );
  INV_X1 U3054 ( .A(n2574), .ZN(n4976) );
  NAND2_X1 U3055 ( .A1(n2978), .A2(n2977), .ZN(n4519) );
  INV_X1 U3056 ( .A(n4519), .ZN(n3093) );
  INV_X1 U3057 ( .A(IR_REG_29__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U3058 ( .A1(n3403), .A2(n3169), .ZN(n3610) );
  NAND2_X1 U3059 ( .A1(n4072), .A2(n4484), .ZN(n2402) );
  INV_X1 U3060 ( .A(n4458), .ZN(n4462) );
  OR2_X1 U3061 ( .A1(n4035), .A2(n4598), .ZN(n2403) );
  INV_X1 U3062 ( .A(n4211), .ZN(n3143) );
  NAND2_X1 U3063 ( .A1(n4681), .A2(n4680), .ZN(n2404) );
  NOR2_X1 U3064 ( .A1(n3130), .A2(n4568), .ZN(n2405) );
  AND2_X1 U3065 ( .A1(n4873), .A2(REG2_REG_5__SCAN_IN), .ZN(n2406) );
  INV_X1 U3066 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2860) );
  AND2_X1 U3067 ( .A1(n4498), .A2(n4115), .ZN(n2407) );
  AND2_X1 U3068 ( .A1(n4249), .A2(n3065), .ZN(n2408) );
  AND2_X1 U3069 ( .A1(n3156), .A2(n4859), .ZN(n4696) );
  NAND2_X1 U3070 ( .A1(n2671), .A2(n2670), .ZN(n4268) );
  AND2_X1 U3071 ( .A1(n4222), .A2(n3144), .ZN(n4661) );
  INV_X1 U3072 ( .A(n4661), .ZN(n3145) );
  XNOR2_X1 U3073 ( .A(n2549), .B(n3213), .ZN(n3211) );
  NAND2_X1 U3074 ( .A1(n3123), .A2(n4355), .ZN(n2409) );
  NAND2_X1 U3075 ( .A1(n3604), .A2(n3616), .ZN(n3065) );
  INV_X1 U3076 ( .A(n4502), .ZN(n3092) );
  AND2_X1 U3077 ( .A1(n3124), .A2(n4690), .ZN(n4310) );
  AND2_X1 U3078 ( .A1(n4225), .A2(n4472), .ZN(n4325) );
  INV_X1 U3079 ( .A(IR_REG_5__SCAN_IN), .ZN(n3668) );
  NAND2_X1 U3080 ( .A1(n2138), .A2(DATAI_1_), .ZN(n2685) );
  NAND2_X1 U3081 ( .A1(n4876), .A2(REG2_REG_1__SCAN_IN), .ZN(n2546) );
  NAND2_X1 U3082 ( .A1(n4868), .A2(REG1_REG_11__SCAN_IN), .ZN(n2499) );
  INV_X1 U3083 ( .A(n3936), .ZN(n2515) );
  NAND2_X1 U3084 ( .A1(n4117), .A2(n4462), .ZN(n3096) );
  INV_X1 U3085 ( .A(IR_REG_26__SCAN_IN), .ZN(n2584) );
  INV_X1 U3086 ( .A(IR_REG_21__SCAN_IN), .ZN(n2432) );
  INV_X1 U3087 ( .A(n3594), .ZN(n2796) );
  INV_X1 U3088 ( .A(n3520), .ZN(n2775) );
  NAND2_X1 U3089 ( .A1(n2135), .A2(n2743), .ZN(n2744) );
  INV_X1 U3090 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3906) );
  OR2_X1 U3091 ( .A1(n2435), .A2(IR_REG_22__SCAN_IN), .ZN(n2419) );
  OR2_X1 U3092 ( .A1(n4871), .A2(REG1_REG_7__SCAN_IN), .ZN(n2477) );
  INV_X1 U3093 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4113) );
  NAND2_X1 U3094 ( .A1(n3419), .A2(n2499), .ZN(n2514) );
  NAND2_X1 U3095 ( .A1(n4976), .A2(n3896), .ZN(n2537) );
  NOR2_X1 U3096 ( .A1(n3155), .A2(n3158), .ZN(n3159) );
  INV_X1 U3097 ( .A(n2135), .ZN(n2854) );
  NAND2_X1 U3098 ( .A1(n4151), .A2(n2971), .ZN(n4024) );
  AOI21_X1 U3099 ( .B1(n2823), .B2(n3551), .A(n2711), .ZN(n2718) );
  NOR2_X1 U3100 ( .A1(n3427), .A2(n3425), .ZN(n3031) );
  INV_X1 U3101 ( .A(n3270), .ZN(n3277) );
  OR2_X1 U3102 ( .A1(n4506), .A2(n2281), .ZN(n2978) );
  NAND2_X1 U3103 ( .A1(n2448), .A2(IR_REG_1__SCAN_IN), .ZN(n2450) );
  INV_X1 U3104 ( .A(n4859), .ZN(n3154) );
  AND2_X1 U3105 ( .A1(n4402), .A2(n4401), .ZN(n4403) );
  INV_X1 U3106 ( .A(n4268), .ZN(n4442) );
  INV_X1 U3107 ( .A(n4351), .ZN(n4536) );
  AND2_X1 U3108 ( .A1(n4637), .A2(n4636), .ZN(n4681) );
  OR2_X1 U3109 ( .A1(n3188), .A2(D_REG_0__SCAN_IN), .ZN(n2626) );
  AND2_X1 U3110 ( .A1(n2138), .A2(DATAI_20_), .ZN(n4559) );
  INV_X1 U3111 ( .A(n4673), .ZN(n4683) );
  INV_X1 U3112 ( .A(n3539), .ZN(n3644) );
  NAND2_X1 U3113 ( .A1(n3156), .A2(n3154), .ZN(n4654) );
  NOR2_X1 U3114 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  OR2_X1 U3115 ( .A1(n2489), .A2(IR_REG_9__SCAN_IN), .ZN(n2494) );
  AND2_X1 U3116 ( .A1(n2666), .A2(n3103), .ZN(n4418) );
  AND2_X1 U3117 ( .A1(n3997), .A2(n4102), .ZN(n3998) );
  NAND2_X1 U3118 ( .A1(n2676), .A2(n4649), .ZN(n4191) );
  OAI21_X1 U3119 ( .B1(n2718), .B2(n2717), .A(n2721), .ZN(n3312) );
  XNOR2_X1 U3120 ( .A(n2604), .B(n2603), .ZN(n2638) );
  INV_X1 U3121 ( .A(n4622), .ZN(n4590) );
  AND4_X1 U3122 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3053)
         );
  INV_X1 U3123 ( .A(n4980), .ZN(n4901) );
  AOI21_X1 U3124 ( .B1(n3950), .B2(n3949), .A(n4908), .ZN(n3955) );
  OR2_X1 U3125 ( .A1(n3165), .A2(n2622), .ZN(n3427) );
  INV_X1 U3126 ( .A(n4089), .ZN(n4631) );
  AND2_X1 U3127 ( .A1(n4955), .A2(n3488), .ZN(n4688) );
  AND2_X1 U3128 ( .A1(n4955), .A2(n3428), .ZN(n4952) );
  NAND2_X1 U3129 ( .A1(n2626), .A2(n2625), .ZN(n3425) );
  INV_X1 U3130 ( .A(n4787), .ZN(n5005) );
  NAND2_X1 U3131 ( .A1(n4704), .A2(n4987), .ZN(n4787) );
  INV_X1 U3132 ( .A(n3162), .ZN(n3302) );
  XNOR2_X1 U3133 ( .A(n2482), .B(n2481), .ZN(n3284) );
  AND2_X1 U3134 ( .A1(n2591), .A2(n2590), .ZN(n4930) );
  NOR2_X1 U3135 ( .A1(n3985), .A2(n3984), .ZN(n4009) );
  INV_X1 U3136 ( .A(n4196), .ZN(n4108) );
  INV_X1 U3137 ( .A(n4102), .ZN(n4199) );
  INV_X1 U3138 ( .A(n4207), .ZN(n4349) );
  NAND2_X1 U3139 ( .A1(n2963), .A2(n2962), .ZN(n4351) );
  OAI211_X1 U3140 ( .C1(n4632), .C2(n2281), .A(n2853), .B(n2852), .ZN(n4608)
         );
  INV_X1 U3141 ( .A(n4940), .ZN(n4905) );
  INV_X1 U3142 ( .A(n4930), .ZN(n4918) );
  INV_X1 U3143 ( .A(n4688), .ZN(n4670) );
  NAND2_X1 U3144 ( .A1(n5022), .A2(n4998), .ZN(n4794) );
  INV_X2 U3145 ( .A(n5019), .ZN(n5022) );
  OR2_X1 U3146 ( .A1(n4010), .A2(n4856), .ZN(n3179) );
  NAND2_X1 U3147 ( .A1(n5013), .A2(n4998), .ZN(n4856) );
  OR2_X1 U31480 ( .A1(n3175), .A2(n3174), .ZN(n5011) );
  INV_X2 U31490 ( .A(n5011), .ZN(n5013) );
  INV_X1 U3150 ( .A(n4972), .ZN(n4971) );
  AND2_X1 U3151 ( .A1(n2587), .A2(n2647), .ZN(n4859) );
  INV_X1 U3152 ( .A(n4341), .ZN(n4864) );
  OR2_X1 U3153 ( .A1(n2521), .A2(n2520), .ZN(n4980) );
  OAI211_X1 U3154 ( .C1(n3034), .C2(n4108), .A(n3033), .B(n2148), .ZN(U3237)
         );
  INV_X2 U3155 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3156 ( .A(n2459), .ZN(n2411) );
  NAND2_X1 U3157 ( .A1(n2411), .A2(n2400), .ZN(n2469) );
  NAND4_X1 U3158 ( .A1(n2485), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n2507)
         );
  NAND4_X1 U3159 ( .A1(n3668), .A2(n2525), .A3(n2518), .A4(n2529), .ZN(n2415)
         );
  NAND2_X1 U3160 ( .A1(n2424), .A2(n2416), .ZN(n2532) );
  NAND3_X1 U3161 ( .A1(n3791), .A2(n2417), .A3(n2630), .ZN(n2418) );
  NOR2_X2 U3162 ( .A1(n2532), .A2(n2418), .ZN(n2429) );
  NOR2_X1 U3163 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2423)
         );
  NAND2_X1 U3164 ( .A1(n2425), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  OR2_X1 U3165 ( .A1(n2638), .A2(U3149), .ZN(n4347) );
  NAND2_X1 U3166 ( .A1(n3162), .A2(n4347), .ZN(n2590) );
  NAND2_X1 U3167 ( .A1(n2435), .A2(IR_REG_31__SCAN_IN), .ZN(n2428) );
  INV_X1 U3168 ( .A(n2429), .ZN(n2430) );
  NAND2_X1 U3169 ( .A1(n2430), .A2(IR_REG_31__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3170 ( .A1(n2431), .A2(IR_REG_21__SCAN_IN), .ZN(n2434) );
  NAND2_X1 U3171 ( .A1(n2434), .A2(n2433), .ZN(n2436) );
  AND2_X2 U3172 ( .A1(n2436), .A2(n2435), .ZN(n4277) );
  INV_X1 U3173 ( .A(n2437), .ZN(n2438) );
  NAND2_X1 U3174 ( .A1(n2438), .A2(n2585), .ZN(n2445) );
  INV_X1 U3175 ( .A(n2446), .ZN(n2443) );
  NOR2_X1 U3176 ( .A1(n2585), .A2(IR_REG_26__SCAN_IN), .ZN(n2442) );
  NAND3_X1 U3177 ( .A1(n2585), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_26__SCAN_IN), .ZN(n2440) );
  OAI211_X1 U3178 ( .C1(IR_REG_31__SCAN_IN), .C2(n2585), .A(n2440), .B(n2439), 
        .ZN(n2441) );
  AOI21_X1 U3179 ( .B1(n3156), .B2(n2638), .A(n2854), .ZN(n2589) );
  OAI21_X1 U3180 ( .B1(n2446), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2447) );
  XNOR2_X1 U3181 ( .A(n2447), .B(IR_REG_27__SCAN_IN), .ZN(n4860) );
  INV_X1 U3182 ( .A(n4860), .ZN(n4359) );
  INV_X1 U3183 ( .A(n2454), .ZN(n2451) );
  AND2_X1 U3184 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3222)
         );
  INV_X1 U3185 ( .A(n3230), .ZN(n4876) );
  NAND2_X1 U3186 ( .A1(n4876), .A2(REG1_REG_1__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3187 ( .A1(n2453), .A2(n2452), .ZN(n4370) );
  INV_X1 U3188 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2456) );
  NAND2_X1 U3189 ( .A1(n2131), .A2(n2456), .ZN(n2457) );
  NAND2_X1 U3190 ( .A1(n4370), .A2(n4371), .ZN(n4369) );
  NAND2_X1 U3191 ( .A1(n2131), .A2(REG1_REG_2__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3192 ( .A1(n2459), .A2(IR_REG_31__SCAN_IN), .ZN(n2461) );
  NAND2_X1 U3193 ( .A1(n2461), .A2(n2460), .ZN(n2466) );
  OR2_X1 U3194 ( .A1(n2461), .A2(n2460), .ZN(n2462) );
  NAND2_X1 U3195 ( .A1(n3210), .A2(REG1_REG_3__SCAN_IN), .ZN(n2465) );
  NAND2_X1 U3196 ( .A1(n2463), .A2(n4874), .ZN(n2464) );
  NAND2_X2 U3197 ( .A1(n2465), .A2(n2464), .ZN(n2468) );
  NAND2_X1 U3198 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2467) );
  XNOR2_X1 U3199 ( .A(n2467), .B(IR_REG_4__SCAN_IN), .ZN(n4884) );
  INV_X1 U3200 ( .A(n4884), .ZN(n2552) );
  XNOR2_X2 U3201 ( .A(n2468), .B(n2552), .ZN(n4879) );
  INV_X1 U3202 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5017) );
  INV_X1 U3203 ( .A(n2509), .ZN(n2472) );
  NAND2_X1 U3204 ( .A1(n2469), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  MUX2_X1 U3205 ( .A(IR_REG_31__SCAN_IN), .B(n2470), .S(IR_REG_5__SCAN_IN), 
        .Z(n2471) );
  NAND2_X1 U3206 ( .A1(n2472), .A2(n2471), .ZN(n3237) );
  MUX2_X1 U3207 ( .A(REG1_REG_5__SCAN_IN), .B(n5017), .S(n3237), .Z(n3231) );
  INV_X1 U3208 ( .A(n3237), .ZN(n4873) );
  OR2_X1 U3209 ( .A1(n2509), .A2(n2517), .ZN(n2473) );
  INV_X1 U32100 ( .A(n2474), .ZN(n2475) );
  NAND2_X1 U32110 ( .A1(n2509), .A2(n2476), .ZN(n2487) );
  NAND2_X1 U32120 ( .A1(n2487), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  INV_X1 U32130 ( .A(n4871), .ZN(n3262) );
  INV_X1 U32140 ( .A(REG1_REG_7__SCAN_IN), .ZN(n5020) );
  INV_X1 U32150 ( .A(n2483), .ZN(n2484) );
  INV_X1 U32160 ( .A(IR_REG_7__SCAN_IN), .ZN(n2478) );
  NAND2_X1 U32170 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  NAND2_X1 U32180 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2482) );
  INV_X1 U32190 ( .A(IR_REG_8__SCAN_IN), .ZN(n2481) );
  INV_X1 U32200 ( .A(n3284), .ZN(n2558) );
  INV_X1 U32210 ( .A(n2485), .ZN(n2486) );
  NAND2_X1 U32220 ( .A1(n2489), .A2(IR_REG_31__SCAN_IN), .ZN(n2488) );
  MUX2_X1 U32230 ( .A(IR_REG_31__SCAN_IN), .B(n2488), .S(IR_REG_9__SCAN_IN), 
        .Z(n2490) );
  NAND2_X1 U32240 ( .A1(n2490), .A2(n2494), .ZN(n3347) );
  XOR2_X1 U32250 ( .A(REG1_REG_9__SCAN_IN), .B(n3347), .Z(n3349) );
  INV_X1 U32260 ( .A(n3347), .ZN(n4870) );
  NAND2_X1 U32270 ( .A1(n2494), .A2(IR_REG_31__SCAN_IN), .ZN(n2491) );
  OR2_X1 U32280 ( .A1(n2492), .A2(n2200), .ZN(n2493) );
  INV_X1 U32290 ( .A(n2494), .ZN(n2496) );
  INV_X1 U32300 ( .A(IR_REG_10__SCAN_IN), .ZN(n2495) );
  NAND2_X1 U32310 ( .A1(n2496), .A2(n2495), .ZN(n2502) );
  NAND2_X1 U32320 ( .A1(n2502), .A2(IR_REG_31__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U32330 ( .A1(n2497), .A2(n3669), .ZN(n2500) );
  OR2_X1 U32340 ( .A1(n2497), .A2(n3669), .ZN(n2498) );
  XOR2_X1 U32350 ( .A(REG1_REG_11__SCAN_IN), .B(n4868), .Z(n3420) );
  NAND2_X1 U32360 ( .A1(n3421), .A2(n3420), .ZN(n3419) );
  INV_X1 U32370 ( .A(n4868), .ZN(n3416) );
  INV_X1 U32380 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U32390 ( .A1(n2500), .A2(IR_REG_31__SCAN_IN), .ZN(n2501) );
  INV_X1 U32400 ( .A(n4867), .ZN(n2564) );
  INV_X1 U32410 ( .A(n2502), .ZN(n2504) );
  NOR2_X1 U32420 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2503) );
  AOI21_X1 U32430 ( .B1(n2504), .B2(n2503), .A(n2517), .ZN(n2505) );
  MUX2_X1 U32440 ( .A(n2517), .B(n2505), .S(IR_REG_13__SCAN_IN), .Z(n2506) );
  INV_X1 U32450 ( .A(n2507), .ZN(n2508) );
  AND2_X1 U32460 ( .A1(n2509), .A2(n2508), .ZN(n2519) );
  INV_X1 U32470 ( .A(n2519), .ZN(n2510) );
  INV_X1 U32480 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4783) );
  XNOR2_X1 U32490 ( .A(n3945), .B(n4783), .ZN(n3939) );
  INV_X1 U32500 ( .A(n3939), .ZN(n2512) );
  AND2_X1 U32510 ( .A1(REG1_REG_12__SCAN_IN), .A2(n2512), .ZN(n2513) );
  NAND2_X1 U32520 ( .A1(n2514), .A2(n4867), .ZN(n3936) );
  NOR2_X1 U32530 ( .A1(n2519), .A2(n2517), .ZN(n2516) );
  MUX2_X1 U32540 ( .A(n2517), .B(n2516), .S(IR_REG_14__SCAN_IN), .Z(n2521) );
  NAND2_X1 U32550 ( .A1(n2519), .A2(n2518), .ZN(n2524) );
  INV_X1 U32560 ( .A(n2524), .ZN(n2520) );
  INV_X1 U32570 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4895) );
  NOR2_X1 U32580 ( .A1(n2522), .A2(n4980), .ZN(n2523) );
  NAND2_X1 U32590 ( .A1(n2524), .A2(IR_REG_31__SCAN_IN), .ZN(n2526) );
  NAND2_X1 U32600 ( .A1(n2526), .A2(n2525), .ZN(n2528) );
  OR2_X1 U32610 ( .A1(n2526), .A2(n2525), .ZN(n2527) );
  XNOR2_X1 U32620 ( .A(n4913), .B(REG1_REG_15__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U32630 ( .A1(n2528), .A2(IR_REG_31__SCAN_IN), .ZN(n2530) );
  XNOR2_X1 U32640 ( .A(n2530), .B(n2529), .ZN(n4978) );
  NAND2_X1 U32650 ( .A1(n2531), .A2(n4978), .ZN(n4932) );
  NAND2_X1 U32660 ( .A1(n2586), .A2(IR_REG_31__SCAN_IN), .ZN(n2533) );
  MUX2_X1 U32670 ( .A(IR_REG_31__SCAN_IN), .B(n2533), .S(IR_REG_17__SCAN_IN), 
        .Z(n2534) );
  AND2_X1 U32680 ( .A1(n2532), .A2(n2534), .ZN(n2574) );
  INV_X1 U32690 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U32700 ( .A1(n2574), .A2(REG1_REG_17__SCAN_IN), .B1(n3896), .B2(
        n4976), .ZN(n4935) );
  INV_X1 U32710 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4920) );
  AND2_X1 U32720 ( .A1(n4920), .A2(n4935), .ZN(n2536) );
  NAND2_X1 U32730 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2538) );
  XNOR2_X1 U32740 ( .A(n2538), .B(IR_REG_18__SCAN_IN), .ZN(n4865) );
  NAND2_X1 U32750 ( .A1(n4865), .A2(REG1_REG_18__SCAN_IN), .ZN(n2539) );
  OAI21_X1 U32760 ( .B1(n4865), .B2(REG1_REG_18__SCAN_IN), .A(n2539), .ZN(
        n3949) );
  INV_X1 U32770 ( .A(n2539), .ZN(n2540) );
  NAND2_X1 U32780 ( .A1(n2541), .A2(n3791), .ZN(n2629) );
  OR2_X1 U32790 ( .A1(n2541), .A2(n3791), .ZN(n2542) );
  XNOR2_X1 U32800 ( .A(n4864), .B(REG1_REG_19__SCAN_IN), .ZN(n2543) );
  INV_X1 U32810 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U32820 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(
        n3224) );
  AOI21_X1 U32830 ( .B1(n3230), .B2(n2544), .A(n3224), .ZN(n2545) );
  INV_X1 U32840 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3449) );
  NAND2_X1 U32850 ( .A1(n2131), .A2(REG2_REG_2__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32860 ( .A1(n3211), .A2(REG2_REG_3__SCAN_IN), .ZN(n2551) );
  NAND2_X1 U32870 ( .A1(n2549), .A2(n4874), .ZN(n2550) );
  INV_X1 U32880 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2555) );
  MUX2_X1 U32890 ( .A(REG2_REG_5__SCAN_IN), .B(n2555), .S(n3237), .Z(n3235) );
  INV_X1 U32900 ( .A(n2556), .ZN(n2557) );
  INV_X1 U32910 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3615) );
  MUX2_X1 U32920 ( .A(n3615), .B(REG2_REG_7__SCAN_IN), .S(n4871), .Z(n3264) );
  INV_X1 U32930 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3493) );
  XNOR2_X1 U32940 ( .A(n3347), .B(REG2_REG_9__SCAN_IN), .ZN(n3344) );
  INV_X1 U32950 ( .A(n2562), .ZN(n2563) );
  INV_X1 U32960 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3854) );
  MUX2_X1 U32970 ( .A(n3854), .B(REG2_REG_11__SCAN_IN), .S(n4868), .Z(n3413)
         );
  NAND2_X1 U32980 ( .A1(n3650), .A2(REG2_REG_12__SCAN_IN), .ZN(n2567) );
  INV_X1 U32990 ( .A(n3945), .ZN(n4866) );
  INV_X1 U33000 ( .A(REG2_REG_13__SCAN_IN), .ZN(n2568) );
  INV_X1 U33010 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4898) );
  NOR2_X1 U33020 ( .A1(n2569), .A2(n4980), .ZN(n2570) );
  XNOR2_X1 U33030 ( .A(n4913), .B(REG2_REG_15__SCAN_IN), .ZN(n4906) );
  INV_X1 U33040 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U33050 ( .A1(n2572), .A2(n4978), .ZN(n2573) );
  NOR2_X1 U33060 ( .A1(n2574), .A2(REG2_REG_17__SCAN_IN), .ZN(n2575) );
  AOI21_X1 U33070 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2574), .A(n2575), .ZN(
        n4938) );
  INV_X1 U33080 ( .A(n2575), .ZN(n2576) );
  XNOR2_X1 U33090 ( .A(n4865), .B(REG2_REG_18__SCAN_IN), .ZN(n3947) );
  XNOR2_X1 U33100 ( .A(n4341), .B(REG2_REG_19__SCAN_IN), .ZN(n2578) );
  XNOR2_X1 U33110 ( .A(n2579), .B(n2578), .ZN(n2588) );
  OR3_X1 U33120 ( .A1(n2446), .A2(IR_REG_27__SCAN_IN), .A3(IR_REG_26__SCAN_IN), 
        .ZN(n2580) );
  NAND2_X1 U33130 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  MUX2_X1 U33140 ( .A(IR_REG_31__SCAN_IN), .B(n2581), .S(IR_REG_28__SCAN_IN), 
        .Z(n2587) );
  AND2_X1 U33150 ( .A1(n4859), .A2(n4860), .ZN(n4360) );
  NAND2_X1 U33160 ( .A1(n2588), .A2(n4940), .ZN(n2595) );
  NAND2_X1 U33170 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4036) );
  INV_X1 U33180 ( .A(n2589), .ZN(n2591) );
  NAND2_X1 U33190 ( .A1(n4930), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2592) );
  OAI211_X1 U33200 ( .C1(n4945), .C2(n4341), .A(n4036), .B(n2592), .ZN(n2593)
         );
  INV_X1 U33210 ( .A(n2593), .ZN(n2594) );
  XNOR2_X1 U33220 ( .A(n2665), .B(REG3_REG_26__SCAN_IN), .ZN(n4447) );
  INV_X1 U33230 ( .A(n4447), .ZN(n3034) );
  NAND2_X1 U33240 ( .A1(n2604), .A2(n2603), .ZN(n2605) );
  NAND3_X1 U33250 ( .A1(n2624), .A2(B_REG_SCAN_IN), .A3(n4861), .ZN(n2610) );
  INV_X1 U33260 ( .A(B_REG_SCAN_IN), .ZN(n2608) );
  NAND2_X1 U33270 ( .A1(n3193), .A2(n2608), .ZN(n2609) );
  OR2_X1 U33280 ( .A1(n3188), .A2(D_REG_1__SCAN_IN), .ZN(n2611) );
  INV_X1 U33290 ( .A(n2602), .ZN(n2623) );
  NAND2_X1 U33300 ( .A1(n2623), .A2(n4861), .ZN(n3189) );
  NAND2_X1 U33310 ( .A1(n2611), .A2(n3189), .ZN(n3165) );
  INV_X1 U33320 ( .A(D_REG_20__SCAN_IN), .ZN(n4964) );
  INV_X1 U33330 ( .A(D_REG_22__SCAN_IN), .ZN(n4962) );
  INV_X1 U33340 ( .A(D_REG_27__SCAN_IN), .ZN(n4959) );
  INV_X1 U33350 ( .A(D_REG_17__SCAN_IN), .ZN(n4965) );
  NAND4_X1 U33360 ( .A1(n4964), .A2(n4962), .A3(n4959), .A4(n4965), .ZN(n2617)
         );
  NOR4_X1 U33370 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_6__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n2615) );
  NOR4_X1 U33380 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_13__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2614) );
  NOR4_X1 U33390 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_18__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2613) );
  NOR4_X1 U33400 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2612) );
  NAND4_X1 U33410 ( .A1(n2615), .A2(n2614), .A3(n2613), .A4(n2612), .ZN(n2616)
         );
  NOR4_X1 U33420 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(n2617), 
        .A4(n2616), .ZN(n2620) );
  NOR4_X1 U33430 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2619) );
  NOR4_X1 U33440 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2618) );
  AND2_X1 U33450 ( .A1(n2619), .A2(n2618), .ZN(n3700) );
  AND2_X1 U33460 ( .A1(n2620), .A2(n3700), .ZN(n2621) );
  INV_X1 U33470 ( .A(n3164), .ZN(n2622) );
  NAND2_X1 U33480 ( .A1(n2624), .A2(n2623), .ZN(n2625) );
  INV_X1 U33490 ( .A(n3031), .ZN(n2644) );
  INV_X1 U33500 ( .A(n3156), .ZN(n2628) );
  INV_X1 U33510 ( .A(n4345), .ZN(n2674) );
  INV_X1 U33520 ( .A(n4277), .ZN(n2675) );
  NAND2_X1 U3353 ( .A1(n3218), .A2(n4864), .ZN(n2627) );
  NAND2_X1 U33540 ( .A1(n2628), .A2(n2627), .ZN(n2633) );
  BUF_X1 U3355 ( .A(n2640), .Z(n2632) );
  INV_X1 U3356 ( .A(n2632), .ZN(n4863) );
  NAND2_X1 U3357 ( .A1(n3029), .A2(n4700), .ZN(n2634) );
  NAND2_X1 U3358 ( .A1(n2644), .A2(n2634), .ZN(n2637) );
  NAND2_X1 U3359 ( .A1(n2632), .A2(n4341), .ZN(n2635) );
  INV_X1 U3360 ( .A(n3161), .ZN(n2636) );
  NAND2_X1 U3361 ( .A1(n2637), .A2(n2636), .ZN(n3300) );
  NAND2_X1 U3362 ( .A1(n2641), .A2(n2638), .ZN(n2639) );
  OAI21_X1 U3363 ( .B1(n3300), .B2(n2639), .A(STATE_REG_SCAN_IN), .ZN(n2645)
         );
  NAND2_X1 U3364 ( .A1(n4345), .A2(n4341), .ZN(n2687) );
  NOR2_X1 U3365 ( .A1(n4973), .A2(n2687), .ZN(n2643) );
  NAND2_X1 U3366 ( .A1(n2643), .A2(n2141), .ZN(n2672) );
  INV_X1 U3367 ( .A(n2672), .ZN(n4343) );
  NAND2_X1 U3368 ( .A1(n2644), .A2(n4343), .ZN(n3301) );
  INV_X1 U3369 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4071) );
  NAND2_X1 U3370 ( .A1(n2991), .A2(n4071), .ZN(n2646) );
  NAND2_X1 U3371 ( .A1(n2665), .A2(n2646), .ZN(n4465) );
  INV_X1 U3372 ( .A(n3962), .ZN(n2650) );
  XNOR2_X2 U3373 ( .A(n2653), .B(n3959), .ZN(n2655) );
  INV_X1 U3374 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U3375 ( .A1(n3270), .A2(REG1_REG_25__SCAN_IN), .ZN(n2657) );
  NAND2_X1 U3376 ( .A1(n2732), .A2(REG0_REG_25__SCAN_IN), .ZN(n2656) );
  OAI211_X1 U3377 ( .C1(n3150), .C2(n4464), .A(n2657), .B(n2656), .ZN(n2658)
         );
  INV_X1 U3378 ( .A(n2658), .ZN(n2659) );
  NOR2_X1 U3379 ( .A1(n2672), .A2(n3154), .ZN(n2661) );
  NAND2_X1 U3380 ( .A1(n3031), .A2(n2661), .ZN(n4169) );
  INV_X1 U3381 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2663) );
  INV_X1 U3382 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2662) );
  OAI21_X1 U3383 ( .B1(n2665), .B2(n2663), .A(n2662), .ZN(n2666) );
  NAND2_X1 U3384 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2664) );
  NAND2_X1 U3385 ( .A1(n4418), .A2(n3014), .ZN(n2671) );
  INV_X1 U3386 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U3387 ( .A1(n3270), .A2(REG1_REG_27__SCAN_IN), .ZN(n2668) );
  NAND2_X1 U3388 ( .A1(n2137), .A2(REG2_REG_27__SCAN_IN), .ZN(n2667) );
  OAI211_X1 U3389 ( .C1(n2680), .C2(n3866), .A(n2668), .B(n2667), .ZN(n2669)
         );
  INV_X1 U3390 ( .A(n2669), .ZN(n2670) );
  NOR2_X1 U3391 ( .A1(n2672), .A2(n4859), .ZN(n2673) );
  NAND2_X1 U3392 ( .A1(n4268), .A2(n4165), .ZN(n2678) );
  NAND3_X1 U3393 ( .A1(n3031), .A2(n4672), .A3(n3302), .ZN(n2676) );
  AND2_X1 U3394 ( .A1(n2632), .A2(n4864), .ZN(n4946) );
  NAND2_X1 U3395 ( .A1(n4995), .A2(n2675), .ZN(n3163) );
  NAND2_X1 U3396 ( .A1(n2138), .A2(DATAI_26_), .ZN(n4445) );
  AOI22_X1 U3397 ( .A1(n4191), .A2(n4439), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n2677) );
  OAI211_X1 U3398 ( .C1(n4117), .C2(n4169), .A(n2678), .B(n2677), .ZN(n2679)
         );
  INV_X1 U3399 ( .A(n2679), .ZN(n3033) );
  NAND2_X1 U3400 ( .A1(n3270), .A2(REG1_REG_1__SCAN_IN), .ZN(n2684) );
  NAND2_X1 U3401 ( .A1(n2139), .A2(REG0_REG_1__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3402 ( .A1(n2875), .A2(REG2_REG_1__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3403 ( .A1(n2769), .A2(REG3_REG_1__SCAN_IN), .ZN(n2681) );
  NAND2_X4 U3404 ( .A1(n2641), .A2(n2686), .ZN(n3989) );
  XNOR2_X1 U3405 ( .A(n2688), .B(n3976), .ZN(n2704) );
  OR2_X4 U3406 ( .A1(n4998), .A2(n3989), .ZN(n2730) );
  XNOR2_X1 U3407 ( .A(n2704), .B(n2705), .ZN(n3299) );
  NAND2_X1 U3408 ( .A1(n3270), .A2(REG1_REG_0__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3409 ( .A1(n2769), .A2(REG3_REG_0__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3410 ( .A1(n2136), .A2(REG2_REG_0__SCAN_IN), .ZN(n2689) );
  AND3_X1 U3411 ( .A1(n2691), .A2(n2690), .A3(n2689), .ZN(n2693) );
  NAND2_X1 U3412 ( .A1(n2732), .A2(REG0_REG_0__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3413 ( .A1(n2141), .A2(n2698), .ZN(n2696) );
  NAND2_X1 U3414 ( .A1(n2726), .A2(n3242), .ZN(n2695) );
  AND2_X1 U3415 ( .A1(n2696), .A2(n2695), .ZN(n2701) );
  NAND2_X1 U3416 ( .A1(n2699), .A2(REG1_REG_0__SCAN_IN), .ZN(n2697) );
  NAND2_X1 U3417 ( .A1(n2701), .A2(n2697), .ZN(n3964) );
  INV_X1 U3418 ( .A(n2698), .ZN(n3111) );
  AOI22_X1 U3419 ( .A1(n2140), .A2(n3242), .B1(IR_REG_0__SCAN_IN), .B2(n2699), 
        .ZN(n2700) );
  OAI21_X1 U3420 ( .B1(n2730), .B2(n3111), .A(n2700), .ZN(n3965) );
  NAND2_X1 U3421 ( .A1(n3964), .A2(n3965), .ZN(n2703) );
  NAND2_X1 U3422 ( .A1(n2701), .A2(n3976), .ZN(n2702) );
  NAND2_X1 U3423 ( .A1(n2703), .A2(n2702), .ZN(n3298) );
  NAND2_X1 U3424 ( .A1(n3299), .A2(n3298), .ZN(n2708) );
  INV_X1 U3425 ( .A(n2704), .ZN(n2706) );
  NAND2_X1 U3426 ( .A1(n2706), .A2(n2705), .ZN(n2707) );
  NAND2_X1 U3427 ( .A1(n2708), .A2(n2707), .ZN(n3309) );
  INV_X1 U3428 ( .A(n3309), .ZN(n2720) );
  NAND2_X1 U3429 ( .A1(n2769), .A2(REG3_REG_2__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3430 ( .A1(n3270), .A2(REG1_REG_2__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U3431 ( .A1(n2137), .A2(REG2_REG_2__SCAN_IN), .ZN(n2713) );
  INV_X1 U3432 ( .A(n2131), .ZN(n2710) );
  NOR2_X1 U3433 ( .A1(n3374), .A2(n2133), .ZN(n2711) );
  AND4_X1 U3434 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2712), .ZN(n3248)
         );
  OAI22_X1 U3435 ( .A1(n3248), .A2(n2133), .B1(n3374), .B2(n3989), .ZN(n2716)
         );
  XNOR2_X1 U3436 ( .A(n2716), .B(n3976), .ZN(n2717) );
  NAND2_X1 U3437 ( .A1(n2717), .A2(n2718), .ZN(n2721) );
  INV_X1 U3438 ( .A(n3312), .ZN(n2719) );
  NAND2_X1 U3439 ( .A1(n2720), .A2(n2719), .ZN(n3310) );
  NAND2_X1 U3440 ( .A1(n3310), .A2(n2721), .ZN(n3355) );
  NAND2_X1 U3441 ( .A1(n3270), .A2(REG1_REG_3__SCAN_IN), .ZN(n2725) );
  INV_X1 U3442 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3556) );
  NAND2_X1 U3443 ( .A1(n2769), .A2(n3556), .ZN(n2724) );
  NAND2_X1 U3444 ( .A1(n2137), .A2(REG2_REG_3__SCAN_IN), .ZN(n2723) );
  NAND2_X1 U3445 ( .A1(n2732), .A2(REG0_REG_3__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3446 ( .A1(n3973), .A2(n3475), .ZN(n2728) );
  MUX2_X1 U3447 ( .A(n4874), .B(DATAI_3_), .S(n2135), .Z(n3550) );
  NAND2_X1 U3448 ( .A1(n2726), .A2(n3550), .ZN(n2727) );
  NAND2_X1 U3449 ( .A1(n2728), .A2(n2727), .ZN(n2729) );
  XNOR2_X1 U3450 ( .A(n2729), .B(n3976), .ZN(n2736) );
  OAI22_X1 U3451 ( .A1(n2730), .A2(n3367), .B1(n3047), .B2(n2134), .ZN(n2735)
         );
  XNOR2_X1 U3452 ( .A(n2736), .B(n2735), .ZN(n3356) );
  NAND2_X1 U3453 ( .A1(n3355), .A2(n3356), .ZN(n3326) );
  NAND2_X1 U3454 ( .A1(n3270), .A2(REG1_REG_4__SCAN_IN), .ZN(n3045) );
  INV_X1 U3455 ( .A(REG3_REG_4__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U3456 ( .A1(n3663), .A2(n3556), .ZN(n2731) );
  AND2_X1 U3457 ( .A1(n2731), .A2(n2751), .ZN(n3483) );
  NAND2_X1 U34580 ( .A1(n2769), .A2(n3483), .ZN(n3044) );
  NAND2_X1 U34590 ( .A1(n2137), .A2(REG2_REG_4__SCAN_IN), .ZN(n3043) );
  NAND2_X1 U3460 ( .A1(n2139), .A2(REG0_REG_4__SCAN_IN), .ZN(n3042) );
  NAND4_X1 U3461 ( .A1(n3045), .A2(n3044), .A3(n3043), .A4(n3042), .ZN(n3040)
         );
  OAI22_X1 U3462 ( .A1(n3053), .A2(n2134), .B1(n3041), .B2(n3989), .ZN(n2734)
         );
  XNOR2_X1 U3463 ( .A(n2734), .B(n3976), .ZN(n2739) );
  OAI22_X1 U3464 ( .A1(n2730), .A2(n3053), .B1(n3041), .B2(n2133), .ZN(n2740)
         );
  XNOR2_X1 U3465 ( .A(n2739), .B(n2740), .ZN(n3327) );
  INV_X1 U3466 ( .A(n2735), .ZN(n2737) );
  NAND2_X1 U34670 ( .A1(n2737), .A2(n2736), .ZN(n3328) );
  AND2_X1 U3468 ( .A1(n3327), .A2(n3328), .ZN(n2738) );
  INV_X1 U34690 ( .A(n2739), .ZN(n2741) );
  NAND2_X1 U3470 ( .A1(n2741), .A2(n2740), .ZN(n2742) );
  XNOR2_X1 U34710 ( .A(n2751), .B(REG3_REG_5__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U3472 ( .A1(n2769), .A2(n3511), .ZN(n3057) );
  NAND2_X1 U34730 ( .A1(n2137), .A2(REG2_REG_5__SCAN_IN), .ZN(n3056) );
  NAND2_X1 U3474 ( .A1(n3270), .A2(REG1_REG_5__SCAN_IN), .ZN(n3055) );
  NAND2_X1 U34750 ( .A1(n2732), .A2(REG0_REG_5__SCAN_IN), .ZN(n3054) );
  INV_X1 U3476 ( .A(DATAI_5_), .ZN(n2743) );
  OAI22_X1 U34770 ( .A1(n3478), .A2(n2134), .B1(n3404), .B2(n3989), .ZN(n2745)
         );
  XNOR2_X1 U3478 ( .A(n2745), .B(n3976), .ZN(n2746) );
  OAI22_X1 U34790 ( .A1(n2730), .A2(n3478), .B1(n3404), .B2(n2133), .ZN(n2747)
         );
  XNOR2_X1 U3480 ( .A(n2746), .B(n2747), .ZN(n3318) );
  INV_X1 U34810 ( .A(n2746), .ZN(n2748) );
  INV_X1 U3482 ( .A(n3334), .ZN(n2761) );
  NAND2_X1 U34830 ( .A1(n3270), .A2(REG1_REG_6__SCAN_IN), .ZN(n2756) );
  INV_X1 U3484 ( .A(n2749), .ZN(n2767) );
  INV_X1 U34850 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2750) );
  INV_X1 U3486 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3693) );
  OAI21_X1 U34870 ( .B1(n2751), .B2(n2750), .A(n3693), .ZN(n2752) );
  AND2_X1 U3488 ( .A1(n2767), .A2(n2752), .ZN(n3564) );
  NAND2_X1 U34890 ( .A1(n3014), .A2(n3564), .ZN(n2755) );
  NAND2_X1 U3490 ( .A1(n2732), .A2(REG0_REG_6__SCAN_IN), .ZN(n2753) );
  NAND2_X1 U34910 ( .A1(n3973), .A2(n4356), .ZN(n2758) );
  MUX2_X1 U3492 ( .A(n4872), .B(DATAI_6_), .S(n2135), .Z(n3406) );
  NAND2_X1 U34930 ( .A1(n2726), .A2(n3406), .ZN(n2757) );
  NAND2_X1 U3494 ( .A1(n2758), .A2(n2757), .ZN(n2759) );
  XNOR2_X1 U34950 ( .A(n2759), .B(n3986), .ZN(n2763) );
  INV_X1 U3496 ( .A(n4356), .ZN(n3604) );
  OAI22_X1 U34970 ( .A1(n2730), .A2(n3604), .B1(n3616), .B2(n2134), .ZN(n2762)
         );
  AND2_X1 U3498 ( .A1(n2763), .A2(n2762), .ZN(n3336) );
  INV_X1 U34990 ( .A(n3336), .ZN(n2760) );
  INV_X1 U3500 ( .A(n2762), .ZN(n2765) );
  INV_X1 U35010 ( .A(n2763), .ZN(n2764) );
  NAND2_X1 U3502 ( .A1(n2765), .A2(n2764), .ZN(n3335) );
  NAND2_X1 U35030 ( .A1(n3270), .A2(REG1_REG_7__SCAN_IN), .ZN(n2773) );
  INV_X1 U3504 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2766) );
  NAND2_X1 U35050 ( .A1(n2767), .A2(n2766), .ZN(n2768) );
  AND2_X1 U35060 ( .A1(n2786), .A2(n2768), .ZN(n3613) );
  NAND2_X1 U35070 ( .A1(n2769), .A2(n3613), .ZN(n2772) );
  NAND2_X1 U35080 ( .A1(n2136), .A2(REG2_REG_7__SCAN_IN), .ZN(n2771) );
  NAND2_X1 U35090 ( .A1(n2732), .A2(REG0_REG_7__SCAN_IN), .ZN(n2770) );
  MUX2_X1 U35100 ( .A(n4871), .B(DATAI_7_), .S(n2135), .Z(n3609) );
  OAI22_X1 U35110 ( .A1(n3392), .A2(n2134), .B1(n3603), .B2(n3989), .ZN(n2774)
         );
  XNOR2_X1 U35120 ( .A(n2774), .B(n3986), .ZN(n2777) );
  OAI22_X1 U35130 ( .A1(n2730), .A2(n3392), .B1(n3603), .B2(n2133), .ZN(n2776)
         );
  XNOR2_X1 U35140 ( .A(n2777), .B(n2776), .ZN(n3520) );
  NAND2_X1 U35150 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  NAND2_X1 U35160 ( .A1(n3270), .A2(REG1_REG_8__SCAN_IN), .ZN(n2782) );
  XNOR2_X1 U35170 ( .A(n2786), .B(REG3_REG_8__SCAN_IN), .ZN(n3491) );
  NAND2_X1 U35180 ( .A1(n3014), .A2(n3491), .ZN(n2781) );
  NAND2_X1 U35190 ( .A1(n2136), .A2(REG2_REG_8__SCAN_IN), .ZN(n2780) );
  NAND2_X1 U35200 ( .A1(n2732), .A2(REG0_REG_8__SCAN_IN), .ZN(n2779) );
  INV_X1 U35210 ( .A(DATAI_8_), .ZN(n3181) );
  MUX2_X1 U35220 ( .A(n3284), .B(n3181), .S(n2135), .Z(n3121) );
  OAI22_X1 U35230 ( .A1(n2730), .A2(n3516), .B1(n3121), .B2(n2134), .ZN(n3437)
         );
  OAI22_X1 U35240 ( .A1(n3516), .A2(n2134), .B1(n3121), .B2(n3989), .ZN(n2783)
         );
  XNOR2_X1 U35250 ( .A(n2783), .B(n3986), .ZN(n3436) );
  NAND2_X1 U35260 ( .A1(n3270), .A2(REG1_REG_9__SCAN_IN), .ZN(n2791) );
  INV_X1 U35270 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2785) );
  INV_X1 U35280 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2784) );
  OAI21_X1 U35290 ( .B1(n2786), .B2(n2785), .A(n2784), .ZN(n2787) );
  AND2_X1 U35300 ( .A1(n2787), .A2(n2797), .ZN(n3598) );
  NAND2_X1 U35310 ( .A1(n3014), .A2(n3598), .ZN(n2790) );
  NAND2_X1 U35320 ( .A1(n2136), .A2(REG2_REG_9__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U35330 ( .A1(n2732), .A2(REG0_REG_9__SCAN_IN), .ZN(n2788) );
  NAND4_X1 U35340 ( .A1(n2791), .A2(n2790), .A3(n2789), .A4(n2788), .ZN(n4355)
         );
  NAND2_X1 U35350 ( .A1(n3973), .A2(n4355), .ZN(n2794) );
  INV_X1 U35360 ( .A(DATAI_9_), .ZN(n2792) );
  MUX2_X1 U35370 ( .A(n3347), .B(n2792), .S(n2135), .Z(n3595) );
  INV_X1 U35380 ( .A(n3595), .ZN(n3123) );
  NAND2_X1 U35390 ( .A1(n2726), .A2(n3123), .ZN(n2793) );
  NAND2_X1 U35400 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  XNOR2_X1 U35410 ( .A(n2795), .B(n3986), .ZN(n2807) );
  OAI22_X1 U35420 ( .A1(n2730), .A2(n3444), .B1(n3595), .B2(n2134), .ZN(n2806)
         );
  XNOR2_X1 U35430 ( .A(n2807), .B(n2806), .ZN(n3594) );
  NAND2_X1 U35440 ( .A1(n3270), .A2(REG1_REG_10__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U35450 ( .A1(n2797), .A2(n3382), .ZN(n2798) );
  NAND2_X1 U35460 ( .A1(n2815), .A2(n2798), .ZN(n3649) );
  INV_X1 U35470 ( .A(n3649), .ZN(n3540) );
  NAND2_X1 U35480 ( .A1(n3014), .A2(n3540), .ZN(n2801) );
  NAND2_X1 U35490 ( .A1(n2136), .A2(REG2_REG_10__SCAN_IN), .ZN(n2800) );
  NAND2_X1 U35500 ( .A1(n2732), .A2(REG0_REG_10__SCAN_IN), .ZN(n2799) );
  NAND4_X1 U35510 ( .A1(n2802), .A2(n2801), .A3(n2800), .A4(n2799), .ZN(n4354)
         );
  NAND2_X1 U35520 ( .A1(n3973), .A2(n4354), .ZN(n2804) );
  MUX2_X1 U35530 ( .A(n4869), .B(DATAI_10_), .S(n4209), .Z(n3539) );
  NAND2_X1 U35540 ( .A1(n2726), .A2(n3539), .ZN(n2803) );
  NAND2_X1 U35550 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  XNOR2_X1 U35560 ( .A(n2805), .B(n3976), .ZN(n2811) );
  OAI22_X1 U35570 ( .A1(n2730), .A2(n4170), .B1(n3644), .B2(n2133), .ZN(n2812)
         );
  XNOR2_X1 U35580 ( .A(n2811), .B(n2812), .ZN(n3642) );
  INV_X1 U35590 ( .A(n2806), .ZN(n2809) );
  INV_X1 U35600 ( .A(n2807), .ZN(n2808) );
  NAND2_X1 U35610 ( .A1(n2809), .A2(n2808), .ZN(n3640) );
  AND2_X1 U35620 ( .A1(n3642), .A2(n3640), .ZN(n2810) );
  NAND2_X1 U35630 ( .A1(n3592), .A2(n2810), .ZN(n3641) );
  INV_X1 U35640 ( .A(n2811), .ZN(n2813) );
  NAND2_X1 U35650 ( .A1(n2813), .A2(n2812), .ZN(n2814) );
  NAND2_X1 U35660 ( .A1(n3641), .A2(n2814), .ZN(n4163) );
  NAND2_X1 U35670 ( .A1(n3270), .A2(REG1_REG_11__SCAN_IN), .ZN(n2820) );
  NAND2_X1 U35680 ( .A1(n2815), .A2(n2225), .ZN(n2816) );
  AND2_X1 U35690 ( .A1(n2828), .A2(n2816), .ZN(n4172) );
  NAND2_X1 U35700 ( .A1(n3014), .A2(n4172), .ZN(n2819) );
  NAND2_X1 U35710 ( .A1(n2137), .A2(REG2_REG_11__SCAN_IN), .ZN(n2818) );
  NAND2_X1 U35720 ( .A1(n2732), .A2(REG0_REG_11__SCAN_IN), .ZN(n2817) );
  MUX2_X1 U35730 ( .A(DATAI_11_), .B(n4868), .S(n2854), .Z(n4166) );
  NAND2_X1 U35740 ( .A1(n4166), .A2(n2726), .ZN(n2821) );
  OAI21_X1 U35750 ( .B1(n4062), .B2(n2134), .A(n2821), .ZN(n2822) );
  XNOR2_X1 U35760 ( .A(n2822), .B(n3976), .ZN(n2824) );
  AOI22_X1 U35770 ( .A1(n2823), .A2(n4353), .B1(n3973), .B2(n4166), .ZN(n2825)
         );
  NAND2_X1 U35780 ( .A1(n2824), .A2(n2825), .ZN(n4161) );
  INV_X1 U35790 ( .A(n2824), .ZN(n2827) );
  INV_X1 U35800 ( .A(n2825), .ZN(n2826) );
  NAND2_X1 U35810 ( .A1(n2827), .A2(n2826), .ZN(n4162) );
  MUX2_X1 U3582 ( .A(DATAI_12_), .B(n4867), .S(n2854), .Z(n4059) );
  NAND2_X1 U3583 ( .A1(n4059), .A2(n2726), .ZN(n2835) );
  NAND2_X1 U3584 ( .A1(n3270), .A2(REG1_REG_12__SCAN_IN), .ZN(n2833) );
  NAND2_X1 U3585 ( .A1(n2828), .A2(n2226), .ZN(n2829) );
  AND2_X1 U3586 ( .A1(n2840), .A2(n2829), .ZN(n4064) );
  NAND2_X1 U3587 ( .A1(n3014), .A2(n4064), .ZN(n2832) );
  NAND2_X1 U3588 ( .A1(n2136), .A2(REG2_REG_12__SCAN_IN), .ZN(n2831) );
  NAND2_X1 U3589 ( .A1(n2732), .A2(REG0_REG_12__SCAN_IN), .ZN(n2830) );
  NAND4_X1 U3590 ( .A1(n2833), .A2(n2832), .A3(n2831), .A4(n2830), .ZN(n4695)
         );
  NAND2_X1 U3591 ( .A1(n3973), .A2(n4695), .ZN(n2834) );
  NAND2_X1 U3592 ( .A1(n2835), .A2(n2834), .ZN(n2836) );
  XNOR2_X1 U3593 ( .A(n2836), .B(n3986), .ZN(n4055) );
  NAND2_X1 U3594 ( .A1(n4059), .A2(n3973), .ZN(n2838) );
  NAND2_X1 U3595 ( .A1(n2823), .A2(n4695), .ZN(n2837) );
  NAND2_X1 U3596 ( .A1(n2838), .A2(n2837), .ZN(n4056) );
  INV_X1 U3597 ( .A(DATAI_13_), .ZN(n2839) );
  MUX2_X1 U3598 ( .A(n3945), .B(n2839), .S(n4209), .Z(n4706) );
  NAND2_X1 U3599 ( .A1(n3270), .A2(REG1_REG_13__SCAN_IN), .ZN(n2845) );
  NAND2_X1 U3600 ( .A1(n2137), .A2(REG2_REG_13__SCAN_IN), .ZN(n2844) );
  NAND2_X1 U3601 ( .A1(n2840), .A2(n3906), .ZN(n2841) );
  AND2_X1 U3602 ( .A1(n2872), .A2(n2841), .ZN(n4709) );
  NAND2_X1 U3603 ( .A1(n3014), .A2(n4709), .ZN(n2843) );
  NAND2_X1 U3604 ( .A1(n2732), .A2(REG0_REG_13__SCAN_IN), .ZN(n2842) );
  OAI22_X1 U3605 ( .A1(n4706), .A2(n3989), .B1(n4677), .B2(n2133), .ZN(n2846)
         );
  XNOR2_X1 U3606 ( .A(n2846), .B(n3986), .ZN(n2847) );
  OAI22_X1 U3607 ( .A1(n4706), .A2(n2134), .B1(n4677), .B2(n2730), .ZN(n2848)
         );
  AND2_X1 U3608 ( .A1(n2847), .A2(n2848), .ZN(n4140) );
  INV_X1 U3609 ( .A(n2847), .ZN(n2850) );
  INV_X1 U3610 ( .A(n2848), .ZN(n2849) );
  NAND2_X1 U3611 ( .A1(n2850), .A2(n2849), .ZN(n4139) );
  NAND2_X1 U3612 ( .A1(n2862), .A2(n4088), .ZN(n2851) );
  NAND2_X1 U3613 ( .A1(n2884), .A2(n2851), .ZN(n4632) );
  AOI22_X1 U3614 ( .A1(n3270), .A2(REG1_REG_16__SCAN_IN), .B1(n2136), .B2(
        REG2_REG_16__SCAN_IN), .ZN(n2853) );
  NAND2_X1 U3615 ( .A1(n2732), .A2(REG0_REG_16__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U3616 ( .A1(n4608), .A2(n2141), .ZN(n2856) );
  INV_X1 U3617 ( .A(DATAI_16_), .ZN(n4977) );
  MUX2_X1 U3618 ( .A(n4977), .B(n4978), .S(n2854), .Z(n4089) );
  OR2_X1 U3619 ( .A1(n4089), .A2(n3989), .ZN(n2855) );
  NAND2_X1 U3620 ( .A1(n2856), .A2(n2855), .ZN(n2857) );
  XNOR2_X1 U3621 ( .A(n2857), .B(n3986), .ZN(n4097) );
  NAND2_X1 U3622 ( .A1(n2823), .A2(n4608), .ZN(n2859) );
  NAND2_X1 U3623 ( .A1(n4631), .A2(n2141), .ZN(n2858) );
  NAND2_X1 U3624 ( .A1(n2859), .A2(n2858), .ZN(n4096) );
  NAND2_X1 U3625 ( .A1(n2874), .A2(n2860), .ZN(n2861) );
  NAND2_X1 U3626 ( .A1(n2862), .A2(n2861), .ZN(n4650) );
  NAND2_X1 U3627 ( .A1(n3270), .A2(REG1_REG_15__SCAN_IN), .ZN(n2864) );
  NAND2_X1 U3628 ( .A1(n2137), .A2(REG2_REG_15__SCAN_IN), .ZN(n2863) );
  AND2_X1 U3629 ( .A1(n2864), .A2(n2863), .ZN(n2866) );
  NAND2_X1 U3630 ( .A1(n2732), .A2(REG0_REG_15__SCAN_IN), .ZN(n2865) );
  NAND2_X1 U3631 ( .A1(n2823), .A2(n4674), .ZN(n2868) );
  MUX2_X1 U3632 ( .A(n4913), .B(DATAI_15_), .S(n2135), .Z(n4629) );
  NAND2_X1 U3633 ( .A1(n2140), .A2(n4629), .ZN(n2867) );
  NAND2_X1 U3634 ( .A1(n2868), .A2(n2867), .ZN(n4189) );
  NAND2_X1 U3635 ( .A1(n4674), .A2(n3973), .ZN(n2870) );
  NAND2_X1 U3636 ( .A1(n2726), .A2(n4629), .ZN(n2869) );
  NAND2_X1 U3637 ( .A1(n2870), .A2(n2869), .ZN(n2871) );
  XNOR2_X1 U3638 ( .A(n2871), .B(n3986), .ZN(n4084) );
  AOI22_X1 U3639 ( .A1(n4097), .A2(n4096), .B1(n4189), .B2(n4084), .ZN(n2882)
         );
  INV_X1 U3640 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3875) );
  NAND2_X1 U3641 ( .A1(n2872), .A2(n3875), .ZN(n2873) );
  AND2_X1 U3642 ( .A1(n2874), .A2(n2873), .ZN(n4685) );
  NAND2_X1 U3643 ( .A1(n4685), .A2(n3014), .ZN(n2879) );
  NAND2_X1 U3644 ( .A1(n3270), .A2(REG1_REG_14__SCAN_IN), .ZN(n2878) );
  NAND2_X1 U3645 ( .A1(n2136), .A2(REG2_REG_14__SCAN_IN), .ZN(n2877) );
  NAND2_X1 U3646 ( .A1(n2732), .A2(REG0_REG_14__SCAN_IN), .ZN(n2876) );
  MUX2_X1 U3647 ( .A(n4901), .B(DATAI_14_), .S(n2138), .Z(n4673) );
  OAI22_X1 U3648 ( .A1(n3076), .A2(n2134), .B1(n4683), .B2(n3989), .ZN(n2880)
         );
  XNOR2_X1 U3649 ( .A(n2880), .B(n3986), .ZN(n4080) );
  OAI22_X1 U3650 ( .A1(n2730), .A2(n3076), .B1(n4683), .B2(n2133), .ZN(n4079)
         );
  NAND2_X1 U3651 ( .A1(n4080), .A2(n4079), .ZN(n2881) );
  NAND2_X1 U3652 ( .A1(n4018), .A2(n2181), .ZN(n2897) );
  INV_X1 U3653 ( .A(n2882), .ZN(n2883) );
  NAND2_X1 U3654 ( .A1(n2884), .A2(n2221), .ZN(n2885) );
  NAND2_X1 U3655 ( .A1(n2899), .A2(n2885), .ZN(n4616) );
  OR2_X1 U3656 ( .A1(n4616), .A2(n2281), .ZN(n2888) );
  AOI22_X1 U3657 ( .A1(n3270), .A2(REG1_REG_17__SCAN_IN), .B1(n2136), .B2(
        REG2_REG_17__SCAN_IN), .ZN(n2887) );
  NAND2_X1 U3658 ( .A1(n2732), .A2(REG0_REG_17__SCAN_IN), .ZN(n2886) );
  INV_X1 U3659 ( .A(DATAI_17_), .ZN(n4975) );
  MUX2_X1 U3660 ( .A(n4976), .B(n4975), .S(n2138), .Z(n4104) );
  OAI22_X1 U3661 ( .A1(n4622), .A2(n2134), .B1(n4104), .B2(n3989), .ZN(n2889)
         );
  XNOR2_X1 U3662 ( .A(n2889), .B(n3986), .ZN(n4098) );
  OAI22_X1 U3663 ( .A1(n4622), .A2(n2730), .B1(n4104), .B2(n2134), .ZN(n4099)
         );
  OAI21_X1 U3664 ( .B1(n4084), .B2(n4189), .A(n4096), .ZN(n2891) );
  INV_X1 U3665 ( .A(n4097), .ZN(n2890) );
  NAND2_X1 U3666 ( .A1(n2891), .A2(n2890), .ZN(n2894) );
  INV_X1 U3667 ( .A(n4084), .ZN(n2892) );
  INV_X1 U3668 ( .A(n4096), .ZN(n4078) );
  INV_X1 U3669 ( .A(n4189), .ZN(n4094) );
  NAND3_X1 U3670 ( .A1(n2892), .A2(n4078), .A3(n4094), .ZN(n2893) );
  OAI211_X1 U3671 ( .C1(n4098), .C2(n4099), .A(n2894), .B(n2893), .ZN(n2895)
         );
  NAND2_X1 U3672 ( .A1(n4098), .A2(n4099), .ZN(n2898) );
  NAND2_X1 U3673 ( .A1(n2899), .A2(n3951), .ZN(n2900) );
  AND2_X1 U3674 ( .A1(n2931), .A2(n2900), .ZN(n4601) );
  NAND2_X1 U3675 ( .A1(n4601), .A2(n3014), .ZN(n2905) );
  INV_X1 U3676 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3900) );
  NAND2_X1 U3677 ( .A1(n2732), .A2(REG0_REG_18__SCAN_IN), .ZN(n2902) );
  NAND2_X1 U3678 ( .A1(n2136), .A2(REG2_REG_18__SCAN_IN), .ZN(n2901) );
  OAI211_X1 U3679 ( .C1(n3277), .C2(n3900), .A(n2902), .B(n2901), .ZN(n2903)
         );
  INV_X1 U3680 ( .A(n2903), .ZN(n2904) );
  MUX2_X1 U3681 ( .A(n4865), .B(DATAI_18_), .S(n2138), .Z(n4598) );
  OAI22_X1 U3682 ( .A1(n4610), .A2(n2133), .B1(n3989), .B2(n4179), .ZN(n2906)
         );
  XNOR2_X1 U3683 ( .A(n2906), .B(n3986), .ZN(n2950) );
  OAI22_X1 U3684 ( .A1(n4610), .A2(n2730), .B1(n2133), .B2(n4179), .ZN(n2951)
         );
  AND2_X1 U3685 ( .A1(n2950), .A2(n2951), .ZN(n4176) );
  NAND2_X1 U3686 ( .A1(n2916), .A2(n4049), .ZN(n2907) );
  AND2_X1 U3687 ( .A1(n2957), .A2(n2907), .ZN(n4539) );
  NAND2_X1 U3688 ( .A1(n4539), .A2(n3014), .ZN(n2912) );
  INV_X1 U3689 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3864) );
  NAND2_X1 U3690 ( .A1(n3270), .A2(REG1_REG_21__SCAN_IN), .ZN(n2909) );
  NAND2_X1 U3691 ( .A1(n2732), .A2(REG0_REG_21__SCAN_IN), .ZN(n2908) );
  OAI211_X1 U3692 ( .C1(n3150), .C2(n3864), .A(n2909), .B(n2908), .ZN(n2910)
         );
  INV_X1 U3693 ( .A(n2910), .ZN(n2911) );
  AND2_X1 U3694 ( .A1(n2135), .A2(DATAI_21_), .ZN(n4533) );
  OAI22_X1 U3695 ( .A1(n4517), .A2(n2133), .B1(n4537), .B2(n3989), .ZN(n2913)
         );
  XNOR2_X1 U3696 ( .A(n2913), .B(n3976), .ZN(n4045) );
  NOR2_X1 U3697 ( .A1(n2133), .A2(n4537), .ZN(n2914) );
  AOI21_X1 U3698 ( .B1(n4555), .B2(n2823), .A(n2914), .ZN(n4044) );
  NAND2_X1 U3699 ( .A1(n4045), .A2(n4044), .ZN(n2945) );
  NAND2_X1 U3700 ( .A1(n2933), .A2(n4133), .ZN(n2915) );
  NAND2_X1 U3701 ( .A1(n2916), .A2(n2915), .ZN(n4132) );
  INV_X1 U3702 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4752) );
  NAND2_X1 U3703 ( .A1(n2732), .A2(REG0_REG_20__SCAN_IN), .ZN(n2918) );
  NAND2_X1 U3704 ( .A1(n2137), .A2(REG2_REG_20__SCAN_IN), .ZN(n2917) );
  OAI211_X1 U3705 ( .C1(n3277), .C2(n4752), .A(n2918), .B(n2917), .ZN(n2919)
         );
  INV_X1 U3706 ( .A(n2919), .ZN(n2920) );
  NAND2_X1 U3707 ( .A1(n4576), .A2(n3973), .ZN(n2923) );
  INV_X1 U3708 ( .A(n4559), .ZN(n4553) );
  OR2_X1 U3709 ( .A1(n3989), .A2(n4553), .ZN(n2922) );
  NAND2_X1 U3710 ( .A1(n2923), .A2(n2922), .ZN(n2924) );
  XNOR2_X1 U3711 ( .A(n2924), .B(n3986), .ZN(n2930) );
  INV_X1 U3712 ( .A(n2930), .ZN(n2928) );
  NAND2_X1 U3713 ( .A1(n4576), .A2(n2823), .ZN(n2926) );
  NAND2_X1 U3714 ( .A1(n3973), .A2(n4559), .ZN(n2925) );
  NAND2_X1 U3715 ( .A1(n2926), .A2(n2925), .ZN(n2929) );
  INV_X1 U3716 ( .A(n2929), .ZN(n2927) );
  NAND2_X1 U3717 ( .A1(n2928), .A2(n2927), .ZN(n4130) );
  NAND2_X1 U3718 ( .A1(n2930), .A2(n2929), .ZN(n4128) );
  INV_X1 U3719 ( .A(n4128), .ZN(n2944) );
  NAND2_X1 U3720 ( .A1(n2931), .A2(n2222), .ZN(n2932) );
  NAND2_X1 U3721 ( .A1(n2933), .A2(n2932), .ZN(n4583) );
  OR2_X1 U3722 ( .A1(n4583), .A2(n2281), .ZN(n2938) );
  INV_X1 U3723 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U3724 ( .A1(n2137), .A2(REG2_REG_19__SCAN_IN), .ZN(n2935) );
  NAND2_X1 U3725 ( .A1(n2732), .A2(REG0_REG_19__SCAN_IN), .ZN(n2934) );
  OAI211_X1 U3726 ( .C1(n4756), .C2(n3277), .A(n2935), .B(n2934), .ZN(n2936)
         );
  INV_X1 U3727 ( .A(n2936), .ZN(n2937) );
  NAND2_X1 U3728 ( .A1(n4352), .A2(n3973), .ZN(n2940) );
  MUX2_X1 U3729 ( .A(n4864), .B(DATAI_19_), .S(n2135), .Z(n4579) );
  NAND2_X1 U3730 ( .A1(n2726), .A2(n4579), .ZN(n2939) );
  NAND2_X1 U3731 ( .A1(n2940), .A2(n2939), .ZN(n2941) );
  XNOR2_X1 U3732 ( .A(n2941), .B(n3986), .ZN(n2947) );
  INV_X1 U3733 ( .A(n2947), .ZN(n2943) );
  INV_X1 U3734 ( .A(n4579), .ZN(n4574) );
  NOR2_X1 U3735 ( .A1(n4574), .A2(n2133), .ZN(n2942) );
  AOI21_X1 U3736 ( .B1(n4352), .B2(n2823), .A(n2942), .ZN(n2946) );
  NAND2_X1 U3737 ( .A1(n2943), .A2(n2946), .ZN(n4125) );
  OR2_X1 U3738 ( .A1(n2944), .A2(n4125), .ZN(n4121) );
  AND2_X1 U3739 ( .A1(n4130), .A2(n4121), .ZN(n4043) );
  AND2_X1 U3740 ( .A1(n2945), .A2(n4043), .ZN(n2954) );
  INV_X1 U3741 ( .A(n2954), .ZN(n2948) );
  XNOR2_X1 U3742 ( .A(n2947), .B(n2946), .ZN(n4123) );
  AND2_X1 U3743 ( .A1(n4123), .A2(n4128), .ZN(n4042) );
  NOR2_X1 U3744 ( .A1(n2948), .A2(n4042), .ZN(n2956) );
  OR2_X1 U3745 ( .A1(n4176), .A2(n2956), .ZN(n2949) );
  INV_X1 U3746 ( .A(n2950), .ZN(n2953) );
  INV_X1 U3747 ( .A(n2951), .ZN(n2952) );
  NAND2_X1 U3748 ( .A1(n2953), .A2(n2952), .ZN(n4175) );
  AND2_X1 U3749 ( .A1(n4175), .A2(n2954), .ZN(n2955) );
  INV_X1 U3750 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U3751 ( .A1(n2957), .A2(n4156), .ZN(n2958) );
  AND2_X1 U3752 ( .A1(n2972), .A2(n2958), .ZN(n4522) );
  NAND2_X1 U3753 ( .A1(n4522), .A2(n3014), .ZN(n2963) );
  INV_X1 U3754 ( .A(REG1_REG_22__SCAN_IN), .ZN(n3862) );
  NAND2_X1 U3755 ( .A1(n2732), .A2(REG0_REG_22__SCAN_IN), .ZN(n2960) );
  NAND2_X1 U3756 ( .A1(n2136), .A2(REG2_REG_22__SCAN_IN), .ZN(n2959) );
  OAI211_X1 U3757 ( .C1(n3277), .C2(n3862), .A(n2960), .B(n2959), .ZN(n2961)
         );
  INV_X1 U3758 ( .A(n2961), .ZN(n2962) );
  NAND2_X1 U3759 ( .A1(n4351), .A2(n3973), .ZN(n2965) );
  NAND2_X1 U3760 ( .A1(n2135), .A2(DATAI_22_), .ZN(n4524) );
  OR2_X1 U3761 ( .A1(n3989), .A2(n4524), .ZN(n2964) );
  NAND2_X1 U3762 ( .A1(n2965), .A2(n2964), .ZN(n2966) );
  XNOR2_X1 U3763 ( .A(n2966), .B(n3976), .ZN(n2984) );
  NOR2_X1 U3764 ( .A1(n2133), .A2(n4524), .ZN(n2967) );
  AOI21_X1 U3765 ( .B1(n4351), .B2(n2823), .A(n2967), .ZN(n2983) );
  XNOR2_X1 U3766 ( .A(n2984), .B(n2983), .ZN(n4154) );
  INV_X1 U3767 ( .A(n4154), .ZN(n2970) );
  INV_X1 U3768 ( .A(n4045), .ZN(n2969) );
  INV_X1 U3769 ( .A(n4044), .ZN(n2968) );
  NAND2_X1 U3770 ( .A1(n2969), .A2(n2968), .ZN(n4150) );
  AND2_X1 U3771 ( .A1(n2970), .A2(n4150), .ZN(n2971) );
  NAND2_X1 U3772 ( .A1(n2972), .A2(n2219), .ZN(n2973) );
  NAND2_X1 U3773 ( .A1(n2989), .A2(n2973), .ZN(n4506) );
  INV_X1 U3774 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U3775 ( .A1(n3270), .A2(REG1_REG_23__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3776 ( .A1(n2732), .A2(REG0_REG_23__SCAN_IN), .ZN(n2974) );
  OAI211_X1 U3777 ( .C1(n3150), .C2(n4505), .A(n2975), .B(n2974), .ZN(n2976)
         );
  INV_X1 U3778 ( .A(n2976), .ZN(n2977) );
  NAND2_X1 U3779 ( .A1(n4519), .A2(n2140), .ZN(n2980) );
  AND2_X1 U3780 ( .A1(n2135), .A2(DATAI_23_), .ZN(n4502) );
  OR2_X1 U3781 ( .A1(n3989), .A2(n3092), .ZN(n2979) );
  NAND2_X1 U3782 ( .A1(n2980), .A2(n2979), .ZN(n2981) );
  XNOR2_X1 U3783 ( .A(n2981), .B(n3986), .ZN(n2988) );
  NOR2_X1 U3784 ( .A1(n2134), .A2(n3092), .ZN(n2982) );
  AOI21_X1 U3785 ( .B1(n4519), .B2(n2823), .A(n2982), .ZN(n2986) );
  XNOR2_X1 U3786 ( .A(n2988), .B(n2986), .ZN(n4027) );
  NAND2_X1 U3787 ( .A1(n2984), .A2(n2983), .ZN(n4025) );
  AND2_X1 U3788 ( .A1(n4027), .A2(n4025), .ZN(n2985) );
  INV_X1 U3789 ( .A(n2986), .ZN(n2987) );
  NAND2_X1 U3790 ( .A1(n2988), .A2(n2987), .ZN(n3002) );
  NAND2_X1 U3791 ( .A1(n2989), .A2(n4113), .ZN(n2990) );
  NAND2_X1 U3792 ( .A1(n4486), .A2(n3014), .ZN(n2996) );
  INV_X1 U3793 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U3794 ( .A1(n2732), .A2(REG0_REG_24__SCAN_IN), .ZN(n2993) );
  NAND2_X1 U3795 ( .A1(n2137), .A2(REG2_REG_24__SCAN_IN), .ZN(n2992) );
  OAI211_X1 U3796 ( .C1(n3277), .C2(n4736), .A(n2993), .B(n2992), .ZN(n2994)
         );
  INV_X1 U3797 ( .A(n2994), .ZN(n2995) );
  AND2_X1 U3798 ( .A1(n2135), .A2(DATAI_24_), .ZN(n4115) );
  INV_X1 U3799 ( .A(n4115), .ZN(n4484) );
  NOR2_X1 U3800 ( .A1(n2134), .A2(n4484), .ZN(n2997) );
  AOI21_X1 U3801 ( .B1(n4498), .B2(n2823), .A(n2997), .ZN(n3003) );
  AND2_X1 U3802 ( .A1(n3002), .A2(n3003), .ZN(n2998) );
  NAND2_X1 U3803 ( .A1(n4498), .A2(n3973), .ZN(n3000) );
  OR2_X1 U3804 ( .A1(n3989), .A2(n4484), .ZN(n2999) );
  NAND2_X1 U3805 ( .A1(n3000), .A2(n2999), .ZN(n3001) );
  XNOR2_X1 U3806 ( .A(n3001), .B(n3986), .ZN(n4112) );
  INV_X1 U3807 ( .A(n3003), .ZN(n3004) );
  NAND2_X1 U3808 ( .A1(n4479), .A2(n2141), .ZN(n3006) );
  AND2_X1 U3809 ( .A1(n2138), .A2(DATAI_25_), .ZN(n4458) );
  OR2_X1 U3810 ( .A1(n3989), .A2(n4462), .ZN(n3005) );
  NAND2_X1 U3811 ( .A1(n3006), .A2(n3005), .ZN(n3007) );
  XNOR2_X1 U3812 ( .A(n3007), .B(n3976), .ZN(n3009) );
  NOR2_X1 U3813 ( .A1(n2133), .A2(n4462), .ZN(n3008) );
  AOI21_X1 U3814 ( .B1(n4479), .B2(n2823), .A(n3008), .ZN(n3010) );
  NAND2_X1 U3815 ( .A1(n3009), .A2(n3010), .ZN(n4067) );
  NAND2_X1 U3816 ( .A1(n4069), .A2(n4067), .ZN(n3013) );
  INV_X1 U3817 ( .A(n3009), .ZN(n3012) );
  INV_X1 U3818 ( .A(n3010), .ZN(n3011) );
  NAND2_X1 U3819 ( .A1(n3012), .A2(n3011), .ZN(n4068) );
  NAND2_X1 U3820 ( .A1(n3013), .A2(n4068), .ZN(n3970) );
  NAND2_X1 U3821 ( .A1(n4447), .A2(n3014), .ZN(n3019) );
  INV_X1 U3822 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U3823 ( .A1(n2732), .A2(REG0_REG_26__SCAN_IN), .ZN(n3016) );
  NAND2_X1 U3824 ( .A1(n2137), .A2(REG2_REG_26__SCAN_IN), .ZN(n3015) );
  OAI211_X1 U3825 ( .C1(n3277), .C2(n4728), .A(n3016), .B(n3015), .ZN(n3017)
         );
  INV_X1 U3826 ( .A(n3017), .ZN(n3018) );
  OAI22_X1 U3827 ( .A1(n4461), .A2(n2133), .B1(n3989), .B2(n4445), .ZN(n3020)
         );
  XNOR2_X1 U3828 ( .A(n3020), .B(n3986), .ZN(n3026) );
  INV_X1 U3829 ( .A(n3026), .ZN(n3024) );
  OR2_X1 U3830 ( .A1(n4461), .A2(n2730), .ZN(n3022) );
  NAND2_X1 U3831 ( .A1(n3973), .A2(n4439), .ZN(n3021) );
  NAND2_X1 U3832 ( .A1(n3022), .A2(n3021), .ZN(n3025) );
  INV_X1 U3833 ( .A(n3025), .ZN(n3023) );
  NAND2_X1 U3834 ( .A1(n3024), .A2(n3023), .ZN(n3971) );
  INV_X1 U3835 ( .A(n3971), .ZN(n3027) );
  AND2_X1 U3836 ( .A1(n3026), .A2(n3025), .ZN(n3969) );
  NOR2_X1 U3837 ( .A1(n3027), .A2(n3969), .ZN(n3028) );
  XNOR2_X1 U3838 ( .A(n3970), .B(n3028), .ZN(n3032) );
  NOR2_X1 U3839 ( .A1(n3029), .A2(n3162), .ZN(n3030) );
  NAND2_X1 U3840 ( .A1(n3110), .A2(n3251), .ZN(n3253) );
  NAND2_X1 U3841 ( .A1(n3253), .A2(n3037), .ZN(n3363) );
  INV_X1 U3842 ( .A(n3363), .ZN(n3039) );
  NAND2_X1 U3843 ( .A1(n3248), .A2(n3365), .ZN(n3115) );
  NAND2_X1 U3844 ( .A1(n3551), .A2(n3374), .ZN(n4281) );
  NAND2_X1 U3845 ( .A1(n3039), .A2(n3038), .ZN(n3362) );
  INV_X1 U3846 ( .A(n3046), .ZN(n3041) );
  NAND2_X1 U3847 ( .A1(n3041), .A2(n3040), .ZN(n3117) );
  NAND2_X1 U3848 ( .A1(n3053), .A2(n3046), .ZN(n3116) );
  AND2_X2 U3849 ( .A1(n3117), .A2(n3116), .ZN(n4239) );
  NAND2_X1 U3850 ( .A1(n3478), .A2(n3404), .ZN(n3052) );
  NAND2_X1 U3851 ( .A1(n3248), .A2(n3374), .ZN(n3546) );
  NAND2_X1 U3852 ( .A1(n3052), .A2(n3469), .ZN(n3048) );
  NOR2_X1 U3853 ( .A1(n4239), .A2(n3048), .ZN(n3049) );
  NAND2_X1 U3854 ( .A1(n3362), .A2(n3049), .ZN(n3064) );
  INV_X1 U3855 ( .A(n4239), .ZN(n3050) );
  NAND2_X1 U3856 ( .A1(n3050), .A2(n3052), .ZN(n3051) );
  NAND2_X1 U3857 ( .A1(n3475), .A2(n3550), .ZN(n3470) );
  NOR2_X1 U3858 ( .A1(n3051), .A2(n3470), .ZN(n3062) );
  INV_X1 U3859 ( .A(n3052), .ZN(n3060) );
  NAND2_X1 U3860 ( .A1(n3040), .A2(n3482), .ZN(n3499) );
  NAND4_X1 U3861 ( .A1(n3057), .A2(n3056), .A3(n3055), .A4(n3054), .ZN(n4357)
         );
  INV_X1 U3862 ( .A(n3404), .ZN(n3507) );
  NAND2_X1 U3863 ( .A1(n4357), .A2(n3507), .ZN(n3058) );
  AND2_X1 U3864 ( .A1(n3499), .A2(n3058), .ZN(n3059) );
  NOR2_X1 U3865 ( .A1(n3060), .A2(n3059), .ZN(n3061) );
  NOR2_X1 U3866 ( .A1(n3062), .A2(n3061), .ZN(n3063) );
  NAND2_X1 U3867 ( .A1(n3392), .A2(n3609), .ZN(n3119) );
  AND2_X1 U3868 ( .A1(n4356), .A2(n3406), .ZN(n3066) );
  AOI22_X1 U3869 ( .A1(n4249), .A2(n3066), .B1(n3609), .B2(n3441), .ZN(n3067)
         );
  NAND2_X1 U3870 ( .A1(n3606), .A2(n3440), .ZN(n3068) );
  INV_X1 U3871 ( .A(n3456), .ZN(n3069) );
  NAND2_X1 U3872 ( .A1(n3444), .A2(n3595), .ZN(n3070) );
  NAND2_X1 U3873 ( .A1(n4166), .A2(n4062), .ZN(n4274) );
  INV_X1 U3874 ( .A(n4166), .ZN(n3573) );
  NAND2_X1 U3875 ( .A1(n3573), .A2(n4353), .ZN(n4309) );
  NAND2_X1 U3876 ( .A1(n4059), .A2(n4695), .ZN(n3072) );
  NAND2_X1 U3877 ( .A1(n3631), .A2(n3072), .ZN(n3074) );
  INV_X1 U3878 ( .A(n4059), .ZN(n3634) );
  INV_X1 U3879 ( .A(n4695), .ZN(n4146) );
  NAND2_X1 U3880 ( .A1(n3634), .A2(n4146), .ZN(n3073) );
  NAND2_X1 U3881 ( .A1(n3074), .A2(n3073), .ZN(n4634) );
  NAND2_X1 U3882 ( .A1(n4706), .A2(n4677), .ZN(n4251) );
  INV_X1 U3883 ( .A(n4251), .ZN(n4635) );
  NAND2_X1 U3884 ( .A1(n4674), .A2(n4629), .ZN(n4639) );
  INV_X1 U3885 ( .A(n4639), .ZN(n3075) );
  NAND2_X1 U3886 ( .A1(n3076), .A2(n4683), .ZN(n4638) );
  NOR2_X1 U3887 ( .A1(n3075), .A2(n4638), .ZN(n3079) );
  OR2_X1 U3888 ( .A1(n4635), .A2(n3079), .ZN(n3081) );
  NAND2_X1 U3889 ( .A1(n3076), .A2(n4673), .ZN(n4657) );
  NAND2_X1 U3890 ( .A1(n4698), .A2(n4683), .ZN(n3128) );
  NAND2_X1 U3891 ( .A1(n4657), .A2(n3128), .ZN(n4680) );
  AND2_X1 U3892 ( .A1(n4680), .A2(n4639), .ZN(n3077) );
  INV_X1 U3893 ( .A(n4706), .ZN(n4143) );
  NAND2_X1 U3894 ( .A1(n4143), .A2(n4058), .ZN(n4636) );
  AND2_X1 U3895 ( .A1(n3077), .A2(n4636), .ZN(n3078) );
  OR2_X1 U3896 ( .A1(n3079), .A2(n3078), .ZN(n3080) );
  NAND2_X1 U3897 ( .A1(n4608), .A2(n4089), .ZN(n4201) );
  OR2_X1 U3898 ( .A1(n4608), .A2(n4089), .ZN(n4317) );
  INV_X1 U3899 ( .A(n4645), .ZN(n3082) );
  INV_X1 U3900 ( .A(n4674), .ZN(n4621) );
  NAND2_X1 U3901 ( .A1(n4621), .A2(n4653), .ZN(n4640) );
  AND2_X1 U3902 ( .A1(n3082), .A2(n4640), .ZN(n3083) );
  NAND2_X1 U3903 ( .A1(n3084), .A2(n3083), .ZN(n4642) );
  NAND2_X1 U3904 ( .A1(n4608), .A2(n4631), .ZN(n3085) );
  NAND2_X1 U3905 ( .A1(n4622), .A2(n4104), .ZN(n3086) );
  NAND2_X1 U3906 ( .A1(n4610), .A2(n4598), .ZN(n4569) );
  NAND2_X1 U3907 ( .A1(n4035), .A2(n4179), .ZN(n4570) );
  NAND2_X1 U3908 ( .A1(n4569), .A2(n4570), .ZN(n4597) );
  NAND2_X1 U3909 ( .A1(n4595), .A2(n4597), .ZN(n4596) );
  NAND2_X1 U3910 ( .A1(n4596), .A2(n2403), .ZN(n4544) );
  NOR2_X1 U3911 ( .A1(n4352), .A2(n4579), .ZN(n4545) );
  NAND2_X1 U3912 ( .A1(n4576), .A2(n4559), .ZN(n4254) );
  NAND2_X1 U3913 ( .A1(n4352), .A2(n4579), .ZN(n4546) );
  OAI211_X1 U3914 ( .C1(n4544), .C2(n4545), .A(n4254), .B(n4546), .ZN(n3087)
         );
  INV_X1 U3915 ( .A(n4576), .ZN(n4048) );
  NAND2_X1 U3916 ( .A1(n4048), .A2(n4553), .ZN(n4255) );
  NAND2_X1 U3917 ( .A1(n3087), .A2(n4255), .ZN(n4529) );
  NAND2_X1 U3918 ( .A1(n4555), .A2(n4533), .ZN(n3089) );
  AOI21_X2 U3919 ( .B1(n4529), .B2(n3089), .A(n3088), .ZN(n4513) );
  NAND2_X1 U3920 ( .A1(n4351), .A2(n4524), .ZN(n3138) );
  NAND2_X1 U3921 ( .A1(n4494), .A2(n3138), .ZN(n4512) );
  INV_X1 U3922 ( .A(n4524), .ZN(n3090) );
  OAI21_X1 U3923 ( .B1(n4470), .B2(n2407), .A(n2402), .ZN(n3095) );
  INV_X1 U3924 ( .A(n3095), .ZN(n4452) );
  NOR2_X1 U3925 ( .A1(n4461), .A2(n4445), .ZN(n3100) );
  NAND2_X1 U3926 ( .A1(n4461), .A2(n4445), .ZN(n3099) );
  NOR2_X1 U3927 ( .A1(n4268), .A2(n4423), .ZN(n3101) );
  INV_X1 U3928 ( .A(n4423), .ZN(n4269) );
  INV_X1 U3929 ( .A(n3103), .ZN(n3102) );
  NAND2_X1 U3930 ( .A1(n3102), .A2(REG3_REG_28__SCAN_IN), .ZN(n4392) );
  INV_X1 U3931 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3832) );
  INV_X1 U3932 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3720) );
  NAND2_X1 U3933 ( .A1(n2732), .A2(REG0_REG_28__SCAN_IN), .ZN(n3105) );
  NAND2_X1 U3934 ( .A1(n2136), .A2(REG2_REG_28__SCAN_IN), .ZN(n3104) );
  OAI211_X1 U3935 ( .C1(n3277), .C2(n3720), .A(n3105), .B(n3104), .ZN(n3106)
         );
  INV_X1 U3936 ( .A(n3106), .ZN(n3107) );
  AND2_X1 U3937 ( .A1(n2138), .A2(DATAI_28_), .ZN(n4405) );
  NAND2_X1 U3938 ( .A1(n4426), .A2(n4405), .ZN(n4393) );
  XNOR2_X1 U3939 ( .A(n2686), .B(n4345), .ZN(n3109) );
  NAND2_X1 U3940 ( .A1(n3109), .A2(n4341), .ZN(n4704) );
  INV_X1 U3941 ( .A(n3110), .ZN(n3112) );
  NAND2_X1 U3942 ( .A1(n3111), .A2(n3242), .ZN(n3244) );
  NAND2_X1 U3943 ( .A1(n3243), .A2(n3113), .ZN(n3114) );
  NAND2_X1 U3944 ( .A1(n3114), .A2(n4238), .ZN(n3369) );
  NAND2_X1 U3945 ( .A1(n3369), .A2(n3115), .ZN(n3549) );
  NAND2_X1 U3946 ( .A1(n3367), .A2(n3550), .ZN(n4283) );
  NAND2_X1 U3947 ( .A1(n3475), .A2(n3047), .ZN(n4280) );
  NAND2_X1 U3948 ( .A1(n3549), .A2(n4245), .ZN(n3548) );
  NAND2_X1 U3949 ( .A1(n3478), .A2(n3507), .ZN(n4297) );
  NAND2_X1 U3950 ( .A1(n4356), .A2(n3616), .ZN(n4301) );
  NAND2_X1 U3951 ( .A1(n3604), .A2(n3406), .ZN(n4286) );
  NAND2_X1 U3952 ( .A1(n3118), .A2(n4286), .ZN(n3602) );
  INV_X1 U3953 ( .A(n3119), .ZN(n3120) );
  NAND2_X1 U3954 ( .A1(n3516), .A2(n3440), .ZN(n4290) );
  NAND2_X1 U3955 ( .A1(n3391), .A2(n4290), .ZN(n3122) );
  NAND2_X1 U3956 ( .A1(n3606), .A2(n3121), .ZN(n4298) );
  NAND2_X1 U3957 ( .A1(n3122), .A2(n4298), .ZN(n3457) );
  AND2_X1 U3958 ( .A1(n4355), .A2(n3595), .ZN(n4303) );
  NAND2_X1 U3959 ( .A1(n3444), .A2(n3123), .ZN(n4291) );
  NAND2_X1 U3960 ( .A1(n4354), .A2(n3644), .ZN(n4308) );
  NAND2_X1 U3961 ( .A1(n4170), .A2(n3539), .ZN(n4305) );
  NAND2_X1 U3962 ( .A1(n4706), .A2(n4058), .ZN(n3124) );
  NAND2_X1 U3963 ( .A1(n3634), .A2(n4695), .ZN(n4690) );
  AND2_X1 U3964 ( .A1(n4310), .A2(n4309), .ZN(n3125) );
  NAND2_X1 U3965 ( .A1(n3627), .A2(n3125), .ZN(n3127) );
  AND2_X1 U3966 ( .A1(n4059), .A2(n4146), .ZN(n4691) );
  NOR2_X1 U3967 ( .A1(n4706), .A2(n4058), .ZN(n3126) );
  AOI21_X1 U3968 ( .B1(n4310), .B2(n4691), .A(n3126), .ZN(n4272) );
  NAND2_X1 U3969 ( .A1(n4621), .A2(n4629), .ZN(n4248) );
  NAND2_X1 U3970 ( .A1(n4248), .A2(n4657), .ZN(n4270) );
  NAND2_X1 U3971 ( .A1(n4674), .A2(n4653), .ZN(n4247) );
  NAND2_X1 U3972 ( .A1(n4247), .A2(n3128), .ZN(n4293) );
  NAND2_X1 U3973 ( .A1(n4293), .A2(n4248), .ZN(n4316) );
  NAND2_X1 U3974 ( .A1(n4352), .A2(n4574), .ZN(n3129) );
  NAND2_X1 U3975 ( .A1(n3129), .A2(n4570), .ZN(n3130) );
  AND2_X1 U3976 ( .A1(n4590), .A2(n4104), .ZN(n4568) );
  AND2_X1 U3977 ( .A1(n4576), .A2(n4553), .ZN(n3137) );
  INV_X1 U3978 ( .A(n3130), .ZN(n3132) );
  NAND2_X1 U3979 ( .A1(n4622), .A2(n2230), .ZN(n4567) );
  NAND2_X1 U3980 ( .A1(n4569), .A2(n4567), .ZN(n3131) );
  NAND2_X1 U3981 ( .A1(n3132), .A2(n3131), .ZN(n3134) );
  INV_X1 U3982 ( .A(n4352), .ZN(n4592) );
  NAND2_X1 U3983 ( .A1(n4592), .A2(n4579), .ZN(n3133) );
  NAND2_X1 U3984 ( .A1(n3134), .A2(n3133), .ZN(n4549) );
  NOR2_X1 U3985 ( .A1(n4576), .A2(n4553), .ZN(n3135) );
  OR2_X1 U3986 ( .A1(n4549), .A2(n3135), .ZN(n3136) );
  INV_X1 U3987 ( .A(n3137), .ZN(n4202) );
  NAND2_X1 U3988 ( .A1(n3136), .A2(n4202), .ZN(n4203) );
  NAND2_X1 U3989 ( .A1(n4494), .A2(n4493), .ZN(n3140) );
  AND2_X1 U3990 ( .A1(n4555), .A2(n4537), .ZN(n4227) );
  NAND2_X1 U3991 ( .A1(n4494), .A2(n4227), .ZN(n3139) );
  NAND2_X1 U3992 ( .A1(n4519), .A2(n3092), .ZN(n4226) );
  AND3_X1 U3993 ( .A1(n3139), .A2(n4226), .A3(n3138), .ZN(n4324) );
  OAI21_X2 U3994 ( .B1(n4492), .B2(n3140), .A(n4324), .ZN(n4473) );
  NAND2_X1 U3995 ( .A1(n4072), .A2(n4115), .ZN(n4225) );
  NAND2_X1 U3996 ( .A1(n3093), .A2(n4502), .ZN(n4472) );
  AND2_X2 U3997 ( .A1(n4473), .A2(n4325), .ZN(n4433) );
  OR2_X1 U3998 ( .A1(n4350), .A2(n4445), .ZN(n3141) );
  NAND2_X1 U3999 ( .A1(n4117), .A2(n4458), .ZN(n4434) );
  NAND2_X1 U4000 ( .A1(n3141), .A2(n4434), .ZN(n4211) );
  NAND2_X1 U4001 ( .A1(n4479), .A2(n4462), .ZN(n4224) );
  NAND2_X1 U4002 ( .A1(n4498), .A2(n4484), .ZN(n4453) );
  NAND2_X1 U4003 ( .A1(n4224), .A2(n4453), .ZN(n4435) );
  AND2_X1 U4004 ( .A1(n4350), .A2(n4445), .ZN(n4214) );
  AOI21_X1 U4005 ( .B1(n3143), .B2(n4435), .A(n4214), .ZN(n4329) );
  XNOR2_X1 U4006 ( .A(n4268), .B(n4423), .ZN(n4422) );
  NAND2_X1 U4007 ( .A1(n4442), .A2(n4423), .ZN(n4206) );
  XNOR2_X1 U4008 ( .A(n4396), .B(n2305), .ZN(n3146) );
  NAND2_X1 U4009 ( .A1(n4863), .A2(n4277), .ZN(n4222) );
  NAND2_X1 U4010 ( .A1(n4345), .A2(n4864), .ZN(n3144) );
  NAND2_X1 U4011 ( .A1(n3146), .A2(n3145), .ZN(n3160) );
  OR2_X1 U4012 ( .A1(n4392), .A2(n2281), .ZN(n3153) );
  INV_X1 U4013 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4014 ( .A1(n3270), .A2(REG1_REG_29__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4015 ( .A1(n2732), .A2(REG0_REG_29__SCAN_IN), .ZN(n3147) );
  OAI211_X1 U4016 ( .C1(n3150), .C2(n3149), .A(n3148), .B(n3147), .ZN(n3151)
         );
  INV_X1 U4017 ( .A(n3151), .ZN(n3152) );
  OAI22_X1 U4018 ( .A1(n4207), .A2(n4654), .B1(n4700), .B2(n3988), .ZN(n3155)
         );
  INV_X1 U4019 ( .A(n4696), .ZN(n3157) );
  OAI21_X1 U4020 ( .B1(n4017), .B2(n5005), .A(n4012), .ZN(n3176) );
  NOR2_X1 U4021 ( .A1(n3162), .A2(n3161), .ZN(n3424) );
  NAND4_X1 U4022 ( .A1(n3165), .A2(n3424), .A3(n3164), .A4(n3163), .ZN(n3175)
         );
  OR2_X1 U4023 ( .A1(n3176), .A2(n5019), .ZN(n3167) );
  OR2_X1 U4024 ( .A1(n5022), .A2(REG1_REG_28__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4025 ( .A1(n3167), .A2(n3166), .ZN(n3173) );
  AND2_X1 U4026 ( .A1(n3616), .A2(n3404), .ZN(n3169) );
  NAND2_X1 U4027 ( .A1(n3461), .A2(n3644), .ZN(n3536) );
  OR2_X2 U4028 ( .A1(n3536), .A2(n4166), .ZN(n3632) );
  NAND2_X1 U4029 ( .A1(n4653), .A2(n4089), .ZN(n3171) );
  NOR2_X4 U4030 ( .A1(n4580), .A2(n4579), .ZN(n4558) );
  OAI21_X1 U4031 ( .B1(n4417), .B2(n3988), .A(n4411), .ZN(n4010) );
  NAND2_X1 U4032 ( .A1(n3173), .A2(n3172), .ZN(U3546) );
  INV_X1 U4033 ( .A(n3425), .ZN(n3174) );
  OR2_X1 U4034 ( .A1(n3176), .A2(n5011), .ZN(n3178) );
  OR2_X1 U4035 ( .A1(n5013), .A2(REG0_REG_28__SCAN_IN), .ZN(n3177) );
  NAND2_X1 U4036 ( .A1(n3178), .A2(n3177), .ZN(n3180) );
  NAND2_X1 U4037 ( .A1(n3180), .A2(n3179), .ZN(U3514) );
  MUX2_X1 U4038 ( .A(n3181), .B(n3284), .S(STATE_REG_SCAN_IN), .Z(n3182) );
  INV_X1 U4039 ( .A(n3182), .ZN(U3344) );
  INV_X1 U4040 ( .A(DATAI_29_), .ZN(n3184) );
  OAI21_X1 U4041 ( .B1(STATE_REG_SCAN_IN), .B2(n3184), .A(n3183), .ZN(U3323)
         );
  INV_X1 U4042 ( .A(DATAI_21_), .ZN(n3751) );
  NAND2_X1 U40430 ( .A1(n4277), .A2(STATE_REG_SCAN_IN), .ZN(n3185) );
  OAI21_X1 U4044 ( .B1(STATE_REG_SCAN_IN), .B2(n3751), .A(n3185), .ZN(U3331)
         );
  INV_X1 U4045 ( .A(DATAI_22_), .ZN(n3732) );
  NAND2_X1 U4046 ( .A1(n4345), .A2(STATE_REG_SCAN_IN), .ZN(n3186) );
  OAI21_X1 U4047 ( .B1(STATE_REG_SCAN_IN), .B2(n3732), .A(n3186), .ZN(U3330)
         );
  INV_X1 U4048 ( .A(DATAI_24_), .ZN(n3735) );
  NAND2_X1 U4049 ( .A1(n3193), .A2(STATE_REG_SCAN_IN), .ZN(n3187) );
  OAI21_X1 U4050 ( .B1(STATE_REG_SCAN_IN), .B2(n3735), .A(n3187), .ZN(U3328)
         );
  INV_X1 U4051 ( .A(D_REG_1__SCAN_IN), .ZN(n3192) );
  INV_X1 U4052 ( .A(n3189), .ZN(n3191) );
  INV_X1 U4053 ( .A(n4973), .ZN(n3190) );
  AOI22_X1 U4054 ( .A1(n4972), .A2(n3192), .B1(n3191), .B2(n3190), .ZN(U3459)
         );
  INV_X1 U4055 ( .A(D_REG_0__SCAN_IN), .ZN(n3195) );
  NOR3_X1 U4056 ( .A1(n3193), .A2(n2602), .A3(n4973), .ZN(n3194) );
  AOI21_X1 U4057 ( .B1(n3195), .B2(n4972), .A(n3194), .ZN(U3458) );
  INV_X1 U4058 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3201) );
  INV_X1 U4059 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U4060 ( .A1(n4860), .A2(n4954), .ZN(n3196) );
  AND2_X1 U4061 ( .A1(n4859), .A2(n3196), .ZN(n4362) );
  OAI21_X1 U4062 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4860), .A(n4362), .ZN(n3197)
         );
  XNOR2_X1 U4063 ( .A(n3197), .B(IR_REG_0__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4064 ( .A1(n3199), .A2(n3198), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3200) );
  OAI21_X1 U4065 ( .B1(n4918), .B2(n3201), .A(n3200), .ZN(U3240) );
  XNOR2_X1 U4066 ( .A(n3202), .B(REG1_REG_6__SCAN_IN), .ZN(n3209) );
  NOR2_X1 U4067 ( .A1(STATE_REG_SCAN_IN), .A2(n3693), .ZN(n3340) );
  INV_X1 U4068 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n3790) );
  XOR2_X1 U4069 ( .A(n3203), .B(REG2_REG_6__SCAN_IN), .Z(n3204) );
  NAND2_X1 U4070 ( .A1(n3204), .A2(n4940), .ZN(n3205) );
  OAI21_X1 U4071 ( .B1(n4918), .B2(n3790), .A(n3205), .ZN(n3206) );
  NOR2_X1 U4072 ( .A1(n3340), .A2(n3206), .ZN(n3208) );
  NAND2_X1 U4073 ( .A1(n4914), .A2(n4872), .ZN(n3207) );
  OAI211_X1 U4074 ( .C1(n3209), .C2(n4908), .A(n3208), .B(n3207), .ZN(U3246)
         );
  XNOR2_X1 U4075 ( .A(n3210), .B(REG1_REG_3__SCAN_IN), .ZN(n3217) );
  XOR2_X1 U4076 ( .A(n3211), .B(REG2_REG_3__SCAN_IN), .Z(n3215) );
  AOI22_X1 U4077 ( .A1(n4930), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3212) );
  OAI21_X1 U4078 ( .B1(n4945), .B2(n3213), .A(n3212), .ZN(n3214) );
  AOI21_X1 U4079 ( .B1(n4940), .B2(n3215), .A(n3214), .ZN(n3216) );
  OAI21_X1 U4080 ( .B1(n3217), .B2(n4908), .A(n3216), .ZN(U3243) );
  NAND2_X1 U4081 ( .A1(n2698), .A2(n3968), .ZN(n4276) );
  AND2_X1 U4082 ( .A1(n3244), .A2(n4276), .ZN(n4234) );
  INV_X1 U4083 ( .A(n4234), .ZN(n4951) );
  INV_X1 U4084 ( .A(n3218), .ZN(n3219) );
  NOR2_X1 U4085 ( .A1(n3968), .A2(n3219), .ZN(n4949) );
  INV_X1 U4086 ( .A(n4704), .ZN(n3474) );
  OAI21_X1 U4087 ( .B1(n3474), .B2(n3145), .A(n4951), .ZN(n3220) );
  OAI21_X1 U4088 ( .B1(n3036), .B2(n4654), .A(n3220), .ZN(n4947) );
  AOI211_X1 U4089 ( .C1(n4995), .C2(n4951), .A(n4949), .B(n4947), .ZN(n4982)
         );
  NAND2_X1 U4090 ( .A1(n5019), .A2(REG1_REG_0__SCAN_IN), .ZN(n3221) );
  OAI21_X1 U4091 ( .B1(n4982), .B2(n5019), .A(n3221), .ZN(U3518) );
  XOR2_X1 U4092 ( .A(n3223), .B(n3222), .Z(n3227) );
  MUX2_X1 U4093 ( .A(REG2_REG_1__SCAN_IN), .B(n2544), .S(n3230), .Z(n3225) );
  AOI211_X1 U4094 ( .C1(n3225), .C2(n3224), .A(n2190), .B(n4905), .ZN(n3226)
         );
  AOI21_X1 U4095 ( .B1(n4942), .B2(n3227), .A(n3226), .ZN(n3229) );
  AOI22_X1 U4096 ( .A1(n4930), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3228) );
  OAI211_X1 U4097 ( .C1(n3230), .C2(n4945), .A(n3229), .B(n3228), .ZN(U3241)
         );
  NOR2_X1 U4098 ( .A1(n4930), .A2(U4043), .ZN(U3148) );
  AOI211_X1 U4099 ( .C1(n3232), .C2(n3231), .A(n2191), .B(n4908), .ZN(n3240)
         );
  AOI211_X1 U4100 ( .C1(n3233), .C2(n3235), .A(n3234), .B(n4905), .ZN(n3239)
         );
  AND2_X1 U4101 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3321) );
  AOI21_X1 U4102 ( .B1(n4930), .B2(ADDR_REG_5__SCAN_IN), .A(n3321), .ZN(n3236)
         );
  OAI21_X1 U4103 ( .B1(n4945), .B2(n3237), .A(n3236), .ZN(n3238) );
  OR3_X1 U4104 ( .A1(n3240), .A2(n3239), .A3(n3238), .ZN(U3245) );
  AOI21_X1 U4105 ( .B1(n3242), .B2(n3035), .A(n3241), .ZN(n3434) );
  NAND2_X1 U4106 ( .A1(n3110), .A2(n3244), .ZN(n3245) );
  NAND2_X1 U4107 ( .A1(n3243), .A2(n3245), .ZN(n3250) );
  NAND2_X1 U4108 ( .A1(n4672), .A2(n3035), .ZN(n3247) );
  NAND2_X1 U4109 ( .A1(n4696), .A2(n2698), .ZN(n3246) );
  OAI211_X1 U4110 ( .C1(n3248), .C2(n4654), .A(n3247), .B(n3246), .ZN(n3249)
         );
  AOI21_X1 U4111 ( .B1(n3250), .B2(n3145), .A(n3249), .ZN(n3255) );
  OR2_X1 U4112 ( .A1(n3251), .A2(n3110), .ZN(n3252) );
  AND2_X1 U4113 ( .A1(n3253), .A2(n3252), .ZN(n3429) );
  NAND2_X1 U4114 ( .A1(n3429), .A2(n3474), .ZN(n3254) );
  NAND2_X1 U4115 ( .A1(n3255), .A2(n3254), .ZN(n3430) );
  INV_X1 U4116 ( .A(n3429), .ZN(n3256) );
  NOR2_X1 U4117 ( .A1(n3256), .A2(n4987), .ZN(n3257) );
  AOI211_X1 U4118 ( .C1(n3434), .C2(n4998), .A(n3430), .B(n3257), .ZN(n4984)
         );
  NAND2_X1 U4119 ( .A1(n5019), .A2(REG1_REG_1__SCAN_IN), .ZN(n3258) );
  OAI21_X1 U4120 ( .B1(n4984), .B2(n5019), .A(n3258), .ZN(U3519) );
  XNOR2_X1 U4121 ( .A(n4871), .B(n5020), .ZN(n3259) );
  XNOR2_X1 U4122 ( .A(n3260), .B(n3259), .ZN(n3268) );
  NAND2_X1 U4123 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3514) );
  NAND2_X1 U4124 ( .A1(n4930), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3261) );
  OAI211_X1 U4125 ( .C1(n4945), .C2(n3262), .A(n3514), .B(n3261), .ZN(n3267)
         );
  AOI211_X1 U4126 ( .C1(n3265), .C2(n3264), .A(n4905), .B(n3263), .ZN(n3266)
         );
  AOI211_X1 U4127 ( .C1(n3268), .C2(n4942), .A(n3267), .B(n3266), .ZN(n3269)
         );
  INV_X1 U4128 ( .A(n3269), .ZN(U3247) );
  INV_X1 U4129 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3815) );
  NAND2_X1 U4130 ( .A1(n3270), .A2(REG1_REG_31__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4131 ( .A1(n2136), .A2(REG2_REG_31__SCAN_IN), .ZN(n3272) );
  NAND2_X1 U4132 ( .A1(n2732), .A2(REG0_REG_31__SCAN_IN), .ZN(n3271) );
  NAND3_X1 U4133 ( .A1(n3273), .A2(n3272), .A3(n3271), .ZN(n4376) );
  NAND2_X1 U4134 ( .A1(U4043), .A2(n4376), .ZN(n3274) );
  OAI21_X1 U4135 ( .B1(U4043), .B2(n3815), .A(n3274), .ZN(U3581) );
  INV_X1 U4136 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3776) );
  INV_X1 U4137 ( .A(REG1_REG_30__SCAN_IN), .ZN(n3716) );
  NAND2_X1 U4138 ( .A1(n2136), .A2(REG2_REG_30__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4139 ( .A1(n2732), .A2(REG0_REG_30__SCAN_IN), .ZN(n3275) );
  OAI211_X1 U4140 ( .C1(n3277), .C2(n3716), .A(n3276), .B(n3275), .ZN(n4399)
         );
  NAND2_X1 U4141 ( .A1(U4043), .A2(n4399), .ZN(n3278) );
  OAI21_X1 U4142 ( .B1(U4043), .B2(n3776), .A(n3278), .ZN(U3580) );
  INV_X1 U4143 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3804) );
  NAND2_X1 U4144 ( .A1(U4043), .A2(n4695), .ZN(n3279) );
  OAI21_X1 U4145 ( .B1(U4043), .B2(n3804), .A(n3279), .ZN(U3562) );
  XNOR2_X1 U4146 ( .A(n3280), .B(n3493), .ZN(n3289) );
  INV_X1 U4147 ( .A(n3281), .ZN(n3282) );
  OAI211_X1 U4148 ( .C1(REG1_REG_8__SCAN_IN), .C2(n3283), .A(n3282), .B(n4942), 
        .ZN(n3288) );
  NAND2_X1 U4149 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3442) );
  INV_X1 U4150 ( .A(n3442), .ZN(n3286) );
  NOR2_X1 U4151 ( .A1(n4945), .A2(n3284), .ZN(n3285) );
  AOI211_X1 U4152 ( .C1(n4930), .C2(ADDR_REG_8__SCAN_IN), .A(n3286), .B(n3285), 
        .ZN(n3287) );
  OAI211_X1 U4153 ( .C1(n3289), .C2(n4905), .A(n3288), .B(n3287), .ZN(U3248)
         );
  INV_X1 U4154 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n3802) );
  NAND2_X1 U4155 ( .A1(n4058), .A2(U4043), .ZN(n3290) );
  OAI21_X1 U4156 ( .B1(U4043), .B2(n3802), .A(n3290), .ZN(U3563) );
  INV_X1 U4157 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4158 ( .A1(n4035), .A2(U4043), .ZN(n3291) );
  OAI21_X1 U4159 ( .B1(U4043), .B2(n3779), .A(n3291), .ZN(U3568) );
  INV_X1 U4160 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n3813) );
  NAND2_X1 U4161 ( .A1(n3441), .A2(U4043), .ZN(n3292) );
  OAI21_X1 U4162 ( .B1(U4043), .B2(n3813), .A(n3292), .ZN(U3557) );
  INV_X1 U4163 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U4164 ( .A1(n4590), .A2(U4043), .ZN(n3293) );
  OAI21_X1 U4165 ( .B1(U4043), .B2(n3805), .A(n3293), .ZN(U3567) );
  INV_X1 U4166 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U4167 ( .A1(n3606), .A2(U4043), .ZN(n3294) );
  OAI21_X1 U4168 ( .B1(U4043), .B2(n3746), .A(n3294), .ZN(U3558) );
  INV_X1 U4169 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n3750) );
  NAND2_X1 U4170 ( .A1(U4043), .A2(n3475), .ZN(n3295) );
  OAI21_X1 U4171 ( .B1(U4043), .B2(n3750), .A(n3295), .ZN(U3553) );
  INV_X1 U4172 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U4173 ( .A1(n3551), .A2(U4043), .ZN(n3296) );
  OAI21_X1 U4174 ( .B1(U4043), .B2(n3749), .A(n3296), .ZN(U3552) );
  INV_X1 U4175 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4176 ( .A1(n4519), .A2(U4043), .ZN(n3297) );
  OAI21_X1 U4177 ( .B1(U4043), .B2(n3744), .A(n3297), .ZN(U3573) );
  XNOR2_X1 U4178 ( .A(n3298), .B(n3299), .ZN(n3308) );
  INV_X1 U4179 ( .A(n3300), .ZN(n3303) );
  NAND3_X1 U4180 ( .A1(n3303), .A2(n3302), .A3(n3301), .ZN(n3963) );
  AOI22_X1 U4181 ( .A1(n4192), .A2(n2698), .B1(n4165), .B2(n3551), .ZN(n3304)
         );
  OAI21_X1 U4182 ( .B1(n4180), .B2(n3305), .A(n3304), .ZN(n3306) );
  AOI21_X1 U4183 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3963), .A(n3306), .ZN(n3307)
         );
  OAI21_X1 U4184 ( .B1(n3308), .B2(n4199), .A(n3307), .ZN(U3219) );
  INV_X1 U4185 ( .A(n3310), .ZN(n3311) );
  AOI21_X1 U4186 ( .B1(n3309), .B2(n3312), .A(n3311), .ZN(n3316) );
  AOI22_X1 U4187 ( .A1(n4192), .A2(n2251), .B1(n4165), .B2(n3475), .ZN(n3313)
         );
  OAI21_X1 U4188 ( .B1(n4180), .B2(n3374), .A(n3313), .ZN(n3314) );
  AOI21_X1 U4189 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3963), .A(n3314), .ZN(n3315)
         );
  OAI21_X1 U4190 ( .B1(n3316), .B2(n4199), .A(n3315), .ZN(U3234) );
  INV_X1 U4191 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n3794) );
  NAND2_X1 U4192 ( .A1(n4498), .A2(U4043), .ZN(n3317) );
  OAI21_X1 U4193 ( .B1(U4043), .B2(n3794), .A(n3317), .ZN(U3574) );
  XNOR2_X1 U4194 ( .A(n3319), .B(n3318), .ZN(n3324) );
  OAI22_X1 U4195 ( .A1(n4180), .A2(n3404), .B1(n3053), .B2(n4169), .ZN(n3320)
         );
  AOI211_X1 U4196 ( .C1(n4165), .C2(n4356), .A(n3321), .B(n3320), .ZN(n3323)
         );
  NAND2_X1 U4197 ( .A1(n4196), .A2(n3511), .ZN(n3322) );
  OAI211_X1 U4198 ( .C1(n3324), .C2(n4199), .A(n3323), .B(n3322), .ZN(U3224)
         );
  NAND2_X1 U4199 ( .A1(n3325), .A2(n4102), .ZN(n3333) );
  AOI21_X1 U4200 ( .B1(n3326), .B2(n3328), .A(n3327), .ZN(n3332) );
  AOI22_X1 U4201 ( .A1(n4192), .A2(n3475), .B1(n4191), .B2(n3482), .ZN(n3329)
         );
  NAND2_X1 U4202 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4885) );
  OAI211_X1 U4203 ( .C1(n3478), .C2(n4194), .A(n3329), .B(n4885), .ZN(n3330)
         );
  AOI21_X1 U4204 ( .B1(n3483), .B2(n4196), .A(n3330), .ZN(n3331) );
  OAI21_X1 U4205 ( .B1(n3333), .B2(n3332), .A(n3331), .ZN(U3227) );
  INV_X1 U4206 ( .A(n3335), .ZN(n3337) );
  NOR2_X1 U4207 ( .A1(n3337), .A2(n3336), .ZN(n3338) );
  XNOR2_X1 U4208 ( .A(n3334), .B(n3338), .ZN(n3343) );
  OAI22_X1 U4209 ( .A1(n4180), .A2(n3616), .B1(n3478), .B2(n4169), .ZN(n3339)
         );
  AOI211_X1 U4210 ( .C1(n4165), .C2(n3441), .A(n3340), .B(n3339), .ZN(n3342)
         );
  NAND2_X1 U4211 ( .A1(n4196), .A2(n3564), .ZN(n3341) );
  OAI211_X1 U4212 ( .C1(n3343), .C2(n4199), .A(n3342), .B(n3341), .ZN(U3236)
         );
  XOR2_X1 U4213 ( .A(n3345), .B(n3344), .Z(n3353) );
  AND2_X1 U4214 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3597) );
  AOI21_X1 U4215 ( .B1(n4930), .B2(ADDR_REG_9__SCAN_IN), .A(n3597), .ZN(n3346)
         );
  OAI21_X1 U4216 ( .B1(n4945), .B2(n3347), .A(n3346), .ZN(n3352) );
  AOI211_X1 U4217 ( .C1(n3350), .C2(n3349), .A(n4908), .B(n3348), .ZN(n3351)
         );
  AOI211_X1 U4218 ( .C1(n4940), .C2(n3353), .A(n3352), .B(n3351), .ZN(n3354)
         );
  INV_X1 U4219 ( .A(n3354), .ZN(U3249) );
  OAI21_X1 U4220 ( .B1(n3356), .B2(n3355), .A(n3326), .ZN(n3360) );
  MUX2_X1 U4221 ( .A(STATE_REG_SCAN_IN), .B(n4108), .S(n3556), .Z(n3358) );
  AOI22_X1 U4222 ( .A1(n4192), .A2(n3551), .B1(n4165), .B2(n3040), .ZN(n3357)
         );
  OAI211_X1 U4223 ( .C1(n4180), .C2(n3047), .A(n3358), .B(n3357), .ZN(n3359)
         );
  AOI21_X1 U4224 ( .B1(n4102), .B2(n3360), .A(n3359), .ZN(n3361) );
  INV_X1 U4225 ( .A(n3361), .ZN(U3215) );
  NAND2_X1 U4226 ( .A1(n3363), .A2(n4238), .ZN(n3364) );
  NAND2_X1 U4227 ( .A1(n3362), .A2(n3364), .ZN(n3453) );
  AOI22_X1 U4228 ( .A1(n2251), .A2(n4696), .B1(n3365), .B2(n4672), .ZN(n3366)
         );
  OAI21_X1 U4229 ( .B1(n3367), .B2(n4654), .A(n3366), .ZN(n3371) );
  NAND3_X1 U4230 ( .A1(n3038), .A2(n3113), .A3(n3243), .ZN(n3368) );
  AOI21_X1 U4231 ( .B1(n3369), .B2(n3368), .A(n4661), .ZN(n3370) );
  AOI211_X1 U4232 ( .C1(n3474), .C2(n3453), .A(n3371), .B(n3370), .ZN(n3450)
         );
  INV_X1 U4233 ( .A(n3450), .ZN(n3372) );
  AOI21_X1 U4234 ( .B1(n4995), .B2(n3453), .A(n3372), .ZN(n3389) );
  OR2_X1 U4235 ( .A1(n3241), .A2(n3374), .ZN(n3375) );
  NAND2_X1 U4236 ( .A1(n3373), .A2(n3375), .ZN(n3455) );
  INV_X1 U4237 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3376) );
  OAI22_X1 U4238 ( .A1(n4856), .A2(n3455), .B1(n5013), .B2(n3376), .ZN(n3377)
         );
  INV_X1 U4239 ( .A(n3377), .ZN(n3378) );
  OAI21_X1 U4240 ( .B1(n3389), .B2(n5011), .A(n3378), .ZN(U3471) );
  XNOR2_X1 U4241 ( .A(n3379), .B(REG2_REG_10__SCAN_IN), .ZN(n3386) );
  OAI211_X1 U4242 ( .C1(n3381), .C2(REG1_REG_10__SCAN_IN), .A(n3380), .B(n4942), .ZN(n3385) );
  NOR2_X1 U4243 ( .A1(STATE_REG_SCAN_IN), .A2(n3382), .ZN(n3646) );
  NOR2_X1 U4244 ( .A1(n4945), .A2(n2200), .ZN(n3383) );
  AOI211_X1 U4245 ( .C1(n4930), .C2(ADDR_REG_10__SCAN_IN), .A(n3646), .B(n3383), .ZN(n3384) );
  OAI211_X1 U4246 ( .C1(n3386), .C2(n4905), .A(n3385), .B(n3384), .ZN(U3250)
         );
  INV_X1 U4247 ( .A(n4794), .ZN(n4766) );
  INV_X1 U4248 ( .A(n3455), .ZN(n3387) );
  AOI22_X1 U4249 ( .A1(n4766), .A2(n3387), .B1(n5019), .B2(REG1_REG_2__SCAN_IN), .ZN(n3388) );
  OAI21_X1 U4250 ( .B1(n3389), .B2(n5019), .A(n3388), .ZN(U3520) );
  AND2_X1 U4251 ( .A1(n4290), .A2(n4298), .ZN(n4233) );
  XNOR2_X1 U4252 ( .A(n3390), .B(n4233), .ZN(n3489) );
  XNOR2_X1 U4253 ( .A(n3391), .B(n4233), .ZN(n3395) );
  OAI22_X1 U4254 ( .A1(n3392), .A2(n3157), .B1(n3444), .B2(n4654), .ZN(n3393)
         );
  AOI21_X1 U4255 ( .B1(n3440), .B2(n4672), .A(n3393), .ZN(n3394) );
  OAI21_X1 U4256 ( .B1(n3395), .B2(n4661), .A(n3394), .ZN(n3490) );
  AOI21_X1 U4257 ( .B1(n3489), .B2(n4787), .A(n3490), .ZN(n3409) );
  AOI21_X1 U4258 ( .B1(n3440), .B2(n3611), .A(n2188), .ZN(n3495) );
  INV_X1 U4259 ( .A(n4856), .ZN(n4836) );
  AOI22_X1 U4260 ( .A1(n3495), .A2(n4836), .B1(REG0_REG_8__SCAN_IN), .B2(n5011), .ZN(n3396) );
  OAI21_X1 U4261 ( .B1(n3409), .B2(n5011), .A(n3396), .ZN(U3483) );
  AND2_X1 U4262 ( .A1(n4286), .A2(n4301), .ZN(n4244) );
  XNOR2_X1 U4263 ( .A(n3397), .B(n4244), .ZN(n3568) );
  XOR2_X1 U4264 ( .A(n3398), .B(n4244), .Z(n3402) );
  OAI22_X1 U4265 ( .A1(n3478), .A2(n3157), .B1(n4700), .B2(n3616), .ZN(n3399)
         );
  AOI21_X1 U4266 ( .B1(n4697), .B2(n3441), .A(n3399), .ZN(n3401) );
  NAND2_X1 U4267 ( .A1(n3568), .A2(n3474), .ZN(n3400) );
  OAI211_X1 U4268 ( .C1(n3402), .C2(n4661), .A(n3401), .B(n3400), .ZN(n3562)
         );
  AOI21_X1 U4269 ( .B1(n4995), .B2(n3568), .A(n3562), .ZN(n3411) );
  AND2_X1 U4270 ( .A1(n3403), .A2(n3404), .ZN(n3510) );
  INV_X1 U4271 ( .A(n3510), .ZN(n3405) );
  AOI21_X1 U4272 ( .B1(n3406), .B2(n3405), .A(n3170), .ZN(n3563) );
  AOI22_X1 U4273 ( .A1(n3563), .A2(n4836), .B1(n5011), .B2(REG0_REG_6__SCAN_IN), .ZN(n3407) );
  OAI21_X1 U4274 ( .B1(n3411), .B2(n5011), .A(n3407), .ZN(U3479) );
  AOI22_X1 U4275 ( .A1(n3495), .A2(n4766), .B1(REG1_REG_8__SCAN_IN), .B2(n5019), .ZN(n3408) );
  OAI21_X1 U4276 ( .B1(n3409), .B2(n5019), .A(n3408), .ZN(U3526) );
  AOI22_X1 U4277 ( .A1(n3563), .A2(n4766), .B1(n5019), .B2(REG1_REG_6__SCAN_IN), .ZN(n3410) );
  OAI21_X1 U4278 ( .B1(n3411), .B2(n5019), .A(n3410), .ZN(U3524) );
  INV_X1 U4279 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4280 ( .A1(n4268), .A2(U4043), .ZN(n3412) );
  OAI21_X1 U4281 ( .B1(U4043), .B2(n3747), .A(n3412), .ZN(U3577) );
  AOI211_X1 U4282 ( .C1(n3414), .C2(n3413), .A(n4905), .B(n2183), .ZN(n3418)
         );
  NAND2_X1 U4283 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4167) );
  NAND2_X1 U4284 ( .A1(n4930), .A2(ADDR_REG_11__SCAN_IN), .ZN(n3415) );
  OAI211_X1 U4285 ( .C1(n4945), .C2(n3416), .A(n4167), .B(n3415), .ZN(n3417)
         );
  NOR2_X1 U4286 ( .A1(n3418), .A2(n3417), .ZN(n3423) );
  OAI211_X1 U4287 ( .C1(n3421), .C2(n3420), .A(n3419), .B(n4942), .ZN(n3422)
         );
  NAND2_X1 U4288 ( .A1(n3423), .A2(n3422), .ZN(U3251) );
  NAND2_X1 U4289 ( .A1(n3425), .A2(n3424), .ZN(n3426) );
  AND2_X1 U4290 ( .A1(n4652), .A2(n4341), .ZN(n4600) );
  OR2_X1 U4291 ( .A1(n2686), .A2(n4341), .ZN(n3487) );
  INV_X1 U4292 ( .A(n3487), .ZN(n3428) );
  NAND2_X1 U4293 ( .A1(n4952), .A2(n3429), .ZN(n3432) );
  AOI22_X1 U4294 ( .A1(n4955), .A2(n3430), .B1(REG3_REG_1__SCAN_IN), .B2(n4950), .ZN(n3431) );
  OAI211_X1 U4295 ( .C1(n4955), .C2(n2544), .A(n3432), .B(n3431), .ZN(n3433)
         );
  AOI21_X1 U4296 ( .B1(n4668), .B2(n3434), .A(n3433), .ZN(n3435) );
  INV_X1 U4297 ( .A(n3435), .ZN(U3289) );
  XOR2_X1 U4298 ( .A(n3437), .B(n3436), .Z(n3438) );
  XNOR2_X1 U4299 ( .A(n3439), .B(n3438), .ZN(n3447) );
  AOI22_X1 U4300 ( .A1(n4192), .A2(n3441), .B1(n4191), .B2(n3440), .ZN(n3443)
         );
  OAI211_X1 U4301 ( .C1(n3444), .C2(n4194), .A(n3443), .B(n3442), .ZN(n3445)
         );
  AOI21_X1 U4302 ( .B1(n3491), .B2(n4196), .A(n3445), .ZN(n3446) );
  OAI21_X1 U4303 ( .B1(n3447), .B2(n4199), .A(n3446), .ZN(U3218) );
  INV_X1 U4304 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3448) );
  OAI22_X1 U4305 ( .A1(n4955), .A2(n3449), .B1(n3448), .B2(n4649), .ZN(n3452)
         );
  NOR2_X1 U4306 ( .A1(n3450), .A2(n2132), .ZN(n3451) );
  AOI211_X1 U4307 ( .C1(n4952), .C2(n3453), .A(n3452), .B(n3451), .ZN(n3454)
         );
  OAI21_X1 U4308 ( .B1(n4711), .B2(n3455), .A(n3454), .ZN(U3288) );
  INV_X1 U4309 ( .A(n4303), .ZN(n4294) );
  AND2_X1 U4310 ( .A1(n4294), .A2(n4291), .ZN(n4246) );
  XNOR2_X1 U4311 ( .A(n3456), .B(n4246), .ZN(n3528) );
  XNOR2_X1 U4312 ( .A(n3457), .B(n4246), .ZN(n3460) );
  OAI22_X1 U4313 ( .A1(n4700), .A2(n3595), .B1(n4170), .B2(n4654), .ZN(n3458)
         );
  AOI21_X1 U4314 ( .B1(n4696), .B2(n3606), .A(n3458), .ZN(n3459) );
  OAI21_X1 U4315 ( .B1(n3460), .B2(n4661), .A(n3459), .ZN(n3524) );
  AOI21_X1 U4316 ( .B1(n3528), .B2(n4787), .A(n3524), .ZN(n3466) );
  NOR2_X1 U4317 ( .A1(n2188), .A2(n3595), .ZN(n3462) );
  OR2_X1 U4318 ( .A1(n3461), .A2(n3462), .ZN(n3526) );
  INV_X1 U4319 ( .A(n3526), .ZN(n3464) );
  AOI22_X1 U4320 ( .A1(n3464), .A2(n4766), .B1(REG1_REG_9__SCAN_IN), .B2(n5019), .ZN(n3463) );
  OAI21_X1 U4321 ( .B1(n3466), .B2(n5019), .A(n3463), .ZN(U3527) );
  AOI22_X1 U4322 ( .A1(n3464), .A2(n4836), .B1(REG0_REG_9__SCAN_IN), .B2(n5011), .ZN(n3465) );
  OAI21_X1 U4323 ( .B1(n3466), .B2(n5011), .A(n3465), .ZN(U3485) );
  INV_X1 U4324 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4325 ( .A1(n4406), .A2(U4043), .ZN(n3467) );
  OAI21_X1 U4326 ( .B1(U4043), .B2(n3801), .A(n3467), .ZN(U3578) );
  XNOR2_X1 U4327 ( .A(n3468), .B(n4239), .ZN(n3480) );
  NAND2_X1 U4328 ( .A1(n3362), .A2(n3469), .ZN(n3471) );
  AND2_X1 U4329 ( .A1(n3471), .A2(n3470), .ZN(n3472) );
  OR2_X1 U4330 ( .A1(n3472), .A2(n4239), .ZN(n3500) );
  NAND2_X1 U4331 ( .A1(n3472), .A2(n4239), .ZN(n3473) );
  AND2_X1 U4332 ( .A1(n3500), .A2(n3473), .ZN(n4996) );
  NAND2_X1 U4333 ( .A1(n4996), .A2(n3474), .ZN(n3477) );
  AOI22_X1 U4334 ( .A1(n4696), .A2(n3475), .B1(n4672), .B2(n3482), .ZN(n3476)
         );
  OAI211_X1 U4335 ( .C1(n3478), .C2(n4654), .A(n3477), .B(n3476), .ZN(n3479)
         );
  AOI21_X1 U4336 ( .B1(n3480), .B2(n3145), .A(n3479), .ZN(n4992) );
  INV_X1 U4337 ( .A(n4998), .ZN(n4986) );
  AOI211_X1 U4338 ( .C1(n3482), .C2(n3481), .A(n4986), .B(n3403), .ZN(n4994)
         );
  AOI22_X1 U4339 ( .A1(n4994), .A2(n4341), .B1(n4950), .B2(n3483), .ZN(n3484)
         );
  AND2_X1 U4340 ( .A1(n4992), .A2(n3484), .ZN(n3486) );
  AOI22_X1 U4341 ( .A1(n4996), .A2(n4952), .B1(REG2_REG_4__SCAN_IN), .B2(n2132), .ZN(n3485) );
  OAI21_X1 U4342 ( .B1(n3486), .B2(n2132), .A(n3485), .ZN(U3286) );
  NAND2_X1 U4343 ( .A1(n4704), .A2(n3487), .ZN(n3488) );
  INV_X1 U4344 ( .A(n3489), .ZN(n3498) );
  NAND2_X1 U4345 ( .A1(n3490), .A2(n4955), .ZN(n3497) );
  INV_X1 U4346 ( .A(n3491), .ZN(n3492) );
  OAI22_X1 U4347 ( .A1(n4652), .A2(n3493), .B1(n3492), .B2(n4649), .ZN(n3494)
         );
  AOI21_X1 U4348 ( .B1(n3495), .B2(n4668), .A(n3494), .ZN(n3496) );
  OAI211_X1 U4349 ( .C1(n4670), .C2(n3498), .A(n3497), .B(n3496), .ZN(U3282)
         );
  NAND2_X1 U4350 ( .A1(n3500), .A2(n3499), .ZN(n3501) );
  NAND2_X1 U4351 ( .A1(n2173), .A2(n4297), .ZN(n4237) );
  XNOR2_X1 U4352 ( .A(n3501), .B(n4237), .ZN(n5002) );
  XNOR2_X1 U4353 ( .A(n3502), .B(n4237), .ZN(n3506) );
  NAND2_X1 U4354 ( .A1(n4672), .A2(n3507), .ZN(n3504) );
  NAND2_X1 U4355 ( .A1(n4697), .A2(n4356), .ZN(n3503) );
  OAI211_X1 U4356 ( .C1(n3157), .C2(n3053), .A(n3504), .B(n3503), .ZN(n3505)
         );
  AOI21_X1 U4357 ( .B1(n3506), .B2(n3145), .A(n3505), .ZN(n5001) );
  MUX2_X1 U4358 ( .A(n5001), .B(n2555), .S(n2132), .Z(n3513) );
  INV_X1 U4359 ( .A(n3403), .ZN(n3508) );
  AND2_X1 U4360 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  NOR2_X1 U4361 ( .A1(n3510), .A2(n3509), .ZN(n4999) );
  AOI22_X1 U4362 ( .A1(n4668), .A2(n4999), .B1(n3511), .B2(n4950), .ZN(n3512)
         );
  OAI211_X1 U4363 ( .C1(n4670), .C2(n5002), .A(n3513), .B(n3512), .ZN(U3285)
         );
  AOI22_X1 U4364 ( .A1(n4192), .A2(n4356), .B1(n4191), .B2(n3609), .ZN(n3515)
         );
  OAI211_X1 U4365 ( .C1(n3516), .C2(n4194), .A(n3515), .B(n3514), .ZN(n3522)
         );
  INV_X1 U4366 ( .A(n3517), .ZN(n3518) );
  AOI211_X1 U4367 ( .C1(n3520), .C2(n3519), .A(n4199), .B(n3518), .ZN(n3521)
         );
  AOI211_X1 U4368 ( .C1(n3613), .C2(n4196), .A(n3522), .B(n3521), .ZN(n3523)
         );
  INV_X1 U4369 ( .A(n3523), .ZN(U3210) );
  INV_X1 U4370 ( .A(n3524), .ZN(n3530) );
  AOI22_X1 U4371 ( .A1(n2132), .A2(REG2_REG_9__SCAN_IN), .B1(n3598), .B2(n4950), .ZN(n3525) );
  OAI21_X1 U4372 ( .B1(n3526), .B2(n4711), .A(n3525), .ZN(n3527) );
  AOI21_X1 U4373 ( .B1(n3528), .B2(n4688), .A(n3527), .ZN(n3529) );
  OAI21_X1 U4374 ( .B1(n3530), .B2(n2132), .A(n3529), .ZN(U3281) );
  AND2_X1 U4375 ( .A1(n4305), .A2(n4308), .ZN(n4232) );
  XNOR2_X1 U4376 ( .A(n3531), .B(n4232), .ZN(n3532) );
  NAND2_X1 U4377 ( .A1(n3532), .A2(n3145), .ZN(n3534) );
  AOI22_X1 U4378 ( .A1(n4353), .A2(n4697), .B1(n4696), .B2(n4355), .ZN(n3533)
         );
  OAI211_X1 U4379 ( .C1(n4700), .C2(n3644), .A(n3534), .B(n3533), .ZN(n3585)
         );
  INV_X1 U4380 ( .A(n3585), .ZN(n3545) );
  XOR2_X1 U4381 ( .A(n3535), .B(n4232), .Z(n3586) );
  INV_X1 U4382 ( .A(n3461), .ZN(n3538) );
  INV_X1 U4383 ( .A(n3536), .ZN(n3537) );
  AOI21_X1 U4384 ( .B1(n3539), .B2(n3538), .A(n3537), .ZN(n3588) );
  INV_X1 U4385 ( .A(n3588), .ZN(n3542) );
  AOI22_X1 U4386 ( .A1(n2132), .A2(REG2_REG_10__SCAN_IN), .B1(n3540), .B2(
        n4950), .ZN(n3541) );
  OAI21_X1 U4387 ( .B1(n3542), .B2(n4711), .A(n3541), .ZN(n3543) );
  AOI21_X1 U4388 ( .B1(n3586), .B2(n4688), .A(n3543), .ZN(n3544) );
  OAI21_X1 U4389 ( .B1(n3545), .B2(n2132), .A(n3544), .ZN(U3280) );
  NAND2_X1 U4390 ( .A1(n3362), .A2(n3546), .ZN(n3547) );
  XNOR2_X1 U4391 ( .A(n3547), .B(n4245), .ZN(n4988) );
  OAI21_X1 U4392 ( .B1(n4245), .B2(n3549), .A(n3548), .ZN(n3554) );
  AOI22_X1 U4393 ( .A1(n3551), .A2(n4696), .B1(n4672), .B2(n3550), .ZN(n3552)
         );
  OAI21_X1 U4394 ( .B1(n3053), .B2(n4654), .A(n3552), .ZN(n3553) );
  AOI21_X1 U4395 ( .B1(n3554), .B2(n3145), .A(n3553), .ZN(n3555) );
  OAI21_X1 U4396 ( .B1(n4988), .B2(n4704), .A(n3555), .ZN(n4990) );
  INV_X1 U4397 ( .A(n4990), .ZN(n3561) );
  INV_X1 U4398 ( .A(n4988), .ZN(n3559) );
  OAI21_X1 U4399 ( .B1(n3168), .B2(n3047), .A(n3481), .ZN(n4985) );
  AOI22_X1 U4400 ( .A1(n2132), .A2(REG2_REG_3__SCAN_IN), .B1(n4950), .B2(n3556), .ZN(n3557) );
  OAI21_X1 U4401 ( .B1(n4711), .B2(n4985), .A(n3557), .ZN(n3558) );
  AOI21_X1 U4402 ( .B1(n4952), .B2(n3559), .A(n3558), .ZN(n3560) );
  OAI21_X1 U4403 ( .B1(n2132), .B2(n3561), .A(n3560), .ZN(U3287) );
  INV_X1 U4404 ( .A(n3562), .ZN(n3570) );
  INV_X1 U4405 ( .A(n3563), .ZN(n3566) );
  AOI22_X1 U4406 ( .A1(n2132), .A2(REG2_REG_6__SCAN_IN), .B1(n3564), .B2(n4950), .ZN(n3565) );
  OAI21_X1 U4407 ( .B1(n3566), .B2(n4711), .A(n3565), .ZN(n3567) );
  AOI21_X1 U4408 ( .B1(n3568), .B2(n4952), .A(n3567), .ZN(n3569) );
  OAI21_X1 U4409 ( .B1(n3570), .B2(n2132), .A(n3569), .ZN(U3284) );
  NAND2_X1 U4410 ( .A1(n3571), .A2(n4305), .ZN(n3572) );
  XOR2_X1 U4411 ( .A(n3572), .B(n4240), .Z(n3578) );
  OAI22_X1 U4412 ( .A1(n3573), .A2(n4700), .B1(n4170), .B2(n3157), .ZN(n3576)
         );
  AOI21_X1 U4413 ( .B1(n4240), .B2(n3574), .A(n2178), .ZN(n3579) );
  NOR2_X1 U4414 ( .A1(n3579), .A2(n4704), .ZN(n3575) );
  AOI211_X1 U4415 ( .C1(n4697), .C2(n4695), .A(n3576), .B(n3575), .ZN(n3577)
         );
  OAI21_X1 U4416 ( .B1(n4661), .B2(n3578), .A(n3577), .ZN(n4790) );
  INV_X1 U4417 ( .A(n4790), .ZN(n3584) );
  INV_X1 U4418 ( .A(n3579), .ZN(n4791) );
  NAND2_X1 U4419 ( .A1(n3536), .A2(n4166), .ZN(n3580) );
  NAND2_X1 U4420 ( .A1(n3632), .A2(n3580), .ZN(n4857) );
  AOI22_X1 U4421 ( .A1(n2132), .A2(REG2_REG_11__SCAN_IN), .B1(n4172), .B2(
        n4950), .ZN(n3581) );
  OAI21_X1 U4422 ( .B1(n4857), .B2(n4711), .A(n3581), .ZN(n3582) );
  AOI21_X1 U4423 ( .B1(n4791), .B2(n4952), .A(n3582), .ZN(n3583) );
  OAI21_X1 U4424 ( .B1(n3584), .B2(n2132), .A(n3583), .ZN(U3279) );
  AOI21_X1 U4425 ( .B1(n4787), .B2(n3586), .A(n3585), .ZN(n3590) );
  AOI22_X1 U4426 ( .A1(n3588), .A2(n4836), .B1(REG0_REG_10__SCAN_IN), .B2(
        n5011), .ZN(n3587) );
  OAI21_X1 U4427 ( .B1(n3590), .B2(n5011), .A(n3587), .ZN(U3487) );
  AOI22_X1 U4428 ( .A1(n3588), .A2(n4766), .B1(REG1_REG_10__SCAN_IN), .B2(
        n5019), .ZN(n3589) );
  OAI21_X1 U4429 ( .B1(n3590), .B2(n5019), .A(n3589), .ZN(U3528) );
  INV_X1 U4430 ( .A(n3592), .ZN(n3593) );
  AOI21_X1 U4431 ( .B1(n3594), .B2(n3591), .A(n3593), .ZN(n3601) );
  OAI22_X1 U4432 ( .A1(n4180), .A2(n3595), .B1(n4194), .B2(n4170), .ZN(n3596)
         );
  AOI211_X1 U4433 ( .C1(n4192), .C2(n3606), .A(n3597), .B(n3596), .ZN(n3600)
         );
  NAND2_X1 U4434 ( .A1(n4196), .A2(n3598), .ZN(n3599) );
  OAI211_X1 U4435 ( .C1(n3601), .C2(n4199), .A(n3600), .B(n3599), .ZN(U3228)
         );
  XNOR2_X1 U4436 ( .A(n3602), .B(n4249), .ZN(n3608) );
  OAI22_X1 U4437 ( .A1(n3604), .A2(n3157), .B1(n4700), .B2(n3603), .ZN(n3605)
         );
  AOI21_X1 U4438 ( .B1(n4697), .B2(n3606), .A(n3605), .ZN(n3607) );
  OAI21_X1 U4439 ( .B1(n3608), .B2(n4661), .A(n3607), .ZN(n5008) );
  INV_X1 U4440 ( .A(n5008), .ZN(n3625) );
  AOI21_X1 U4441 ( .B1(n3610), .B2(n3609), .A(n4986), .ZN(n3612) );
  AND2_X1 U4442 ( .A1(n3612), .A2(n3611), .ZN(n5009) );
  INV_X1 U4443 ( .A(n3613), .ZN(n3614) );
  OAI22_X1 U4444 ( .A1(n4955), .A2(n3615), .B1(n3614), .B2(n4649), .ZN(n3623)
         );
  OR2_X1 U4445 ( .A1(n3397), .A2(n4356), .ZN(n3619) );
  NAND2_X1 U4446 ( .A1(n3397), .A2(n4356), .ZN(n3617) );
  NAND2_X1 U4447 ( .A1(n3617), .A2(n3616), .ZN(n3618) );
  AND2_X1 U4448 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  NOR2_X1 U4449 ( .A1(n3620), .A2(n4249), .ZN(n5007) );
  INV_X1 U4450 ( .A(n3620), .ZN(n3621) );
  INV_X1 U4451 ( .A(n4249), .ZN(n4287) );
  NOR2_X1 U4452 ( .A1(n3621), .A2(n4287), .ZN(n5006) );
  NOR3_X1 U4453 ( .A1(n5007), .A2(n5006), .A3(n4670), .ZN(n3622) );
  AOI211_X1 U4454 ( .C1(n4600), .C2(n5009), .A(n3623), .B(n3622), .ZN(n3624)
         );
  OAI21_X1 U4455 ( .B1(n2132), .B2(n3625), .A(n3624), .ZN(U3283) );
  INV_X1 U4456 ( .A(n4691), .ZN(n3626) );
  AND2_X1 U4457 ( .A1(n3626), .A2(n4690), .ZN(n4257) );
  AND2_X1 U4458 ( .A1(n3627), .A2(n4309), .ZN(n4692) );
  XOR2_X1 U4459 ( .A(n4257), .B(n4692), .Z(n3630) );
  OAI22_X1 U4460 ( .A1(n4062), .A2(n3157), .B1(n4677), .B2(n4654), .ZN(n3628)
         );
  AOI21_X1 U4461 ( .B1(n4059), .B2(n4672), .A(n3628), .ZN(n3629) );
  OAI21_X1 U4462 ( .B1(n3630), .B2(n4661), .A(n3629), .ZN(n4785) );
  INV_X1 U4463 ( .A(n4785), .ZN(n3639) );
  XOR2_X1 U4464 ( .A(n3631), .B(n4257), .Z(n4786) );
  INV_X1 U4465 ( .A(n3632), .ZN(n3635) );
  INV_X1 U4466 ( .A(n4707), .ZN(n3633) );
  OAI21_X1 U4467 ( .B1(n3635), .B2(n3634), .A(n3633), .ZN(n4852) );
  AOI22_X1 U4468 ( .A1(n2132), .A2(REG2_REG_12__SCAN_IN), .B1(n4064), .B2(
        n4950), .ZN(n3636) );
  OAI21_X1 U4469 ( .B1(n4852), .B2(n4711), .A(n3636), .ZN(n3637) );
  AOI21_X1 U4470 ( .B1(n4786), .B2(n4688), .A(n3637), .ZN(n3638) );
  OAI21_X1 U4471 ( .B1(n3639), .B2(n2132), .A(n3638), .ZN(U3278) );
  AND2_X1 U4472 ( .A1(n3592), .A2(n3640), .ZN(n3643) );
  OAI211_X1 U4473 ( .C1(n3643), .C2(n3642), .A(n4102), .B(n3641), .ZN(n3648)
         );
  OAI22_X1 U4474 ( .A1(n4180), .A2(n3644), .B1(n4194), .B2(n4062), .ZN(n3645)
         );
  AOI211_X1 U4475 ( .C1(n4192), .C2(n4355), .A(n3646), .B(n3645), .ZN(n3647)
         );
  OAI211_X1 U4476 ( .C1(n4108), .C2(n3649), .A(n3648), .B(n3647), .ZN(U3214)
         );
  XNOR2_X1 U4477 ( .A(n3650), .B(REG2_REG_12__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4478 ( .A1(n3651), .A2(REG1_REG_12__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4479 ( .C1(n3651), .C2(REG1_REG_12__SCAN_IN), .A(n3937), .B(n4942), .ZN(n3654) );
  INV_X1 U4480 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4481 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4060) );
  OAI21_X1 U4482 ( .B1(n4918), .B2(n3726), .A(n4060), .ZN(n3652) );
  AOI21_X1 U4483 ( .B1(n4867), .B2(n4914), .A(n3652), .ZN(n3653) );
  OAI211_X1 U4484 ( .C1(n3655), .C2(n4905), .A(n3654), .B(n3653), .ZN(n3932)
         );
  INV_X1 U4485 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4826) );
  INV_X1 U4486 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3847) );
  NAND4_X1 U4487 ( .A1(REG0_REG_18__SCAN_IN), .A2(n4826), .A3(n3847), .A4(
        n4920), .ZN(n3656) );
  NOR3_X1 U4488 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG0_REG_11__SCAN_IN), .A3(
        n3656), .ZN(n3657) );
  INV_X1 U4489 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4846) );
  NAND3_X1 U4490 ( .A1(n3657), .A2(REG2_REG_11__SCAN_IN), .A3(n4846), .ZN(
        n3660) );
  NAND4_X1 U4491 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(n2792), .ZN(n3659) );
  INV_X1 U4492 ( .A(REG0_REG_16__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4493 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_17__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(n3842), .ZN(n3658) );
  NOR3_X1 U4494 ( .A1(n3660), .A2(n3659), .A3(n3658), .ZN(n3683) );
  NAND4_X1 U4495 ( .A1(REG1_REG_17__SCAN_IN), .A2(REG2_REG_2__SCAN_IN), .A3(
        n2860), .A4(n4898), .ZN(n3666) );
  INV_X1 U4496 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4497 ( .A1(n3875), .A2(n3906), .A3(n3493), .A4(n3922), .ZN(n3665)
         );
  INV_X1 U4498 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5004) );
  INV_X1 U4499 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4997) );
  NAND4_X1 U4500 ( .A1(REG2_REG_1__SCAN_IN), .A2(REG0_REG_12__SCAN_IN), .A3(
        REG2_REG_0__SCAN_IN), .A4(n4997), .ZN(n3661) );
  NOR2_X1 U4501 ( .A1(REG0_REG_6__SCAN_IN), .A2(n3661), .ZN(n3662) );
  NAND4_X1 U4502 ( .A1(n3663), .A2(REG1_REG_7__SCAN_IN), .A3(n5004), .A4(n3662), .ZN(n3664) );
  NOR3_X1 U4503 ( .A1(n3666), .A2(n3665), .A3(n3664), .ZN(n3682) );
  AND3_X1 U4504 ( .A1(n2585), .A2(n3735), .A3(n3732), .ZN(n3667) );
  NAND4_X1 U4505 ( .A1(n3669), .A2(n3668), .A3(IR_REG_9__SCAN_IN), .A4(n3667), 
        .ZN(n3672) );
  INV_X1 U4506 ( .A(IR_REG_22__SCAN_IN), .ZN(n3670) );
  NAND4_X1 U4507 ( .A1(n3670), .A2(DATAI_27_), .A3(DATAI_26_), .A4(DATAI_21_), 
        .ZN(n3671) );
  NOR2_X1 U4508 ( .A1(n3672), .A2(n3671), .ZN(n3675) );
  INV_X1 U4509 ( .A(DATAI_0_), .ZN(n3673) );
  AND4_X1 U4510 ( .A1(n3673), .A2(DATAO_REG_23__SCAN_IN), .A3(
        DATAO_REG_2__SCAN_IN), .A4(DATAO_REG_3__SCAN_IN), .ZN(n3674) );
  AND4_X1 U4511 ( .A1(n3675), .A2(n3747), .A3(n3746), .A4(n3674), .ZN(n3681)
         );
  INV_X1 U4512 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4805) );
  NAND4_X1 U4513 ( .A1(REG0_REG_24__SCAN_IN), .A2(n4805), .A3(n4728), .A4(
        n4736), .ZN(n3679) );
  INV_X1 U4514 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4822) );
  NAND4_X1 U4515 ( .A1(REG2_REG_21__SCAN_IN), .A2(n3862), .A3(n4822), .A4(
        n4752), .ZN(n3678) );
  INV_X1 U4516 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4517 ( .A1(REG1_REG_1__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .A3(
        ADDR_REG_12__SCAN_IN), .A4(n3715), .ZN(n3677) );
  NAND4_X1 U4518 ( .A1(REG0_REG_28__SCAN_IN), .A2(REG0_REG_27__SCAN_IN), .A3(
        n3720), .A4(n3716), .ZN(n3676) );
  NOR4_X1 U4519 ( .A1(n3679), .A2(n3678), .A3(n3677), .A4(n3676), .ZN(n3680)
         );
  NAND4_X1 U4520 ( .A1(n3683), .A2(n3682), .A3(n3681), .A4(n3680), .ZN(n3713)
         );
  NAND4_X1 U4521 ( .A1(REG1_REG_18__SCAN_IN), .A2(ADDR_REG_19__SCAN_IN), .A3(
        n4071), .A4(n4756), .ZN(n3684) );
  NOR4_X1 U4522 ( .A1(IR_REG_2__SCAN_IN), .A2(REG2_REG_28__SCAN_IN), .A3(
        REG2_REG_25__SCAN_IN), .A4(n3684), .ZN(n3707) );
  INV_X1 U4523 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3834) );
  NOR4_X1 U4524 ( .A1(REG2_REG_23__SCAN_IN), .A2(REG2_REG_22__SCAN_IN), .A3(
        n4975), .A4(n3834), .ZN(n3706) );
  NOR4_X1 U4525 ( .A1(ADDR_REG_6__SCAN_IN), .A2(ADDR_REG_13__SCAN_IN), .A3(
        ADDR_REG_0__SCAN_IN), .A4(n2226), .ZN(n3685) );
  NAND3_X1 U4526 ( .A1(IR_REG_19__SCAN_IN), .A2(DATAI_14_), .A3(n3685), .ZN(
        n3699) );
  INV_X1 U4527 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4904) );
  NOR4_X1 U4528 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .A3(
        REG3_REG_19__SCAN_IN), .A4(n4904), .ZN(n3686) );
  AND3_X1 U4529 ( .A1(IR_REG_18__SCAN_IN), .A2(n3686), .A3(DATAI_3_), .ZN(
        n3688) );
  NOR2_X1 U4530 ( .A1(DATAO_REG_18__SCAN_IN), .A2(DATAO_REG_30__SCAN_IN), .ZN(
        n3687) );
  NAND4_X1 U4531 ( .A1(n3688), .A2(n3687), .A3(IR_REG_12__SCAN_IN), .A4(
        IR_REG_30__SCAN_IN), .ZN(n3691) );
  INV_X1 U4532 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n3689) );
  INV_X1 U4533 ( .A(REG1_REG_31__SCAN_IN), .ZN(n3778) );
  NAND4_X1 U4534 ( .A1(n3689), .A2(n3805), .A3(n3778), .A4(IR_REG_15__SCAN_IN), 
        .ZN(n3690) );
  NOR2_X1 U4535 ( .A1(n3691), .A2(n3690), .ZN(n3697) );
  NAND4_X1 U4536 ( .A1(n3832), .A2(n4113), .A3(n4088), .A4(REG3_REG_3__SCAN_IN), .ZN(n3695) );
  INV_X1 U4537 ( .A(DATAI_25_), .ZN(n3692) );
  NAND4_X1 U4538 ( .A1(n3693), .A2(n3692), .A3(REG1_REG_0__SCAN_IN), .A4(
        REG2_REG_6__SCAN_IN), .ZN(n3694) );
  NOR2_X1 U4539 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  NAND4_X1 U4540 ( .A1(n3697), .A2(n3696), .A3(DATAO_REG_31__SCAN_IN), .A4(
        DATAO_REG_13__SCAN_IN), .ZN(n3698) );
  NOR2_X1 U4541 ( .A1(n3699), .A2(n3698), .ZN(n3705) );
  INV_X1 U4542 ( .A(n3700), .ZN(n3703) );
  NOR4_X1 U4543 ( .A1(REG2_REG_27__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .A3(
        REG2_REG_30__SCAN_IN), .A4(n4156), .ZN(n3701) );
  NAND3_X1 U4544 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG2_REG_19__SCAN_IN), .A3(
        n3701), .ZN(n3702) );
  NOR2_X1 U4545 ( .A1(n3703), .A2(n3702), .ZN(n3704) );
  AND4_X1 U4546 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3711)
         );
  INV_X1 U4547 ( .A(DATAI_12_), .ZN(n3708) );
  NOR4_X1 U4548 ( .A1(DATAO_REG_28__SCAN_IN), .A2(DATAI_31_), .A3(
        DATAO_REG_7__SCAN_IN), .A4(n3708), .ZN(n3710) );
  INV_X1 U4549 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4917) );
  NOR4_X1 U4550 ( .A1(REG3_REG_27__SCAN_IN), .A2(DATAO_REG_24__SCAN_IN), .A3(
        n4917), .A4(n3804), .ZN(n3709) );
  NAND3_X1 U4551 ( .A1(n3711), .A2(n3710), .A3(n3709), .ZN(n3712) );
  OAI21_X1 U4552 ( .B1(n3713), .B2(n3712), .A(IR_REG_26__SCAN_IN), .ZN(n3829)
         );
  AOI22_X1 U4553 ( .A1(n3716), .A2(keyinput47), .B1(keyinput51), .B2(n3715), 
        .ZN(n3714) );
  OAI221_X1 U4554 ( .B1(n3716), .B2(keyinput47), .C1(n3715), .C2(keyinput51), 
        .A(n3714), .ZN(n3717) );
  INV_X1 U4555 ( .A(n3717), .ZN(n3730) );
  INV_X1 U4556 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4557 ( .A1(n3720), .A2(keyinput117), .B1(n3719), .B2(keyinput109), 
        .ZN(n3718) );
  OAI221_X1 U4558 ( .B1(n3720), .B2(keyinput117), .C1(n3719), .C2(keyinput109), 
        .A(n3718), .ZN(n3721) );
  INV_X1 U4559 ( .A(n3721), .ZN(n3729) );
  XNOR2_X1 U4560 ( .A(IR_REG_11__SCAN_IN), .B(keyinput38), .ZN(n3724) );
  XNOR2_X1 U4561 ( .A(REG1_REG_1__SCAN_IN), .B(keyinput69), .ZN(n3723) );
  XNOR2_X1 U4562 ( .A(IR_REG_3__SCAN_IN), .B(keyinput42), .ZN(n3722) );
  AND3_X1 U4563 ( .A1(n3724), .A2(n3723), .A3(n3722), .ZN(n3728) );
  INV_X1 U4564 ( .A(keyinput71), .ZN(n3725) );
  XNOR2_X1 U4565 ( .A(n3726), .B(n3725), .ZN(n3727) );
  AND4_X1 U4566 ( .A1(n3730), .A2(n3729), .A3(n3728), .A4(n3727), .ZN(n3774)
         );
  INV_X1 U4567 ( .A(DATAI_27_), .ZN(n3733) );
  AOI22_X1 U4568 ( .A1(n3733), .A2(keyinput15), .B1(keyinput31), .B2(n3732), 
        .ZN(n3731) );
  OAI221_X1 U4569 ( .B1(n3733), .B2(keyinput15), .C1(n3732), .C2(keyinput31), 
        .A(n3731), .ZN(n3742) );
  INV_X1 U4570 ( .A(D_REG_24__SCAN_IN), .ZN(n4961) );
  INV_X1 U4571 ( .A(D_REG_30__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U4572 ( .A1(n4961), .A2(keyinput19), .B1(keyinput3), .B2(n4957), 
        .ZN(n3734) );
  OAI221_X1 U4573 ( .B1(n4961), .B2(keyinput19), .C1(n4957), .C2(keyinput3), 
        .A(n3734), .ZN(n3741) );
  XOR2_X1 U4574 ( .A(n3735), .B(keyinput39), .Z(n3739) );
  XNOR2_X1 U4575 ( .A(keyinput116), .B(IR_REG_27__SCAN_IN), .ZN(n3738) );
  XNOR2_X1 U4576 ( .A(IR_REG_5__SCAN_IN), .B(keyinput23), .ZN(n3737) );
  XNOR2_X1 U4577 ( .A(IR_REG_9__SCAN_IN), .B(keyinput11), .ZN(n3736) );
  NAND4_X1 U4578 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  NOR3_X1 U4579 ( .A1(n3742), .A2(n3741), .A3(n3740), .ZN(n3773) );
  INV_X1 U4580 ( .A(D_REG_12__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U4581 ( .A1(n4968), .A2(keyinput29), .B1(keyinput28), .B2(n3744), 
        .ZN(n3743) );
  OAI221_X1 U4582 ( .B1(n4968), .B2(keyinput29), .C1(n3744), .C2(keyinput28), 
        .A(n3743), .ZN(n3757) );
  AOI22_X1 U4583 ( .A1(n3747), .A2(keyinput63), .B1(keyinput103), .B2(n3746), 
        .ZN(n3745) );
  OAI221_X1 U4584 ( .B1(n3747), .B2(keyinput63), .C1(n3746), .C2(keyinput103), 
        .A(n3745), .ZN(n3756) );
  AOI22_X1 U4585 ( .A1(n3750), .A2(keyinput119), .B1(keyinput107), .B2(n3749), 
        .ZN(n3748) );
  OAI221_X1 U4586 ( .B1(n3750), .B2(keyinput119), .C1(n3749), .C2(keyinput107), 
        .A(n3748), .ZN(n3755) );
  XOR2_X1 U4587 ( .A(n3751), .B(keyinput55), .Z(n3753) );
  XNOR2_X1 U4588 ( .A(DATAI_0_), .B(keyinput123), .ZN(n3752) );
  NAND2_X1 U4589 ( .A1(n3753), .A2(n3752), .ZN(n3754) );
  NOR4_X1 U4590 ( .A1(n3757), .A2(n3756), .A3(n3755), .A4(n3754), .ZN(n3772)
         );
  INV_X1 U4591 ( .A(D_REG_21__SCAN_IN), .ZN(n4963) );
  INV_X1 U4592 ( .A(DATAI_26_), .ZN(n3759) );
  AOI22_X1 U4593 ( .A1(n4963), .A2(keyinput20), .B1(keyinput24), .B2(n3759), 
        .ZN(n3758) );
  OAI221_X1 U4594 ( .B1(n4963), .B2(keyinput20), .C1(n3759), .C2(keyinput24), 
        .A(n3758), .ZN(n3760) );
  INV_X1 U4595 ( .A(n3760), .ZN(n3770) );
  INV_X1 U4596 ( .A(keyinput0), .ZN(n3761) );
  XNOR2_X1 U4597 ( .A(n4904), .B(n3761), .ZN(n3769) );
  INV_X1 U4598 ( .A(D_REG_10__SCAN_IN), .ZN(n4969) );
  INV_X1 U4599 ( .A(keyinput34), .ZN(n3762) );
  XNOR2_X1 U4600 ( .A(n4969), .B(n3762), .ZN(n3768) );
  XNOR2_X1 U4601 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput37), .ZN(n3766) );
  XNOR2_X1 U4602 ( .A(IR_REG_22__SCAN_IN), .B(keyinput33), .ZN(n3765) );
  XNOR2_X1 U4603 ( .A(IR_REG_13__SCAN_IN), .B(keyinput17), .ZN(n3764) );
  XNOR2_X1 U4604 ( .A(IR_REG_6__SCAN_IN), .B(keyinput9), .ZN(n3763) );
  AND4_X1 U4605 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3767)
         );
  AND4_X1 U4606 ( .A1(n3770), .A2(n3769), .A3(n3768), .A4(n3767), .ZN(n3771)
         );
  NAND4_X1 U4607 ( .A1(n3774), .A2(n3773), .A3(n3772), .A4(n3771), .ZN(n3828)
         );
  INV_X1 U4608 ( .A(D_REG_5__SCAN_IN), .ZN(n4970) );
  AOI22_X1 U4609 ( .A1(n4970), .A2(keyinput122), .B1(keyinput125), .B2(n3776), 
        .ZN(n3775) );
  OAI221_X1 U4610 ( .B1(n4970), .B2(keyinput122), .C1(n3776), .C2(keyinput125), 
        .A(n3775), .ZN(n3787) );
  AOI22_X1 U4611 ( .A1(n3779), .A2(keyinput18), .B1(n3778), .B2(keyinput21), 
        .ZN(n3777) );
  OAI221_X1 U4612 ( .B1(n3779), .B2(keyinput18), .C1(n3778), .C2(keyinput21), 
        .A(n3777), .ZN(n3786) );
  INV_X1 U4613 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n3780) );
  XOR2_X1 U4614 ( .A(n3780), .B(keyinput114), .Z(n3784) );
  XNOR2_X1 U4615 ( .A(DATAI_25_), .B(keyinput13), .ZN(n3783) );
  XNOR2_X1 U4616 ( .A(IR_REG_18__SCAN_IN), .B(keyinput124), .ZN(n3782) );
  XNOR2_X1 U4617 ( .A(IR_REG_30__SCAN_IN), .B(keyinput118), .ZN(n3781) );
  NAND4_X1 U4618 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3785)
         );
  NOR3_X1 U4619 ( .A1(n3787), .A2(n3786), .A3(n3785), .ZN(n3826) );
  INV_X1 U4620 ( .A(DATAI_14_), .ZN(n4979) );
  AOI22_X1 U4621 ( .A1(n2226), .A2(keyinput113), .B1(keyinput108), .B2(n4979), 
        .ZN(n3788) );
  OAI221_X1 U4622 ( .B1(n2226), .B2(keyinput113), .C1(n4979), .C2(keyinput108), 
        .A(n3788), .ZN(n3798) );
  AOI22_X1 U4623 ( .A1(n3791), .A2(keyinput110), .B1(keyinput105), .B2(n3790), 
        .ZN(n3789) );
  OAI221_X1 U4624 ( .B1(n3791), .B2(keyinput110), .C1(n3790), .C2(keyinput105), 
        .A(n3789), .ZN(n3797) );
  AOI22_X1 U4625 ( .A1(n3201), .A2(keyinput98), .B1(n4917), .B2(keyinput101), 
        .ZN(n3792) );
  OAI221_X1 U4626 ( .B1(n3201), .B2(keyinput98), .C1(n4917), .C2(keyinput101), 
        .A(n3792), .ZN(n3796) );
  AOI22_X1 U4627 ( .A1(n2662), .A2(keyinput96), .B1(keyinput84), .B2(n3794), 
        .ZN(n3793) );
  OAI221_X1 U4628 ( .B1(n2662), .B2(keyinput96), .C1(n3794), .C2(keyinput84), 
        .A(n3793), .ZN(n3795) );
  NOR4_X1 U4629 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3825)
         );
  INV_X1 U4630 ( .A(DATAI_31_), .ZN(n3960) );
  INV_X1 U4631 ( .A(D_REG_16__SCAN_IN), .ZN(n4966) );
  AOI22_X1 U4632 ( .A1(n3960), .A2(keyinput66), .B1(n4966), .B2(keyinput64), 
        .ZN(n3799) );
  OAI221_X1 U4633 ( .B1(n3960), .B2(keyinput66), .C1(n4966), .C2(keyinput64), 
        .A(n3799), .ZN(n3811) );
  AOI22_X1 U4634 ( .A1(n3802), .A2(keyinput72), .B1(keyinput68), .B2(n3801), 
        .ZN(n3800) );
  OAI221_X1 U4635 ( .B1(n3802), .B2(keyinput72), .C1(n3801), .C2(keyinput68), 
        .A(n3800), .ZN(n3810) );
  AOI22_X1 U4636 ( .A1(n3804), .A2(keyinput86), .B1(n4088), .B2(keyinput81), 
        .ZN(n3803) );
  OAI221_X1 U4637 ( .B1(n3804), .B2(keyinput86), .C1(n4088), .C2(keyinput81), 
        .A(n3803), .ZN(n3809) );
  XOR2_X1 U4638 ( .A(n3805), .B(keyinput74), .Z(n3807) );
  XNOR2_X1 U4639 ( .A(IR_REG_12__SCAN_IN), .B(keyinput76), .ZN(n3806) );
  NAND2_X1 U4640 ( .A1(n3807), .A2(n3806), .ZN(n3808) );
  NOR4_X1 U4641 ( .A1(n3811), .A2(n3810), .A3(n3809), .A4(n3808), .ZN(n3824)
         );
  INV_X1 U4642 ( .A(D_REG_26__SCAN_IN), .ZN(n4960) );
  AOI22_X1 U4643 ( .A1(n4960), .A2(keyinput60), .B1(keyinput58), .B2(n3813), 
        .ZN(n3812) );
  OAI221_X1 U4644 ( .B1(n4960), .B2(keyinput60), .C1(n3813), .C2(keyinput58), 
        .A(n3812), .ZN(n3822) );
  AOI22_X1 U4645 ( .A1(n3815), .A2(keyinput52), .B1(n3693), .B2(keyinput50), 
        .ZN(n3814) );
  OAI221_X1 U4646 ( .B1(n3815), .B2(keyinput52), .C1(n3693), .C2(keyinput50), 
        .A(n3814), .ZN(n3821) );
  XNOR2_X1 U4647 ( .A(IR_REG_15__SCAN_IN), .B(keyinput56), .ZN(n3819) );
  XNOR2_X1 U4648 ( .A(IR_REG_2__SCAN_IN), .B(keyinput44), .ZN(n3818) );
  XNOR2_X1 U4649 ( .A(keyinput57), .B(DATAI_12_), .ZN(n3817) );
  XNOR2_X1 U4650 ( .A(keyinput49), .B(DATAI_3_), .ZN(n3816) );
  NAND4_X1 U4651 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  NOR3_X1 U4652 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3823) );
  NAND4_X1 U4653 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3827)
         );
  AOI211_X1 U4654 ( .C1(keyinput102), .C2(n3829), .A(n3828), .B(n3827), .ZN(
        n3930) );
  AOI22_X1 U4655 ( .A1(n4113), .A2(keyinput61), .B1(keyinput53), .B2(n4133), 
        .ZN(n3830) );
  OAI221_X1 U4656 ( .B1(n4113), .B2(keyinput61), .C1(n4133), .C2(keyinput53), 
        .A(n3830), .ZN(n3840) );
  AOI22_X1 U4657 ( .A1(n3149), .A2(keyinput115), .B1(keyinput97), .B2(n3832), 
        .ZN(n3831) );
  OAI221_X1 U4658 ( .B1(n3149), .B2(keyinput115), .C1(n3832), .C2(keyinput97), 
        .A(n3831), .ZN(n3839) );
  INV_X1 U4659 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4660 ( .A1(n3835), .A2(keyinput46), .B1(keyinput40), .B2(n3834), 
        .ZN(n3833) );
  OAI221_X1 U4661 ( .B1(n3835), .B2(keyinput46), .C1(n3834), .C2(keyinput40), 
        .A(n3833), .ZN(n3838) );
  INV_X1 U4662 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U4663 ( .A1(n4156), .A2(keyinput70), .B1(keyinput12), .B2(n4391), 
        .ZN(n3836) );
  OAI221_X1 U4664 ( .B1(n4156), .B2(keyinput70), .C1(n4391), .C2(keyinput12), 
        .A(n3836), .ZN(n3837) );
  NOR4_X1 U4665 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3929)
         );
  AOI22_X1 U4666 ( .A1(n3842), .A2(keyinput111), .B1(n4920), .B2(keyinput89), 
        .ZN(n3841) );
  OAI221_X1 U4667 ( .B1(n3842), .B2(keyinput111), .C1(n4920), .C2(keyinput89), 
        .A(n3841), .ZN(n3851) );
  INV_X1 U4668 ( .A(D_REG_28__SCAN_IN), .ZN(n4958) );
  INV_X1 U4669 ( .A(D_REG_13__SCAN_IN), .ZN(n4967) );
  AOI22_X1 U4670 ( .A1(n4958), .A2(keyinput75), .B1(keyinput54), .B2(n4967), 
        .ZN(n3843) );
  OAI221_X1 U4671 ( .B1(n4958), .B2(keyinput75), .C1(n4967), .C2(keyinput54), 
        .A(n3843), .ZN(n3850) );
  AOI22_X1 U4672 ( .A1(n4826), .A2(keyinput6), .B1(keyinput121), .B2(n4752), 
        .ZN(n3844) );
  OAI221_X1 U4673 ( .B1(n4826), .B2(keyinput6), .C1(n4752), .C2(keyinput121), 
        .A(n3844), .ZN(n3849) );
  INV_X1 U4674 ( .A(REG0_REG_18__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4675 ( .A1(n3847), .A2(keyinput10), .B1(keyinput2), .B2(n3846), 
        .ZN(n3845) );
  OAI221_X1 U4676 ( .B1(n3847), .B2(keyinput10), .C1(n3846), .C2(keyinput2), 
        .A(n3845), .ZN(n3848) );
  NOR4_X1 U4677 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3928)
         );
  AOI22_X1 U4678 ( .A1(n4846), .A2(keyinput94), .B1(keyinput45), .B2(n2792), 
        .ZN(n3852) );
  OAI221_X1 U4679 ( .B1(n4846), .B2(keyinput94), .C1(n2792), .C2(keyinput45), 
        .A(n3852), .ZN(n3860) );
  INV_X1 U4680 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4854) );
  AOI22_X1 U4681 ( .A1(n4854), .A2(keyinput65), .B1(n3854), .B2(keyinput32), 
        .ZN(n3853) );
  OAI221_X1 U4682 ( .B1(n4854), .B2(keyinput65), .C1(n3854), .C2(keyinput32), 
        .A(n3853), .ZN(n3859) );
  AOI22_X1 U4683 ( .A1(n4959), .A2(keyinput41), .B1(keyinput59), .B2(n4965), 
        .ZN(n3855) );
  OAI221_X1 U4684 ( .B1(n4959), .B2(keyinput41), .C1(n4965), .C2(keyinput59), 
        .A(n3855), .ZN(n3858) );
  AOI22_X1 U4685 ( .A1(n4964), .A2(keyinput80), .B1(keyinput48), .B2(n4962), 
        .ZN(n3856) );
  OAI221_X1 U4686 ( .B1(n4964), .B2(keyinput80), .C1(n4962), .C2(keyinput48), 
        .A(n3856), .ZN(n3857) );
  NOR4_X1 U4687 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3926)
         );
  AOI22_X1 U4688 ( .A1(n3862), .A2(keyinput88), .B1(keyinput85), .B2(n4736), 
        .ZN(n3861) );
  OAI221_X1 U4689 ( .B1(n3862), .B2(keyinput88), .C1(n4736), .C2(keyinput85), 
        .A(n3861), .ZN(n3871) );
  AOI22_X1 U4690 ( .A1(n4822), .A2(keyinput91), .B1(n3864), .B2(keyinput82), 
        .ZN(n3863) );
  OAI221_X1 U4691 ( .B1(n4822), .B2(keyinput91), .C1(n3864), .C2(keyinput82), 
        .A(n3863), .ZN(n3870) );
  AOI22_X1 U4692 ( .A1(n4805), .A2(keyinput126), .B1(n3866), .B2(keyinput27), 
        .ZN(n3865) );
  OAI221_X1 U4693 ( .B1(n4805), .B2(keyinput126), .C1(n3866), .C2(keyinput27), 
        .A(n3865), .ZN(n3869) );
  INV_X1 U4694 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4813) );
  AOI22_X1 U4695 ( .A1(n4813), .A2(keyinput22), .B1(n4728), .B2(keyinput99), 
        .ZN(n3867) );
  OAI221_X1 U4696 ( .B1(n4813), .B2(keyinput22), .C1(n4728), .C2(keyinput99), 
        .A(n3867), .ZN(n3868) );
  NOR4_X1 U4697 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3925)
         );
  INV_X1 U4698 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4699 ( .A1(n5004), .A2(keyinput127), .B1(n3873), .B2(keyinput106), 
        .ZN(n3872) );
  OAI221_X1 U4700 ( .B1(n5004), .B2(keyinput127), .C1(n3873), .C2(keyinput106), 
        .A(n3872), .ZN(n3888) );
  AOI22_X1 U4701 ( .A1(n3875), .A2(keyinput104), .B1(n2860), .B2(keyinput95), 
        .ZN(n3874) );
  OAI221_X1 U4702 ( .B1(n3875), .B2(keyinput104), .C1(n2860), .C2(keyinput95), 
        .A(n3874), .ZN(n3887) );
  XNOR2_X1 U4703 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput83), .ZN(n3879) );
  XNOR2_X1 U4704 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput62), .ZN(n3878) );
  XNOR2_X1 U4705 ( .A(REG1_REG_0__SCAN_IN), .B(keyinput43), .ZN(n3877) );
  XNOR2_X1 U4706 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput14), .ZN(n3876) );
  AND4_X1 U4707 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  XNOR2_X1 U4708 ( .A(keyinput26), .B(REG0_REG_4__SCAN_IN), .ZN(n3884) );
  XNOR2_X1 U4709 ( .A(keyinput87), .B(n3689), .ZN(n3881) );
  XNOR2_X1 U4710 ( .A(keyinput1), .B(n2544), .ZN(n3880) );
  NOR2_X1 U4711 ( .A1(n3881), .A2(n3880), .ZN(n3883) );
  XNOR2_X1 U4712 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput8), .ZN(n3882) );
  NAND4_X1 U4713 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  NOR3_X1 U4714 ( .A1(n3888), .A2(n3887), .A3(n3886), .ZN(n3920) );
  INV_X1 U4715 ( .A(REG2_REG_22__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4716 ( .A1(n4505), .A2(keyinput7), .B1(keyinput92), .B2(n3890), 
        .ZN(n3889) );
  OAI221_X1 U4717 ( .B1(n4505), .B2(keyinput7), .C1(n3890), .C2(keyinput92), 
        .A(n3889), .ZN(n3894) );
  INV_X1 U4718 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4719 ( .A1(n3892), .A2(keyinput4), .B1(keyinput78), .B2(n4464), 
        .ZN(n3891) );
  OAI221_X1 U4720 ( .B1(n3892), .B2(keyinput4), .C1(n4464), .C2(keyinput78), 
        .A(n3891), .ZN(n3893) );
  NOR2_X1 U4721 ( .A1(n3894), .A2(n3893), .ZN(n3919) );
  AOI22_X1 U4722 ( .A1(n3896), .A2(keyinput79), .B1(keyinput93), .B2(n4898), 
        .ZN(n3895) );
  OAI221_X1 U4723 ( .B1(n3896), .B2(keyinput79), .C1(n4898), .C2(keyinput93), 
        .A(n3895), .ZN(n3903) );
  INV_X1 U4724 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4725 ( .A1(n3898), .A2(keyinput112), .B1(n4756), .B2(keyinput35), 
        .ZN(n3897) );
  OAI221_X1 U4726 ( .B1(n3898), .B2(keyinput112), .C1(n4756), .C2(keyinput35), 
        .A(n3897), .ZN(n3902) );
  INV_X1 U4727 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4584) );
  AOI22_X1 U4728 ( .A1(n3900), .A2(keyinput90), .B1(n4584), .B2(keyinput73), 
        .ZN(n3899) );
  OAI221_X1 U4729 ( .B1(n3900), .B2(keyinput90), .C1(n4584), .C2(keyinput73), 
        .A(n3899), .ZN(n3901) );
  NOR3_X1 U4730 ( .A1(n3903), .A2(n3902), .A3(n3901), .ZN(n3918) );
  INV_X1 U4731 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4850) );
  AOI22_X1 U4732 ( .A1(n4850), .A2(keyinput100), .B1(keyinput67), .B2(n4954), 
        .ZN(n3904) );
  OAI221_X1 U4733 ( .B1(n4850), .B2(keyinput100), .C1(n4954), .C2(keyinput67), 
        .A(n3904), .ZN(n3916) );
  AOI22_X1 U4734 ( .A1(n3493), .A2(keyinput25), .B1(n3906), .B2(keyinput36), 
        .ZN(n3905) );
  OAI221_X1 U4735 ( .B1(n3493), .B2(keyinput25), .C1(n3906), .C2(keyinput36), 
        .A(n3905), .ZN(n3915) );
  INV_X1 U4736 ( .A(keyinput102), .ZN(n3908) );
  AND2_X1 U4737 ( .A1(n4071), .A2(keyinput77), .ZN(n3907) );
  AOI21_X1 U4738 ( .B1(n3908), .B2(IR_REG_26__SCAN_IN), .A(n3907), .ZN(n3913)
         );
  XNOR2_X1 U4739 ( .A(keyinput5), .B(REG1_REG_7__SCAN_IN), .ZN(n3912) );
  XNOR2_X1 U4740 ( .A(DATAI_17_), .B(keyinput30), .ZN(n3911) );
  INV_X1 U4741 ( .A(keyinput77), .ZN(n3909) );
  NAND2_X1 U4742 ( .A1(n3909), .A2(REG3_REG_25__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4743 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  NOR3_X1 U4744 ( .A1(n3916), .A2(n3915), .A3(n3914), .ZN(n3917) );
  AND4_X1 U4745 ( .A1(n3920), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3924)
         );
  OAI22_X1 U4746 ( .A1(n2331), .A2(keyinput120), .B1(n3922), .B2(keyinput16), 
        .ZN(n3921) );
  AOI221_X1 U4747 ( .B1(n2331), .B2(keyinput120), .C1(keyinput16), .C2(n3922), 
        .A(n3921), .ZN(n3923) );
  AND4_X1 U4748 ( .A1(n3926), .A2(n3925), .A3(n3924), .A4(n3923), .ZN(n3927)
         );
  NAND4_X1 U4749 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  XNOR2_X1 U4750 ( .A(n3932), .B(n3931), .ZN(U3252) );
  XNOR2_X1 U4751 ( .A(n3945), .B(REG2_REG_13__SCAN_IN), .ZN(n3935) );
  AOI21_X1 U4752 ( .B1(n3935), .B2(n3933), .A(n4905), .ZN(n3934) );
  OAI21_X1 U4753 ( .B1(n3933), .B2(n3935), .A(n3934), .ZN(n3944) );
  NAND2_X1 U4754 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4144) );
  INV_X1 U4755 ( .A(n4144), .ZN(n3942) );
  AND2_X1 U4756 ( .A1(n3937), .A2(n3936), .ZN(n3940) );
  AOI211_X1 U4757 ( .C1(n3940), .C2(n3939), .A(n3938), .B(n4908), .ZN(n3941)
         );
  AOI211_X1 U4758 ( .C1(n4930), .C2(ADDR_REG_13__SCAN_IN), .A(n3942), .B(n3941), .ZN(n3943) );
  OAI211_X1 U4759 ( .C1(n4945), .C2(n3945), .A(n3944), .B(n3943), .ZN(U3253)
         );
  INV_X1 U4760 ( .A(n4865), .ZN(n3958) );
  AOI21_X1 U4761 ( .B1(n3947), .B2(n3946), .A(n2167), .ZN(n3948) );
  NAND2_X1 U4762 ( .A1(n4940), .A2(n3948), .ZN(n3957) );
  NAND2_X1 U4763 ( .A1(n4930), .A2(ADDR_REG_18__SCAN_IN), .ZN(n3953) );
  NOR2_X1 U4764 ( .A1(n3951), .A2(STATE_REG_SCAN_IN), .ZN(n4182) );
  INV_X1 U4765 ( .A(n4182), .ZN(n3952) );
  NAND2_X1 U4766 ( .A1(n3953), .A2(n3952), .ZN(n3954) );
  OAI211_X1 U4767 ( .C1(n3958), .C2(n4945), .A(n3957), .B(n3956), .ZN(U3258)
         );
  NAND3_X1 U4768 ( .A1(n3959), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3961) );
  OAI22_X1 U4769 ( .A1(n3962), .A2(n3961), .B1(STATE_REG_SCAN_IN), .B2(n3960), 
        .ZN(U3321) );
  NAND2_X1 U4770 ( .A1(n3963), .A2(REG3_REG_0__SCAN_IN), .ZN(n3967) );
  XOR2_X1 U4771 ( .A(n3965), .B(n3964), .Z(n4365) );
  AOI22_X1 U4772 ( .A1(n4365), .A2(n4102), .B1(n4165), .B2(n2251), .ZN(n3966)
         );
  OAI211_X1 U4773 ( .C1(n4180), .C2(n3968), .A(n3967), .B(n3966), .ZN(U3229)
         );
  OR2_X2 U4774 ( .A1(n3970), .A2(n3969), .ZN(n3972) );
  NAND2_X1 U4775 ( .A1(n4268), .A2(n2140), .ZN(n3975) );
  OR2_X1 U4776 ( .A1(n3989), .A2(n4269), .ZN(n3974) );
  NAND2_X1 U4777 ( .A1(n3975), .A2(n3974), .ZN(n3977) );
  XNOR2_X1 U4778 ( .A(n3977), .B(n3976), .ZN(n3993) );
  NOR2_X1 U4779 ( .A1(n2134), .A2(n4269), .ZN(n3978) );
  AOI21_X1 U4780 ( .B1(n4268), .B2(n2823), .A(n3978), .ZN(n3994) );
  XNOR2_X1 U4781 ( .A(n3993), .B(n3994), .ZN(n3984) );
  XNOR2_X1 U4782 ( .A(n3985), .B(n3984), .ZN(n3983) );
  NOR2_X1 U4783 ( .A1(n4461), .A2(n4169), .ZN(n3981) );
  AOI22_X1 U4784 ( .A1(n4191), .A2(n4423), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3979) );
  OAI21_X1 U4785 ( .B1(n4426), .B2(n4194), .A(n3979), .ZN(n3980) );
  AOI211_X1 U4786 ( .C1(n4418), .C2(n4196), .A(n3981), .B(n3980), .ZN(n3982)
         );
  OAI21_X1 U4787 ( .B1(n3983), .B2(n4199), .A(n3982), .ZN(U3211) );
  OAI22_X1 U4788 ( .A1(n4426), .A2(n2730), .B1(n2134), .B2(n3988), .ZN(n3987)
         );
  XNOR2_X1 U4789 ( .A(n3987), .B(n3986), .ZN(n3992) );
  OAI22_X1 U4790 ( .A1(n4426), .A2(n2133), .B1(n3989), .B2(n3988), .ZN(n3991)
         );
  XNOR2_X1 U4791 ( .A(n3992), .B(n3991), .ZN(n3997) );
  INV_X1 U4792 ( .A(n3997), .ZN(n4002) );
  INV_X1 U4793 ( .A(n3993), .ZN(n3996) );
  INV_X1 U4794 ( .A(n3994), .ZN(n3995) );
  NAND2_X1 U4795 ( .A1(n3996), .A2(n3995), .ZN(n4001) );
  NAND3_X1 U4796 ( .A1(n4002), .A2(n4102), .A3(n4001), .ZN(n4008) );
  NAND2_X1 U4797 ( .A1(n4009), .A2(n3998), .ZN(n4007) );
  INV_X1 U4798 ( .A(n4011), .ZN(n4005) );
  NAND2_X1 U4799 ( .A1(n4349), .A2(n4165), .ZN(n4000) );
  AOI22_X1 U4800 ( .A1(n4191), .A2(n4405), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3999) );
  OAI211_X1 U4801 ( .C1(n4442), .C2(n4169), .A(n4000), .B(n3999), .ZN(n4004)
         );
  NOR3_X1 U4802 ( .A1(n4002), .A2(n4199), .A3(n4001), .ZN(n4003) );
  AOI211_X1 U4803 ( .C1(n4005), .C2(n4196), .A(n4004), .B(n4003), .ZN(n4006)
         );
  OAI211_X1 U4804 ( .C1(n4009), .C2(n4008), .A(n4007), .B(n4006), .ZN(U3217)
         );
  INV_X1 U4805 ( .A(n4010), .ZN(n4015) );
  OAI22_X1 U4806 ( .A1(n4011), .A2(n4649), .B1(n3892), .B2(n4955), .ZN(n4014)
         );
  NOR2_X1 U4807 ( .A1(n4012), .A2(n2132), .ZN(n4013) );
  AOI211_X1 U4808 ( .C1(n4668), .C2(n4015), .A(n4014), .B(n4013), .ZN(n4016)
         );
  OAI21_X1 U4809 ( .B1(n4017), .B2(n4670), .A(n4016), .ZN(U3262) );
  XNOR2_X1 U4810 ( .A(n4080), .B(n4079), .ZN(n4019) );
  XNOR2_X1 U4811 ( .A(n4018), .B(n4019), .ZN(n4023) );
  AOI22_X1 U4812 ( .A1(n4191), .A2(n4673), .B1(n4165), .B2(n4674), .ZN(n4020)
         );
  NAND2_X1 U4813 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4902) );
  OAI211_X1 U4814 ( .C1(n4677), .C2(n4169), .A(n4020), .B(n4902), .ZN(n4021)
         );
  AOI21_X1 U4815 ( .B1(n4685), .B2(n4196), .A(n4021), .ZN(n4022) );
  OAI21_X1 U4816 ( .B1(n4023), .B2(n4199), .A(n4022), .ZN(U3212) );
  AND2_X1 U4817 ( .A1(n4024), .A2(n4025), .ZN(n4028) );
  OAI211_X1 U4818 ( .C1(n4028), .C2(n4027), .A(n4102), .B(n4026), .ZN(n4032)
         );
  OAI22_X1 U4819 ( .A1(n4536), .A2(n4169), .B1(n4180), .B2(n3092), .ZN(n4030)
         );
  NOR2_X1 U4820 ( .A1(n4072), .A2(n4194), .ZN(n4029) );
  AOI211_X1 U4821 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n4030), .B(n4029), .ZN(n4031) );
  OAI211_X1 U4822 ( .C1(n4108), .C2(n4506), .A(n4032), .B(n4031), .ZN(U3213)
         );
  OR2_X1 U4823 ( .A1(n4033), .A2(n4176), .ZN(n4034) );
  NAND2_X1 U4824 ( .A1(n4034), .A2(n4175), .ZN(n4124) );
  XOR2_X1 U4825 ( .A(n4123), .B(n4124), .Z(n4041) );
  INV_X1 U4826 ( .A(n4583), .ZN(n4039) );
  AOI22_X1 U4827 ( .A1(n4192), .A2(n4035), .B1(n4191), .B2(n4579), .ZN(n4037)
         );
  OAI211_X1 U4828 ( .C1(n4048), .C2(n4194), .A(n4037), .B(n4036), .ZN(n4038)
         );
  AOI21_X1 U4829 ( .B1(n4039), .B2(n4196), .A(n4038), .ZN(n4040) );
  OAI21_X1 U4830 ( .B1(n4041), .B2(n4199), .A(n4040), .ZN(U3216) );
  NAND2_X1 U4831 ( .A1(n4124), .A2(n4042), .ZN(n4122) );
  NAND2_X1 U4832 ( .A1(n4122), .A2(n4043), .ZN(n4047) );
  XNOR2_X1 U4833 ( .A(n4045), .B(n4044), .ZN(n4046) );
  XNOR2_X1 U4834 ( .A(n4047), .B(n4046), .ZN(n4053) );
  OAI22_X1 U4835 ( .A1(n4180), .A2(n4537), .B1(n4048), .B2(n4169), .ZN(n4051)
         );
  OAI22_X1 U4836 ( .A1(n4536), .A2(n4194), .B1(STATE_REG_SCAN_IN), .B2(n4049), 
        .ZN(n4050) );
  AOI211_X1 U4837 ( .C1(n4539), .C2(n4196), .A(n4051), .B(n4050), .ZN(n4052)
         );
  OAI21_X1 U4838 ( .B1(n4053), .B2(n4199), .A(n4052), .ZN(U3220) );
  XOR2_X1 U4839 ( .A(n4056), .B(n4055), .Z(n4057) );
  XNOR2_X1 U4840 ( .A(n4054), .B(n4057), .ZN(n4066) );
  AOI22_X1 U4841 ( .A1(n4191), .A2(n4059), .B1(n4165), .B2(n4058), .ZN(n4061)
         );
  OAI211_X1 U4842 ( .C1(n4062), .C2(n4169), .A(n4061), .B(n4060), .ZN(n4063)
         );
  AOI21_X1 U4843 ( .B1(n4064), .B2(n4196), .A(n4063), .ZN(n4065) );
  OAI21_X1 U4844 ( .B1(n4066), .B2(n4199), .A(n4065), .ZN(U3221) );
  NAND2_X1 U4845 ( .A1(n4068), .A2(n4067), .ZN(n4070) );
  XOR2_X1 U4846 ( .A(n4070), .B(n4069), .Z(n4077) );
  OAI22_X1 U4847 ( .A1(n4072), .A2(n4169), .B1(STATE_REG_SCAN_IN), .B2(n4071), 
        .ZN(n4073) );
  AOI21_X1 U4848 ( .B1(n4458), .B2(n4191), .A(n4073), .ZN(n4074) );
  OAI21_X1 U4849 ( .B1(n4108), .B2(n4465), .A(n4074), .ZN(n4075) );
  AOI21_X1 U4850 ( .B1(n4165), .B2(n4350), .A(n4075), .ZN(n4076) );
  OAI21_X1 U4851 ( .B1(n4077), .B2(n4199), .A(n4076), .ZN(U3222) );
  XNOR2_X1 U4852 ( .A(n4097), .B(n4078), .ZN(n4093) );
  INV_X1 U4853 ( .A(n4080), .ZN(n4083) );
  INV_X1 U4854 ( .A(n4018), .ZN(n4081) );
  OAI21_X1 U4855 ( .B1(n4081), .B2(n4080), .A(n4079), .ZN(n4082) );
  OAI21_X1 U4856 ( .B1(n4083), .B2(n4018), .A(n4082), .ZN(n4085) );
  NAND2_X1 U4857 ( .A1(n4085), .A2(n4084), .ZN(n4186) );
  NOR2_X1 U4858 ( .A1(n4085), .A2(n4084), .ZN(n4188) );
  AOI21_X1 U4859 ( .B1(n4094), .B2(n4186), .A(n4188), .ZN(n4086) );
  XOR2_X1 U4860 ( .A(n4093), .B(n4086), .Z(n4087) );
  NAND2_X1 U4861 ( .A1(n4087), .A2(n4102), .ZN(n4092) );
  NOR2_X1 U4862 ( .A1(n4088), .A2(STATE_REG_SCAN_IN), .ZN(n4919) );
  OAI22_X1 U4863 ( .A1(n4180), .A2(n4089), .B1(n4621), .B2(n4169), .ZN(n4090)
         );
  AOI211_X1 U4864 ( .C1(n4165), .C2(n4590), .A(n4919), .B(n4090), .ZN(n4091)
         );
  OAI211_X1 U4865 ( .C1(n4108), .C2(n4632), .A(n4092), .B(n4091), .ZN(U3223)
         );
  OAI211_X1 U4866 ( .C1(n4188), .C2(n4094), .A(n4093), .B(n4186), .ZN(n4095)
         );
  OAI21_X1 U4867 ( .B1(n4097), .B2(n4096), .A(n4095), .ZN(n4101) );
  XOR2_X1 U4868 ( .A(n4099), .B(n4098), .Z(n4100) );
  XNOR2_X1 U4869 ( .A(n4101), .B(n4100), .ZN(n4103) );
  NAND2_X1 U4870 ( .A1(n4103), .A2(n4102), .ZN(n4107) );
  AND2_X1 U4871 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4929) );
  OAI22_X1 U4872 ( .A1(n4180), .A2(n4104), .B1(n4194), .B2(n4610), .ZN(n4105)
         );
  AOI211_X1 U4873 ( .C1(n4192), .C2(n4608), .A(n4929), .B(n4105), .ZN(n4106)
         );
  OAI211_X1 U4874 ( .C1(n4108), .C2(n4616), .A(n4107), .B(n4106), .ZN(U3225)
         );
  NAND2_X1 U4875 ( .A1(n4109), .A2(n4110), .ZN(n4111) );
  XOR2_X1 U4876 ( .A(n4112), .B(n4111), .Z(n4120) );
  OAI22_X1 U4877 ( .A1(n3093), .A2(n4169), .B1(STATE_REG_SCAN_IN), .B2(n4113), 
        .ZN(n4114) );
  AOI21_X1 U4878 ( .B1(n4115), .B2(n4191), .A(n4114), .ZN(n4116) );
  OAI21_X1 U4879 ( .B1(n4117), .B2(n4194), .A(n4116), .ZN(n4118) );
  AOI21_X1 U4880 ( .B1(n4486), .B2(n4196), .A(n4118), .ZN(n4119) );
  OAI21_X1 U4881 ( .B1(n4120), .B2(n4199), .A(n4119), .ZN(U3226) );
  NAND2_X1 U4882 ( .A1(n4122), .A2(n4121), .ZN(n4131) );
  NAND2_X1 U4883 ( .A1(n4124), .A2(n4123), .ZN(n4126) );
  NAND2_X1 U4884 ( .A1(n4126), .A2(n4125), .ZN(n4127) );
  AOI21_X1 U4885 ( .B1(n4130), .B2(n4128), .A(n4127), .ZN(n4129) );
  AOI21_X1 U4886 ( .B1(n4131), .B2(n4130), .A(n4129), .ZN(n4137) );
  INV_X1 U4887 ( .A(n4132), .ZN(n4562) );
  OAI22_X1 U4888 ( .A1(n4194), .A2(n4517), .B1(STATE_REG_SCAN_IN), .B2(n4133), 
        .ZN(n4135) );
  OAI22_X1 U4889 ( .A1(n4180), .A2(n4553), .B1(n4592), .B2(n4169), .ZN(n4134)
         );
  AOI211_X1 U4890 ( .C1(n4562), .C2(n4196), .A(n4135), .B(n4134), .ZN(n4136)
         );
  OAI21_X1 U4891 ( .B1(n4137), .B2(n4199), .A(n4136), .ZN(U3230) );
  INV_X1 U4892 ( .A(n4139), .ZN(n4141) );
  NOR2_X1 U4893 ( .A1(n4141), .A2(n4140), .ZN(n4142) );
  XNOR2_X1 U4894 ( .A(n4138), .B(n4142), .ZN(n4149) );
  AOI22_X1 U4895 ( .A1(n4191), .A2(n4143), .B1(n4165), .B2(n4698), .ZN(n4145)
         );
  OAI211_X1 U4896 ( .C1(n4146), .C2(n4169), .A(n4145), .B(n4144), .ZN(n4147)
         );
  AOI21_X1 U4897 ( .B1(n4709), .B2(n4196), .A(n4147), .ZN(n4148) );
  OAI21_X1 U4898 ( .B1(n4149), .B2(n4199), .A(n4148), .ZN(U3231) );
  NAND2_X1 U4899 ( .A1(n4151), .A2(n4150), .ZN(n4153) );
  INV_X1 U4900 ( .A(n4024), .ZN(n4152) );
  AOI21_X1 U4901 ( .B1(n4154), .B2(n4153), .A(n4152), .ZN(n4160) );
  OAI22_X1 U4902 ( .A1(n4180), .A2(n4524), .B1(n4517), .B2(n4169), .ZN(n4158)
         );
  NAND2_X1 U4903 ( .A1(n4519), .A2(n4165), .ZN(n4155) );
  OAI21_X1 U4904 ( .B1(STATE_REG_SCAN_IN), .B2(n4156), .A(n4155), .ZN(n4157)
         );
  AOI211_X1 U4905 ( .C1(n4522), .C2(n4196), .A(n4158), .B(n4157), .ZN(n4159)
         );
  OAI21_X1 U4906 ( .B1(n4160), .B2(n4199), .A(n4159), .ZN(U3232) );
  NAND2_X1 U4907 ( .A1(n4162), .A2(n4161), .ZN(n4164) );
  XOR2_X1 U4908 ( .A(n4164), .B(n4163), .Z(n4174) );
  AOI22_X1 U4909 ( .A1(n4191), .A2(n4166), .B1(n4165), .B2(n4695), .ZN(n4168)
         );
  OAI211_X1 U4910 ( .C1(n4170), .C2(n4169), .A(n4168), .B(n4167), .ZN(n4171)
         );
  AOI21_X1 U4911 ( .B1(n4172), .B2(n4196), .A(n4171), .ZN(n4173) );
  OAI21_X1 U4912 ( .B1(n4174), .B2(n4199), .A(n4173), .ZN(U3233) );
  INV_X1 U4913 ( .A(n4175), .ZN(n4177) );
  NOR2_X1 U4914 ( .A1(n4177), .A2(n4176), .ZN(n4178) );
  XNOR2_X1 U4915 ( .A(n4033), .B(n4178), .ZN(n4185) );
  OAI22_X1 U4916 ( .A1(n4180), .A2(n4179), .B1(n4194), .B2(n4592), .ZN(n4181)
         );
  AOI211_X1 U4917 ( .C1(n4192), .C2(n4590), .A(n4182), .B(n4181), .ZN(n4184)
         );
  NAND2_X1 U4918 ( .A1(n4196), .A2(n4601), .ZN(n4183) );
  OAI211_X1 U4919 ( .C1(n4185), .C2(n4199), .A(n4184), .B(n4183), .ZN(U3235)
         );
  INV_X1 U4920 ( .A(n4186), .ZN(n4187) );
  NOR2_X1 U4921 ( .A1(n4188), .A2(n4187), .ZN(n4190) );
  XNOR2_X1 U4922 ( .A(n4190), .B(n4189), .ZN(n4200) );
  INV_X1 U4923 ( .A(n4650), .ZN(n4197) );
  INV_X1 U4924 ( .A(n4608), .ZN(n4655) );
  AOI22_X1 U4925 ( .A1(n4192), .A2(n4698), .B1(n4191), .B2(n4629), .ZN(n4193)
         );
  NAND2_X1 U4926 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4915) );
  OAI211_X1 U4927 ( .C1(n4655), .C2(n4194), .A(n4193), .B(n4915), .ZN(n4195)
         );
  AOI21_X1 U4928 ( .B1(n4197), .B2(n4196), .A(n4195), .ZN(n4198) );
  OAI21_X1 U4929 ( .B1(n4200), .B2(n4199), .A(n4198), .ZN(U3238) );
  INV_X1 U4930 ( .A(n4201), .ZN(n4318) );
  NAND2_X1 U4931 ( .A1(n2405), .A2(n4202), .ZN(n4320) );
  AOI211_X1 U4932 ( .C1(n4624), .C2(n4317), .A(n4318), .B(n4320), .ZN(n4204)
         );
  NAND3_X1 U4933 ( .A1(n4494), .A2(n4203), .A3(n4493), .ZN(n4321) );
  OAI21_X1 U4934 ( .B1(n4204), .B2(n4321), .A(n4324), .ZN(n4205) );
  AOI21_X1 U4935 ( .B1(n4205), .B2(n4325), .A(n4435), .ZN(n4212) );
  NAND2_X1 U4936 ( .A1(n4393), .A2(n4206), .ZN(n4215) );
  AND2_X1 U4937 ( .A1(n2138), .A2(DATAI_29_), .ZN(n4412) );
  NAND2_X1 U4938 ( .A1(n4207), .A2(n4412), .ZN(n4264) );
  INV_X1 U4939 ( .A(n4399), .ZN(n4208) );
  NAND2_X1 U4940 ( .A1(n2138), .A2(DATAI_30_), .ZN(n4383) );
  INV_X1 U4941 ( .A(n4383), .ZN(n4386) );
  NAND2_X1 U4942 ( .A1(n4208), .A2(n4386), .ZN(n4210) );
  NAND2_X1 U4943 ( .A1(n4209), .A2(DATAI_31_), .ZN(n4377) );
  NAND2_X1 U4944 ( .A1(n4376), .A2(n4377), .ZN(n4333) );
  AND2_X1 U4945 ( .A1(n4210), .A2(n4333), .ZN(n4235) );
  NAND2_X1 U4946 ( .A1(n4264), .A2(n4235), .ZN(n4216) );
  NOR4_X1 U4947 ( .A1(n4212), .A2(n4211), .A3(n4215), .A4(n4216), .ZN(n4221)
         );
  INV_X1 U4948 ( .A(n4412), .ZN(n4213) );
  NAND2_X1 U4949 ( .A1(n4349), .A2(n4213), .ZN(n4263) );
  NAND2_X1 U4950 ( .A1(n4395), .A2(n4263), .ZN(n4267) );
  NOR2_X1 U4951 ( .A1(n4267), .A2(n4214), .ZN(n4219) );
  INV_X1 U4952 ( .A(n4215), .ZN(n4218) );
  INV_X1 U4953 ( .A(n4216), .ZN(n4217) );
  OAI21_X1 U4954 ( .B1(n4218), .B2(n4267), .A(n4217), .ZN(n4331) );
  AOI21_X1 U4955 ( .B1(n4422), .B2(n4219), .A(n4331), .ZN(n4220) );
  OAI22_X1 U4956 ( .A1(n4221), .A2(n4220), .B1(n4376), .B2(n4383), .ZN(n4340)
         );
  NAND2_X1 U4957 ( .A1(n4399), .A2(n4383), .ZN(n4230) );
  AOI21_X1 U4958 ( .B1(n4230), .B2(n4376), .A(n4377), .ZN(n4223) );
  NOR2_X1 U4959 ( .A1(n4223), .A2(n4222), .ZN(n4339) );
  XNOR2_X1 U4960 ( .A(n4461), .B(n4445), .ZN(n4436) );
  NAND2_X1 U4961 ( .A1(n4434), .A2(n4224), .ZN(n4455) );
  INV_X1 U4962 ( .A(n4455), .ZN(n4262) );
  NAND2_X1 U4963 ( .A1(n4225), .A2(n4453), .ZN(n4471) );
  INV_X1 U4964 ( .A(n4471), .ZN(n4474) );
  NAND2_X1 U4965 ( .A1(n4472), .A2(n4226), .ZN(n4495) );
  INV_X1 U4966 ( .A(n4495), .ZN(n4261) );
  INV_X1 U4967 ( .A(n4227), .ZN(n4228) );
  INV_X1 U4968 ( .A(n4568), .ZN(n4229) );
  AND2_X1 U4969 ( .A1(n4229), .A2(n4567), .ZN(n4613) );
  OAI21_X1 U4970 ( .B1(n4376), .B2(n4377), .A(n4230), .ZN(n4332) );
  NOR2_X1 U4971 ( .A1(n4332), .A2(n4277), .ZN(n4231) );
  AND4_X1 U4972 ( .A1(n4234), .A2(n4233), .A3(n4232), .A4(n4231), .ZN(n4243)
         );
  INV_X1 U4973 ( .A(n4235), .ZN(n4236) );
  NOR2_X1 U4974 ( .A1(n4237), .A2(n4236), .ZN(n4242) );
  INV_X1 U4975 ( .A(n4680), .ZN(n4671) );
  AND4_X1 U4976 ( .A1(n4671), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(n4241)
         );
  AND4_X1 U4977 ( .A1(n4613), .A2(n4243), .A3(n4242), .A4(n4241), .ZN(n4253)
         );
  NAND4_X1 U4978 ( .A1(n3112), .A2(n4246), .A3(n4245), .A4(n4244), .ZN(n4250)
         );
  NAND2_X1 U4979 ( .A1(n4248), .A2(n4247), .ZN(n4662) );
  NOR4_X1 U4980 ( .A1(n4597), .A2(n4250), .A3(n4249), .A4(n4662), .ZN(n4252)
         );
  NAND2_X1 U4981 ( .A1(n4636), .A2(n4251), .ZN(n4694) );
  NAND4_X1 U4982 ( .A1(n4531), .A2(n4253), .A3(n4252), .A4(n4694), .ZN(n4259)
         );
  NAND2_X1 U4983 ( .A1(n4255), .A2(n4254), .ZN(n4551) );
  INV_X1 U4984 ( .A(n4546), .ZN(n4256) );
  OR2_X1 U4985 ( .A1(n4256), .A2(n4545), .ZN(n4572) );
  NAND4_X1 U4986 ( .A1(n4551), .A2(n4645), .A3(n4257), .A4(n4572), .ZN(n4258)
         );
  NOR3_X1 U4987 ( .A1(n4259), .A2(n4512), .A3(n4258), .ZN(n4260) );
  NAND4_X1 U4988 ( .A1(n4262), .A2(n4474), .A3(n4261), .A4(n4260), .ZN(n4265)
         );
  NAND2_X1 U4989 ( .A1(n4264), .A2(n4263), .ZN(n4409) );
  NOR2_X1 U4990 ( .A1(n4265), .A2(n4409), .ZN(n4266) );
  AND4_X1 U4991 ( .A1(n2305), .A2(n4422), .A3(n4436), .A4(n4266), .ZN(n4337)
         );
  AOI21_X1 U4992 ( .B1(n4269), .B2(n4268), .A(n4267), .ZN(n4330) );
  INV_X1 U4993 ( .A(n4310), .ZN(n4273) );
  INV_X1 U4994 ( .A(n4270), .ZN(n4271) );
  OAI211_X1 U4995 ( .C1(n4274), .C2(n4273), .A(n4272), .B(n4271), .ZN(n4315)
         );
  OAI211_X1 U4996 ( .C1(n4278), .C2(n4277), .A(n4276), .B(n4275), .ZN(n4279)
         );
  NAND3_X1 U4997 ( .A1(n4279), .A2(n3115), .A3(n3113), .ZN(n4282) );
  NAND3_X1 U4998 ( .A1(n4282), .A2(n4281), .A3(n4280), .ZN(n4284) );
  NAND3_X1 U4999 ( .A1(n4284), .A2(n3116), .A3(n4283), .ZN(n4285) );
  NAND4_X1 U5000 ( .A1(n4285), .A2(n3117), .A3(n4301), .A4(n2173), .ZN(n4288)
         );
  NAND3_X1 U5001 ( .A1(n4288), .A2(n4287), .A3(n4286), .ZN(n4289) );
  NAND3_X1 U5002 ( .A1(n4289), .A2(n4299), .A3(n4298), .ZN(n4292) );
  NAND3_X1 U5003 ( .A1(n4292), .A2(n4291), .A3(n4290), .ZN(n4296) );
  INV_X1 U5004 ( .A(n4293), .ZN(n4295) );
  NAND3_X1 U5005 ( .A1(n4296), .A2(n4295), .A3(n4294), .ZN(n4313) );
  INV_X1 U5006 ( .A(n4297), .ZN(n4300) );
  NAND3_X1 U5007 ( .A1(n4300), .A2(n4299), .A3(n4298), .ZN(n4304) );
  INV_X1 U5008 ( .A(n4301), .ZN(n4302) );
  NOR3_X1 U5009 ( .A1(n4304), .A2(n4303), .A3(n4302), .ZN(n4307) );
  INV_X1 U5010 ( .A(n4305), .ZN(n4306) );
  OAI21_X1 U5011 ( .B1(n4307), .B2(n4306), .A(n4316), .ZN(n4312) );
  NAND3_X1 U5012 ( .A1(n4310), .A2(n4309), .A3(n4308), .ZN(n4311) );
  AOI21_X1 U5013 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(n4314) );
  AOI21_X1 U5014 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4319) );
  OAI21_X1 U5015 ( .B1(n4319), .B2(n4318), .A(n4317), .ZN(n4323) );
  INV_X1 U5016 ( .A(n4320), .ZN(n4322) );
  AOI21_X1 U5017 ( .B1(n4323), .B2(n4322), .A(n4321), .ZN(n4327) );
  INV_X1 U5018 ( .A(n4324), .ZN(n4326) );
  OAI211_X1 U5019 ( .C1(n4327), .C2(n4326), .A(n3143), .B(n4325), .ZN(n4328)
         );
  NAND3_X1 U5020 ( .A1(n4330), .A2(n4329), .A3(n4328), .ZN(n4335) );
  INV_X1 U5021 ( .A(n4331), .ZN(n4334) );
  AOI22_X1 U5022 ( .A1(n4335), .A2(n4334), .B1(n4333), .B2(n4332), .ZN(n4336)
         );
  MUX2_X1 U5023 ( .A(n4337), .B(n4336), .S(n2640), .Z(n4338) );
  AOI21_X1 U5024 ( .B1(n4340), .B2(n4339), .A(n4338), .ZN(n4342) );
  XNOR2_X1 U5025 ( .A(n4342), .B(n4341), .ZN(n4348) );
  NAND2_X1 U5026 ( .A1(n4343), .A2(n4360), .ZN(n4344) );
  OAI211_X1 U5027 ( .C1(n4345), .C2(n4347), .A(n4344), .B(B_REG_SCAN_IN), .ZN(
        n4346) );
  OAI21_X1 U5028 ( .B1(n4348), .B2(n4347), .A(n4346), .ZN(U3239) );
  MUX2_X1 U5029 ( .A(n4349), .B(DATAO_REG_29__SCAN_IN), .S(n4358), .Z(U3579)
         );
  MUX2_X1 U5030 ( .A(n4350), .B(DATAO_REG_26__SCAN_IN), .S(n4358), .Z(U3576)
         );
  MUX2_X1 U5031 ( .A(n4479), .B(DATAO_REG_25__SCAN_IN), .S(n4358), .Z(U3575)
         );
  MUX2_X1 U5032 ( .A(n4351), .B(DATAO_REG_22__SCAN_IN), .S(n4358), .Z(U3572)
         );
  MUX2_X1 U5033 ( .A(n4555), .B(DATAO_REG_21__SCAN_IN), .S(n4358), .Z(U3571)
         );
  MUX2_X1 U5034 ( .A(n4576), .B(DATAO_REG_20__SCAN_IN), .S(n4358), .Z(U3570)
         );
  MUX2_X1 U5035 ( .A(n4352), .B(DATAO_REG_19__SCAN_IN), .S(n4358), .Z(U3569)
         );
  MUX2_X1 U5036 ( .A(n4608), .B(DATAO_REG_16__SCAN_IN), .S(n4358), .Z(U3566)
         );
  MUX2_X1 U5037 ( .A(n4674), .B(DATAO_REG_15__SCAN_IN), .S(n4358), .Z(U3565)
         );
  MUX2_X1 U5038 ( .A(n4698), .B(DATAO_REG_14__SCAN_IN), .S(n4358), .Z(U3564)
         );
  MUX2_X1 U5039 ( .A(n4353), .B(DATAO_REG_11__SCAN_IN), .S(n4358), .Z(U3561)
         );
  MUX2_X1 U5040 ( .A(n4354), .B(DATAO_REG_10__SCAN_IN), .S(n4358), .Z(U3560)
         );
  MUX2_X1 U5041 ( .A(n4355), .B(DATAO_REG_9__SCAN_IN), .S(n4358), .Z(U3559) );
  MUX2_X1 U5042 ( .A(n4356), .B(DATAO_REG_6__SCAN_IN), .S(n4358), .Z(U3556) );
  MUX2_X1 U5043 ( .A(n4357), .B(DATAO_REG_5__SCAN_IN), .S(n4358), .Z(U3555) );
  MUX2_X1 U5044 ( .A(n3040), .B(DATAO_REG_4__SCAN_IN), .S(n4358), .Z(U3554) );
  MUX2_X1 U5045 ( .A(n2251), .B(DATAO_REG_1__SCAN_IN), .S(n4358), .Z(U3551) );
  MUX2_X1 U5046 ( .A(n2698), .B(DATAO_REG_0__SCAN_IN), .S(n4358), .Z(U3550) );
  NAND2_X1 U5047 ( .A1(n4859), .A2(n4359), .ZN(n4364) );
  NAND2_X1 U5048 ( .A1(n4360), .A2(REG2_REG_0__SCAN_IN), .ZN(n4361) );
  MUX2_X1 U5049 ( .A(n4362), .B(n4361), .S(IR_REG_0__SCAN_IN), .Z(n4363) );
  OAI211_X1 U5050 ( .C1(n4365), .C2(n4364), .A(U4043), .B(n4363), .ZN(n4891)
         );
  AOI22_X1 U5051 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4930), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4374) );
  XOR2_X1 U5052 ( .A(n4366), .B(n4367), .Z(n4368) );
  AOI22_X1 U5053 ( .A1(n2131), .A2(n4914), .B1(n4940), .B2(n4368), .ZN(n4373)
         );
  OAI211_X1 U5054 ( .C1(n4371), .C2(n4370), .A(n4942), .B(n4369), .ZN(n4372)
         );
  NAND4_X1 U5055 ( .A1(n4891), .A2(n4374), .A3(n4373), .A4(n4372), .ZN(U3242)
         );
  NAND2_X1 U5056 ( .A1(n4384), .A2(n4383), .ZN(n4382) );
  AND2_X1 U5057 ( .A1(n4860), .A2(B_REG_SCAN_IN), .ZN(n4375) );
  NOR2_X1 U5058 ( .A1(n4654), .A2(n4375), .ZN(n4400) );
  NAND2_X1 U5059 ( .A1(n4400), .A2(n4376), .ZN(n4388) );
  INV_X1 U5060 ( .A(n4377), .ZN(n4378) );
  NAND2_X1 U5061 ( .A1(n4672), .A2(n4378), .ZN(n4379) );
  NAND2_X1 U5062 ( .A1(n4388), .A2(n4379), .ZN(n4795) );
  NAND2_X1 U5063 ( .A1(n4652), .A2(n4795), .ZN(n4381) );
  NAND2_X1 U5064 ( .A1(n2132), .A2(REG2_REG_31__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U5065 ( .C1(n4798), .C2(n4711), .A(n4381), .B(n4380), .ZN(U3260)
         );
  OAI21_X1 U5066 ( .B1(n4384), .B2(n4383), .A(n4382), .ZN(n4802) );
  INV_X1 U5067 ( .A(n4802), .ZN(n4385) );
  NAND2_X1 U5068 ( .A1(n4385), .A2(n4668), .ZN(n4390) );
  NAND2_X1 U5069 ( .A1(n4672), .A2(n4386), .ZN(n4387) );
  NAND2_X1 U5070 ( .A1(n4388), .A2(n4387), .ZN(n4799) );
  NAND2_X1 U5071 ( .A1(n4652), .A2(n4799), .ZN(n4389) );
  OAI211_X1 U5072 ( .C1(n4652), .C2(n4391), .A(n4390), .B(n4389), .ZN(U3261)
         );
  INV_X1 U5073 ( .A(n4392), .ZN(n4404) );
  INV_X1 U5074 ( .A(n4393), .ZN(n4394) );
  NAND2_X1 U5075 ( .A1(n4406), .A2(n4696), .ZN(n4402) );
  AOI22_X1 U5076 ( .A1(n4400), .A2(n4399), .B1(n4412), .B2(n4672), .ZN(n4401)
         );
  AOI21_X1 U5077 ( .B1(n4404), .B2(n4950), .A(n4720), .ZN(n4415) );
  NAND2_X1 U5078 ( .A1(n4721), .A2(n4688), .ZN(n4414) );
  AOI21_X1 U5079 ( .B1(n4412), .B2(n4411), .A(n4384), .ZN(n4719) );
  AOI22_X1 U5080 ( .A1(n4719), .A2(n4668), .B1(REG2_REG_29__SCAN_IN), .B2(
        n2132), .ZN(n4413) );
  OAI211_X1 U5081 ( .C1(n2132), .C2(n4415), .A(n4414), .B(n4413), .ZN(U3354)
         );
  XNOR2_X1 U5082 ( .A(n4416), .B(n4422), .ZN(n4725) );
  AOI21_X1 U5083 ( .B1(n4423), .B2(n4444), .A(n4417), .ZN(n4722) );
  INV_X1 U5084 ( .A(n4418), .ZN(n4419) );
  OAI22_X1 U5085 ( .A1(n4419), .A2(n4649), .B1(n3835), .B2(n4955), .ZN(n4430)
         );
  OAI21_X1 U5086 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n4428) );
  NAND2_X1 U5087 ( .A1(n4672), .A2(n4423), .ZN(n4425) );
  OR2_X1 U5088 ( .A1(n4461), .A2(n3157), .ZN(n4424) );
  OAI211_X1 U5089 ( .C1(n4426), .C2(n4654), .A(n4425), .B(n4424), .ZN(n4427)
         );
  AOI21_X1 U5090 ( .B1(n4428), .B2(n3145), .A(n4427), .ZN(n4724) );
  NOR2_X1 U5091 ( .A1(n4724), .A2(n2132), .ZN(n4429) );
  AOI211_X1 U5092 ( .C1(n4668), .C2(n4722), .A(n4430), .B(n4429), .ZN(n4431)
         );
  OAI21_X1 U5093 ( .B1(n4725), .B2(n4670), .A(n4431), .ZN(U3263) );
  XNOR2_X1 U5094 ( .A(n4432), .B(n4436), .ZN(n4727) );
  INV_X1 U5095 ( .A(n4727), .ZN(n4451) );
  OAI21_X1 U5096 ( .B1(n4433), .B2(n4435), .A(n4434), .ZN(n4437) );
  XNOR2_X1 U5097 ( .A(n4437), .B(n4436), .ZN(n4438) );
  NAND2_X1 U5098 ( .A1(n4438), .A2(n3145), .ZN(n4441) );
  AOI22_X1 U5099 ( .A1(n4479), .A2(n4696), .B1(n4439), .B2(n4672), .ZN(n4440)
         );
  OAI211_X1 U5100 ( .C1(n4442), .C2(n4654), .A(n4441), .B(n4440), .ZN(n4726)
         );
  INV_X1 U5101 ( .A(n4443), .ZN(n4446) );
  OAI21_X1 U5102 ( .B1(n4446), .B2(n4445), .A(n4444), .ZN(n4807) );
  AOI22_X1 U5103 ( .A1(n4447), .A2(n4950), .B1(REG2_REG_26__SCAN_IN), .B2(
        n2132), .ZN(n4448) );
  OAI21_X1 U5104 ( .B1(n4807), .B2(n4711), .A(n4448), .ZN(n4449) );
  AOI21_X1 U5105 ( .B1(n4726), .B2(n4955), .A(n4449), .ZN(n4450) );
  OAI21_X1 U5106 ( .B1(n4451), .B2(n4670), .A(n4450), .ZN(U3264) );
  XOR2_X1 U5107 ( .A(n4455), .B(n4452), .Z(n4731) );
  INV_X1 U5108 ( .A(n4731), .ZN(n4469) );
  NAND2_X1 U5109 ( .A1(n4454), .A2(n4453), .ZN(n4456) );
  XNOR2_X1 U5110 ( .A(n4456), .B(n4455), .ZN(n4457) );
  NAND2_X1 U5111 ( .A1(n4457), .A2(n3145), .ZN(n4460) );
  AOI22_X1 U5112 ( .A1(n4498), .A2(n4696), .B1(n4458), .B2(n4672), .ZN(n4459)
         );
  OAI211_X1 U5113 ( .C1(n4461), .C2(n4654), .A(n4460), .B(n4459), .ZN(n4730)
         );
  OR2_X1 U5114 ( .A1(n4482), .A2(n4462), .ZN(n4463) );
  NAND2_X1 U5115 ( .A1(n4443), .A2(n4463), .ZN(n4811) );
  NOR2_X1 U5116 ( .A1(n4811), .A2(n4711), .ZN(n4467) );
  OAI22_X1 U5117 ( .A1(n4465), .A2(n4649), .B1(n4464), .B2(n4955), .ZN(n4466)
         );
  AOI211_X1 U5118 ( .C1(n4730), .C2(n4955), .A(n4467), .B(n4466), .ZN(n4468)
         );
  OAI21_X1 U5119 ( .B1(n4469), .B2(n4670), .A(n4468), .ZN(U3265) );
  XOR2_X1 U5120 ( .A(n4471), .B(n4470), .Z(n4735) );
  INV_X1 U5121 ( .A(n4735), .ZN(n4490) );
  NAND2_X1 U5122 ( .A1(n4473), .A2(n4472), .ZN(n4475) );
  XNOR2_X1 U5123 ( .A(n4475), .B(n4474), .ZN(n4476) );
  NAND2_X1 U5124 ( .A1(n4476), .A2(n3145), .ZN(n4481) );
  NAND2_X1 U5125 ( .A1(n4519), .A2(n4696), .ZN(n4477) );
  OAI21_X1 U5126 ( .B1(n4700), .B2(n4484), .A(n4477), .ZN(n4478) );
  AOI21_X1 U5127 ( .B1(n4479), .B2(n4697), .A(n4478), .ZN(n4480) );
  NAND2_X1 U5128 ( .A1(n4481), .A2(n4480), .ZN(n4734) );
  INV_X1 U5129 ( .A(n4504), .ZN(n4485) );
  INV_X1 U5130 ( .A(n4482), .ZN(n4483) );
  OAI21_X1 U5131 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(n4815) );
  AOI22_X1 U5132 ( .A1(n4486), .A2(n4950), .B1(REG2_REG_24__SCAN_IN), .B2(
        n2132), .ZN(n4487) );
  OAI21_X1 U5133 ( .B1(n4815), .B2(n4711), .A(n4487), .ZN(n4488) );
  AOI21_X1 U5134 ( .B1(n4734), .B2(n4955), .A(n4488), .ZN(n4489) );
  OAI21_X1 U5135 ( .B1(n4490), .B2(n4670), .A(n4489), .ZN(U3266) );
  XOR2_X1 U5136 ( .A(n4495), .B(n4491), .Z(n4739) );
  INV_X1 U5137 ( .A(n4739), .ZN(n4510) );
  NAND2_X1 U5138 ( .A1(n4492), .A2(n4531), .ZN(n4530) );
  NAND2_X1 U5139 ( .A1(n4530), .A2(n4493), .ZN(n4515) );
  NAND2_X1 U5140 ( .A1(n4515), .A2(n2293), .ZN(n4514) );
  NAND2_X1 U5141 ( .A1(n4514), .A2(n4494), .ZN(n4496) );
  XNOR2_X1 U5142 ( .A(n4496), .B(n4495), .ZN(n4500) );
  OAI22_X1 U5143 ( .A1(n4536), .A2(n3157), .B1(n4700), .B2(n3092), .ZN(n4497)
         );
  AOI21_X1 U5144 ( .B1(n4697), .B2(n4498), .A(n4497), .ZN(n4499) );
  OAI21_X1 U5145 ( .B1(n4500), .B2(n4661), .A(n4499), .ZN(n4738) );
  NAND2_X1 U5146 ( .A1(n4501), .A2(n4502), .ZN(n4503) );
  NAND2_X1 U5147 ( .A1(n4504), .A2(n4503), .ZN(n4819) );
  NOR2_X1 U5148 ( .A1(n4819), .A2(n4711), .ZN(n4508) );
  OAI22_X1 U5149 ( .A1(n4506), .A2(n4649), .B1(n4505), .B2(n4955), .ZN(n4507)
         );
  AOI211_X1 U5150 ( .C1(n4738), .C2(n4955), .A(n4508), .B(n4507), .ZN(n4509)
         );
  OAI21_X1 U5151 ( .B1(n4510), .B2(n4670), .A(n4509), .ZN(U3267) );
  OAI21_X1 U5152 ( .B1(n4513), .B2(n4512), .A(n4511), .ZN(n4745) );
  OAI21_X1 U5153 ( .B1(n2293), .B2(n4515), .A(n4514), .ZN(n4516) );
  NAND2_X1 U5154 ( .A1(n4516), .A2(n3145), .ZN(n4521) );
  OAI22_X1 U5155 ( .A1(n4517), .A2(n3157), .B1(n4524), .B2(n4700), .ZN(n4518)
         );
  AOI21_X1 U5156 ( .B1(n4697), .B2(n4519), .A(n4518), .ZN(n4520) );
  AOI22_X1 U5157 ( .A1(n4522), .A2(n4950), .B1(n2132), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4526) );
  OR2_X1 U5158 ( .A1(n4523), .A2(n4524), .ZN(n4742) );
  NAND3_X1 U5159 ( .A1(n4742), .A2(n4501), .A3(n4668), .ZN(n4525) );
  OAI211_X1 U5160 ( .C1(n4744), .C2(n2132), .A(n4526), .B(n4525), .ZN(n4527)
         );
  INV_X1 U5161 ( .A(n4527), .ZN(n4528) );
  OAI21_X1 U5162 ( .B1(n4745), .B2(n4670), .A(n4528), .ZN(U3268) );
  XOR2_X1 U5163 ( .A(n4531), .B(n4529), .Z(n4747) );
  INV_X1 U5164 ( .A(n4747), .ZN(n4543) );
  OAI21_X1 U5165 ( .B1(n4531), .B2(n4492), .A(n4530), .ZN(n4532) );
  NAND2_X1 U5166 ( .A1(n4532), .A2(n3145), .ZN(n4535) );
  AOI22_X1 U5167 ( .A1(n4576), .A2(n4696), .B1(n4672), .B2(n4533), .ZN(n4534)
         );
  OAI211_X1 U5168 ( .C1(n4536), .C2(n4654), .A(n4535), .B(n4534), .ZN(n4746)
         );
  NOR2_X1 U5169 ( .A1(n4560), .A2(n4537), .ZN(n4538) );
  OR2_X1 U5170 ( .A1(n4523), .A2(n4538), .ZN(n4824) );
  AOI22_X1 U5171 ( .A1(n2132), .A2(REG2_REG_21__SCAN_IN), .B1(n4539), .B2(
        n4950), .ZN(n4540) );
  OAI21_X1 U5172 ( .B1(n4824), .B2(n4711), .A(n4540), .ZN(n4541) );
  AOI21_X1 U5173 ( .B1(n4746), .B2(n4652), .A(n4541), .ZN(n4542) );
  OAI21_X1 U5174 ( .B1(n4543), .B2(n4670), .A(n4542), .ZN(U3269) );
  AOI21_X1 U5175 ( .B1(n4544), .B2(n4546), .A(n4545), .ZN(n4547) );
  XNOR2_X1 U5176 ( .A(n4547), .B(n4551), .ZN(n4751) );
  INV_X1 U5177 ( .A(n4751), .ZN(n4566) );
  INV_X1 U5178 ( .A(n4549), .ZN(n4550) );
  NAND2_X1 U5179 ( .A1(n4548), .A2(n4550), .ZN(n4552) );
  XOR2_X1 U5180 ( .A(n4552), .B(n4551), .Z(n4557) );
  OAI22_X1 U5181 ( .A1(n4592), .A2(n3157), .B1(n4553), .B2(n4700), .ZN(n4554)
         );
  AOI21_X1 U5182 ( .B1(n4555), .B2(n4697), .A(n4554), .ZN(n4556) );
  OAI21_X1 U5183 ( .B1(n4557), .B2(n4661), .A(n4556), .ZN(n4750) );
  INV_X1 U5184 ( .A(n4558), .ZN(n4582) );
  AND2_X1 U5185 ( .A1(n4582), .A2(n4559), .ZN(n4561) );
  OR2_X1 U5186 ( .A1(n4561), .A2(n4560), .ZN(n4828) );
  AOI22_X1 U5187 ( .A1(n2132), .A2(REG2_REG_20__SCAN_IN), .B1(n4562), .B2(
        n4950), .ZN(n4563) );
  OAI21_X1 U5188 ( .B1(n4828), .B2(n4711), .A(n4563), .ZN(n4564) );
  AOI21_X1 U5189 ( .B1(n4750), .B2(n4652), .A(n4564), .ZN(n4565) );
  OAI21_X1 U5190 ( .B1(n4566), .B2(n4670), .A(n4565), .ZN(U3270) );
  XOR2_X1 U5191 ( .A(n4572), .B(n4544), .Z(n4755) );
  INV_X1 U5192 ( .A(n4755), .ZN(n4588) );
  OAI21_X1 U5193 ( .B1(n4607), .B2(n4568), .A(n4567), .ZN(n4589) );
  INV_X1 U5194 ( .A(n4569), .ZN(n4571) );
  OAI21_X1 U5195 ( .B1(n4589), .B2(n4571), .A(n4570), .ZN(n4573) );
  XNOR2_X1 U5196 ( .A(n4573), .B(n4572), .ZN(n4578) );
  OAI22_X1 U5197 ( .A1(n4610), .A2(n3157), .B1(n4574), .B2(n4700), .ZN(n4575)
         );
  AOI21_X1 U5198 ( .B1(n4697), .B2(n4576), .A(n4575), .ZN(n4577) );
  OAI21_X1 U5199 ( .B1(n4578), .B2(n4661), .A(n4577), .ZN(n4754) );
  NAND2_X1 U5200 ( .A1(n4580), .A2(n4579), .ZN(n4581) );
  NAND2_X1 U5201 ( .A1(n4582), .A2(n4581), .ZN(n4832) );
  NOR2_X1 U5202 ( .A1(n4832), .A2(n4711), .ZN(n4586) );
  OAI22_X1 U5203 ( .A1(n4652), .A2(n4584), .B1(n4583), .B2(n4649), .ZN(n4585)
         );
  AOI211_X1 U5204 ( .C1(n4754), .C2(n4652), .A(n4586), .B(n4585), .ZN(n4587)
         );
  OAI21_X1 U5205 ( .B1(n4588), .B2(n4670), .A(n4587), .ZN(U3271) );
  XOR2_X1 U5206 ( .A(n4597), .B(n4589), .Z(n4594) );
  AOI22_X1 U5207 ( .A1(n4590), .A2(n4696), .B1(n4598), .B2(n4672), .ZN(n4591)
         );
  OAI21_X1 U5208 ( .B1(n4592), .B2(n4654), .A(n4591), .ZN(n4593) );
  AOI21_X1 U5209 ( .B1(n4594), .B2(n3145), .A(n4593), .ZN(n4760) );
  OAI21_X1 U5210 ( .B1(n4595), .B2(n4597), .A(n4596), .ZN(n4758) );
  XNOR2_X1 U5211 ( .A(n2401), .B(n4598), .ZN(n4599) );
  NAND2_X1 U5212 ( .A1(n4599), .A2(n4998), .ZN(n4759) );
  INV_X1 U5213 ( .A(n4600), .ZN(n4603) );
  AOI22_X1 U5214 ( .A1(n2132), .A2(REG2_REG_18__SCAN_IN), .B1(n4601), .B2(
        n4950), .ZN(n4602) );
  OAI21_X1 U5215 ( .B1(n4759), .B2(n4603), .A(n4602), .ZN(n4604) );
  AOI21_X1 U5216 ( .B1(n4758), .B2(n4688), .A(n4604), .ZN(n4605) );
  OAI21_X1 U5217 ( .B1(n4760), .B2(n2132), .A(n4605), .ZN(U3272) );
  INV_X1 U5218 ( .A(n4613), .ZN(n4606) );
  XNOR2_X1 U5219 ( .A(n4607), .B(n4606), .ZN(n4612) );
  AOI22_X1 U5220 ( .A1(n4608), .A2(n4696), .B1(n4672), .B2(n2230), .ZN(n4609)
         );
  OAI21_X1 U5221 ( .B1(n4610), .B2(n4654), .A(n4609), .ZN(n4611) );
  AOI21_X1 U5222 ( .B1(n4612), .B2(n3145), .A(n4611), .ZN(n4763) );
  XNOR2_X1 U5223 ( .A(n4614), .B(n4613), .ZN(n4762) );
  NAND2_X1 U5224 ( .A1(n4762), .A2(n4688), .ZN(n4620) );
  AOI21_X1 U5225 ( .B1(n2230), .B2(n2231), .A(n2401), .ZN(n4837) );
  INV_X1 U5226 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4617) );
  OAI22_X1 U5227 ( .A1(n4652), .A2(n4617), .B1(n4616), .B2(n4649), .ZN(n4618)
         );
  AOI21_X1 U5228 ( .B1(n4837), .B2(n4668), .A(n4618), .ZN(n4619) );
  OAI211_X1 U5229 ( .C1(n4763), .C2(n2132), .A(n4620), .B(n4619), .ZN(U3273)
         );
  OAI22_X1 U5230 ( .A1(n4622), .A2(n4654), .B1(n4621), .B2(n3157), .ZN(n4627)
         );
  OAI211_X1 U5231 ( .C1(n4624), .C2(n4645), .A(n4623), .B(n3145), .ZN(n4625)
         );
  INV_X1 U5232 ( .A(n4625), .ZN(n4626) );
  AOI211_X1 U5233 ( .C1(n4672), .C2(n4631), .A(n4627), .B(n4626), .ZN(n4770)
         );
  OR2_X1 U5234 ( .A1(n4628), .A2(n4629), .ZN(n4630) );
  AOI21_X1 U5235 ( .B1(n4631), .B2(n4630), .A(n4615), .ZN(n4768) );
  OAI22_X1 U5236 ( .A1(n4955), .A2(n4923), .B1(n4632), .B2(n4649), .ZN(n4633)
         );
  AOI21_X1 U5237 ( .B1(n4768), .B2(n4668), .A(n4633), .ZN(n4647) );
  OR2_X1 U5238 ( .A1(n4634), .A2(n4635), .ZN(n4637) );
  NAND2_X1 U5239 ( .A1(n2404), .A2(n4638), .ZN(n4648) );
  NAND2_X1 U5240 ( .A1(n4648), .A2(n4639), .ZN(n4641) );
  NAND2_X1 U5241 ( .A1(n4641), .A2(n4640), .ZN(n4644) );
  INV_X1 U5242 ( .A(n4642), .ZN(n4643) );
  AOI21_X1 U5243 ( .B1(n4645), .B2(n4644), .A(n4643), .ZN(n4769) );
  NAND2_X1 U5244 ( .A1(n4769), .A2(n4688), .ZN(n4646) );
  OAI211_X1 U5245 ( .C1(n4770), .C2(n2132), .A(n4647), .B(n4646), .ZN(U3274)
         );
  XOR2_X1 U5246 ( .A(n4662), .B(n4648), .Z(n4775) );
  XNOR2_X1 U5247 ( .A(n4628), .B(n4653), .ZN(n4772) );
  INV_X1 U5248 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4651) );
  OAI22_X1 U5249 ( .A1(n4652), .A2(n4651), .B1(n4650), .B2(n4649), .ZN(n4667)
         );
  OAI22_X1 U5250 ( .A1(n4655), .A2(n4654), .B1(n4700), .B2(n4653), .ZN(n4665)
         );
  NAND2_X1 U5251 ( .A1(n4656), .A2(n4671), .ZN(n4658) );
  NAND2_X1 U5252 ( .A1(n4658), .A2(n4657), .ZN(n4663) );
  INV_X1 U5253 ( .A(n4663), .ZN(n4660) );
  INV_X1 U5254 ( .A(n4662), .ZN(n4659) );
  AOI211_X1 U5255 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n2394), .ZN(n4664)
         );
  AOI211_X1 U5256 ( .C1(n4696), .C2(n4698), .A(n4665), .B(n4664), .ZN(n4774)
         );
  NOR2_X1 U5257 ( .A1(n4774), .A2(n2132), .ZN(n4666) );
  AOI211_X1 U5258 ( .C1(n4668), .C2(n4772), .A(n4667), .B(n4666), .ZN(n4669)
         );
  OAI21_X1 U5259 ( .B1(n4775), .B2(n4670), .A(n4669), .ZN(U3275) );
  XNOR2_X1 U5260 ( .A(n4656), .B(n4671), .ZN(n4679) );
  NAND2_X1 U5261 ( .A1(n4673), .A2(n4672), .ZN(n4676) );
  NAND2_X1 U5262 ( .A1(n4674), .A2(n4697), .ZN(n4675) );
  OAI211_X1 U5263 ( .C1(n4677), .C2(n3157), .A(n4676), .B(n4675), .ZN(n4678)
         );
  AOI21_X1 U5264 ( .B1(n4679), .B2(n3145), .A(n4678), .ZN(n4777) );
  OAI21_X1 U5265 ( .B1(n4681), .B2(n4680), .A(n2404), .ZN(n4776) );
  OR2_X1 U5266 ( .A1(n4682), .A2(n4683), .ZN(n4684) );
  NAND2_X1 U5267 ( .A1(n4628), .A2(n4684), .ZN(n4844) );
  AOI22_X1 U5268 ( .A1(n2132), .A2(REG2_REG_14__SCAN_IN), .B1(n4685), .B2(
        n4950), .ZN(n4686) );
  OAI21_X1 U5269 ( .B1(n4844), .B2(n4711), .A(n4686), .ZN(n4687) );
  AOI21_X1 U5270 ( .B1(n4776), .B2(n4688), .A(n4687), .ZN(n4689) );
  OAI21_X1 U5271 ( .B1(n2132), .B2(n4777), .A(n4689), .ZN(U3276) );
  XNOR2_X1 U5272 ( .A(n4634), .B(n4694), .ZN(n4705) );
  OAI21_X1 U5273 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(n4693) );
  XOR2_X1 U5274 ( .A(n4694), .B(n4693), .Z(n4702) );
  AOI22_X1 U5275 ( .A1(n4698), .A2(n4697), .B1(n4696), .B2(n4695), .ZN(n4699)
         );
  OAI21_X1 U5276 ( .B1(n4706), .B2(n4700), .A(n4699), .ZN(n4701) );
  AOI21_X1 U5277 ( .B1(n4702), .B2(n3145), .A(n4701), .ZN(n4703) );
  OAI21_X1 U5278 ( .B1(n4704), .B2(n4705), .A(n4703), .ZN(n4781) );
  INV_X1 U5279 ( .A(n4781), .ZN(n4714) );
  INV_X1 U5280 ( .A(n4705), .ZN(n4782) );
  NOR2_X1 U5281 ( .A1(n4707), .A2(n4706), .ZN(n4708) );
  OR2_X1 U5282 ( .A1(n4682), .A2(n4708), .ZN(n4848) );
  AOI22_X1 U5283 ( .A1(n2132), .A2(REG2_REG_13__SCAN_IN), .B1(n4709), .B2(
        n4950), .ZN(n4710) );
  OAI21_X1 U5284 ( .B1(n4848), .B2(n4711), .A(n4710), .ZN(n4712) );
  AOI21_X1 U5285 ( .B1(n4782), .B2(n4952), .A(n4712), .ZN(n4713) );
  OAI21_X1 U5286 ( .B1(n4714), .B2(n2132), .A(n4713), .ZN(U3277) );
  NAND2_X1 U5287 ( .A1(n5022), .A2(n4795), .ZN(n4716) );
  NAND2_X1 U5288 ( .A1(n5019), .A2(REG1_REG_31__SCAN_IN), .ZN(n4715) );
  OAI211_X1 U5289 ( .C1(n4798), .C2(n4794), .A(n4716), .B(n4715), .ZN(U3549)
         );
  NAND2_X1 U5290 ( .A1(n5022), .A2(n4799), .ZN(n4718) );
  NAND2_X1 U5291 ( .A1(n5019), .A2(REG1_REG_30__SCAN_IN), .ZN(n4717) );
  OAI211_X1 U5292 ( .C1(n4802), .C2(n4794), .A(n4718), .B(n4717), .ZN(U3548)
         );
  NAND2_X1 U5293 ( .A1(n4722), .A2(n4998), .ZN(n4723) );
  OAI211_X1 U5294 ( .C1(n4725), .C2(n5005), .A(n4724), .B(n4723), .ZN(n4803)
         );
  MUX2_X1 U5295 ( .A(REG1_REG_27__SCAN_IN), .B(n4803), .S(n5022), .Z(U3545) );
  AOI21_X1 U5296 ( .B1(n4727), .B2(n4787), .A(n4726), .ZN(n4804) );
  MUX2_X1 U5297 ( .A(n4728), .B(n4804), .S(n5022), .Z(n4729) );
  OAI21_X1 U5298 ( .B1(n4794), .B2(n4807), .A(n4729), .ZN(U3544) );
  INV_X1 U5299 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4732) );
  AOI21_X1 U5300 ( .B1(n4731), .B2(n4787), .A(n4730), .ZN(n4808) );
  MUX2_X1 U5301 ( .A(n4732), .B(n4808), .S(n5022), .Z(n4733) );
  OAI21_X1 U5302 ( .B1(n4794), .B2(n4811), .A(n4733), .ZN(U3543) );
  AOI21_X1 U5303 ( .B1(n4735), .B2(n4787), .A(n4734), .ZN(n4812) );
  MUX2_X1 U5304 ( .A(n4736), .B(n4812), .S(n5022), .Z(n4737) );
  OAI21_X1 U5305 ( .B1(n4794), .B2(n4815), .A(n4737), .ZN(U3542) );
  INV_X1 U5306 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4740) );
  AOI21_X1 U5307 ( .B1(n4739), .B2(n4787), .A(n4738), .ZN(n4816) );
  MUX2_X1 U5308 ( .A(n4740), .B(n4816), .S(n5022), .Z(n4741) );
  OAI21_X1 U5309 ( .B1(n4794), .B2(n4819), .A(n4741), .ZN(U3541) );
  NAND3_X1 U5310 ( .A1(n4742), .A2(n4998), .A3(n4501), .ZN(n4743) );
  OAI211_X1 U5311 ( .C1(n4745), .C2(n5005), .A(n4744), .B(n4743), .ZN(n4820)
         );
  MUX2_X1 U5312 ( .A(REG1_REG_22__SCAN_IN), .B(n4820), .S(n5022), .Z(U3540) );
  INV_X1 U5313 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4748) );
  AOI21_X1 U5314 ( .B1(n4747), .B2(n4787), .A(n4746), .ZN(n4821) );
  MUX2_X1 U5315 ( .A(n4748), .B(n4821), .S(n5022), .Z(n4749) );
  OAI21_X1 U5316 ( .B1(n4794), .B2(n4824), .A(n4749), .ZN(U3539) );
  AOI21_X1 U5317 ( .B1(n4751), .B2(n4787), .A(n4750), .ZN(n4825) );
  MUX2_X1 U5318 ( .A(n4752), .B(n4825), .S(n5022), .Z(n4753) );
  OAI21_X1 U5319 ( .B1(n4794), .B2(n4828), .A(n4753), .ZN(U3538) );
  AOI21_X1 U5320 ( .B1(n4755), .B2(n4787), .A(n4754), .ZN(n4829) );
  MUX2_X1 U5321 ( .A(n4756), .B(n4829), .S(n5022), .Z(n4757) );
  OAI21_X1 U5322 ( .B1(n4794), .B2(n4832), .A(n4757), .ZN(U3537) );
  INV_X1 U5323 ( .A(n4758), .ZN(n4761) );
  OAI211_X1 U5324 ( .C1(n4761), .C2(n5005), .A(n4760), .B(n4759), .ZN(n4833)
         );
  MUX2_X1 U5325 ( .A(REG1_REG_18__SCAN_IN), .B(n4833), .S(n5022), .Z(U3536) );
  NAND2_X1 U5326 ( .A1(n4762), .A2(n4787), .ZN(n4764) );
  NAND2_X1 U5327 ( .A1(n4764), .A2(n4763), .ZN(n4834) );
  MUX2_X1 U5328 ( .A(REG1_REG_17__SCAN_IN), .B(n4834), .S(n5022), .Z(n4765) );
  AOI21_X1 U5329 ( .B1(n4766), .B2(n4837), .A(n4765), .ZN(n4767) );
  INV_X1 U5330 ( .A(n4767), .ZN(U3535) );
  AOI22_X1 U5331 ( .A1(n4769), .A2(n4787), .B1(n4768), .B2(n4998), .ZN(n4771)
         );
  NAND2_X1 U5332 ( .A1(n4771), .A2(n4770), .ZN(n4839) );
  MUX2_X1 U5333 ( .A(REG1_REG_16__SCAN_IN), .B(n4839), .S(n5022), .Z(U3534) );
  NAND2_X1 U5334 ( .A1(n4772), .A2(n4998), .ZN(n4773) );
  OAI211_X1 U5335 ( .C1(n5005), .C2(n4775), .A(n4774), .B(n4773), .ZN(n4840)
         );
  MUX2_X1 U5336 ( .A(REG1_REG_15__SCAN_IN), .B(n4840), .S(n5022), .Z(U3533) );
  NAND2_X1 U5337 ( .A1(n4776), .A2(n4787), .ZN(n4778) );
  NAND2_X1 U5338 ( .A1(n4778), .A2(n4777), .ZN(n4841) );
  MUX2_X1 U5339 ( .A(REG1_REG_14__SCAN_IN), .B(n4841), .S(n5022), .Z(n4779) );
  INV_X1 U5340 ( .A(n4779), .ZN(n4780) );
  OAI21_X1 U5341 ( .B1(n4794), .B2(n4844), .A(n4780), .ZN(U3532) );
  AOI21_X1 U5342 ( .B1(n4995), .B2(n4782), .A(n4781), .ZN(n4845) );
  MUX2_X1 U5343 ( .A(n4783), .B(n4845), .S(n5022), .Z(n4784) );
  OAI21_X1 U5344 ( .B1(n4794), .B2(n4848), .A(n4784), .ZN(U3531) );
  INV_X1 U5345 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4788) );
  AOI21_X1 U5346 ( .B1(n4787), .B2(n4786), .A(n4785), .ZN(n4849) );
  MUX2_X1 U5347 ( .A(n4788), .B(n4849), .S(n5022), .Z(n4789) );
  OAI21_X1 U5348 ( .B1(n4794), .B2(n4852), .A(n4789), .ZN(U3530) );
  AOI21_X1 U5349 ( .B1(n4995), .B2(n4791), .A(n4790), .ZN(n4853) );
  MUX2_X1 U5350 ( .A(n4792), .B(n4853), .S(n5022), .Z(n4793) );
  OAI21_X1 U5351 ( .B1(n4794), .B2(n4857), .A(n4793), .ZN(U3529) );
  NAND2_X1 U5352 ( .A1(n5013), .A2(n4795), .ZN(n4797) );
  NAND2_X1 U5353 ( .A1(n5011), .A2(REG0_REG_31__SCAN_IN), .ZN(n4796) );
  OAI211_X1 U5354 ( .C1(n4798), .C2(n4856), .A(n4797), .B(n4796), .ZN(U3517)
         );
  NAND2_X1 U5355 ( .A1(n5013), .A2(n4799), .ZN(n4801) );
  NAND2_X1 U5356 ( .A1(n5011), .A2(REG0_REG_30__SCAN_IN), .ZN(n4800) );
  OAI211_X1 U5357 ( .C1(n4802), .C2(n4856), .A(n4801), .B(n4800), .ZN(U3516)
         );
  MUX2_X1 U5358 ( .A(REG0_REG_27__SCAN_IN), .B(n4803), .S(n5013), .Z(U3513) );
  MUX2_X1 U5359 ( .A(n4805), .B(n4804), .S(n5013), .Z(n4806) );
  OAI21_X1 U5360 ( .B1(n4807), .B2(n4856), .A(n4806), .ZN(U3512) );
  INV_X1 U5361 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4809) );
  MUX2_X1 U5362 ( .A(n4809), .B(n4808), .S(n5013), .Z(n4810) );
  OAI21_X1 U5363 ( .B1(n4811), .B2(n4856), .A(n4810), .ZN(U3511) );
  MUX2_X1 U5364 ( .A(n4813), .B(n4812), .S(n5013), .Z(n4814) );
  OAI21_X1 U5365 ( .B1(n4815), .B2(n4856), .A(n4814), .ZN(U3510) );
  INV_X1 U5366 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4817) );
  MUX2_X1 U5367 ( .A(n4817), .B(n4816), .S(n5013), .Z(n4818) );
  OAI21_X1 U5368 ( .B1(n4819), .B2(n4856), .A(n4818), .ZN(U3509) );
  MUX2_X1 U5369 ( .A(REG0_REG_22__SCAN_IN), .B(n4820), .S(n5013), .Z(U3508) );
  MUX2_X1 U5370 ( .A(n4822), .B(n4821), .S(n5013), .Z(n4823) );
  OAI21_X1 U5371 ( .B1(n4824), .B2(n4856), .A(n4823), .ZN(U3507) );
  MUX2_X1 U5372 ( .A(n4826), .B(n4825), .S(n5013), .Z(n4827) );
  OAI21_X1 U5373 ( .B1(n4828), .B2(n4856), .A(n4827), .ZN(U3506) );
  INV_X1 U5374 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4830) );
  MUX2_X1 U5375 ( .A(n4830), .B(n4829), .S(n5013), .Z(n4831) );
  OAI21_X1 U5376 ( .B1(n4832), .B2(n4856), .A(n4831), .ZN(U3505) );
  MUX2_X1 U5377 ( .A(REG0_REG_18__SCAN_IN), .B(n4833), .S(n5013), .Z(U3503) );
  MUX2_X1 U5378 ( .A(n4834), .B(REG0_REG_17__SCAN_IN), .S(n5011), .Z(n4835) );
  AOI21_X1 U5379 ( .B1(n4837), .B2(n4836), .A(n4835), .ZN(n4838) );
  INV_X1 U5380 ( .A(n4838), .ZN(U3501) );
  MUX2_X1 U5381 ( .A(REG0_REG_16__SCAN_IN), .B(n4839), .S(n5013), .Z(U3499) );
  MUX2_X1 U5382 ( .A(REG0_REG_15__SCAN_IN), .B(n4840), .S(n5013), .Z(U3497) );
  MUX2_X1 U5383 ( .A(REG0_REG_14__SCAN_IN), .B(n4841), .S(n5013), .Z(n4842) );
  INV_X1 U5384 ( .A(n4842), .ZN(n4843) );
  OAI21_X1 U5385 ( .B1(n4844), .B2(n4856), .A(n4843), .ZN(U3495) );
  MUX2_X1 U5386 ( .A(n4846), .B(n4845), .S(n5013), .Z(n4847) );
  OAI21_X1 U5387 ( .B1(n4848), .B2(n4856), .A(n4847), .ZN(U3493) );
  MUX2_X1 U5388 ( .A(n4850), .B(n4849), .S(n5013), .Z(n4851) );
  OAI21_X1 U5389 ( .B1(n4852), .B2(n4856), .A(n4851), .ZN(U3491) );
  MUX2_X1 U5390 ( .A(n4854), .B(n4853), .S(n5013), .Z(n4855) );
  OAI21_X1 U5391 ( .B1(n4857), .B2(n4856), .A(n4855), .ZN(U3489) );
  MUX2_X1 U5392 ( .A(DATAI_30_), .B(n4858), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5393 ( .A(n4859), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5394 ( .A(DATAI_27_), .B(n4860), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5395 ( .A(DATAI_26_), .B(n2602), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  INV_X1 U5396 ( .A(n4861), .ZN(n4862) );
  MUX2_X1 U5397 ( .A(DATAI_25_), .B(n4862), .S(STATE_REG_SCAN_IN), .Z(U3327)
         );
  MUX2_X1 U5398 ( .A(DATAI_20_), .B(n4863), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5399 ( .A(n4864), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5400 ( .A(n4865), .B(DATAI_18_), .S(U3149), .Z(U3334) );
  MUX2_X1 U5401 ( .A(n4913), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5402 ( .A(n4866), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5403 ( .A(DATAI_12_), .B(n4867), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5404 ( .A(DATAI_11_), .B(n4868), .S(STATE_REG_SCAN_IN), .Z(U3341)
         );
  MUX2_X1 U5405 ( .A(n4869), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5406 ( .A(n4870), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5407 ( .A(DATAI_7_), .B(n4871), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5408 ( .A(n4872), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5409 ( .A(n4873), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5410 ( .A(DATAI_4_), .B(n4884), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5411 ( .A(n4874), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5412 ( .A(n2131), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5413 ( .A(n4876), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5414 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5415 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4878) );
  XNOR2_X1 U5416 ( .A(n4879), .B(n4878), .ZN(n4880) );
  NAND2_X1 U5417 ( .A1(n4942), .A2(n4880), .ZN(n4890) );
  INV_X1 U5418 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4881) );
  XNOR2_X1 U5419 ( .A(n4882), .B(n4881), .ZN(n4883) );
  NAND2_X1 U5420 ( .A1(n4940), .A2(n4883), .ZN(n4889) );
  NAND2_X1 U5421 ( .A1(n4914), .A2(n4884), .ZN(n4888) );
  INV_X1 U5422 ( .A(n4885), .ZN(n4886) );
  AOI21_X1 U5423 ( .B1(n4930), .B2(ADDR_REG_4__SCAN_IN), .A(n4886), .ZN(n4887)
         );
  AND4_X1 U5424 ( .A1(n4890), .A2(n4889), .A3(n4888), .A4(n4887), .ZN(n4892)
         );
  NAND2_X1 U5425 ( .A1(n4892), .A2(n4891), .ZN(U3244) );
  AOI211_X1 U5426 ( .C1(n4895), .C2(n4894), .A(n4893), .B(n4908), .ZN(n4900)
         );
  AOI211_X1 U5427 ( .C1(n4898), .C2(n4897), .A(n4896), .B(n4905), .ZN(n4899)
         );
  AOI211_X1 U5428 ( .C1(n4914), .C2(n4901), .A(n4900), .B(n4899), .ZN(n4903)
         );
  OAI211_X1 U5429 ( .C1(n4918), .C2(n4904), .A(n4903), .B(n4902), .ZN(U3254)
         );
  AOI211_X1 U5430 ( .C1(n4907), .C2(n4906), .A(n4905), .B(n2155), .ZN(n4912)
         );
  AOI211_X1 U5431 ( .C1(n4910), .C2(n4909), .A(n4908), .B(n2156), .ZN(n4911)
         );
  AOI211_X1 U5432 ( .C1(n4914), .C2(n4913), .A(n4912), .B(n4911), .ZN(n4916)
         );
  OAI211_X1 U5433 ( .C1(n4918), .C2(n4917), .A(n4916), .B(n4915), .ZN(U3255)
         );
  AOI21_X1 U5434 ( .B1(n4930), .B2(ADDR_REG_16__SCAN_IN), .A(n4919), .ZN(n4928) );
  NAND2_X1 U5435 ( .A1(n4921), .A2(n4920), .ZN(n4931) );
  OAI21_X1 U5436 ( .B1(n4921), .B2(n4920), .A(n4931), .ZN(n4926) );
  OAI21_X1 U5437 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4925) );
  AOI22_X1 U5438 ( .A1(n4942), .A2(n4926), .B1(n4940), .B2(n4925), .ZN(n4927)
         );
  OAI211_X1 U5439 ( .C1(n4978), .C2(n4945), .A(n4928), .B(n4927), .ZN(U3256)
         );
  AOI21_X1 U5440 ( .B1(n4930), .B2(ADDR_REG_17__SCAN_IN), .A(n4929), .ZN(n4944) );
  NAND2_X1 U5441 ( .A1(n4932), .A2(n4931), .ZN(n4934) );
  OAI21_X1 U5442 ( .B1(n4935), .B2(n4934), .A(n4933), .ZN(n4941) );
  OAI21_X1 U5443 ( .B1(n4938), .B2(n4937), .A(n4936), .ZN(n4939) );
  AOI22_X1 U5444 ( .A1(n4942), .A2(n4941), .B1(n4940), .B2(n4939), .ZN(n4943)
         );
  OAI211_X1 U5445 ( .C1(n4976), .C2(n4945), .A(n4944), .B(n4943), .ZN(U3257)
         );
  INV_X1 U5446 ( .A(n4946), .ZN(n4948) );
  AOI21_X1 U5447 ( .B1(n4949), .B2(n4948), .A(n4947), .ZN(n4956) );
  AOI22_X1 U5448 ( .A1(n4952), .A2(n4951), .B1(REG3_REG_0__SCAN_IN), .B2(n4950), .ZN(n4953) );
  OAI221_X1 U5449 ( .B1(n2132), .B2(n4956), .C1(n4955), .C2(n4954), .A(n4953), 
        .ZN(U3290) );
  AND2_X1 U5450 ( .A1(D_REG_31__SCAN_IN), .A2(n4972), .ZN(U3291) );
  NOR2_X1 U5451 ( .A1(n4971), .A2(n4957), .ZN(U3292) );
  AND2_X1 U5452 ( .A1(D_REG_29__SCAN_IN), .A2(n4972), .ZN(U3293) );
  NOR2_X1 U5453 ( .A1(n4971), .A2(n4958), .ZN(U3294) );
  NOR2_X1 U5454 ( .A1(n4971), .A2(n4959), .ZN(U3295) );
  NOR2_X1 U5455 ( .A1(n4971), .A2(n4960), .ZN(U3296) );
  AND2_X1 U5456 ( .A1(D_REG_25__SCAN_IN), .A2(n4972), .ZN(U3297) );
  NOR2_X1 U5457 ( .A1(n4971), .A2(n4961), .ZN(U3298) );
  AND2_X1 U5458 ( .A1(D_REG_23__SCAN_IN), .A2(n4972), .ZN(U3299) );
  NOR2_X1 U5459 ( .A1(n4971), .A2(n4962), .ZN(U3300) );
  NOR2_X1 U5460 ( .A1(n4971), .A2(n4963), .ZN(U3301) );
  NOR2_X1 U5461 ( .A1(n4971), .A2(n4964), .ZN(U3302) );
  AND2_X1 U5462 ( .A1(D_REG_19__SCAN_IN), .A2(n4972), .ZN(U3303) );
  AND2_X1 U5463 ( .A1(D_REG_18__SCAN_IN), .A2(n4972), .ZN(U3304) );
  NOR2_X1 U5464 ( .A1(n4971), .A2(n4965), .ZN(U3305) );
  NOR2_X1 U5465 ( .A1(n4971), .A2(n4966), .ZN(U3306) );
  AND2_X1 U5466 ( .A1(D_REG_15__SCAN_IN), .A2(n4972), .ZN(U3307) );
  AND2_X1 U5467 ( .A1(D_REG_14__SCAN_IN), .A2(n4972), .ZN(U3308) );
  NOR2_X1 U5468 ( .A1(n4971), .A2(n4967), .ZN(U3309) );
  NOR2_X1 U5469 ( .A1(n4971), .A2(n4968), .ZN(U3310) );
  AND2_X1 U5470 ( .A1(D_REG_11__SCAN_IN), .A2(n4972), .ZN(U3311) );
  NOR2_X1 U5471 ( .A1(n4971), .A2(n4969), .ZN(U3312) );
  AND2_X1 U5472 ( .A1(D_REG_9__SCAN_IN), .A2(n4972), .ZN(U3313) );
  AND2_X1 U5473 ( .A1(D_REG_8__SCAN_IN), .A2(n4972), .ZN(U3314) );
  AND2_X1 U5474 ( .A1(D_REG_7__SCAN_IN), .A2(n4972), .ZN(U3315) );
  AND2_X1 U5475 ( .A1(D_REG_6__SCAN_IN), .A2(n4972), .ZN(U3316) );
  NOR2_X1 U5476 ( .A1(n4971), .A2(n4970), .ZN(U3317) );
  AND2_X1 U5477 ( .A1(D_REG_4__SCAN_IN), .A2(n4972), .ZN(U3318) );
  AND2_X1 U5478 ( .A1(D_REG_3__SCAN_IN), .A2(n4972), .ZN(U3319) );
  AND2_X1 U5479 ( .A1(D_REG_2__SCAN_IN), .A2(n4972), .ZN(U3320) );
  OAI21_X1 U5480 ( .B1(STATE_REG_SCAN_IN), .B2(DATAI_23_), .A(n4973), .ZN(
        n4974) );
  INV_X1 U5481 ( .A(n4974), .ZN(U3329) );
  AOI22_X1 U5482 ( .A1(STATE_REG_SCAN_IN), .A2(n4976), .B1(n4975), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5483 ( .A1(STATE_REG_SCAN_IN), .A2(n4978), .B1(n4977), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5484 ( .A1(STATE_REG_SCAN_IN), .A2(n4980), .B1(n4979), .B2(U3149), 
        .ZN(U3338) );
  INV_X1 U5485 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4981) );
  AOI22_X1 U5486 ( .A1(n5013), .A2(n4982), .B1(n4981), .B2(n5011), .ZN(U3467)
         );
  INV_X1 U5487 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4983) );
  AOI22_X1 U5488 ( .A1(n5013), .A2(n4984), .B1(n4983), .B2(n5011), .ZN(U3469)
         );
  OAI22_X1 U5489 ( .A1(n4988), .A2(n4987), .B1(n4986), .B2(n4985), .ZN(n4989)
         );
  NOR2_X1 U5490 ( .A1(n4990), .A2(n4989), .ZN(n5015) );
  INV_X1 U5491 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4991) );
  AOI22_X1 U5492 ( .A1(n5013), .A2(n5015), .B1(n4991), .B2(n5011), .ZN(U3473)
         );
  INV_X1 U5493 ( .A(n4992), .ZN(n4993) );
  AOI211_X1 U5494 ( .C1(n4996), .C2(n4995), .A(n4994), .B(n4993), .ZN(n5016)
         );
  AOI22_X1 U5495 ( .A1(n5013), .A2(n5016), .B1(n4997), .B2(n5011), .ZN(U3475)
         );
  NAND2_X1 U5496 ( .A1(n4999), .A2(n4998), .ZN(n5000) );
  OAI211_X1 U5497 ( .C1(n5002), .C2(n5005), .A(n5001), .B(n5000), .ZN(n5003)
         );
  INV_X1 U5498 ( .A(n5003), .ZN(n5018) );
  AOI22_X1 U5499 ( .A1(n5013), .A2(n5018), .B1(n5004), .B2(n5011), .ZN(U3477)
         );
  NOR3_X1 U5500 ( .A1(n5007), .A2(n5006), .A3(n5005), .ZN(n5010) );
  NOR3_X1 U5501 ( .A1(n5010), .A2(n5009), .A3(n5008), .ZN(n5021) );
  INV_X1 U5502 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5012) );
  AOI22_X1 U5503 ( .A1(n5013), .A2(n5021), .B1(n5012), .B2(n5011), .ZN(U3481)
         );
  INV_X1 U5504 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5014) );
  AOI22_X1 U5505 ( .A1(n5022), .A2(n5015), .B1(n5014), .B2(n5019), .ZN(U3521)
         );
  AOI22_X1 U5506 ( .A1(n5022), .A2(n5016), .B1(n4878), .B2(n5019), .ZN(U3522)
         );
  AOI22_X1 U5507 ( .A1(n5022), .A2(n5018), .B1(n5017), .B2(n5019), .ZN(U3523)
         );
  AOI22_X1 U5508 ( .A1(n5022), .A2(n5021), .B1(n5020), .B2(n5019), .ZN(U3525)
         );
  CLKBUF_X3 U2373 ( .A(n3990), .Z(n2134) );
  CLKBUF_X1 U2411 ( .A(n4652), .Z(n4955) );
endmodule

