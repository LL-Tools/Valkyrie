

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput63, keyinput62, keyinput61, keyinput60, keyinput59, keyinput58, 
        keyinput57, keyinput56, keyinput55, keyinput54, keyinput53, keyinput52, 
        keyinput51, keyinput50, keyinput49, keyinput48, keyinput47, keyinput46, 
        keyinput45, keyinput44, keyinput43, keyinput42, keyinput41, keyinput40, 
        keyinput39, keyinput38, keyinput37, keyinput36, keyinput35, keyinput34, 
        keyinput33, keyinput32, keyinput31, keyinput30, keyinput29, keyinput28, 
        keyinput27, keyinput26, keyinput25, keyinput24, keyinput23, keyinput22, 
        keyinput21, keyinput20, keyinput19, keyinput18, keyinput17, keyinput16, 
        keyinput15, keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, 
        keyinput9, keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, 
        keyinput3, keyinput2, keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135;

  OAI21_X1 U4796 ( .B1(n5366), .B2(n5365), .A(n5364), .ZN(n5372) );
  BUF_X2 U4797 ( .A(n6572), .Z(n4295) );
  CLKBUF_X2 U4798 ( .A(n5704), .Z(n8729) );
  AND2_X1 U4799 ( .A1(n8737), .A2(n8868), .ZN(n6784) );
  BUF_X1 U4800 ( .A(n8616), .Z(n4307) );
  AND2_X1 U4801 ( .A1(n6516), .A2(n6515), .ZN(n7571) );
  NOR2_X1 U4802 ( .A1(n9964), .A2(n9963), .ZN(n9962) );
  INV_X1 U4803 ( .A(n4292), .ZN(n4293) );
  OR2_X1 U4804 ( .A1(n7154), .A2(n7058), .ZN(n8653) );
  BUF_X1 U4806 ( .A(n7210), .Z(n7583) );
  NOR2_X1 U4807 ( .A1(n9962), .A2(n4407), .ZN(n8063) );
  OR2_X1 U4808 ( .A1(n8109), .A2(n8110), .ZN(n4693) );
  OAI22_X1 U4809 ( .A1(n8186), .A2(n5456), .B1(n7968), .B2(n5499), .ZN(n5561)
         );
  INV_X1 U4810 ( .A(n7903), .ZN(n7907) );
  CLKBUF_X3 U4811 ( .A(n5058), .Z(n7739) );
  NAND2_X1 U4812 ( .A1(n4591), .A2(n4383), .ZN(n8482) );
  INV_X1 U4813 ( .A(n6139), .ZN(n7620) );
  INV_X1 U4814 ( .A(n4307), .ZN(n5736) );
  NAND2_X1 U4815 ( .A1(n8803), .A2(n8662), .ZN(n8763) );
  INV_X1 U4816 ( .A(n6995), .ZN(n9799) );
  NAND2_X1 U4817 ( .A1(n8789), .A2(n6753), .ZN(n6772) );
  NAND2_X1 U4818 ( .A1(n5802), .A2(n5801), .ZN(n7339) );
  NAND2_X1 U4819 ( .A1(n6164), .A2(n6163), .ZN(n9228) );
  INV_X2 U4820 ( .A(n5642), .ZN(n7747) );
  AND4_X1 U4821 ( .A1(n4741), .A2(n5165), .A3(n4740), .A4(n5149), .ZN(n4290)
         );
  INV_X1 U4822 ( .A(n5687), .ZN(n4292) );
  XNOR2_X1 U4823 ( .A(n5087), .B(P2_IR_REG_2__SCAN_IN), .ZN(n6572) );
  AND2_X2 U4824 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9565) );
  NAND2_X2 U4826 ( .A1(n6777), .A2(n8791), .ZN(n9747) );
  AOI211_X2 U4827 ( .C1(n9959), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8128), .B(
        n8127), .ZN(n8135) );
  OAI21_X2 U4828 ( .B1(n6934), .B2(n6936), .A(n6935), .ZN(n5777) );
  NOR2_X2 U4829 ( .A1(n9892), .A2(n6551), .ZN(n9891) );
  NAND2_X1 U4830 ( .A1(n7611), .A2(n9677), .ZN(n4310) );
  NAND2_X1 U4831 ( .A1(n7611), .A2(n9677), .ZN(n4311) );
  NAND2_X1 U4832 ( .A1(n5606), .A2(n5605), .ZN(n4291) );
  INV_X2 U4833 ( .A(n4292), .ZN(n4294) );
  NAND4_X2 U4834 ( .A1(n5715), .A2(n5714), .A3(n5713), .A4(n5712), .ZN(n8896)
         );
  NOR4_X2 U4835 ( .A1(n8863), .A2(n8862), .A3(n8861), .A4(n8860), .ZN(n8883)
         );
  NAND2_X2 U4836 ( .A1(n5646), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5648) );
  NOR2_X1 U4837 ( .A1(n8898), .A2(n9775), .ZN(n6776) );
  NAND4_X2 U4838 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(n8898)
         );
  OAI22_X2 U4839 ( .A1(n8235), .A2(n7922), .B1(n7972), .B2(n7703), .ZN(n8225)
         );
  AOI22_X2 U4840 ( .A1(n8245), .A2(n8251), .B1(n8426), .B2(n8261), .ZN(n8235)
         );
  NAND2_X2 U4841 ( .A1(n5840), .A2(n5839), .ZN(n7154) );
  OAI211_X2 U4842 ( .C1(n4311), .C2(n6657), .A(n5686), .B(n5685), .ZN(n6767)
         );
  OR2_X1 U4843 ( .A1(n5797), .A2(n6251), .ZN(n5686) );
  NAND2_X2 U4844 ( .A1(n5877), .A2(n5876), .ZN(n7510) );
  INV_X1 U4845 ( .A(n6449), .ZN(n8145) );
  XNOR2_X1 U4846 ( .A(n9172), .B(n9195), .ZN(n9431) );
  NAND2_X1 U4847 ( .A1(n6019), .A2(n8573), .ZN(n8501) );
  NAND2_X1 U4848 ( .A1(n5956), .A2(n5955), .ZN(n5960) );
  NAND2_X1 U4849 ( .A1(n4735), .A2(n4982), .ZN(n5204) );
  INV_X1 U4850 ( .A(n9656), .ZN(n9808) );
  INV_X1 U4851 ( .A(n9671), .ZN(n9789) );
  NAND2_X1 U4852 ( .A1(n5073), .A2(n6794), .ZN(n5489) );
  CLKBUF_X1 U4853 ( .A(n5086), .Z(n5169) );
  CLKBUF_X2 U4854 ( .A(n8616), .Z(n4306) );
  OR2_X2 U4856 ( .A1(n7603), .A2(n8455), .ZN(n5076) );
  NAND2_X1 U4857 ( .A1(n5606), .A2(n9555), .ZN(n8620) );
  AND2_X1 U4858 ( .A1(n4560), .A2(n4559), .ZN(n5028) );
  AND2_X1 U4859 ( .A1(n5798), .A2(n5598), .ZN(n4685) );
  AND2_X1 U4860 ( .A1(n4875), .A2(n4873), .ZN(n6183) );
  NAND2_X1 U4861 ( .A1(n9206), .A2(n9171), .ZN(n9172) );
  AND2_X1 U4862 ( .A1(n8736), .A2(n8867), .ZN(n8864) );
  NAND2_X1 U4863 ( .A1(n4660), .A2(n4361), .ZN(n9206) );
  NOR3_X1 U4864 ( .A1(n8871), .A2(n8832), .A3(n8775), .ZN(n8857) );
  NOR2_X1 U4865 ( .A1(n7900), .A2(n7899), .ZN(n7908) );
  INV_X1 U4866 ( .A(n8740), .ZN(n9500) );
  INV_X1 U4867 ( .A(n9195), .ZN(n4447) );
  OR2_X1 U4868 ( .A1(n9428), .A2(n8725), .ZN(n8778) );
  NAND2_X1 U4869 ( .A1(n8723), .A2(n8722), .ZN(n9428) );
  NAND2_X1 U4870 ( .A1(n7614), .A2(n7613), .ZN(n9212) );
  AOI21_X1 U4871 ( .B1(n4567), .B2(n5960), .A(n4568), .ZN(n4566) );
  NAND2_X1 U4872 ( .A1(n5567), .A2(n5566), .ZN(n7593) );
  AND2_X1 U4873 ( .A1(n5960), .A2(n5959), .ZN(n4570) );
  NAND2_X1 U4874 ( .A1(n8257), .A2(n5333), .ZN(n8245) );
  XNOR2_X1 U4875 ( .A(n5458), .B(n5457), .ZN(n8463) );
  OR2_X1 U4876 ( .A1(n5956), .A2(n5955), .ZN(n4906) );
  OR2_X1 U4877 ( .A1(n9275), .A2(n8697), .ZN(n9185) );
  INV_X1 U4878 ( .A(n7880), .ZN(n4296) );
  NAND2_X1 U4879 ( .A1(n9146), .A2(n9145), .ZN(n9373) );
  AOI21_X2 U4880 ( .B1(n7365), .B2(n7753), .A(n4404), .ZN(n8415) );
  OR2_X1 U4881 ( .A1(n8038), .A2(n8039), .ZN(n4597) );
  NAND2_X1 U4882 ( .A1(n5393), .A2(n5404), .ZN(n7365) );
  NAND2_X1 U4883 ( .A1(n6041), .A2(n6040), .ZN(n9471) );
  NAND2_X1 U4884 ( .A1(n6023), .A2(n6022), .ZN(n9356) );
  NAND2_X1 U4885 ( .A1(n8744), .A2(n8838), .ZN(n4674) );
  OR2_X1 U4886 ( .A1(n9411), .A2(n8645), .ZN(n8744) );
  NAND2_X1 U4887 ( .A1(n9411), .A2(n8645), .ZN(n8838) );
  NAND2_X1 U4888 ( .A1(n5941), .A2(n5940), .ZN(n9139) );
  NAND2_X1 U4889 ( .A1(n8658), .A2(n8656), .ZN(n7371) );
  NAND2_X1 U4890 ( .A1(n8653), .A2(n8650), .ZN(n8758) );
  NAND2_X1 U4891 ( .A1(n5173), .A2(n5172), .ZN(n7042) );
  NAND2_X1 U4892 ( .A1(n5859), .A2(n5858), .ZN(n7305) );
  INV_X1 U4893 ( .A(n7031), .ZN(n9813) );
  XNOR2_X1 U4894 ( .A(n5204), .B(n5203), .ZN(n6294) );
  NAND2_X1 U4895 ( .A1(n7074), .A2(n7082), .ZN(n7073) );
  OR2_X1 U4896 ( .A1(n7072), .A2(n7071), .ZN(n7074) );
  NAND2_X1 U4897 ( .A1(n5094), .A2(n5093), .ZN(n6719) );
  OAI21_X1 U4898 ( .B1(n5183), .B2(n5184), .A(n4977), .ZN(n5196) );
  INV_X2 U4899 ( .A(n10016), .ZN(n8334) );
  NAND2_X1 U4900 ( .A1(n4698), .A2(n9942), .ZN(n6886) );
  NAND2_X2 U4901 ( .A1(n6764), .A2(n9741), .ZN(n9394) );
  INV_X1 U4902 ( .A(n8497), .ZN(n9783) );
  NAND2_X1 U4903 ( .A1(n5705), .A2(n4466), .ZN(n8497) );
  NAND2_X1 U4904 ( .A1(n4962), .A2(n4961), .ZN(n5136) );
  NAND2_X1 U4905 ( .A1(n5083), .A2(n5082), .ZN(n5092) );
  OR2_X1 U4906 ( .A1(n4601), .A2(n6567), .ZN(n9926) );
  INV_X1 U4907 ( .A(n5655), .ZN(n6139) );
  NAND4_X1 U4908 ( .A1(n5665), .A2(n5664), .A3(n5663), .A4(n5662), .ZN(n6771)
         );
  INV_X2 U4909 ( .A(n5169), .ZN(n7753) );
  AND2_X2 U4910 ( .A1(n6244), .A2(n6279), .ZN(P1_U3973) );
  CLKBUF_X1 U4911 ( .A(n7739), .Z(n5460) );
  INV_X2 U4912 ( .A(n5078), .ZN(n6839) );
  NAND3_X1 U4913 ( .A1(n8870), .A2(n5651), .A3(n6785), .ZN(n5652) );
  CLKBUF_X3 U4914 ( .A(n8620), .Z(n4309) );
  INV_X1 U4915 ( .A(n8615), .ZN(n6218) );
  OR2_X1 U4916 ( .A1(n4291), .A2(n6626), .ZN(n5608) );
  NAND2_X1 U4917 ( .A1(n6185), .A2(n5621), .ZN(n6243) );
  NAND2_X2 U4918 ( .A1(n7635), .A2(n5605), .ZN(n8615) );
  NAND2_X2 U4919 ( .A1(n4584), .A2(n4582), .ZN(n8868) );
  CLKBUF_X2 U4920 ( .A(n5604), .Z(n7635) );
  INV_X1 U4921 ( .A(n9555), .ZN(n5605) );
  XNOR2_X1 U4922 ( .A(n4920), .B(n4919), .ZN(n7603) );
  OR2_X1 U4923 ( .A1(n5631), .A2(n5838), .ZN(n5633) );
  XNOR2_X1 U4924 ( .A(n5603), .B(n5602), .ZN(n9555) );
  NAND2_X1 U4925 ( .A1(n5634), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U4926 ( .A1(n5645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6002) );
  INV_X2 U4927 ( .A(n8465), .ZN(n8456) );
  XNOR2_X1 U4928 ( .A(n4956), .B(SI_3_), .ZN(n5104) );
  OAI21_X1 U4929 ( .B1(n6249), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4459), .ZN(
        n4953) );
  XNOR2_X1 U4930 ( .A(n5102), .B(n4820), .ZN(n9888) );
  AND2_X2 U4931 ( .A1(n4685), .A2(n4871), .ZN(n5617) );
  INV_X2 U4932 ( .A(n5642), .ZN(n6249) );
  OR2_X1 U4933 ( .A1(n4917), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4765) );
  NOR2_X1 U4934 ( .A1(n4915), .A2(n4914), .ZN(n4916) );
  NOR2_X1 U4935 ( .A1(n4893), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4892) );
  AND2_X2 U4936 ( .A1(n4702), .A2(n4703), .ZN(n5642) );
  AND2_X1 U4937 ( .A1(n6430), .A2(n4907), .ZN(n4908) );
  NAND2_X1 U4938 ( .A1(n9565), .A2(n4946), .ZN(n4702) );
  AND2_X2 U4939 ( .A1(n5638), .A2(n5684), .ZN(n5702) );
  AND4_X1 U4940 ( .A1(n5589), .A2(n5762), .A3(n5764), .A4(n5716), .ZN(n4571)
         );
  NOR2_X1 U4941 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5034) );
  INV_X1 U4942 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5716) );
  INV_X1 U4943 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5684) );
  INV_X1 U4944 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5647) );
  NOR2_X2 U4945 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5638) );
  INV_X4 U4946 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U4947 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U4948 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6430) );
  INV_X1 U4949 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5149) );
  INV_X1 U4950 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5764) );
  INV_X1 U4951 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5762) );
  NOR2_X1 U4952 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5590) );
  NOR2_X1 U4953 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5591) );
  NOR2_X1 U4954 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5592) );
  NOR2_X1 U4955 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5593) );
  NOR2_X1 U4956 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n5589) );
  INV_X1 U4957 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5632) );
  AOI21_X2 U4958 ( .B1(n8294), .B2(n8297), .A(n5315), .ZN(n8281) );
  XNOR2_X1 U4959 ( .A(n5285), .B(n5284), .ZN(n6703) );
  OAI21_X1 U4960 ( .B1(n5642), .B2(n4461), .A(n4460), .ZN(n4950) );
  XNOR2_X1 U4961 ( .A(n4950), .B(SI_1_), .ZN(n5060) );
  CLKBUF_X1 U4962 ( .A(n9637), .Z(n4297) );
  CLKBUF_X1 U4963 ( .A(n7301), .Z(n4298) );
  INV_X1 U4964 ( .A(n6874), .ZN(n4300) );
  NAND2_X1 U4965 ( .A1(n4664), .A2(n4666), .ZN(n7301) );
  AND2_X2 U4966 ( .A1(n4571), .A2(n5702), .ZN(n5798) );
  INV_X1 U4967 ( .A(n6874), .ZN(n9769) );
  NAND2_X2 U4968 ( .A1(n4663), .A2(n4661), .ZN(n4660) );
  CLKBUF_X1 U4969 ( .A(n9373), .Z(n4301) );
  CLKBUF_X1 U4970 ( .A(n6991), .Z(n4302) );
  CLKBUF_X1 U4971 ( .A(n6852), .Z(n4303) );
  CLKBUF_X1 U4972 ( .A(n9385), .Z(n4304) );
  AND2_X1 U4974 ( .A1(n4684), .A2(n4685), .ZN(n5631) );
  AND2_X1 U4975 ( .A1(n7635), .A2(n9555), .ZN(n8616) );
  NAND2_X1 U4976 ( .A1(n7611), .A2(n9677), .ZN(n6281) );
  INV_X2 U4977 ( .A(n5797), .ZN(n8730) );
  OR2_X1 U4978 ( .A1(n6267), .A2(n5797), .ZN(n5789) );
  OAI21_X2 U4979 ( .B1(n9314), .B2(n4354), .A(n9156), .ZN(n9305) );
  OAI21_X2 U4980 ( .B1(n9330), .B2(n4390), .A(n9154), .ZN(n9314) );
  OAI21_X2 U4981 ( .B1(n9373), .B2(n4373), .A(n9148), .ZN(n9352) );
  OAI222_X1 U4982 ( .A1(P1_U3086), .A2(n9677), .B1(n9562), .B2(n9557), .C1(
        n9556), .C2(n9559), .ZN(P1_U3328) );
  NAND2_X1 U4983 ( .A1(n7684), .A2(n8237), .ZN(n4502) );
  XNOR2_X1 U4984 ( .A(n8415), .B(n7571), .ZN(n7572) );
  NOR2_X1 U4985 ( .A1(n7093), .A2(n5208), .ZN(n4766) );
  AOI21_X1 U4986 ( .B1(n4838), .B2(n4836), .A(n4369), .ZN(n4835) );
  INV_X1 U4987 ( .A(n4840), .ZN(n4836) );
  NAND2_X1 U4988 ( .A1(n5539), .A2(n7962), .ZN(n7903) );
  INV_X1 U4989 ( .A(n5343), .ZN(n6844) );
  INV_X1 U4990 ( .A(n5378), .ZN(n6840) );
  NAND2_X1 U4991 ( .A1(n6882), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U4992 ( .A1(n6900), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4699) );
  AND2_X1 U4993 ( .A1(n4768), .A2(n4767), .ZN(n7233) );
  INV_X1 U4994 ( .A(n7084), .ZN(n4767) );
  OR2_X1 U4995 ( .A1(n6692), .A2(n6691), .ZN(n4525) );
  MUX2_X1 U4996 ( .A(n8693), .B(n8692), .S(n8738), .Z(n8696) );
  OR2_X1 U4997 ( .A1(n5584), .A2(n7585), .ZN(n7898) );
  NAND2_X1 U4998 ( .A1(n5318), .A2(n5317), .ZN(n4733) );
  NAND2_X1 U4999 ( .A1(n5000), .A2(n4999), .ZN(n5003) );
  INV_X1 U5000 ( .A(SI_9_), .ZN(n4978) );
  NAND2_X1 U5001 ( .A1(n7684), .A2(n7569), .ZN(n4796) );
  INV_X1 U5002 ( .A(n4338), .ZN(n4804) );
  INV_X1 U5003 ( .A(n7715), .ZN(n4805) );
  NOR2_X1 U5004 ( .A1(n7663), .A2(n7577), .ZN(n7579) );
  NAND2_X1 U5005 ( .A1(n7744), .A2(n7902), .ZN(n7951) );
  OR2_X1 U5006 ( .A1(n7744), .A2(n7902), .ZN(n7952) );
  INV_X1 U5007 ( .A(n7897), .ZN(n7954) );
  AND2_X1 U5008 ( .A1(n7578), .A2(n8208), .ZN(n7884) );
  AND2_X1 U5009 ( .A1(n7889), .A2(n7888), .ZN(n7919) );
  NAND2_X1 U5010 ( .A1(n8412), .A2(n8218), .ZN(n4843) );
  INV_X1 U5011 ( .A(n8415), .ZN(n5497) );
  OR2_X1 U5012 ( .A1(n7575), .A2(n8218), .ZN(n7885) );
  OR2_X1 U5013 ( .A1(n7562), .A2(n8261), .ZN(n7869) );
  NAND2_X1 U5014 ( .A1(n5316), .A2(n4846), .ZN(n4849) );
  NOR2_X1 U5015 ( .A1(n8274), .A2(n4847), .ZN(n4846) );
  INV_X1 U5016 ( .A(n4850), .ZN(n4847) );
  OR2_X1 U5017 ( .A1(n7692), .A2(n8271), .ZN(n7863) );
  OR2_X1 U5018 ( .A1(n7644), .A2(n8283), .ZN(n7857) );
  OR2_X1 U5019 ( .A1(n7547), .A2(n8325), .ZN(n7846) );
  NOR2_X1 U5020 ( .A1(n5255), .A2(n4854), .ZN(n4853) );
  INV_X1 U5021 ( .A(n5242), .ZN(n4854) );
  AND2_X1 U5022 ( .A1(n5197), .A2(n4858), .ZN(n4560) );
  AND2_X1 U5023 ( .A1(n4916), .A2(n4560), .ZN(n5534) );
  INV_X1 U5024 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4909) );
  INV_X1 U5025 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n4740) );
  NOR2_X1 U5026 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n4741) );
  AND2_X1 U5027 ( .A1(n6243), .A2(n5630), .ZN(n5655) );
  NOR2_X1 U5028 ( .A1(n9207), .A2(n4617), .ZN(n4613) );
  INV_X1 U5029 ( .A(n9180), .ZN(n4608) );
  NAND2_X1 U5030 ( .A1(n9471), .A2(n8678), .ZN(n9179) );
  NAND2_X1 U5031 ( .A1(n4649), .A2(n9828), .ZN(n4648) );
  OAI21_X1 U5032 ( .B1(n7595), .B2(n9118), .A(n7594), .ZN(n7601) );
  OR2_X1 U5033 ( .A1(n7593), .A2(n7592), .ZN(n7594) );
  OR2_X1 U5034 ( .A1(n7601), .A2(n7600), .ZN(n7746) );
  XNOR2_X1 U5035 ( .A(n7593), .B(n7592), .ZN(n7595) );
  AND2_X1 U5036 ( .A1(n4871), .A2(n5798), .ZN(n5644) );
  NAND2_X1 U5037 ( .A1(n4726), .A2(n5008), .ZN(n4725) );
  INV_X1 U5038 ( .A(n5284), .ZN(n5008) );
  NAND2_X1 U5039 ( .A1(n5007), .A2(n5006), .ZN(n4726) );
  OAI21_X1 U5040 ( .B1(n4295), .B2(P2_REG1_REG_2__SCAN_IN), .A(n4505), .ZN(
        n4504) );
  NAND2_X1 U5041 ( .A1(n4295), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U5042 ( .A1(n6885), .A2(n6886), .ZN(n9941) );
  INV_X1 U5043 ( .A(n4698), .ZN(n6884) );
  NAND2_X1 U5044 ( .A1(n4512), .A2(n4513), .ZN(n4768) );
  NAND2_X1 U5045 ( .A1(n4427), .A2(n4426), .ZN(n4596) );
  INV_X1 U5046 ( .A(n7076), .ZN(n4426) );
  AND2_X1 U5047 ( .A1(n4509), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4506) );
  XNOR2_X1 U5048 ( .A(n7743), .B(n7954), .ZN(n5583) );
  NAND2_X1 U5049 ( .A1(n5573), .A2(n5572), .ZN(n7743) );
  NAND2_X1 U5050 ( .A1(n4833), .A2(n4832), .ZN(n8186) );
  AOI21_X1 U5051 ( .B1(n4835), .B2(n4837), .A(n4368), .ZN(n4832) );
  INV_X1 U5052 ( .A(n4756), .ZN(n4755) );
  OAI21_X1 U5053 ( .B1(n4759), .B2(n4327), .A(n7891), .ZN(n4756) );
  AND2_X1 U5054 ( .A1(n5455), .A2(n5454), .ZN(n8199) );
  NAND2_X1 U5055 ( .A1(n7575), .A2(n8218), .ZN(n7886) );
  OR2_X1 U5056 ( .A1(n5497), .A2(n8227), .ZN(n7880) );
  NAND2_X1 U5057 ( .A1(n7644), .A2(n7975), .ZN(n4848) );
  AND2_X1 U5058 ( .A1(n8299), .A2(n7977), .ZN(n5315) );
  AOI21_X1 U5059 ( .B1(n7536), .B2(n7535), .A(n5270), .ZN(n8322) );
  AOI21_X1 U5060 ( .B1(n7115), .B2(n7802), .A(n7806), .ZN(n7177) );
  NAND2_X1 U5061 ( .A1(n9989), .A2(n7793), .ZN(n4751) );
  AND2_X1 U5062 ( .A1(n7756), .A2(n5540), .ZN(n10013) );
  AND2_X1 U5063 ( .A1(n5506), .A2(n6504), .ZN(n10010) );
  OR2_X1 U5064 ( .A1(n7989), .A2(n6604), .ZN(n7763) );
  INV_X1 U5065 ( .A(n9984), .ZN(n10007) );
  NAND2_X1 U5066 ( .A1(n5446), .A2(n5445), .ZN(n5499) );
  INV_X1 U5067 ( .A(n5460), .ZN(n7752) );
  NOR2_X1 U5069 ( .A1(n4765), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5070 ( .A1(n4311), .A2(n5642), .ZN(n5704) );
  AND2_X1 U5071 ( .A1(n6208), .A2(n8786), .ZN(n6465) );
  OR2_X1 U5072 ( .A1(n9257), .A2(n9165), .ZN(n4456) );
  NAND2_X1 U5073 ( .A1(n9188), .A2(n9187), .ZN(n9237) );
  NOR2_X1 U5074 ( .A1(n9405), .A2(n9392), .ZN(n9391) );
  NOR2_X1 U5075 ( .A1(n4332), .A2(n4670), .ZN(n4669) );
  AND3_X1 U5076 ( .A1(n6243), .A2(P1_STATE_REG_SCAN_IN), .A3(n6279), .ZN(n8877) );
  NAND2_X1 U5077 ( .A1(n5617), .A2(n4891), .ZN(n5615) );
  INV_X1 U5078 ( .A(n4893), .ZN(n4891) );
  NAND2_X1 U5079 ( .A1(n5372), .A2(n5371), .ZN(n5386) );
  INV_X1 U5080 ( .A(n7969), .ZN(n8208) );
  OR2_X1 U5081 ( .A1(n8857), .A2(n8776), .ZN(n4437) );
  NAND2_X1 U5082 ( .A1(n4525), .A2(n4524), .ZN(n4523) );
  NAND2_X1 U5083 ( .A1(n6331), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4524) );
  MUX2_X1 U5084 ( .A(n7841), .B(n7840), .S(n7907), .Z(n7843) );
  NAND2_X1 U5085 ( .A1(n4422), .A2(n4419), .ZN(n7855) );
  NAND2_X1 U5086 ( .A1(n7851), .A2(n7907), .ZN(n4422) );
  OAI21_X1 U5087 ( .B1(n4421), .B2(n7842), .A(n4420), .ZN(n4419) );
  AND2_X1 U5088 ( .A1(n7876), .A2(n7878), .ZN(n4416) );
  NAND2_X1 U5089 ( .A1(n4423), .A2(n7866), .ZN(n7871) );
  AND2_X1 U5090 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  NAND2_X1 U5091 ( .A1(n8782), .A2(n8704), .ZN(n4442) );
  NAND2_X1 U5092 ( .A1(n8816), .A2(n8738), .ZN(n4443) );
  OR2_X1 U5093 ( .A1(n7205), .A2(n4814), .ZN(n4813) );
  INV_X1 U5094 ( .A(n7131), .ZN(n4814) );
  INV_X1 U5095 ( .A(n4813), .ZN(n4810) );
  NAND2_X1 U5096 ( .A1(n4491), .A2(n6967), .ZN(n4488) );
  INV_X1 U5097 ( .A(n6967), .ZN(n4489) );
  NAND2_X1 U5098 ( .A1(n4440), .A2(n8711), .ZN(n8716) );
  OR2_X1 U5099 ( .A1(n9212), .A2(n9170), .ZN(n8777) );
  NOR2_X1 U5100 ( .A1(n9257), .A2(n9275), .ZN(n4658) );
  INV_X1 U5101 ( .A(n5302), .ZN(n4722) );
  NAND2_X1 U5102 ( .A1(n5012), .A2(n5011), .ZN(n5015) );
  AND2_X1 U5103 ( .A1(n7014), .A2(n8154), .ZN(n6514) );
  AOI21_X1 U5104 ( .B1(n5500), .B2(n4347), .A(n4553), .ZN(n7755) );
  OR2_X1 U5105 ( .A1(n7906), .A2(n4554), .ZN(n4553) );
  AND2_X1 U5106 ( .A1(n7898), .A2(n4555), .ZN(n4554) );
  NAND2_X1 U5107 ( .A1(n5343), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5055) );
  OR2_X1 U5108 ( .A1(n6437), .A2(n6793), .ZN(n6451) );
  NAND2_X1 U5109 ( .A1(n6563), .A2(n6562), .ZN(n6564) );
  OAI21_X1 U5110 ( .B1(n9891), .B2(n4696), .A(n4695), .ZN(n6566) );
  NAND2_X1 U5111 ( .A1(n9908), .A2(n4334), .ZN(n4695) );
  NAND2_X1 U5112 ( .A1(n4334), .A2(n4697), .ZN(n4696) );
  OR2_X1 U5113 ( .A1(n6905), .A2(n6904), .ZN(n4773) );
  NOR2_X1 U5114 ( .A1(n8013), .A2(n4403), .ZN(n8014) );
  OR2_X1 U5115 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  NAND2_X1 U5116 ( .A1(n4771), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4770) );
  OR2_X1 U5117 ( .A1(n7578), .A2(n8208), .ZN(n7891) );
  AND2_X1 U5118 ( .A1(n8418), .A2(n7971), .ZN(n7921) );
  INV_X1 U5119 ( .A(n7856), .ZN(n4762) );
  NOR2_X1 U5120 ( .A1(n7185), .A2(n7984), .ZN(n4829) );
  INV_X1 U5121 ( .A(n7790), .ZN(n4745) );
  AND2_X1 U5122 ( .A1(n5519), .A2(n5518), .ZN(n6594) );
  AND2_X1 U5123 ( .A1(n9111), .A2(n4817), .ZN(n4816) );
  INV_X1 U5124 ( .A(n4880), .ZN(n4879) );
  OAI21_X1 U5125 ( .B1(n5836), .B2(n4881), .A(n5835), .ZN(n4880) );
  AND2_X1 U5126 ( .A1(n8512), .A2(n4888), .ZN(n4887) );
  NAND2_X1 U5127 ( .A1(n8557), .A2(n6057), .ZN(n4888) );
  INV_X1 U5128 ( .A(n6057), .ZN(n4885) );
  NOR2_X1 U5129 ( .A1(n4886), .A2(n4593), .ZN(n4592) );
  INV_X1 U5130 ( .A(n8503), .ZN(n4593) );
  INV_X1 U5131 ( .A(n4887), .ZN(n4886) );
  NAND2_X1 U5132 ( .A1(n4592), .A2(n8502), .ZN(n4590) );
  OAI21_X1 U5133 ( .B1(n9317), .B2(n4608), .A(n9181), .ZN(n4607) );
  NOR2_X1 U5134 ( .A1(n9356), .A2(n9377), .ZN(n4651) );
  NAND2_X1 U5135 ( .A1(n4467), .A2(n5963), .ZN(n9411) );
  NOR2_X1 U5136 ( .A1(n7400), .A2(n8476), .ZN(n4653) );
  INV_X1 U5137 ( .A(n7371), .ZN(n8762) );
  AND2_X1 U5138 ( .A1(n4635), .A2(n8658), .ZN(n4634) );
  AND2_X1 U5139 ( .A1(n7025), .A2(n9730), .ZN(n4680) );
  NAND2_X1 U5140 ( .A1(n9722), .A2(n8623), .ZN(n7053) );
  INV_X1 U5141 ( .A(n6998), .ZN(n4623) );
  AND2_X1 U5142 ( .A1(n4351), .A2(n6802), .ZN(n4626) );
  INV_X1 U5143 ( .A(n6271), .ZN(n6201) );
  NOR2_X1 U5144 ( .A1(n9192), .A2(n4618), .ZN(n4617) );
  INV_X1 U5145 ( .A(n9189), .ZN(n4618) );
  AOI22_X1 U5146 ( .A1(n4616), .A2(n9191), .B1(n4617), .B2(n9190), .ZN(n4615)
         );
  INV_X1 U5147 ( .A(n9221), .ZN(n4616) );
  NOR2_X1 U5148 ( .A1(n7306), .A2(n7510), .ZN(n7397) );
  NOR2_X1 U5149 ( .A1(n7339), .A2(n7031), .ZN(n4649) );
  OR2_X1 U5150 ( .A1(n8738), .A2(n8853), .ZN(n9767) );
  NAND2_X1 U5151 ( .A1(n5423), .A2(n5422), .ZN(n5438) );
  AOI21_X1 U5152 ( .B1(n4708), .B2(n4711), .A(n4706), .ZN(n4705) );
  AND2_X1 U5153 ( .A1(n5403), .A2(n5390), .ZN(n5391) );
  AOI21_X1 U5154 ( .B1(n4732), .B2(n4730), .A(n4729), .ZN(n4728) );
  INV_X1 U5155 ( .A(n5336), .ZN(n4729) );
  INV_X1 U5156 ( .A(n5317), .ZN(n4730) );
  NAND2_X1 U5157 ( .A1(n4412), .A2(n4732), .ZN(n4727) );
  AND2_X1 U5158 ( .A1(n5336), .A2(n5323), .ZN(n5334) );
  INV_X1 U5159 ( .A(n4724), .ZN(n4723) );
  OAI21_X1 U5160 ( .B1(n4725), .B2(n5006), .A(n5010), .ZN(n4724) );
  INV_X1 U5161 ( .A(n5271), .ZN(n5007) );
  XNOR2_X1 U5162 ( .A(n5004), .B(SI_15_), .ZN(n5271) );
  NAND2_X1 U5163 ( .A1(n4734), .A2(n4998), .ZN(n5256) );
  INV_X1 U5164 ( .A(n5243), .ZN(n4996) );
  NAND2_X1 U5165 ( .A1(n5003), .A2(n5002), .ZN(n5257) );
  XNOR2_X1 U5166 ( .A(n4997), .B(SI_13_), .ZN(n5243) );
  XNOR2_X1 U5167 ( .A(n4993), .B(SI_12_), .ZN(n5229) );
  NAND2_X1 U5168 ( .A1(n4985), .A2(SI_10_), .ZN(n4986) );
  INV_X1 U5169 ( .A(n5203), .ZN(n4983) );
  NAND2_X1 U5170 ( .A1(n4977), .A2(n4976), .ZN(n5184) );
  AND2_X1 U5171 ( .A1(n4477), .A2(n4319), .ZN(n4474) );
  NAND2_X1 U5172 ( .A1(n4312), .A2(n4329), .ZN(n4477) );
  OR2_X1 U5173 ( .A1(n7579), .A2(n7581), .ZN(n7582) );
  NAND2_X1 U5174 ( .A1(n4795), .A2(n7569), .ZN(n4503) );
  INV_X1 U5175 ( .A(n4502), .ZN(n4795) );
  INV_X1 U5176 ( .A(n7660), .ZN(n4500) );
  INV_X1 U5177 ( .A(n7661), .ZN(n4499) );
  AOI21_X1 U5178 ( .B1(n4807), .B2(n7487), .A(n4370), .ZN(n4487) );
  AND2_X1 U5179 ( .A1(n7660), .A2(n7574), .ZN(n7684) );
  NOR2_X1 U5180 ( .A1(n6713), .A2(n4819), .ZN(n4818) );
  INV_X1 U5181 ( .A(n6709), .ZN(n4819) );
  NAND2_X1 U5182 ( .A1(n4936), .A2(n4935), .ZN(n5328) );
  INV_X1 U5183 ( .A(n5049), .ZN(n4936) );
  NAND2_X1 U5184 ( .A1(n4480), .A2(n4478), .ZN(n7652) );
  AOI21_X1 U5185 ( .B1(n4482), .B2(n4801), .A(n4479), .ZN(n4478) );
  INV_X1 U5186 ( .A(n7651), .ZN(n4479) );
  OR2_X1 U5187 ( .A1(n5359), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U5188 ( .A1(n7484), .A2(n7483), .ZN(n7524) );
  NOR3_X1 U5189 ( .A1(n7949), .A2(n7950), .A3(n4452), .ZN(n7953) );
  INV_X1 U5190 ( .A(n7951), .ZN(n4452) );
  NAND2_X1 U5191 ( .A1(n7917), .A2(n7918), .ZN(n4738) );
  INV_X1 U5192 ( .A(n7916), .ZN(n4739) );
  OR2_X1 U5193 ( .A1(n7905), .A2(n7904), .ZN(n7914) );
  INV_X1 U5194 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4910) );
  OR2_X1 U5195 ( .A1(n5076), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5095) );
  OR2_X1 U5196 ( .A1(n5028), .A2(n8452), .ZN(n5030) );
  NAND2_X1 U5197 ( .A1(n6456), .A2(n4504), .ZN(n6570) );
  XNOR2_X1 U5198 ( .A(n6564), .B(n9888), .ZN(n9892) );
  OR2_X1 U5199 ( .A1(n9889), .A2(n6575), .ZN(n4520) );
  NAND2_X1 U5200 ( .A1(n4520), .A2(n4519), .ZN(n6578) );
  INV_X1 U5201 ( .A(n9906), .ZN(n4519) );
  XNOR2_X1 U5202 ( .A(n6577), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n9908) );
  AND2_X1 U5203 ( .A1(n4596), .A2(n4595), .ZN(n7260) );
  NAND2_X1 U5204 ( .A1(n7234), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4595) );
  OR2_X1 U5205 ( .A1(n7233), .A2(n4400), .ZN(n4508) );
  NOR2_X1 U5206 ( .A1(n7265), .A2(n7264), .ZN(n8025) );
  NAND2_X1 U5207 ( .A1(n8014), .A2(n8019), .ZN(n4771) );
  OR2_X1 U5208 ( .A1(n8014), .A2(n8019), .ZN(n4772) );
  INV_X1 U5209 ( .A(n4770), .ZN(n4769) );
  AND3_X1 U5210 ( .A1(n4690), .A2(P2_REG2_REG_13__SCAN_IN), .A3(n8034), .ZN(
        n8035) );
  OR2_X1 U5211 ( .A1(n8091), .A2(n8383), .ZN(n4788) );
  NAND2_X1 U5212 ( .A1(n4693), .A2(n4692), .ZN(n8138) );
  INV_X1 U5213 ( .A(n8112), .ZN(n4692) );
  INV_X1 U5214 ( .A(n7886), .ZN(n4757) );
  INV_X1 U5215 ( .A(n7919), .ZN(n8190) );
  OR2_X1 U5216 ( .A1(n4841), .A2(n4839), .ZN(n4838) );
  INV_X1 U5217 ( .A(n4843), .ZN(n4839) );
  AND2_X1 U5218 ( .A1(n4842), .A2(n8209), .ZN(n4841) );
  NAND2_X1 U5219 ( .A1(n4336), .A2(n4844), .ZN(n4842) );
  INV_X1 U5220 ( .A(n8200), .ZN(n8196) );
  AND2_X1 U5221 ( .A1(n4843), .A2(n4844), .ZN(n4840) );
  NOR2_X1 U5222 ( .A1(n5498), .A2(n4296), .ZN(n4759) );
  AND2_X1 U5223 ( .A1(n7890), .A2(n7891), .ZN(n8200) );
  OR2_X1 U5224 ( .A1(n5497), .A2(n7970), .ZN(n4844) );
  OAI21_X1 U5225 ( .B1(n8238), .B2(n4748), .A(n4746), .ZN(n8222) );
  AOI21_X1 U5226 ( .B1(n4749), .B2(n4747), .A(n7920), .ZN(n4746) );
  INV_X1 U5227 ( .A(n4749), .ZN(n4748) );
  INV_X1 U5228 ( .A(n7874), .ZN(n4747) );
  OR2_X1 U5229 ( .A1(n5376), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5396) );
  AND2_X1 U5230 ( .A1(n5402), .A2(n5401), .ZN(n8227) );
  OR2_X1 U5231 ( .A1(n7921), .A2(n7920), .ZN(n8228) );
  AND3_X1 U5232 ( .A1(n5346), .A2(n5345), .A3(n5344), .ZN(n8261) );
  NAND2_X1 U5233 ( .A1(n4849), .A2(n4348), .ZN(n8257) );
  OAI21_X1 U5234 ( .B1(n8296), .B2(n8438), .A(n8281), .ZN(n5316) );
  NAND2_X1 U5235 ( .A1(n8438), .A2(n8296), .ZN(n4850) );
  OR2_X1 U5236 ( .A1(n7722), .A2(n8296), .ZN(n7856) );
  AND2_X1 U5237 ( .A1(n7857), .A2(n7859), .ZN(n8274) );
  OR2_X1 U5238 ( .A1(n5310), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5239 ( .A1(n4541), .A2(n7847), .ZN(n5493) );
  INV_X1 U5240 ( .A(n8298), .ZN(n4541) );
  NAND2_X1 U5241 ( .A1(n5493), .A2(n4315), .ZN(n8284) );
  OR2_X1 U5242 ( .A1(n5292), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5308) );
  AND2_X1 U5243 ( .A1(n7846), .A2(n7849), .ZN(n8314) );
  OAI21_X1 U5244 ( .B1(n8328), .B2(n7840), .A(n7839), .ZN(n8313) );
  NAND2_X1 U5245 ( .A1(n8322), .A2(n8321), .ZN(n8320) );
  OR2_X1 U5246 ( .A1(n5264), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5277) );
  AND2_X1 U5247 ( .A1(n4548), .A2(n7832), .ZN(n4547) );
  NAND2_X1 U5248 ( .A1(n4549), .A2(n7831), .ZN(n4548) );
  INV_X1 U5249 ( .A(n7828), .ZN(n4549) );
  INV_X1 U5250 ( .A(n7831), .ZN(n4550) );
  AND4_X1 U5251 ( .A1(n5282), .A2(n5281), .A3(n5280), .A4(n5279), .ZN(n8308)
         );
  NAND2_X1 U5252 ( .A1(n4852), .A2(n4851), .ZN(n7536) );
  AOI21_X1 U5253 ( .B1(n4853), .B2(n5241), .A(n4359), .ZN(n4851) );
  NAND2_X1 U5254 ( .A1(n4929), .A2(n7273), .ZN(n5248) );
  INV_X1 U5255 ( .A(n5235), .ZN(n4929) );
  AND2_X1 U5256 ( .A1(n7832), .A2(n7831), .ZN(n7923) );
  NAND2_X1 U5257 ( .A1(n4537), .A2(n4535), .ZN(n7455) );
  AOI21_X1 U5258 ( .B1(n4339), .B2(n4540), .A(n4536), .ZN(n4535) );
  INV_X1 U5259 ( .A(n7822), .ZN(n4536) );
  INV_X1 U5260 ( .A(n7983), .ZN(n7431) );
  NAND2_X1 U5261 ( .A1(n4831), .A2(n4330), .ZN(n4830) );
  INV_X1 U5262 ( .A(n7178), .ZN(n4831) );
  INV_X1 U5263 ( .A(n4829), .ZN(n4827) );
  OR2_X1 U5264 ( .A1(n5174), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5189) );
  INV_X1 U5265 ( .A(n7984), .ZN(n7316) );
  NAND2_X1 U5266 ( .A1(n4751), .A2(n4349), .ZN(n7115) );
  NAND2_X1 U5267 ( .A1(n4551), .A2(n5490), .ZN(n9989) );
  INV_X1 U5268 ( .A(n6981), .ZN(n4551) );
  NOR2_X1 U5269 ( .A1(n5123), .A2(n10030), .ZN(n4857) );
  NAND2_X1 U5270 ( .A1(n6725), .A2(n4924), .ZN(n5125) );
  INV_X1 U5271 ( .A(n6284), .ZN(n6503) );
  AOI21_X1 U5272 ( .B1(n5583), .B2(n10010), .A(n5580), .ZN(n5581) );
  OR2_X1 U5273 ( .A1(n5582), .A2(n10013), .ZN(n4823) );
  NAND2_X1 U5274 ( .A1(n5410), .A2(n5409), .ZN(n7575) );
  NAND2_X1 U5275 ( .A1(n5358), .A2(n5357), .ZN(n7703) );
  NAND2_X1 U5276 ( .A1(n5338), .A2(n5337), .ZN(n7562) );
  NAND2_X1 U5277 ( .A1(n5039), .A2(n5038), .ZN(n7644) );
  NAND2_X1 U5278 ( .A1(n5291), .A2(n5290), .ZN(n7547) );
  OR2_X1 U5279 ( .A1(n5533), .A2(n7418), .ZN(n6496) );
  NAND2_X1 U5280 ( .A1(n5534), .A2(n5536), .ZN(n5508) );
  NAND2_X1 U5281 ( .A1(n6286), .A2(n5516), .ZN(n6283) );
  AND2_X1 U5282 ( .A1(n5534), .A2(n4764), .ZN(n5025) );
  NOR2_X1 U5283 ( .A1(n4765), .A2(n4371), .ZN(n4764) );
  INV_X1 U5284 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5509) );
  INV_X1 U5285 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9109) );
  NAND2_X1 U5286 ( .A1(n5475), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  OAI21_X1 U5287 ( .B1(n5471), .B2(P2_IR_REG_19__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5474) );
  INV_X1 U5288 ( .A(n5218), .ZN(n5031) );
  INV_X1 U5289 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5165) );
  OR2_X1 U5290 ( .A1(n5164), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5181) );
  NAND2_X1 U5291 ( .A1(n4908), .A2(n4820), .ZN(n5117) );
  NOR2_X1 U5292 ( .A1(n5117), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5133) );
  OR2_X1 U5293 ( .A1(n6430), .A2(n8452), .ZN(n5087) );
  INV_X1 U5294 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4945) );
  INV_X1 U5295 ( .A(n8470), .ZN(n4865) );
  INV_X1 U5296 ( .A(n4576), .ZN(n7356) );
  AOI21_X1 U5297 ( .B1(n6771), .B2(n7620), .A(n5670), .ZN(n5675) );
  NAND2_X1 U5298 ( .A1(n6125), .A2(n8519), .ZN(n4876) );
  AND2_X1 U5299 ( .A1(n8547), .A2(n8519), .ZN(n4877) );
  INV_X1 U5300 ( .A(n8530), .ZN(n4568) );
  NAND2_X1 U5301 ( .A1(n8546), .A2(n8547), .ZN(n8545) );
  XNOR2_X1 U5302 ( .A(n6096), .B(n6173), .ZN(n8484) );
  NAND2_X1 U5303 ( .A1(n4570), .A2(n4906), .ZN(n8595) );
  INV_X1 U5304 ( .A(n7017), .ZN(n8853) );
  NOR2_X1 U5305 ( .A1(n7142), .A2(n4533), .ZN(n8920) );
  AND2_X1 U5306 ( .A1(n7143), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U5307 ( .A1(n8956), .A2(n4527), .ZN(n8962) );
  OR2_X1 U5308 ( .A1(n8957), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4527) );
  AND2_X1 U5309 ( .A1(n9178), .A2(n9214), .ZN(n9173) );
  NAND2_X1 U5310 ( .A1(n9289), .A2(n4654), .ZN(n9226) );
  NOR2_X1 U5311 ( .A1(n4655), .A2(n9228), .ZN(n4654) );
  INV_X1 U5312 ( .A(n4656), .ZN(n4655) );
  NOR2_X1 U5313 ( .A1(n9226), .A2(n9212), .ZN(n9214) );
  AND2_X1 U5314 ( .A1(n9306), .A2(n9522), .ZN(n9289) );
  NAND2_X1 U5315 ( .A1(n8684), .A2(n8844), .ZN(n9180) );
  NOR2_X1 U5316 ( .A1(n9321), .A2(n9307), .ZN(n9306) );
  NAND2_X1 U5317 ( .A1(n9339), .A2(n9179), .ZN(n9316) );
  AND2_X1 U5318 ( .A1(n8844), .A2(n8742), .ZN(n9317) );
  NAND2_X1 U5319 ( .A1(n9316), .A2(n9317), .ZN(n9315) );
  NAND2_X1 U5320 ( .A1(n4642), .A2(n4640), .ZN(n9340) );
  AOI21_X1 U5321 ( .B1(n4340), .B2(n8840), .A(n4641), .ZN(n4640) );
  INV_X1 U5322 ( .A(n8843), .ZN(n4641) );
  AND2_X1 U5323 ( .A1(n4643), .A2(n8842), .ZN(n9347) );
  OR2_X1 U5324 ( .A1(n9387), .A2(n8840), .ZN(n4643) );
  OR2_X1 U5325 ( .A1(n9139), .A2(n8885), .ZN(n4676) );
  AND2_X1 U5326 ( .A1(n9139), .A2(n8885), .ZN(n4677) );
  CLKBUF_X1 U5327 ( .A(n9411), .Z(n4457) );
  INV_X1 U5328 ( .A(n4674), .ZN(n9414) );
  NAND2_X1 U5329 ( .A1(n7374), .A2(n7373), .ZN(n7401) );
  NAND2_X1 U5330 ( .A1(n9701), .A2(n7055), .ZN(n7025) );
  NAND2_X1 U5331 ( .A1(n4351), .A2(n4625), .ZN(n4624) );
  INV_X1 U5332 ( .A(n8790), .ZN(n4625) );
  NAND2_X1 U5333 ( .A1(n6803), .A2(n4626), .ZN(n4622) );
  NAND2_X1 U5334 ( .A1(n4432), .A2(n4409), .ZN(n8735) );
  NAND2_X1 U5335 ( .A1(n8731), .A2(n8730), .ZN(n4432) );
  NAND2_X1 U5336 ( .A1(n5984), .A2(n5983), .ZN(n9392) );
  AND2_X1 U5337 ( .A1(n7004), .A2(n9767), .ZN(n9632) );
  NAND2_X1 U5338 ( .A1(n7746), .A2(n7602), .ZN(n8607) );
  AND2_X1 U5339 ( .A1(n5598), .A2(n5632), .ZN(n4683) );
  NAND2_X1 U5340 ( .A1(n5438), .A2(n5437), .ZN(n5440) );
  NAND2_X1 U5341 ( .A1(n5617), .A2(n4892), .ZN(n5634) );
  AND2_X1 U5342 ( .A1(n5385), .A2(n5370), .ZN(n5371) );
  AOI21_X1 U5343 ( .B1(n4586), .B2(P1_IR_REG_31__SCAN_IN), .A(
        P1_IR_REG_22__SCAN_IN), .ZN(n4585) );
  XNOR2_X1 U5344 ( .A(n5366), .B(n5365), .ZN(n7188) );
  AND2_X1 U5345 ( .A1(n5644), .A2(n5622), .ZN(n5626) );
  XNOR2_X1 U5346 ( .A(n5256), .B(n5257), .ZN(n6619) );
  NAND2_X1 U5347 ( .A1(n5375), .A2(n5374), .ZN(n7641) );
  INV_X1 U5348 ( .A(n5092), .ZN(n6641) );
  AND3_X1 U5349 ( .A1(n5332), .A2(n5331), .A3(n5330), .ZN(n8271) );
  AND4_X1 U5350 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n8309)
         );
  NAND2_X1 U5351 ( .A1(n5307), .A2(n5306), .ZN(n8299) );
  AND4_X1 U5352 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), .ZN(n8283)
         );
  INV_X1 U5353 ( .A(n7988), .ZN(n10008) );
  AND4_X1 U5354 ( .A1(n5269), .A2(n5268), .A3(n5267), .A4(n5266), .ZN(n8326)
         );
  NAND2_X1 U5355 ( .A1(n5436), .A2(n5435), .ZN(n7969) );
  AND2_X1 U5356 ( .A1(n5419), .A2(n5418), .ZN(n8218) );
  INV_X1 U5357 ( .A(n8227), .ZN(n7970) );
  INV_X1 U5358 ( .A(n8283), .ZN(n7975) );
  NAND2_X1 U5359 ( .A1(n5071), .A2(n5070), .ZN(n7989) );
  AND2_X1 U5360 ( .A1(n5343), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5068) );
  INV_X1 U5361 ( .A(n6577), .ZN(n9915) );
  NAND2_X1 U5362 ( .A1(n4599), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4600) );
  INV_X1 U5363 ( .A(n9941), .ZN(n4599) );
  OR2_X1 U5364 ( .A1(n6887), .A2(n6890), .ZN(n4598) );
  OR2_X1 U5365 ( .A1(n7990), .A2(n7075), .ZN(n4427) );
  INV_X1 U5366 ( .A(n4768), .ZN(n7085) );
  INV_X1 U5367 ( .A(n4596), .ZN(n7231) );
  NAND2_X1 U5368 ( .A1(n4597), .A2(n4337), .ZN(n4688) );
  INV_X1 U5369 ( .A(n8080), .ZN(n4516) );
  AND2_X1 U5370 ( .A1(n4688), .A2(n4687), .ZN(n8087) );
  INV_X1 U5371 ( .A(n8066), .ZN(n4687) );
  NAND2_X1 U5372 ( .A1(n4789), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U5373 ( .A1(n8131), .A2(n4789), .ZN(n4785) );
  INV_X1 U5374 ( .A(n8132), .ZN(n4789) );
  AND2_X1 U5375 ( .A1(n9885), .A2(n9882), .ZN(n9951) );
  NAND2_X1 U5376 ( .A1(n8138), .A2(n8137), .ZN(n4691) );
  NAND2_X1 U5377 ( .A1(n5500), .A2(n7889), .ZN(n5501) );
  AOI21_X1 U5378 ( .B1(n5485), .B2(n9987), .A(n5484), .ZN(n8185) );
  AND2_X1 U5379 ( .A1(n4861), .A2(n4858), .ZN(n4558) );
  AND2_X1 U5380 ( .A1(n4345), .A2(n4922), .ZN(n4861) );
  NOR2_X1 U5381 ( .A1(n7421), .A2(n7370), .ZN(n5621) );
  NAND2_X1 U5382 ( .A1(n6076), .A2(n6075), .ZN(n9291) );
  NAND2_X1 U5383 ( .A1(n4429), .A2(n4428), .ZN(n8862) );
  NAND2_X1 U5384 ( .A1(n4431), .A2(n8834), .ZN(n4428) );
  OR2_X1 U5385 ( .A1(n4431), .A2(n4430), .ZN(n4429) );
  OAI21_X1 U5386 ( .B1(n8833), .B2(n8832), .A(n8831), .ZN(n4431) );
  INV_X1 U5387 ( .A(n6390), .ZN(n4522) );
  AOI21_X1 U5388 ( .B1(n4444), .B2(n9738), .A(n4453), .ZN(n9426) );
  INV_X1 U5389 ( .A(n9201), .ZN(n4453) );
  XNOR2_X1 U5390 ( .A(n9194), .B(n4447), .ZN(n4444) );
  NAND2_X1 U5391 ( .A1(n4663), .A2(n9168), .ZN(n9220) );
  OAI21_X1 U5392 ( .B1(n9237), .B2(n9190), .A(n9189), .ZN(n9222) );
  OR2_X1 U5393 ( .A1(n9758), .A2(n8980), .ZN(n9413) );
  INV_X1 U5394 ( .A(n9489), .ZN(n4435) );
  MUX2_X1 U5395 ( .A(n7764), .B(n7763), .S(n7762), .Z(n7770) );
  NOR2_X1 U5396 ( .A1(n7843), .A2(n7842), .ZN(n7844) );
  INV_X1 U5397 ( .A(n7850), .ZN(n4421) );
  NOR2_X1 U5398 ( .A1(n7848), .A2(n7907), .ZN(n4420) );
  NAND2_X1 U5399 ( .A1(n4425), .A2(n4424), .ZN(n4423) );
  AOI21_X1 U5400 ( .B1(n7862), .B2(n7903), .A(n7867), .ZN(n4424) );
  NAND2_X1 U5401 ( .A1(n7861), .A2(n7907), .ZN(n4425) );
  AND2_X1 U5402 ( .A1(n4416), .A2(n8221), .ZN(n4415) );
  INV_X1 U5403 ( .A(n8701), .ZN(n4438) );
  AND2_X1 U5404 ( .A1(n8699), .A2(n8698), .ZN(n4439) );
  OAI21_X1 U5405 ( .B1(n8696), .B2(n9299), .A(n4441), .ZN(n8700) );
  AOI21_X1 U5406 ( .B1(n4715), .B2(n4718), .A(n4713), .ZN(n4712) );
  INV_X1 U5407 ( .A(n5562), .ZN(n4713) );
  INV_X1 U5408 ( .A(n5572), .ZN(n4555) );
  INV_X1 U5409 ( .A(n4897), .ZN(n4697) );
  OR2_X1 U5410 ( .A1(n9651), .A2(n4882), .ZN(n4881) );
  INV_X1 U5411 ( .A(n5796), .ZN(n4882) );
  INV_X1 U5412 ( .A(n5836), .ZN(n4883) );
  INV_X1 U5413 ( .A(n5420), .ZN(n4706) );
  NAND2_X1 U5414 ( .A1(n4988), .A2(n4987), .ZN(n4991) );
  NAND2_X1 U5415 ( .A1(n4974), .A2(n4973), .ZN(n4977) );
  AOI21_X1 U5416 ( .B1(n4800), .B2(n4803), .A(n4483), .ZN(n4482) );
  INV_X1 U5417 ( .A(n4812), .ZN(n4811) );
  OAI211_X1 U5418 ( .C1(n4492), .C2(n4489), .A(n4810), .B(n4488), .ZN(n4809)
         );
  OAI21_X1 U5419 ( .B1(n4813), .B2(n6970), .A(n7204), .ZN(n4812) );
  NAND2_X1 U5420 ( .A1(n7954), .A2(n4418), .ZN(n4417) );
  INV_X1 U5421 ( .A(n7899), .ZN(n4418) );
  OR2_X1 U5422 ( .A1(n4780), .A2(n10080), .ZN(n4778) );
  NAND2_X1 U5423 ( .A1(n4773), .A2(n7081), .ZN(n7083) );
  NAND2_X1 U5424 ( .A1(n7083), .A2(n7082), .ZN(n4513) );
  NOR2_X1 U5425 ( .A1(n7950), .A2(n4557), .ZN(n4556) );
  INV_X1 U5426 ( .A(n7889), .ZN(n4557) );
  INV_X1 U5427 ( .A(n4838), .ZN(n4837) );
  NOR2_X1 U5428 ( .A1(n7921), .A2(n7873), .ZN(n4749) );
  AND2_X1 U5429 ( .A1(n7872), .A2(n7874), .ZN(n7922) );
  OR2_X1 U5430 ( .A1(n7525), .A2(n8308), .ZN(n7839) );
  OR2_X1 U5431 ( .A1(n7813), .A2(n4540), .ZN(n4539) );
  INV_X1 U5432 ( .A(n7816), .ZN(n4540) );
  NAND2_X1 U5433 ( .A1(n7898), .A2(n7742), .ZN(n7897) );
  INV_X1 U5434 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5026) );
  INV_X1 U5435 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4946) );
  NOR2_X1 U5436 ( .A1(n5964), .A2(n8927), .ZN(n5986) );
  NOR2_X1 U5437 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  INV_X1 U5438 ( .A(n7357), .ZN(n4581) );
  INV_X1 U5439 ( .A(n7438), .ZN(n4580) );
  AND2_X1 U5440 ( .A1(n5986), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6005) );
  INV_X1 U5441 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4907) );
  AND2_X1 U5442 ( .A1(n4658), .A2(n4657), .ZN(n4656) );
  OR2_X1 U5443 ( .A1(n9228), .A2(n8706), .ZN(n8779) );
  OR2_X1 U5444 ( .A1(n9291), .A2(n8695), .ZN(n8741) );
  INV_X1 U5445 ( .A(n7376), .ZN(n4670) );
  NAND2_X1 U5446 ( .A1(n6773), .A2(n6874), .ZN(n6753) );
  NAND2_X1 U5447 ( .A1(n9289), .A2(n4658), .ZN(n9255) );
  NAND2_X1 U5448 ( .A1(n9289), .A2(n9518), .ZN(n9272) );
  NAND2_X1 U5449 ( .A1(n9749), .A2(n9783), .ZN(n6809) );
  AND2_X1 U5450 ( .A1(n5439), .A2(n5427), .ZN(n5437) );
  NAND2_X1 U5451 ( .A1(n5599), .A2(n4894), .ZN(n4893) );
  INV_X1 U5452 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4894) );
  INV_X1 U5453 ( .A(n5391), .ZN(n4711) );
  AOI21_X1 U5454 ( .B1(n5391), .B2(n4710), .A(n4709), .ZN(n4708) );
  INV_X1 U5455 ( .A(n5403), .ZN(n4709) );
  INV_X1 U5456 ( .A(n5385), .ZN(n4710) );
  AOI21_X1 U5457 ( .B1(n5272), .B2(n4395), .A(n4720), .ZN(n4719) );
  NAND2_X1 U5458 ( .A1(n4721), .A2(n5015), .ZN(n4720) );
  NAND2_X1 U5459 ( .A1(n4723), .A2(n4397), .ZN(n4721) );
  OR2_X1 U5460 ( .A1(n5899), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U5461 ( .A(n4984), .B(SI_10_), .ZN(n5203) );
  AND2_X1 U5462 ( .A1(n4982), .A2(n4981), .ZN(n5195) );
  NAND2_X1 U5463 ( .A1(n4926), .A2(n6973), .ZN(n5174) );
  INV_X1 U5464 ( .A(n5158), .ZN(n4926) );
  INV_X1 U5465 ( .A(n6969), .ZN(n4815) );
  NAND2_X1 U5466 ( .A1(n4496), .A2(n4503), .ZN(n4497) );
  NAND2_X1 U5467 ( .A1(n7132), .A2(n7131), .ZN(n7206) );
  INV_X1 U5468 ( .A(n5341), .ZN(n5340) );
  XNOR2_X1 U5469 ( .A(n7571), .B(n6794), .ZN(n6526) );
  NAND2_X1 U5470 ( .A1(n4806), .A2(n4805), .ZN(n4802) );
  NAND2_X1 U5471 ( .A1(n6832), .A2(n4318), .ZN(n4491) );
  OR2_X1 U5472 ( .A1(n5430), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5449) );
  OAI21_X1 U5473 ( .B1(n6435), .B2(n6434), .A(n6450), .ZN(n6437) );
  NAND2_X1 U5474 ( .A1(n6447), .A2(n4790), .ZN(n6431) );
  NAND2_X1 U5475 ( .A1(n4791), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4790) );
  AND2_X1 U5476 ( .A1(n6566), .A2(n6565), .ZN(n4601) );
  NAND2_X1 U5477 ( .A1(n6578), .A2(n4780), .ZN(n4782) );
  NAND2_X1 U5478 ( .A1(n6578), .A2(n4783), .ZN(n4775) );
  OAI21_X1 U5479 ( .B1(n6578), .B2(n4779), .A(n4776), .ZN(n6580) );
  NOR2_X1 U5480 ( .A1(n9928), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4779) );
  AND2_X1 U5481 ( .A1(n4778), .A2(n4777), .ZN(n4776) );
  NAND2_X1 U5482 ( .A1(n9928), .A2(n4784), .ZN(n4777) );
  OR2_X1 U5483 ( .A1(n8001), .A2(n10085), .ZN(n4512) );
  OAI21_X1 U5484 ( .B1(n7083), .B2(n7082), .A(n4513), .ZN(n8001) );
  NAND2_X1 U5485 ( .A1(n4766), .A2(n4511), .ZN(n4509) );
  AND2_X1 U5486 ( .A1(n4510), .A2(n4341), .ZN(n7272) );
  NOR2_X1 U5487 ( .A1(n7261), .A2(n7262), .ZN(n7265) );
  OAI21_X1 U5488 ( .B1(n8042), .B2(n4515), .A(n4514), .ZN(n8089) );
  NAND2_X1 U5489 ( .A1(n4518), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n4515) );
  NAND2_X1 U5490 ( .A1(n8080), .A2(n4518), .ZN(n4514) );
  INV_X1 U5491 ( .A(n8081), .ZN(n4518) );
  OR2_X1 U5492 ( .A1(n8042), .A2(n8392), .ZN(n4517) );
  AND2_X1 U5493 ( .A1(n8090), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4686) );
  OR2_X1 U5494 ( .A1(n5463), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8164) );
  AOI21_X1 U5495 ( .B1(n4755), .B2(n4327), .A(n4754), .ZN(n4753) );
  NAND2_X1 U5496 ( .A1(n4313), .A2(n4755), .ZN(n4752) );
  INV_X1 U5497 ( .A(n7888), .ZN(n4754) );
  OR2_X1 U5498 ( .A1(n8199), .A2(n5499), .ZN(n7889) );
  INV_X1 U5499 ( .A(n7967), .ZN(n8188) );
  AND2_X1 U5500 ( .A1(n5496), .A2(n7880), .ZN(n8221) );
  NAND2_X1 U5501 ( .A1(n5395), .A2(n5394), .ZN(n5413) );
  INV_X1 U5502 ( .A(n5396), .ZN(n5395) );
  NAND2_X1 U5503 ( .A1(n7869), .A2(n7868), .ZN(n8251) );
  OAI21_X1 U5504 ( .B1(n5493), .B2(n4333), .A(n4760), .ZN(n8262) );
  INV_X1 U5505 ( .A(n4761), .ZN(n4760) );
  OAI21_X1 U5506 ( .B1(n4315), .B2(n4333), .A(n7859), .ZN(n4761) );
  INV_X1 U5507 ( .A(n5308), .ZN(n4934) );
  NAND2_X1 U5508 ( .A1(n8311), .A2(n5300), .ZN(n8294) );
  OAI21_X1 U5509 ( .B1(n4542), .B2(n7842), .A(n7846), .ZN(n8298) );
  INV_X1 U5510 ( .A(n8313), .ZN(n4542) );
  INV_X1 U5511 ( .A(n8314), .ZN(n5298) );
  NAND2_X1 U5512 ( .A1(n4933), .A2(n4932), .ZN(n5292) );
  NAND2_X1 U5513 ( .A1(n4545), .A2(n4543), .ZN(n8328) );
  AOI21_X1 U5514 ( .B1(n4320), .B2(n4550), .A(n4544), .ZN(n4543) );
  INV_X1 U5515 ( .A(n7835), .ZN(n4544) );
  NAND2_X1 U5516 ( .A1(n4931), .A2(n4930), .ZN(n5264) );
  INV_X1 U5517 ( .A(n5248), .ZN(n4931) );
  OR2_X1 U5518 ( .A1(n5222), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5235) );
  AOI21_X1 U5519 ( .B1(n4826), .B2(n4828), .A(n4375), .ZN(n4825) );
  INV_X1 U5520 ( .A(n4330), .ZN(n4826) );
  OR2_X1 U5521 ( .A1(n5209), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U5522 ( .A1(n4928), .A2(n4927), .ZN(n5209) );
  INV_X1 U5523 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n4927) );
  INV_X1 U5524 ( .A(n5189), .ZN(n4928) );
  INV_X1 U5525 ( .A(n7804), .ZN(n5491) );
  OAI21_X1 U5526 ( .B1(n6983), .B2(n5141), .A(n5140), .ZN(n9981) );
  INV_X1 U5527 ( .A(n5125), .ZN(n4925) );
  NAND2_X1 U5528 ( .A1(n4552), .A2(n4742), .ZN(n6981) );
  AND2_X1 U5529 ( .A1(n4743), .A2(n7784), .ZN(n4742) );
  NAND2_X1 U5530 ( .A1(n4745), .A2(n7792), .ZN(n4743) );
  CLKBUF_X1 U5531 ( .A(n5073), .Z(n10006) );
  NAND2_X1 U5532 ( .A1(n5570), .A2(n5569), .ZN(n5584) );
  NAND2_X1 U5533 ( .A1(n5429), .A2(n5428), .ZN(n7578) );
  NAND2_X1 U5534 ( .A1(n5325), .A2(n5324), .ZN(n7692) );
  OR2_X1 U5535 ( .A1(n5460), .A2(n6255), .ZN(n5121) );
  OR2_X1 U5536 ( .A1(n7903), .A2(n5505), .ZN(n6504) );
  AND2_X1 U5537 ( .A1(n6722), .A2(n7761), .ZN(n10046) );
  INV_X1 U5538 ( .A(n10013), .ZN(n9987) );
  NOR2_X1 U5539 ( .A1(n4859), .A2(P2_IR_REG_22__SCAN_IN), .ZN(n4858) );
  INV_X1 U5540 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5036) );
  NAND2_X1 U5541 ( .A1(n5031), .A2(n4321), .ZN(n5258) );
  INV_X1 U5542 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U5543 ( .A(n4792), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U5544 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4792) );
  NAND2_X1 U5545 ( .A1(n9652), .A2(n9651), .ZN(n9650) );
  AND2_X1 U5546 ( .A1(n5829), .A2(n5828), .ZN(n7285) );
  NAND2_X1 U5547 ( .A1(n5687), .A2(n6874), .ZN(n4572) );
  INV_X1 U5548 ( .A(n7505), .ZN(n4578) );
  NAND2_X1 U5549 ( .A1(n4904), .A2(n7437), .ZN(n4576) );
  NAND2_X1 U5550 ( .A1(n8528), .A2(n5980), .ZN(n8537) );
  NAND2_X1 U5551 ( .A1(n8537), .A2(n8538), .ZN(n8536) );
  OR2_X1 U5552 ( .A1(n6089), .A2(n8488), .ZN(n6111) );
  NAND2_X1 U5553 ( .A1(n4890), .A2(n4889), .ZN(n8554) );
  INV_X1 U5554 ( .A(n8557), .ZN(n4889) );
  INV_X1 U5555 ( .A(n8556), .ZN(n4890) );
  AOI21_X1 U5556 ( .B1(n4887), .B2(n4885), .A(n4362), .ZN(n4884) );
  AND3_X1 U5557 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5755) );
  NOR2_X1 U5558 ( .A1(n5751), .A2(n4869), .ZN(n4868) );
  INV_X1 U5559 ( .A(n5734), .ZN(n4869) );
  NOR2_X1 U5560 ( .A1(n6158), .A2(n4874), .ZN(n4873) );
  OR2_X1 U5561 ( .A1(n8584), .A2(n8585), .ZN(n6158) );
  INV_X1 U5562 ( .A(n4876), .ZN(n4874) );
  INV_X1 U5563 ( .A(n8835), .ZN(n4430) );
  OR2_X1 U5564 ( .A1(n8829), .A2(n4445), .ZN(n8775) );
  NAND2_X1 U5565 ( .A1(n4447), .A2(n4446), .ZN(n4445) );
  NOR2_X1 U5566 ( .A1(n8774), .A2(n9207), .ZN(n4446) );
  XNOR2_X1 U5567 ( .A(n6657), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6655) );
  NAND2_X1 U5568 ( .A1(n6654), .A2(n6655), .ZN(n6653) );
  NOR2_X1 U5569 ( .A1(n6378), .A2(n4391), .ZN(n6353) );
  NAND2_X1 U5570 ( .A1(n6353), .A2(n6354), .ZN(n6408) );
  NOR2_X1 U5571 ( .A1(n8922), .A2(n8921), .ZN(n8925) );
  NOR2_X1 U5572 ( .A1(n8962), .A2(n8961), .ZN(n8969) );
  INV_X1 U5573 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9081) );
  AOI21_X1 U5574 ( .B1(n4615), .B2(n4613), .A(n4612), .ZN(n4611) );
  INV_X1 U5575 ( .A(n9193), .ZN(n4612) );
  OR2_X1 U5576 ( .A1(n9228), .A2(n9169), .ZN(n4662) );
  NOR2_X1 U5577 ( .A1(n9221), .A2(n8772), .ZN(n4661) );
  OAI21_X1 U5578 ( .B1(n9264), .B2(n9164), .A(n9163), .ZN(n9248) );
  AND2_X1 U5579 ( .A1(n8741), .A2(n9265), .ZN(n9295) );
  AOI21_X1 U5580 ( .B1(n4606), .B2(n4608), .A(n4605), .ZN(n4604) );
  INV_X1 U5581 ( .A(n9182), .ZN(n4605) );
  NAND2_X1 U5582 ( .A1(n9391), .A2(n4322), .ZN(n9321) );
  NAND2_X1 U5583 ( .A1(n9391), .A2(n4317), .ZN(n9331) );
  AND2_X1 U5584 ( .A1(n8845), .A2(n9179), .ZN(n9341) );
  AND2_X1 U5585 ( .A1(n8743), .A2(n8843), .ZN(n9353) );
  AND2_X1 U5586 ( .A1(n9391), .A2(n4651), .ZN(n9354) );
  AND2_X1 U5587 ( .A1(n9391), .A2(n9538), .ZN(n9375) );
  NAND2_X1 U5588 ( .A1(n8839), .A2(n8838), .ZN(n9387) );
  NAND2_X1 U5589 ( .A1(n9637), .A2(n9142), .ZN(n9385) );
  NAND2_X1 U5590 ( .A1(n7397), .A2(n4323), .ZN(n9405) );
  NAND2_X1 U5591 ( .A1(n7397), .A2(n4316), .ZN(n9404) );
  NAND2_X1 U5592 ( .A1(n8837), .A2(n8836), .ZN(n9400) );
  AOI21_X1 U5593 ( .B1(n4630), .B2(n4629), .A(n4632), .ZN(n4628) );
  INV_X1 U5594 ( .A(n4634), .ZN(n4630) );
  OR2_X1 U5595 ( .A1(n7464), .A2(n7463), .ZN(n8837) );
  AND2_X1 U5596 ( .A1(n7397), .A2(n9847), .ZN(n7395) );
  NAND2_X1 U5597 ( .A1(n7397), .A2(n4653), .ZN(n7470) );
  NAND2_X1 U5598 ( .A1(n7390), .A2(n8799), .ZN(n7462) );
  OR2_X1 U5599 ( .A1(n7510), .A2(n7296), .ZN(n8658) );
  NAND2_X1 U5600 ( .A1(n7379), .A2(n4634), .ZN(n7390) );
  AOI21_X1 U5601 ( .B1(n8758), .B2(n4667), .A(n4364), .ZN(n4666) );
  INV_X1 U5602 ( .A(n7067), .ZN(n4667) );
  NAND2_X1 U5603 ( .A1(n4637), .A2(n4357), .ZN(n8785) );
  INV_X1 U5604 ( .A(n7053), .ZN(n4637) );
  NAND3_X1 U5605 ( .A1(n8785), .A2(n8794), .A3(n4636), .ZN(n7294) );
  INV_X1 U5606 ( .A(n8729), .ZN(n6021) );
  NOR2_X1 U5607 ( .A1(n9714), .A2(n7031), .ZN(n9715) );
  INV_X1 U5608 ( .A(n6997), .ZN(n4681) );
  NAND2_X1 U5609 ( .A1(n4621), .A2(n4619), .ZN(n9722) );
  INV_X1 U5610 ( .A(n4620), .ZN(n4619) );
  OAI21_X1 U5611 ( .B1(n4623), .B2(n4624), .A(n8792), .ZN(n4620) );
  INV_X1 U5612 ( .A(n6939), .ZN(n8988) );
  NAND2_X1 U5613 ( .A1(n4610), .A2(n4615), .ZN(n9208) );
  NAND2_X1 U5614 ( .A1(n9237), .A2(n4617), .ZN(n4610) );
  NAND2_X1 U5615 ( .A1(n6141), .A2(n6140), .ZN(n9241) );
  NAND2_X1 U5616 ( .A1(n6128), .A2(n6127), .ZN(n9257) );
  NOR2_X1 U5617 ( .A1(n9714), .A2(n4647), .ZN(n7063) );
  INV_X1 U5618 ( .A(n4649), .ZN(n4647) );
  NOR2_X1 U5619 ( .A1(n6474), .A2(n6760), .ZN(n9491) );
  XNOR2_X1 U5620 ( .A(n7751), .B(n7750), .ZN(n8731) );
  NAND2_X1 U5621 ( .A1(n7746), .A2(n7745), .ZN(n7751) );
  XNOR2_X1 U5622 ( .A(n5600), .B(n9546), .ZN(n5604) );
  OR2_X1 U5623 ( .A1(n9545), .A2(n5838), .ZN(n5600) );
  XNOR2_X1 U5624 ( .A(n7595), .B(SI_29_), .ZN(n8720) );
  AOI21_X1 U5625 ( .B1(n5457), .B2(n4717), .A(n4716), .ZN(n4715) );
  INV_X1 U5626 ( .A(n5459), .ZN(n4716) );
  INV_X1 U5627 ( .A(n5439), .ZN(n4717) );
  INV_X1 U5628 ( .A(n5457), .ZN(n4718) );
  INV_X1 U5629 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n4872) );
  NAND2_X1 U5630 ( .A1(n5440), .A2(n5439), .ZN(n5458) );
  XNOR2_X1 U5631 ( .A(n5438), .B(n5437), .ZN(n7459) );
  XNOR2_X1 U5632 ( .A(n5421), .B(n5420), .ZN(n7416) );
  NAND2_X1 U5633 ( .A1(n4704), .A2(n4708), .ZN(n5421) );
  OR2_X1 U5634 ( .A1(n5386), .A2(n4711), .ZN(n4704) );
  NAND2_X1 U5635 ( .A1(n5392), .A2(n5391), .ZN(n5404) );
  OR2_X1 U5636 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  NAND2_X1 U5637 ( .A1(n5386), .A2(n5385), .ZN(n5392) );
  NAND2_X1 U5638 ( .A1(n4727), .A2(n4728), .ZN(n5348) );
  XNOR2_X1 U5639 ( .A(n5335), .B(n5334), .ZN(n7012) );
  NAND2_X1 U5640 ( .A1(n4731), .A2(n5317), .ZN(n5335) );
  OR2_X1 U5641 ( .A1(n5319), .A2(n5318), .ZN(n4731) );
  AND2_X1 U5642 ( .A1(n5594), .A2(n5595), .ZN(n4870) );
  OAI21_X1 U5643 ( .B1(n5272), .B2(n4725), .A(n4723), .ZN(n5301) );
  OAI21_X1 U5644 ( .B1(n5272), .B2(n5007), .A(n5006), .ZN(n5285) );
  XNOR2_X1 U5645 ( .A(n4963), .B(SI_5_), .ZN(n5137) );
  XNOR2_X1 U5646 ( .A(n4959), .B(SI_4_), .ZN(n5115) );
  NOR2_X1 U5647 ( .A1(n5717), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5763) );
  NAND2_X1 U5648 ( .A1(n4798), .A2(n4797), .ZN(n7637) );
  NAND2_X1 U5649 ( .A1(n6639), .A2(n6638), .ZN(n6710) );
  NAND2_X1 U5650 ( .A1(n4802), .A2(n4799), .ZN(n7697) );
  OAI21_X1 U5651 ( .B1(n4475), .B2(n4472), .A(n4473), .ZN(n4471) );
  NAND2_X1 U5652 ( .A1(n4376), .A2(n4477), .ZN(n4473) );
  NAND2_X1 U5653 ( .A1(n7582), .A2(n4474), .ZN(n4472) );
  INV_X1 U5654 ( .A(n4449), .ZN(n4475) );
  NAND2_X1 U5655 ( .A1(n7582), .A2(n4353), .ZN(n4476) );
  NAND2_X1 U5656 ( .A1(n5462), .A2(n5461), .ZN(n7589) );
  NAND2_X1 U5657 ( .A1(n7763), .A2(n6517), .ZN(n6524) );
  NAND2_X1 U5658 ( .A1(n4495), .A2(n4450), .ZN(n4494) );
  NAND2_X1 U5659 ( .A1(n4486), .A2(n4484), .ZN(n7669) );
  AOI21_X1 U5660 ( .B1(n4487), .B2(n4808), .A(n4485), .ZN(n4484) );
  INV_X1 U5661 ( .A(n7670), .ZN(n4485) );
  OAI21_X1 U5662 ( .B1(n7484), .B2(n4808), .A(n4487), .ZN(n7671) );
  INV_X1 U5663 ( .A(n4798), .ZN(n7685) );
  NAND2_X1 U5664 ( .A1(n6710), .A2(n6709), .ZN(n6712) );
  NAND2_X1 U5665 ( .A1(n7714), .A2(n4799), .ZN(n4481) );
  NOR2_X1 U5666 ( .A1(n7704), .A2(n4794), .ZN(n4793) );
  INV_X1 U5667 ( .A(n7565), .ZN(n4794) );
  NAND2_X1 U5668 ( .A1(n7652), .A2(n7565), .ZN(n7705) );
  AND4_X1 U5669 ( .A1(n5163), .A2(n5162), .A3(n5161), .A4(n5160), .ZN(n7129)
         );
  OR2_X1 U5670 ( .A1(n6519), .A2(n6491), .ZN(n7731) );
  NAND2_X1 U5671 ( .A1(n4492), .A2(n4490), .ZN(n6968) );
  INV_X1 U5672 ( .A(n4491), .ZN(n4490) );
  AND2_X1 U5673 ( .A1(n4492), .A2(n4318), .ZN(n6833) );
  NAND2_X1 U5674 ( .A1(n6507), .A2(n6506), .ZN(n7734) );
  OR2_X1 U5675 ( .A1(n6519), .A2(n6518), .ZN(n7730) );
  NAND2_X1 U5676 ( .A1(n7524), .A2(n7523), .ZN(n7526) );
  NAND2_X1 U5677 ( .A1(n7524), .A2(n4807), .ZN(n7546) );
  NAND2_X1 U5678 ( .A1(n4342), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U5679 ( .A1(n7955), .A2(n4326), .ZN(n4736) );
  XNOR2_X1 U5680 ( .A(n5477), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7962) );
  AND2_X1 U5681 ( .A1(n6842), .A2(n5483), .ZN(n7585) );
  INV_X1 U5682 ( .A(n8199), .ZN(n7968) );
  INV_X1 U5683 ( .A(n8247), .ZN(n7972) );
  NAND4_X1 U5684 ( .A1(n5180), .A2(n5179), .A3(n5178), .A4(n5177), .ZN(n7985)
         );
  INV_X1 U5685 ( .A(n7129), .ZN(n9985) );
  NAND2_X1 U5686 ( .A1(n5100), .A2(n5099), .ZN(n7988) );
  NOR2_X1 U5687 ( .A1(n5098), .A2(n4902), .ZN(n5099) );
  AND3_X1 U5688 ( .A1(n5081), .A2(n5080), .A3(n5079), .ZN(n5082) );
  INV_X1 U5689 ( .A(P2_U3893), .ZN(n8122) );
  OAI21_X1 U5690 ( .B1(n6456), .B2(n4504), .A(n6570), .ZN(n6457) );
  INV_X1 U5691 ( .A(n4520), .ZN(n9907) );
  INV_X1 U5692 ( .A(n6578), .ZN(n9905) );
  NOR2_X1 U5693 ( .A1(n9891), .A2(n4897), .ZN(n9909) );
  NAND2_X1 U5694 ( .A1(n4411), .A2(n4781), .ZN(n9934) );
  INV_X1 U5695 ( .A(n4600), .ZN(n9940) );
  INV_X1 U5696 ( .A(n4512), .ZN(n8003) );
  XNOR2_X1 U5697 ( .A(n7260), .B(n7268), .ZN(n7232) );
  NOR2_X1 U5698 ( .A1(n7232), .A2(n7433), .ZN(n7261) );
  NAND2_X1 U5699 ( .A1(n4772), .A2(n4771), .ZN(n8015) );
  NAND2_X1 U5700 ( .A1(n4690), .A2(n8034), .ZN(n8028) );
  INV_X1 U5701 ( .A(n4597), .ZN(n8064) );
  INV_X1 U5702 ( .A(n4517), .ZN(n8079) );
  AOI21_X1 U5703 ( .B1(n4521), .B2(n9951), .A(n4355), .ZN(n8104) );
  NAND2_X1 U5704 ( .A1(n4788), .A2(n8092), .ZN(n4521) );
  INV_X1 U5705 ( .A(n4693), .ZN(n8113) );
  INV_X1 U5706 ( .A(n8131), .ZN(n4787) );
  AOI22_X1 U5707 ( .A1(n8731), .A2(n7753), .B1(n7752), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8166) );
  NAND2_X1 U5708 ( .A1(n4823), .A2(n5581), .ZN(n8170) );
  OAI21_X1 U5709 ( .B1(n4313), .B2(n4327), .A(n4755), .ZN(n8189) );
  NAND2_X1 U5710 ( .A1(n4834), .A2(n4838), .ZN(n8197) );
  NAND2_X1 U5711 ( .A1(n4758), .A2(n7886), .ZN(n8201) );
  NAND2_X1 U5712 ( .A1(n4313), .A2(n4759), .ZN(n4758) );
  XNOR2_X1 U5713 ( .A(n4455), .B(n4454), .ZN(n8207) );
  INV_X1 U5714 ( .A(n8209), .ZN(n4454) );
  OAI21_X1 U5715 ( .B1(n8216), .B2(n4336), .A(n4844), .ZN(n4455) );
  NAND2_X1 U5716 ( .A1(n4313), .A2(n7880), .ZN(n8210) );
  NAND2_X1 U5717 ( .A1(n4750), .A2(n7872), .ZN(n8229) );
  NAND2_X1 U5718 ( .A1(n8238), .A2(n7874), .ZN(n4750) );
  AND2_X1 U5719 ( .A1(n4845), .A2(n4848), .ZN(n8258) );
  NAND2_X1 U5720 ( .A1(n5316), .A2(n4850), .ZN(n8269) );
  NAND2_X1 U5721 ( .A1(n8284), .A2(n7856), .ZN(n8275) );
  NAND2_X1 U5722 ( .A1(n5493), .A2(n7854), .ZN(n8287) );
  NAND2_X1 U5723 ( .A1(n8320), .A2(n5283), .ZN(n8306) );
  NAND2_X1 U5724 ( .A1(n4546), .A2(n4547), .ZN(n7534) );
  OR2_X1 U5725 ( .A1(n10069), .A2(n4550), .ZN(n4546) );
  NAND2_X1 U5726 ( .A1(n5262), .A2(n5261), .ZN(n9619) );
  NAND2_X1 U5727 ( .A1(n10069), .A2(n7828), .ZN(n7493) );
  NAND2_X1 U5728 ( .A1(n5247), .A2(n5246), .ZN(n9627) );
  NAND2_X1 U5729 ( .A1(n4855), .A2(n5242), .ZN(n7494) );
  OR2_X1 U5730 ( .A1(n7450), .A2(n5241), .ZN(n4855) );
  OR2_X1 U5731 ( .A1(n7455), .A2(n7938), .ZN(n10069) );
  NAND2_X1 U5732 ( .A1(n5234), .A2(n5233), .ZN(n10072) );
  NAND2_X1 U5733 ( .A1(n4538), .A2(n7816), .ZN(n7423) );
  NAND2_X1 U5734 ( .A1(n7313), .A2(n7813), .ZN(n4538) );
  NAND2_X1 U5735 ( .A1(n5221), .A2(n5220), .ZN(n10065) );
  NAND2_X1 U5736 ( .A1(n4830), .A2(n4827), .ZN(n7315) );
  NAND2_X1 U5737 ( .A1(n4751), .A2(n7928), .ZN(n7117) );
  NAND2_X1 U5738 ( .A1(n4744), .A2(n7790), .ZN(n6913) );
  NAND2_X1 U5739 ( .A1(n6721), .A2(n7926), .ZN(n4744) );
  OAI211_X1 U5740 ( .C1(n6246), .C2(n9888), .A(n5106), .B(n5105), .ZN(n6726)
         );
  OR2_X1 U5741 ( .A1(n5169), .A2(n6256), .ZN(n5105) );
  AND2_X1 U5742 ( .A1(n10016), .A2(n6724), .ZN(n9996) );
  OR2_X1 U5743 ( .A1(n10054), .A2(n6722), .ZN(n10003) );
  OR2_X1 U5744 ( .A1(n6481), .A2(n6503), .ZN(n10002) );
  INV_X1 U5745 ( .A(n10002), .ZN(n9994) );
  INV_X1 U5746 ( .A(n5584), .ZN(n8171) );
  AND2_X1 U5747 ( .A1(n5581), .A2(n10092), .ZN(n4822) );
  INV_X1 U5748 ( .A(n7589), .ZN(n8181) );
  INV_X1 U5749 ( .A(n8166), .ZN(n8395) );
  NAND2_X1 U5750 ( .A1(n7741), .A2(n7740), .ZN(n7744) );
  NAND2_X1 U5751 ( .A1(n8183), .A2(n10068), .ZN(n5507) );
  INV_X1 U5752 ( .A(n5499), .ZN(n8404) );
  INV_X1 U5753 ( .A(n7578), .ZN(n8408) );
  INV_X1 U5754 ( .A(n7575), .ZN(n8412) );
  INV_X1 U5755 ( .A(n7641), .ZN(n8418) );
  INV_X1 U5756 ( .A(n7562), .ZN(n8426) );
  NAND2_X1 U5757 ( .A1(n5186), .A2(n5185), .ZN(n7139) );
  OR2_X1 U5758 ( .A1(n10076), .A2(n10054), .ZN(n8450) );
  INV_X2 U5759 ( .A(n10076), .ZN(n10074) );
  XNOR2_X1 U5760 ( .A(n5515), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5761 ( .A1(n4862), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4920) );
  NAND2_X1 U5762 ( .A1(n5513), .A2(n5512), .ZN(n7366) );
  INV_X1 U5763 ( .A(n5539), .ZN(n7762) );
  OR2_X1 U5764 ( .A1(n5474), .A2(n5472), .ZN(n5476) );
  INV_X1 U5765 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U5766 ( .A1(n5031), .A2(n9111), .ZN(n5231) );
  INV_X1 U5767 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9103) );
  INV_X1 U5768 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6295) );
  INV_X1 U5769 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6289) );
  INV_X1 U5770 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6265) );
  INV_X1 U5771 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6264) );
  INV_X1 U5772 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6260) );
  NAND2_X1 U5773 ( .A1(n5118), .A2(n5119), .ZN(n6577) );
  INV_X1 U5774 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6255) );
  INV_X1 U5775 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6257) );
  INV_X1 U5776 ( .A(n6447), .ZN(n6435) );
  INV_X1 U5777 ( .A(n4867), .ZN(n4863) );
  INV_X1 U5778 ( .A(n6623), .ZN(n4565) );
  NAND2_X1 U5779 ( .A1(n8554), .A2(n6057), .ZN(n8511) );
  NAND2_X1 U5780 ( .A1(n8545), .A2(n6126), .ZN(n8520) );
  NAND2_X1 U5781 ( .A1(n4875), .A2(n4876), .ZN(n8518) );
  NAND2_X1 U5782 ( .A1(n8595), .A2(n5960), .ZN(n8529) );
  NAND2_X1 U5783 ( .A1(n4594), .A2(n8503), .ZN(n8556) );
  NAND2_X1 U5784 ( .A1(n4589), .A2(n4588), .ZN(n4594) );
  INV_X1 U5785 ( .A(n8501), .ZN(n4589) );
  XNOR2_X1 U5786 ( .A(n8482), .B(n8484), .ZN(n8566) );
  NAND2_X1 U5787 ( .A1(n6085), .A2(n6084), .ZN(n9307) );
  INV_X1 U5788 ( .A(n9660), .ZN(n8599) );
  AND2_X1 U5789 ( .A1(n6230), .A2(n6209), .ZN(n9649) );
  INV_X1 U5790 ( .A(n9649), .ZN(n9665) );
  OR2_X1 U5791 ( .A1(n6542), .A2(n5661), .ZN(n5662) );
  NOR2_X1 U5792 ( .A1(n6330), .A2(n4526), .ZN(n6692) );
  NOR2_X1 U5793 ( .A1(n6329), .A2(n6766), .ZN(n4526) );
  INV_X1 U5794 ( .A(n4525), .ZN(n6690) );
  NOR2_X1 U5795 ( .A1(n6361), .A2(n4532), .ZN(n6380) );
  AND2_X1 U5796 ( .A1(n6350), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4532) );
  NOR2_X1 U5797 ( .A1(n6380), .A2(n6379), .ZN(n6378) );
  NOR2_X1 U5798 ( .A1(n6605), .A2(n4529), .ZN(n6609) );
  AND2_X1 U5799 ( .A1(n6606), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4529) );
  NOR2_X1 U5800 ( .A1(n6608), .A2(n6609), .ZN(n6732) );
  NOR2_X1 U5801 ( .A1(n4530), .A2(n6732), .ZN(n9684) );
  AND2_X1 U5802 ( .A1(n6733), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U5803 ( .A1(n9684), .A2(n9685), .ZN(n9683) );
  NOR2_X1 U5804 ( .A1(n6957), .A2(n4534), .ZN(n6961) );
  AND2_X1 U5805 ( .A1(n6958), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4534) );
  NOR2_X1 U5806 ( .A1(n6961), .A2(n6960), .ZN(n7142) );
  XNOR2_X1 U5807 ( .A(n8920), .B(n8919), .ZN(n7144) );
  NOR2_X1 U5808 ( .A1(n7469), .A2(n7144), .ZN(n8921) );
  NOR2_X1 U5809 ( .A1(n8933), .A2(n4528), .ZN(n8936) );
  AND2_X1 U5810 ( .A1(n8934), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5811 ( .A1(n8936), .A2(n8935), .ZN(n8956) );
  OR3_X1 U5812 ( .A1(n9214), .A2(n9213), .A3(n9403), .ZN(n9432) );
  NAND2_X1 U5813 ( .A1(n9315), .A2(n9180), .ZN(n9300) );
  INV_X1 U5814 ( .A(n4297), .ZN(n9140) );
  INV_X1 U5815 ( .A(n4676), .ZN(n4672) );
  NAND2_X1 U5816 ( .A1(n4671), .A2(n7376), .ZN(n7474) );
  NAND2_X1 U5817 ( .A1(n4668), .A2(n7067), .ZN(n7153) );
  NAND2_X1 U5818 ( .A1(n7066), .A2(n8753), .ZN(n4668) );
  NAND2_X1 U5819 ( .A1(n4682), .A2(n6997), .ZN(n7026) );
  NAND2_X1 U5820 ( .A1(n4622), .A2(n4624), .ZN(n6999) );
  NAND2_X1 U5821 ( .A1(n6803), .A2(n6802), .ZN(n6847) );
  NAND2_X1 U5822 ( .A1(n8877), .A2(n6471), .ZN(n9741) );
  INV_X1 U5823 ( .A(n9744), .ZN(n9410) );
  NAND2_X1 U5824 ( .A1(n9877), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n4464) );
  AND2_X1 U5825 ( .A1(n9426), .A2(n9429), .ZN(n9430) );
  INV_X1 U5826 ( .A(n9291), .ZN(n9522) );
  NAND2_X1 U5827 ( .A1(n5615), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U5828 ( .A1(n5386), .A2(n5373), .ZN(n7193) );
  NOR2_X1 U5829 ( .A1(n6202), .A2(n5838), .ZN(n4583) );
  INV_X1 U5830 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6376) );
  INV_X1 U5831 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6296) );
  INV_X1 U5832 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6290) );
  INV_X1 U5833 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6276) );
  INV_X1 U5834 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6266) );
  INV_X1 U5835 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6262) );
  INV_X1 U5836 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6258) );
  INV_X1 U5837 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9102) );
  INV_X1 U5838 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6252) );
  XNOR2_X1 U5839 ( .A(n4531), .B(n5684), .ZN(n6657) );
  OR2_X1 U5840 ( .A1(n5638), .A2(n5838), .ZN(n4531) );
  NOR2_X2 U5841 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9566) );
  AND2_X1 U5842 ( .A1(n4600), .A2(n6886), .ZN(n6888) );
  INV_X1 U5843 ( .A(n4427), .ZN(n7077) );
  INV_X1 U5844 ( .A(n4688), .ZN(n8067) );
  XNOR2_X1 U5845 ( .A(n4691), .B(n8139), .ZN(n8161) );
  INV_X1 U5846 ( .A(n4523), .ZN(n6391) );
  INV_X1 U5847 ( .A(n4638), .ZN(n9203) );
  OAI21_X1 U5848 ( .B1(n9426), .B2(n9758), .A(n4639), .ZN(n4638) );
  AOI21_X1 U5849 ( .B1(n9427), .B2(n9754), .A(n9202), .ZN(n4639) );
  NAND2_X1 U5850 ( .A1(n4465), .A2(n4462), .ZN(P1_U3550) );
  INV_X1 U5851 ( .A(n4463), .ZN(n4462) );
  NAND2_X1 U5852 ( .A1(n9502), .A2(n9879), .ZN(n4465) );
  OAI21_X1 U5853 ( .B1(n9503), .B2(n9489), .A(n4464), .ZN(n4463) );
  AOI21_X1 U5854 ( .B1(n9228), .B2(n4435), .A(n4434), .ZN(n4433) );
  NOR2_X1 U5855 ( .A1(n9879), .A2(n9439), .ZN(n4434) );
  NAND2_X1 U5856 ( .A1(n4470), .A2(n4468), .ZN(P1_U3518) );
  AOI22_X1 U5857 ( .A1(n9212), .A2(n4469), .B1(P1_REG0_REG_28__SCAN_IN), .B2(
        n9860), .ZN(n4468) );
  NAND2_X1 U5858 ( .A1(n9502), .A2(n9862), .ZN(n4470) );
  NAND2_X1 U5859 ( .A1(n9228), .A2(n4469), .ZN(n4451) );
  XOR2_X1 U5860 ( .A(n7950), .B(n7210), .Z(n4312) );
  OAI21_X1 U5861 ( .B1(n7356), .B2(n7439), .A(n4579), .ZN(n7441) );
  NAND2_X1 U5862 ( .A1(n4450), .A2(n7569), .ZN(n4798) );
  OR2_X1 U5863 ( .A1(n8222), .A2(n7879), .ZN(n4313) );
  AND2_X1 U5864 ( .A1(n4374), .A2(n4798), .ZN(n4314) );
  AND2_X1 U5865 ( .A1(n4763), .A2(n7854), .ZN(n4315) );
  AND2_X1 U5866 ( .A1(n4653), .A2(n9641), .ZN(n4316) );
  AND2_X1 U5867 ( .A1(n9338), .A2(n4651), .ZN(n4317) );
  INV_X1 U5868 ( .A(n8438), .ZN(n7722) );
  AND2_X1 U5869 ( .A1(n5047), .A2(n5046), .ZN(n8438) );
  NAND2_X1 U5870 ( .A1(n6829), .A2(n6828), .ZN(n4318) );
  XOR2_X1 U5871 ( .A(n7584), .B(n7968), .Z(n4319) );
  AND2_X1 U5872 ( .A1(n4547), .A2(n7836), .ZN(n4320) );
  AND2_X1 U5873 ( .A1(n4816), .A2(n5032), .ZN(n4321) );
  NAND2_X1 U5874 ( .A1(n6004), .A2(n6003), .ZN(n9377) );
  AND2_X1 U5875 ( .A1(n4317), .A2(n4650), .ZN(n4322) );
  AND2_X1 U5876 ( .A1(n4316), .A2(n4652), .ZN(n4323) );
  AND3_X1 U5877 ( .A1(n5122), .A2(n5121), .A3(n5120), .ZN(n10030) );
  INV_X1 U5878 ( .A(n10030), .ZN(n4856) );
  NAND3_X1 U5879 ( .A1(n4916), .A2(n5197), .A3(n4860), .ZN(n4324) );
  NAND2_X1 U5880 ( .A1(n5383), .A2(n5382), .ZN(n7971) );
  INV_X1 U5881 ( .A(n7971), .ZN(n8237) );
  INV_X1 U5882 ( .A(n9228), .ZN(n9507) );
  AND2_X1 U5883 ( .A1(n4565), .A2(n5678), .ZN(n4325) );
  INV_X1 U5884 ( .A(n8758), .ZN(n4636) );
  NAND2_X1 U5885 ( .A1(n4815), .A2(n6970), .ZN(n7132) );
  NAND2_X1 U5886 ( .A1(n4775), .A2(n9928), .ZN(n4781) );
  INV_X1 U5887 ( .A(n7268), .ZN(n4511) );
  NOR2_X1 U5888 ( .A1(n5539), .A2(n7014), .ZN(n4326) );
  NAND2_X1 U5889 ( .A1(n4496), .A2(n7570), .ZN(n4797) );
  OR2_X1 U5890 ( .A1(n7884), .A2(n4757), .ZN(n4327) );
  AND2_X1 U5891 ( .A1(n4481), .A2(n4800), .ZN(n4328) );
  INV_X1 U5892 ( .A(n4808), .ZN(n4807) );
  NAND2_X1 U5893 ( .A1(n7528), .A2(n7523), .ZN(n4808) );
  AND2_X1 U5894 ( .A1(n7584), .A2(n7968), .ZN(n4329) );
  INV_X1 U5895 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n4820) );
  OR2_X1 U5896 ( .A1(n7316), .A2(n10049), .ZN(n4330) );
  OR2_X1 U5897 ( .A1(n8177), .A2(n10056), .ZN(n4331) );
  NOR2_X1 U5898 ( .A1(n8476), .A2(n8886), .ZN(n4332) );
  OR2_X1 U5899 ( .A1(n5494), .A2(n4762), .ZN(n4333) );
  NAND2_X1 U5900 ( .A1(n6577), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4334) );
  OR2_X1 U5901 ( .A1(n4310), .A2(n6305), .ZN(n4335) );
  NOR2_X1 U5902 ( .A1(n8415), .A2(n8227), .ZN(n4336) );
  NAND2_X1 U5903 ( .A1(n4501), .A2(n4497), .ZN(n7659) );
  NAND2_X1 U5904 ( .A1(n4939), .A2(n8455), .ZN(n5078) );
  OR2_X1 U5905 ( .A1(n8078), .A2(n8063), .ZN(n4337) );
  INV_X1 U5906 ( .A(n9275), .ZN(n9518) );
  AND2_X1 U5907 ( .A1(n7555), .A2(n8296), .ZN(n4338) );
  AND2_X1 U5908 ( .A1(n4539), .A2(n7422), .ZN(n4339) );
  AND2_X1 U5909 ( .A1(n9353), .A2(n8842), .ZN(n4340) );
  OR2_X1 U5910 ( .A1(n7268), .A2(n7267), .ZN(n4341) );
  OR2_X1 U5911 ( .A1(n8395), .A2(n8163), .ZN(n4342) );
  AND2_X1 U5912 ( .A1(n9291), .A2(n9160), .ZN(n4343) );
  OR2_X1 U5913 ( .A1(n4310), .A2(n6329), .ZN(n4344) );
  AND2_X1 U5914 ( .A1(n7706), .A2(n7568), .ZN(n4450) );
  NAND2_X1 U5915 ( .A1(n7726), .A2(n8208), .ZN(n4449) );
  AND2_X1 U5916 ( .A1(n5029), .A2(n5026), .ZN(n4345) );
  NAND2_X1 U5917 ( .A1(n5599), .A2(n5617), .ZN(n5613) );
  AND2_X1 U5918 ( .A1(n4772), .A2(n4770), .ZN(n4346) );
  XNOR2_X1 U5919 ( .A(n7641), .B(n7210), .ZN(n7569) );
  INV_X1 U5920 ( .A(n4802), .ZN(n7713) );
  XNOR2_X1 U5921 ( .A(n7589), .B(n8188), .ZN(n7950) );
  AND2_X1 U5922 ( .A1(n4556), .A2(n7898), .ZN(n4347) );
  INV_X1 U5923 ( .A(n4908), .ZN(n5101) );
  AND2_X1 U5924 ( .A1(n8263), .A2(n4848), .ZN(n4348) );
  INV_X1 U5925 ( .A(n4801), .ZN(n4800) );
  OAI21_X1 U5926 ( .B1(n4805), .B2(n4803), .A(n7561), .ZN(n4801) );
  INV_X1 U5927 ( .A(n8296), .ZN(n7976) );
  AND4_X1 U5928 ( .A1(n5053), .A2(n5052), .A3(n5051), .A4(n5050), .ZN(n8296)
         );
  AND2_X1 U5929 ( .A1(n5202), .A2(n5201), .ZN(n10049) );
  OR2_X1 U5930 ( .A1(n7703), .A2(n8247), .ZN(n7872) );
  INV_X1 U5931 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8452) );
  AND2_X1 U5932 ( .A1(n5491), .A2(n7928), .ZN(n4349) );
  AND2_X1 U5933 ( .A1(n4523), .A2(n4522), .ZN(n4350) );
  INV_X1 U5934 ( .A(n4784), .ZN(n4783) );
  OR2_X1 U5935 ( .A1(n8896), .A2(n9789), .ZN(n4351) );
  AND2_X1 U5936 ( .A1(n4883), .A2(n5796), .ZN(n4352) );
  NAND2_X1 U5937 ( .A1(n9289), .A2(n4656), .ZN(n4659) );
  OR2_X1 U5938 ( .A1(n5135), .A2(n5134), .ZN(n9928) );
  AND2_X1 U5939 ( .A1(n4312), .A2(n4319), .ZN(n4353) );
  NOR2_X1 U5940 ( .A1(n9323), .A2(n9155), .ZN(n4354) );
  AND2_X1 U5941 ( .A1(n8101), .A2(n9970), .ZN(n4355) );
  NOR2_X1 U5942 ( .A1(n7713), .A2(n4338), .ZN(n4356) );
  AND2_X1 U5943 ( .A1(n8754), .A2(n8638), .ZN(n4357) );
  AND2_X1 U5944 ( .A1(n4517), .A2(n4516), .ZN(n4358) );
  OR2_X1 U5945 ( .A1(n9257), .A2(n8702), .ZN(n9187) );
  AND2_X1 U5946 ( .A1(n9627), .A2(n7980), .ZN(n4359) );
  AND2_X1 U5947 ( .A1(n4614), .A2(n9187), .ZN(n4360) );
  AND2_X1 U5948 ( .A1(n9207), .A2(n4662), .ZN(n4361) );
  AND2_X1 U5949 ( .A1(n6074), .A2(n6073), .ZN(n4362) );
  AND2_X1 U5950 ( .A1(n4449), .A2(n7582), .ZN(n4363) );
  NOR2_X1 U5951 ( .A1(n7154), .A2(n8890), .ZN(n4364) );
  OR2_X1 U5952 ( .A1(n8299), .A2(n8309), .ZN(n7847) );
  NAND2_X1 U5953 ( .A1(n8778), .A2(n8826), .ZN(n9195) );
  OR2_X1 U5954 ( .A1(n9619), .A2(n8326), .ZN(n7836) );
  AND2_X1 U5955 ( .A1(n7582), .A2(n4319), .ZN(n4365) );
  AND2_X1 U5956 ( .A1(n5034), .A2(n5033), .ZN(n4366) );
  OR2_X1 U5957 ( .A1(n5508), .A2(n4917), .ZN(n4367) );
  AND2_X1 U5958 ( .A1(n5497), .A2(n8227), .ZN(n7879) );
  INV_X1 U5959 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5032) );
  INV_X1 U5960 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U5961 ( .A1(n8408), .A2(n8208), .ZN(n4368) );
  NOR2_X1 U5962 ( .A1(n7578), .A2(n7969), .ZN(n4369) );
  INV_X1 U5963 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5536) );
  AND2_X1 U5964 ( .A1(n7545), .A2(n7978), .ZN(n4370) );
  OR2_X1 U5965 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4371) );
  AND2_X1 U5966 ( .A1(n4892), .A2(n5635), .ZN(n4372) );
  NOR2_X1 U5967 ( .A1(n6124), .A2(n6123), .ZN(n6125) );
  AND2_X1 U5968 ( .A1(n9377), .A2(n9147), .ZN(n4373) );
  AND2_X1 U5969 ( .A1(n4797), .A2(n8237), .ZN(n4374) );
  INV_X1 U5970 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6248) );
  NOR2_X1 U5971 ( .A1(n10055), .A2(n7431), .ZN(n4375) );
  INV_X1 U5972 ( .A(n8286), .ZN(n4763) );
  OR2_X1 U5973 ( .A1(n4312), .A2(n4329), .ZN(n4376) );
  AND2_X1 U5974 ( .A1(n7505), .A2(n4581), .ZN(n4377) );
  AND2_X1 U5975 ( .A1(n7027), .A2(n9808), .ZN(n4378) );
  AND2_X1 U5976 ( .A1(n4788), .A2(n4787), .ZN(n4379) );
  AND2_X1 U5977 ( .A1(n5595), .A2(n4872), .ZN(n4380) );
  NOR2_X1 U5978 ( .A1(n5215), .A2(n4829), .ZN(n4828) );
  AND2_X1 U5979 ( .A1(n6001), .A2(n6015), .ZN(n4381) );
  AND2_X1 U5980 ( .A1(n4626), .A2(n6998), .ZN(n4382) );
  AND2_X1 U5981 ( .A1(n4590), .A2(n4884), .ZN(n4383) );
  AND2_X1 U5982 ( .A1(n5623), .A2(n5624), .ZN(n4384) );
  AND2_X1 U5983 ( .A1(n5298), .A2(n5283), .ZN(n4385) );
  AND2_X1 U5984 ( .A1(n4321), .A2(n4366), .ZN(n4386) );
  AND2_X1 U5985 ( .A1(n5931), .A2(n5919), .ZN(n4387) );
  INV_X1 U5986 ( .A(n4860), .ZN(n4859) );
  AND2_X1 U5987 ( .A1(n4909), .A2(n4910), .ZN(n4860) );
  AND2_X1 U5988 ( .A1(n4820), .A2(n4860), .ZN(n4388) );
  INV_X1 U5989 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5635) );
  NAND2_X1 U5990 ( .A1(n7660), .A2(n4503), .ZN(n4389) );
  AND2_X1 U5991 ( .A1(n9471), .A2(n9153), .ZN(n4390) );
  INV_X1 U5992 ( .A(n9241), .ZN(n4657) );
  NAND2_X1 U5993 ( .A1(n6059), .A2(n6058), .ZN(n9323) );
  INV_X1 U5994 ( .A(n9323), .ZN(n4650) );
  NAND2_X1 U5995 ( .A1(n9650), .A2(n5796), .ZN(n7282) );
  NAND2_X1 U5996 ( .A1(n7356), .A2(n7357), .ZN(n7355) );
  INV_X1 U5997 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4461) );
  INV_X1 U5998 ( .A(n4457), .ZN(n4652) );
  INV_X1 U5999 ( .A(n8799), .ZN(n4633) );
  INV_X1 U6000 ( .A(n9212), .ZN(n9503) );
  AND2_X1 U6001 ( .A1(n6352), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4391) );
  INV_X1 U6002 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4817) );
  AND2_X1 U6003 ( .A1(n5197), .A2(n4909), .ZN(n5199) );
  AND2_X1 U6004 ( .A1(n9783), .A2(n9789), .ZN(n4392) );
  INV_X1 U6005 ( .A(n7650), .ZN(n4483) );
  OR2_X1 U6006 ( .A1(n8412), .A2(n8394), .ZN(n4393) );
  AND4_X1 U6007 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n8325)
         );
  AND2_X1 U6008 ( .A1(n7379), .A2(n8658), .ZN(n4394) );
  NAND2_X1 U6009 ( .A1(n5594), .A2(n4299), .ZN(n5961) );
  OR2_X1 U6010 ( .A1(n8476), .A2(n7377), .ZN(n8803) );
  INV_X1 U6011 ( .A(n8803), .ZN(n4632) );
  NAND2_X1 U6012 ( .A1(n7645), .A2(n4804), .ZN(n4803) );
  INV_X1 U6013 ( .A(n4803), .ZN(n4799) );
  AND2_X1 U6014 ( .A1(n4723), .A2(n4722), .ZN(n4395) );
  NOR2_X1 U6015 ( .A1(n4864), .A2(n4863), .ZN(n4396) );
  AND2_X1 U6016 ( .A1(n4725), .A2(n4722), .ZN(n4397) );
  AND2_X1 U6017 ( .A1(n6036), .A2(n6037), .ZN(n8502) );
  INV_X1 U6018 ( .A(n8502), .ZN(n4588) );
  AND2_X1 U6019 ( .A1(n5031), .A2(n4386), .ZN(n5042) );
  AND2_X1 U6020 ( .A1(n4733), .A2(n5334), .ZN(n4732) );
  AND2_X1 U6021 ( .A1(n4728), .A2(n5347), .ZN(n4398) );
  AND2_X1 U6022 ( .A1(n5031), .A2(n4816), .ZN(n4399) );
  OR2_X1 U6023 ( .A1(n4766), .A2(n4511), .ZN(n4400) );
  AND2_X1 U6024 ( .A1(n4769), .A2(n4772), .ZN(n4401) );
  OR2_X1 U6025 ( .A1(n4675), .A2(n4672), .ZN(n4402) );
  INV_X1 U6026 ( .A(n9542), .ZN(n4469) );
  AND2_X1 U6027 ( .A1(n8023), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n4403) );
  NOR2_X1 U6028 ( .A1(n7739), .A2(n7367), .ZN(n4404) );
  OR2_X1 U6029 ( .A1(n9714), .A2(n4648), .ZN(n4405) );
  NAND2_X1 U6030 ( .A1(n8868), .A2(n8980), .ZN(n8738) );
  NAND2_X1 U6031 ( .A1(n4870), .A2(n4299), .ZN(n5981) );
  AND2_X1 U6032 ( .A1(n8785), .A2(n8794), .ZN(n4406) );
  NOR3_X1 U6033 ( .A1(n9714), .A2(n7305), .A3(n4648), .ZN(n4646) );
  NAND2_X1 U6034 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  OR2_X1 U6035 ( .A1(n6518), .A2(n7903), .ZN(n8307) );
  INV_X1 U6036 ( .A(n9879), .ZN(n9877) );
  AND2_X1 U6037 ( .A1(n9979), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4407) );
  AND2_X1 U6038 ( .A1(n4781), .A2(n4782), .ZN(n4408) );
  OR2_X1 U6039 ( .A1(n8729), .A2(n6846), .ZN(n4409) );
  NOR2_X1 U6040 ( .A1(n9909), .A2(n9908), .ZN(n4410) );
  AND2_X1 U6041 ( .A1(n4782), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4411) );
  INV_X1 U6042 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4791) );
  XNOR2_X1 U6043 ( .A(n5037), .B(n5036), .ZN(n8154) );
  NOR2_X1 U6044 ( .A1(n5601), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U6045 ( .A1(n4495), .A2(n4389), .ZN(n4493) );
  INV_X1 U6046 ( .A(n5319), .ZN(n4412) );
  OAI21_X1 U6047 ( .B1(n4501), .B2(n4500), .A(n4499), .ZN(n4498) );
  OAI21_X2 U6048 ( .B1(n5256), .B2(n5257), .A(n5003), .ZN(n5272) );
  OAI21_X2 U6049 ( .B1(n5230), .B2(n4992), .A(n4995), .ZN(n5244) );
  OAI21_X2 U6050 ( .B1(n5204), .B2(n4983), .A(n4986), .ZN(n5217) );
  OAI21_X2 U6051 ( .B1(n5217), .B2(n5216), .A(n4991), .ZN(n5230) );
  NAND2_X1 U6052 ( .A1(n4413), .A2(n4955), .ZN(n5103) );
  NAND2_X1 U6053 ( .A1(n5084), .A2(n5085), .ZN(n4413) );
  AOI21_X1 U6054 ( .B1(n4414), .B2(n7883), .A(n8209), .ZN(n7894) );
  NAND2_X1 U6055 ( .A1(n7877), .A2(n4415), .ZN(n4414) );
  NAND2_X1 U6056 ( .A1(n7900), .A2(n4417), .ZN(n7909) );
  XNOR2_X1 U6057 ( .A(n8063), .B(n8078), .ZN(n8038) );
  XNOR2_X1 U6058 ( .A(n8108), .B(n8130), .ZN(n8088) );
  NOR2_X2 U6059 ( .A1(n8087), .A2(n4686), .ZN(n8108) );
  NOR2_X2 U6060 ( .A1(n9926), .A2(n5124), .ZN(n9925) );
  OAI22_X1 U6061 ( .A1(n9941), .A2(n4598), .B1(n6886), .B2(n6887), .ZN(n7072)
         );
  NOR2_X1 U6062 ( .A1(n6566), .A2(n6565), .ZN(n6567) );
  INV_X1 U6063 ( .A(n8735), .ZN(n9496) );
  NAND2_X1 U6064 ( .A1(n5020), .A2(n5019), .ZN(n5319) );
  INV_X1 U6065 ( .A(n4607), .ZN(n4606) );
  NAND2_X1 U6066 ( .A1(n9251), .A2(n9186), .ZN(n9188) );
  NAND2_X1 U6067 ( .A1(n9283), .A2(n9184), .ZN(n9268) );
  NAND2_X1 U6068 ( .A1(n4436), .A2(n4433), .ZN(P1_U3549) );
  OR2_X1 U6069 ( .A1(n9504), .A2(n9877), .ZN(n4436) );
  OAI211_X1 U6070 ( .C1(n4739), .C2(n4737), .A(n7956), .B(n4736), .ZN(n7958)
         );
  OR2_X1 U6071 ( .A1(n8726), .A2(n9195), .ZN(n8728) );
  NAND2_X1 U6072 ( .A1(n8709), .A2(n9186), .ZN(n4440) );
  AOI21_X1 U6073 ( .B1(n8864), .B2(n8786), .A(n4437), .ZN(n8863) );
  AND4_X1 U6074 ( .A1(n8716), .A2(n8777), .A3(n8715), .A4(n8714), .ZN(n8718)
         );
  AOI21_X1 U6075 ( .B1(n8700), .B2(n4439), .A(n4438), .ZN(n8709) );
  NAND3_X1 U6076 ( .A1(n8732), .A2(n8733), .A3(n8831), .ZN(n8736) );
  INV_X1 U6077 ( .A(n9207), .ZN(n4614) );
  XNOR2_X1 U6078 ( .A(n5563), .B(n5562), .ZN(n8459) );
  AOI21_X2 U6079 ( .B1(n8484), .B2(n4587), .A(n8564), .ZN(n8485) );
  NAND2_X1 U6080 ( .A1(n5659), .A2(n6668), .ZN(n6623) );
  NAND2_X1 U6081 ( .A1(n9664), .A2(n5730), .ZN(n9661) );
  OAI21_X2 U6082 ( .B1(n9248), .B2(n9166), .A(n4456), .ZN(n9235) );
  OAI21_X2 U6083 ( .B1(n4569), .B2(n4570), .A(n4566), .ZN(n8528) );
  NAND2_X1 U6084 ( .A1(n8493), .A2(n8494), .ZN(n9664) );
  NOR2_X1 U6085 ( .A1(n7439), .A2(n4578), .ZN(n4577) );
  OAI21_X1 U6086 ( .B1(n8827), .B2(n8828), .A(n8826), .ZN(n8847) );
  NAND3_X1 U6087 ( .A1(n7895), .A2(n7954), .A3(n7896), .ZN(n7900) );
  NAND2_X1 U6088 ( .A1(n4502), .A2(n4796), .ZN(n4501) );
  INV_X1 U6089 ( .A(n4498), .ZN(n4495) );
  OAI21_X1 U6090 ( .B1(n7915), .B2(n7914), .A(n7913), .ZN(n7916) );
  OAI211_X1 U6091 ( .C1(n4363), .C2(n4319), .A(n7727), .B(n4448), .ZN(n7609)
         );
  NAND2_X1 U6092 ( .A1(n4365), .A2(n4449), .ZN(n4448) );
  NAND2_X1 U6093 ( .A1(n4714), .A2(n4712), .ZN(n5567) );
  NAND2_X1 U6094 ( .A1(n6703), .A2(n8730), .ZN(n4467) );
  NAND2_X1 U6095 ( .A1(n4966), .A2(n4965), .ZN(n5151) );
  NAND2_X1 U6096 ( .A1(n7401), .A2(n7402), .ZN(n4671) );
  NAND2_X1 U6097 ( .A1(n7372), .A2(n7371), .ZN(n7374) );
  OAI21_X2 U6098 ( .B1(n9294), .B2(n4343), .A(n9161), .ZN(n9264) );
  NAND2_X1 U6099 ( .A1(n9152), .A2(n9151), .ZN(n9330) );
  OR2_X2 U6100 ( .A1(n9235), .A2(n9167), .ZN(n4663) );
  NAND2_X1 U6101 ( .A1(n5642), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4460) );
  NAND2_X1 U6102 ( .A1(n9506), .A2(n4451), .ZN(P1_U3517) );
  NOR2_X1 U6103 ( .A1(n8763), .A2(n4633), .ZN(n4629) );
  OAI21_X1 U6104 ( .B1(n7379), .B2(n4631), .A(n4628), .ZN(n7464) );
  INV_X1 U6105 ( .A(n9563), .ZN(n6185) );
  NAND2_X1 U6106 ( .A1(n4727), .A2(n4398), .ZN(n5352) );
  NAND3_X1 U6107 ( .A1(n9188), .A2(n4615), .A3(n4360), .ZN(n4609) );
  NAND2_X1 U6108 ( .A1(n4719), .A2(n5040), .ZN(n5020) );
  NAND2_X1 U6109 ( .A1(n8353), .A2(n4393), .ZN(P2_U3484) );
  OR2_X1 U6110 ( .A1(n5642), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4459) );
  NAND2_X1 U6111 ( .A1(n4674), .A2(n4676), .ZN(n4673) );
  NAND2_X1 U6112 ( .A1(n4866), .A2(n4865), .ZN(n4864) );
  NAND2_X1 U6113 ( .A1(n4575), .A2(n4574), .ZN(n4573) );
  NAND2_X1 U6114 ( .A1(n7513), .A2(n7514), .ZN(n7512) );
  NAND2_X1 U6115 ( .A1(n4700), .A2(n4972), .ZN(n5183) );
  NAND2_X1 U6116 ( .A1(n4458), .A2(n4958), .ZN(n5114) );
  NAND2_X1 U6117 ( .A1(n4952), .A2(n4951), .ZN(n5084) );
  AND2_X1 U6118 ( .A1(n8758), .A2(n8753), .ZN(n4665) );
  NAND2_X1 U6119 ( .A1(n5103), .A2(n5104), .ZN(n4458) );
  NOR2_X1 U6120 ( .A1(n8088), .A2(n8301), .ZN(n8109) );
  INV_X1 U6121 ( .A(n8026), .ZN(n4689) );
  OR2_X2 U6122 ( .A1(n4675), .A2(n4673), .ZN(n9637) );
  NAND2_X1 U6123 ( .A1(n9566), .A2(n4945), .ZN(n4703) );
  OAI211_X2 U6124 ( .C1(n6281), .C2(n6372), .A(n5789), .B(n5788), .ZN(n9656)
         );
  NAND2_X1 U6125 ( .A1(n4707), .A2(n4705), .ZN(n5423) );
  NAND2_X1 U6126 ( .A1(n4701), .A2(n4969), .ZN(n5167) );
  OAI21_X1 U6127 ( .B1(n5440), .B2(n4718), .A(n4715), .ZN(n5563) );
  NAND2_X1 U6128 ( .A1(n6798), .A2(n8746), .ZN(n6801) );
  NAND2_X1 U6129 ( .A1(n8788), .A2(n6802), .ZN(n8746) );
  AND2_X1 U6130 ( .A1(n5706), .A2(n4344), .ZN(n4466) );
  NAND2_X1 U6131 ( .A1(n5136), .A2(n5137), .ZN(n4966) );
  NAND2_X1 U6132 ( .A1(n5244), .A2(n4996), .ZN(n4734) );
  NAND2_X1 U6133 ( .A1(n4660), .A2(n4662), .ZN(n9204) );
  NAND2_X1 U6134 ( .A1(n9159), .A2(n9158), .ZN(n9294) );
  NAND2_X1 U6135 ( .A1(n5196), .A2(n5195), .ZN(n4735) );
  INV_X1 U6136 ( .A(n9352), .ZN(n9149) );
  OAI21_X1 U6137 ( .B1(n4476), .B2(n4475), .A(n4471), .ZN(n7591) );
  NAND2_X1 U6138 ( .A1(n7714), .A2(n4482), .ZN(n4480) );
  NAND2_X1 U6139 ( .A1(n7484), .A2(n4487), .ZN(n4486) );
  NAND2_X1 U6140 ( .A1(n6831), .A2(n6830), .ZN(n4492) );
  AND3_X2 U6141 ( .A1(n4908), .A2(n4820), .A3(n4290), .ZN(n5197) );
  NAND2_X1 U6142 ( .A1(n7706), .A2(n7568), .ZN(n4496) );
  NAND2_X1 U6143 ( .A1(n4494), .A2(n4493), .ZN(n7663) );
  NAND3_X1 U6144 ( .A1(n6286), .A2(n5516), .A3(n5517), .ZN(n5519) );
  NAND2_X1 U6145 ( .A1(n7233), .A2(n4511), .ZN(n4507) );
  NOR2_X1 U6146 ( .A1(n7233), .A2(n4766), .ZN(n7267) );
  NAND3_X1 U6147 ( .A1(n4508), .A2(n4507), .A3(n4509), .ZN(n7235) );
  NAND3_X1 U6148 ( .A1(n4508), .A2(n4507), .A3(n4506), .ZN(n4510) );
  INV_X1 U6149 ( .A(n4510), .ZN(n7269) );
  XNOR2_X1 U6150 ( .A(n8077), .B(n8078), .ZN(n8042) );
  NAND2_X1 U6151 ( .A1(n7313), .A2(n4339), .ZN(n4537) );
  AND2_X2 U6152 ( .A1(n7603), .A2(n8455), .ZN(n5343) );
  NAND2_X1 U6153 ( .A1(n10069), .A2(n4320), .ZN(n4545) );
  NAND3_X1 U6154 ( .A1(n6721), .A2(n7792), .A3(n7926), .ZN(n4552) );
  NAND2_X1 U6155 ( .A1(n5500), .A2(n4556), .ZN(n5573) );
  AND2_X1 U6156 ( .A1(n4916), .A2(n4561), .ZN(n4559) );
  NAND4_X1 U6157 ( .A1(n4561), .A2(n4916), .A3(n5197), .A4(n4558), .ZN(n4862)
         );
  NAND3_X1 U6158 ( .A1(n4563), .A2(n6669), .A3(n4562), .ZN(n6670) );
  NAND2_X1 U6159 ( .A1(n6624), .A2(n6668), .ZN(n4562) );
  NAND2_X1 U6160 ( .A1(n6668), .A2(n6623), .ZN(n4563) );
  INV_X1 U6161 ( .A(n6668), .ZN(n4564) );
  INV_X1 U6162 ( .A(n4906), .ZN(n4567) );
  INV_X1 U6163 ( .A(n5960), .ZN(n4569) );
  AND2_X2 U6164 ( .A1(n5594), .A2(n4380), .ZN(n4871) );
  AND4_X2 U6165 ( .A1(n5590), .A2(n5591), .A3(n5592), .A4(n5593), .ZN(n5594)
         );
  NAND2_X2 U6166 ( .A1(n7618), .A2(n6138), .ZN(n5687) );
  NAND2_X4 U6167 ( .A1(n5652), .A2(n6243), .ZN(n7618) );
  NAND2_X1 U6168 ( .A1(n5653), .A2(n4572), .ZN(n5654) );
  AOI21_X1 U6169 ( .B1(n7437), .B2(n4581), .A(n4580), .ZN(n4579) );
  AOI21_X1 U6170 ( .B1(n4577), .B2(n4576), .A(n4573), .ZN(n5897) );
  NAND2_X1 U6171 ( .A1(n4580), .A2(n7505), .ZN(n4574) );
  NAND2_X1 U6172 ( .A1(n7437), .A2(n4377), .ZN(n4575) );
  NAND2_X1 U6173 ( .A1(n7512), .A2(n5919), .ZN(n5933) );
  NAND2_X1 U6174 ( .A1(n7512), .A2(n4387), .ZN(n4866) );
  NAND2_X1 U6175 ( .A1(n5626), .A2(n5623), .ZN(n5643) );
  NAND2_X1 U6176 ( .A1(n4586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U6177 ( .A1(n4586), .A2(n4583), .ZN(n4582) );
  INV_X1 U6178 ( .A(n4585), .ZN(n4584) );
  NAND2_X1 U6179 ( .A1(n5626), .A2(n4384), .ZN(n4586) );
  CLKBUF_X1 U6180 ( .A(n8482), .Z(n4587) );
  NAND2_X1 U6181 ( .A1(n8501), .A2(n4592), .ZN(n4591) );
  NOR2_X2 U6182 ( .A1(n8566), .A2(n8565), .ZN(n8564) );
  OAI211_X2 U6183 ( .C1(n6261), .C2(n5797), .A(n4335), .B(n4602), .ZN(n6874)
         );
  OR2_X1 U6184 ( .A1(n5704), .A2(n4461), .ZN(n4602) );
  NAND2_X1 U6185 ( .A1(n6752), .A2(n4300), .ZN(n8789) );
  NAND2_X1 U6186 ( .A1(n9316), .A2(n4606), .ZN(n4603) );
  NAND2_X1 U6187 ( .A1(n4603), .A2(n4604), .ZN(n9284) );
  NAND2_X1 U6188 ( .A1(n4609), .A2(n4611), .ZN(n9194) );
  NAND2_X1 U6189 ( .A1(n6803), .A2(n4382), .ZN(n4621) );
  NAND2_X1 U6190 ( .A1(n4627), .A2(n8799), .ZN(n4631) );
  INV_X1 U6191 ( .A(n8763), .ZN(n4627) );
  INV_X1 U6192 ( .A(n7402), .ZN(n4635) );
  NAND2_X1 U6193 ( .A1(n9387), .A2(n4340), .ZN(n4642) );
  AND3_X1 U6194 ( .A1(n9799), .A2(n9794), .A3(n9749), .ZN(n4644) );
  NAND2_X1 U6195 ( .A1(n4392), .A2(n4644), .ZN(n9731) );
  AND2_X1 U6196 ( .A1(n4392), .A2(n4645), .ZN(n9732) );
  AND2_X1 U6197 ( .A1(n9794), .A2(n9749), .ZN(n4645) );
  NAND2_X1 U6198 ( .A1(n4392), .A2(n9749), .ZN(n6857) );
  INV_X1 U6199 ( .A(n4646), .ZN(n7306) );
  INV_X1 U6200 ( .A(n4659), .ZN(n9240) );
  NAND2_X1 U6201 ( .A1(n7066), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U6202 ( .A1(n4671), .A2(n4669), .ZN(n7476) );
  NOR2_X2 U6203 ( .A1(n9138), .A2(n4677), .ZN(n4675) );
  NAND2_X1 U6204 ( .A1(n4679), .A2(n4678), .ZN(n9700) );
  AOI21_X1 U6205 ( .B1(n7025), .B2(n4681), .A(n4378), .ZN(n4678) );
  NAND2_X1 U6206 ( .A1(n9729), .A2(n4680), .ZN(n4679) );
  NAND2_X1 U6207 ( .A1(n9729), .A2(n9730), .ZN(n4682) );
  AND2_X1 U6208 ( .A1(n4871), .A2(n4372), .ZN(n4684) );
  NAND4_X1 U6209 ( .A1(n4871), .A2(n4372), .A3(n5798), .A4(n4683), .ZN(n5601)
         );
  NAND2_X1 U6210 ( .A1(n7476), .A2(n7475), .ZN(n9138) );
  NAND2_X1 U6211 ( .A1(n6801), .A2(n6800), .ZN(n6852) );
  INV_X1 U6212 ( .A(n6752), .ZN(n6773) );
  NAND2_X1 U6213 ( .A1(n6855), .A2(n6854), .ZN(n6991) );
  NAND2_X1 U6214 ( .A1(n4689), .A2(n8019), .ZN(n4690) );
  NAND2_X1 U6215 ( .A1(n8026), .A2(n8050), .ZN(n8034) );
  NOR2_X2 U6216 ( .A1(n8035), .A2(n8036), .ZN(n9964) );
  NAND2_X1 U6217 ( .A1(n6572), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4694) );
  OAI21_X1 U6218 ( .B1(n6572), .B2(P2_REG2_REG_2__SCAN_IN), .A(n4694), .ZN(
        n6453) );
  NAND2_X1 U6219 ( .A1(n6452), .A2(n6453), .ZN(n6563) );
  NAND2_X1 U6220 ( .A1(n5114), .A2(n5115), .ZN(n4962) );
  NAND2_X1 U6221 ( .A1(n5167), .A2(n5168), .ZN(n4700) );
  NAND2_X1 U6222 ( .A1(n5151), .A2(n5152), .ZN(n4701) );
  NAND2_X1 U6223 ( .A1(n5386), .A2(n4708), .ZN(n4707) );
  NAND2_X1 U6224 ( .A1(n5440), .A2(n4715), .ZN(n4714) );
  INV_X1 U6225 ( .A(n4719), .ZN(n5041) );
  NAND2_X1 U6226 ( .A1(n4752), .A2(n4753), .ZN(n5500) );
  INV_X1 U6227 ( .A(n4773), .ZN(n7080) );
  NOR2_X1 U6228 ( .A1(n9953), .A2(n4774), .ZN(n6905) );
  AND2_X1 U6229 ( .A1(n6903), .A2(n9942), .ZN(n4774) );
  AND2_X1 U6230 ( .A1(n6565), .A2(n4783), .ZN(n4780) );
  NOR2_X1 U6231 ( .A1(n9915), .A2(n6579), .ZN(n4784) );
  XNOR2_X1 U6232 ( .A(n8129), .B(n8130), .ZN(n8091) );
  OAI21_X1 U6233 ( .B1(n4786), .B2(n8091), .A(n4785), .ZN(n8142) );
  NAND2_X1 U6234 ( .A1(n7652), .A2(n4793), .ZN(n7706) );
  INV_X1 U6235 ( .A(n7714), .ZN(n4806) );
  NAND2_X1 U6236 ( .A1(n4809), .A2(n4811), .ZN(n7208) );
  NAND2_X1 U6237 ( .A1(n6710), .A2(n4818), .ZN(n6819) );
  NAND3_X1 U6238 ( .A1(n4908), .A2(n4388), .A3(n4290), .ZN(n5218) );
  NAND2_X1 U6239 ( .A1(n4821), .A2(n6240), .ZN(n6242) );
  NAND3_X1 U6240 ( .A1(n4331), .A2(n4823), .A3(n4822), .ZN(n4821) );
  NAND3_X1 U6241 ( .A1(n4331), .A2(n5581), .A3(n4823), .ZN(n6241) );
  NAND2_X1 U6242 ( .A1(n7178), .A2(n4828), .ZN(n4824) );
  NAND2_X1 U6243 ( .A1(n4824), .A2(n4825), .ZN(n7428) );
  NAND2_X1 U6244 ( .A1(n8320), .A2(n4385), .ZN(n8311) );
  NAND2_X1 U6245 ( .A1(n8216), .A2(n4835), .ZN(n4833) );
  NAND2_X1 U6246 ( .A1(n8216), .A2(n4840), .ZN(n4834) );
  CLKBUF_X1 U6247 ( .A(n4849), .Z(n4845) );
  INV_X1 U6248 ( .A(n4845), .ZN(n8270) );
  NAND2_X1 U6249 ( .A1(n7450), .A2(n4853), .ZN(n4852) );
  OAI22_X2 U6250 ( .A1(n6914), .A2(n4857), .B1(n7987), .B2(n4856), .ZN(n6983)
         );
  NAND2_X1 U6251 ( .A1(n5028), .A2(n4345), .ZN(n4921) );
  NAND2_X1 U6252 ( .A1(n4906), .A2(n5960), .ZN(n8598) );
  NAND2_X1 U6253 ( .A1(n4864), .A2(n4867), .ZN(n5956) );
  NAND2_X1 U6254 ( .A1(n5933), .A2(n5932), .ZN(n4867) );
  NAND2_X1 U6255 ( .A1(n4866), .A2(n4867), .ZN(n8469) );
  NAND2_X1 U6256 ( .A1(n9661), .A2(n5734), .ZN(n5752) );
  NAND2_X1 U6257 ( .A1(n9661), .A2(n4868), .ZN(n6922) );
  NAND2_X1 U6258 ( .A1(n8536), .A2(n6001), .ZN(n6018) );
  NAND2_X1 U6259 ( .A1(n8536), .A2(n4381), .ZN(n8574) );
  NAND2_X1 U6260 ( .A1(n8546), .A2(n4877), .ZN(n4875) );
  INV_X1 U6261 ( .A(n5777), .ZN(n9652) );
  NAND2_X1 U6262 ( .A1(n4878), .A2(n4879), .ZN(n5852) );
  NAND2_X1 U6263 ( .A1(n5777), .A2(n4352), .ZN(n4878) );
  NAND2_X1 U6264 ( .A1(n5557), .A2(n10074), .ZN(n5547) );
  NAND2_X1 U6265 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  INV_X1 U6266 ( .A(n8455), .ZN(n4938) );
  OAI21_X1 U6267 ( .B1(n9435), .B2(n9632), .A(n9434), .ZN(n9502) );
  XNOR2_X1 U6268 ( .A(n7958), .B(n8154), .ZN(n7965) );
  INV_X1 U6269 ( .A(n7763), .ZN(n5488) );
  AND3_X2 U6270 ( .A1(n5091), .A2(n5090), .A3(n5089), .ZN(n10018) );
  OR2_X1 U6271 ( .A1(n5025), .A2(n8452), .ZN(n5027) );
  NAND2_X1 U6272 ( .A1(n7211), .A2(n7342), .ZN(n7345) );
  OR2_X1 U6273 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  OAI21_X1 U6274 ( .B1(n7755), .B2(n7754), .A(n8395), .ZN(n7758) );
  NAND2_X1 U6275 ( .A1(n7347), .A2(n7346), .ZN(n7408) );
  NAND2_X2 U6276 ( .A1(n7765), .A2(n5489), .ZN(n5486) );
  NAND2_X1 U6277 ( .A1(n4921), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4923) );
  OAI21_X2 U6278 ( .B1(n7042), .B2(n5188), .A(n5187), .ZN(n7178) );
  INV_X1 U6279 ( .A(n5604), .ZN(n5606) );
  OAI22_X2 U6280 ( .A1(n8225), .A2(n5384), .B1(n8418), .B2(n8237), .ZN(n8216)
         );
  AND3_X2 U6281 ( .A1(n6592), .A2(n5556), .A3(n5555), .ZN(n10092) );
  INV_X1 U6282 ( .A(n7724), .ZN(n7727) );
  OR2_X1 U6283 ( .A1(n10074), .A2(n5467), .ZN(n4895) );
  OR2_X1 U6284 ( .A1(n8181), .A2(n8450), .ZN(n4896) );
  INV_X1 U6285 ( .A(n7987), .ZN(n5123) );
  AND2_X1 U6286 ( .A1(n6564), .A2(n9888), .ZN(n4897) );
  OR2_X1 U6287 ( .A1(n9507), .A2(n8594), .ZN(n4898) );
  OR2_X1 U6288 ( .A1(n8181), .A2(n8394), .ZN(n4899) );
  OR2_X1 U6289 ( .A1(n8171), .A2(n8394), .ZN(n4900) );
  AND2_X1 U6290 ( .A1(n4896), .A2(n4895), .ZN(n4901) );
  NOR2_X1 U6291 ( .A1(n5378), .A2(n5097), .ZN(n4902) );
  OR2_X1 U6292 ( .A1(n9356), .A2(n9150), .ZN(n4903) );
  INV_X1 U6293 ( .A(n8329), .ZN(n9993) );
  INV_X1 U6294 ( .A(n7783), .ZN(n5490) );
  OR2_X1 U6295 ( .A1(n5852), .A2(n5851), .ZN(n4904) );
  AND2_X1 U6296 ( .A1(n5559), .A2(n5558), .ZN(n4905) );
  INV_X2 U6297 ( .A(n9394), .ZN(n9758) );
  NOR2_X1 U6298 ( .A1(n7966), .A2(n7907), .ZN(n7904) );
  AOI21_X1 U6299 ( .B1(n7912), .B2(n7911), .A(n7910), .ZN(n7913) );
  INV_X1 U6300 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9111) );
  AND2_X1 U6301 ( .A1(n7576), .A2(n8218), .ZN(n7577) );
  INV_X1 U6302 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5595) );
  NOR2_X1 U6303 ( .A1(n8484), .A2(n8483), .ZN(n6100) );
  AND4_X1 U6304 ( .A1(n5597), .A2(n5596), .A3(n6205), .A4(n5647), .ZN(n5598)
         );
  AOI21_X1 U6305 ( .B1(n5539), .B2(n7014), .A(n6514), .ZN(n6515) );
  INV_X1 U6306 ( .A(n5413), .ZN(n5412) );
  INV_X1 U6307 ( .A(n5449), .ZN(n5448) );
  OR2_X1 U6308 ( .A1(n7692), .A2(n7974), .ZN(n5333) );
  INV_X1 U6309 ( .A(n5277), .ZN(n4933) );
  OR2_X1 U6310 ( .A1(n6103), .A2(n8481), .ZN(n6106) );
  INV_X2 U6311 ( .A(n6139), .ZN(n6097) );
  NOR2_X1 U6312 ( .A1(n6044), .A2(n6043), .ZN(n6060) );
  AND2_X1 U6313 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  NAND2_X1 U6314 ( .A1(n9284), .A2(n9295), .ZN(n9283) );
  NOR2_X1 U6315 ( .A1(n5881), .A2(n5878), .ZN(n5903) );
  INV_X1 U6316 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5599) );
  INV_X1 U6317 ( .A(n5229), .ZN(n4992) );
  INV_X1 U6318 ( .A(SI_8_), .ZN(n4973) );
  INV_X1 U6319 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5029) );
  INV_X1 U6320 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n4924) );
  NAND2_X1 U6321 ( .A1(n5412), .A2(n5411), .ZN(n5430) );
  OR2_X1 U6322 ( .A1(n5078), .A2(n6793), .ZN(n5057) );
  NAND2_X1 U6323 ( .A1(n5448), .A2(n5447), .ZN(n5463) );
  NAND2_X1 U6324 ( .A1(n4934), .A2(n9097), .ZN(n5310) );
  OR2_X1 U6325 ( .A1(n6829), .A2(n10034), .ZN(n5140) );
  INV_X1 U6326 ( .A(n5486), .ZN(n5487) );
  XNOR2_X1 U6327 ( .A(n5092), .B(n10018), .ZN(n7929) );
  AND2_X1 U6328 ( .A1(n6060), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6077) );
  AND2_X1 U6329 ( .A1(n6106), .A2(n6105), .ZN(n6107) );
  INV_X1 U6330 ( .A(n8597), .ZN(n5959) );
  OR2_X1 U6331 ( .A1(n5816), .A2(n5805), .ZN(n5842) );
  AOI21_X1 U6332 ( .B1(n9200), .B2(n9199), .A(n9198), .ZN(n9201) );
  OR2_X1 U6333 ( .A1(n6025), .A2(n6024), .ZN(n6044) );
  OR2_X1 U6334 ( .A1(n5945), .A2(n5944), .ZN(n5964) );
  OR2_X1 U6335 ( .A1(n5842), .A2(n5841), .ZN(n5881) );
  OAI21_X1 U6336 ( .B1(n9736), .B2(n6776), .A(n8791), .ZN(n6754) );
  AND2_X1 U6337 ( .A1(n9433), .A2(n9432), .ZN(n9434) );
  INV_X1 U6338 ( .A(n6281), .ZN(n6020) );
  OR2_X1 U6339 ( .A1(n9731), .A2(n9656), .ZN(n9714) );
  INV_X1 U6340 ( .A(n6784), .ZN(n6785) );
  NAND2_X1 U6341 ( .A1(n4994), .A2(SI_12_), .ZN(n4995) );
  NAND2_X1 U6342 ( .A1(n4979), .A2(n4978), .ZN(n4982) );
  NAND2_X1 U6343 ( .A1(n5340), .A2(n5339), .ZN(n5359) );
  INV_X1 U6344 ( .A(n7986), .ZN(n7119) );
  INV_X1 U6345 ( .A(n8154), .ZN(n7957) );
  INV_X1 U6346 ( .A(n9928), .ZN(n6565) );
  INV_X1 U6347 ( .A(n9951), .ZN(n9974) );
  NAND2_X1 U6348 ( .A1(n7885), .A2(n7886), .ZN(n8209) );
  NAND2_X1 U6349 ( .A1(n5488), .A2(n5487), .ZN(n6678) );
  AND2_X1 U6350 ( .A1(n7903), .A2(n5552), .ZN(n6593) );
  INV_X1 U6351 ( .A(n7981), .ZN(n7826) );
  AND2_X1 U6352 ( .A1(n7790), .A2(n7782), .ZN(n7926) );
  NOR2_X1 U6353 ( .A1(n10010), .A2(n10046), .ZN(n10061) );
  AND2_X1 U6354 ( .A1(n5755), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5778) );
  AND2_X1 U6355 ( .A1(n6162), .A2(n6161), .ZN(n6180) );
  OR2_X1 U6356 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  OR2_X1 U6357 ( .A1(n6111), .A2(n8550), .ZN(n6129) );
  AND2_X1 U6358 ( .A1(n6099), .A2(n6098), .ZN(n8483) );
  OR2_X1 U6359 ( .A1(n6235), .A2(n6231), .ZN(n9660) );
  NOR2_X1 U6360 ( .A1(n8925), .A2(n8924), .ZN(n8933) );
  NAND2_X1 U6361 ( .A1(n9149), .A2(n4903), .ZN(n9152) );
  AND2_X1 U6362 ( .A1(n9367), .A2(n9366), .ZN(n9386) );
  NAND2_X1 U6363 ( .A1(n7295), .A2(n8652), .ZN(n7378) );
  OR2_X1 U6364 ( .A1(n9758), .A2(n6765), .ZN(n9744) );
  INV_X1 U6365 ( .A(n9738), .ZN(n9706) );
  AND2_X1 U6366 ( .A1(n5422), .A2(n5408), .ZN(n5420) );
  NAND2_X1 U6367 ( .A1(n4991), .A2(n4990), .ZN(n5216) );
  NAND2_X2 U6368 ( .A1(n6423), .A2(n6449), .ZN(n6246) );
  NAND2_X1 U6369 ( .A1(n4925), .A2(n9081), .ZN(n5142) );
  OR2_X1 U6370 ( .A1(n5142), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5158) );
  AND3_X1 U6371 ( .A1(n5363), .A2(n5362), .A3(n5361), .ZN(n8247) );
  INV_X1 U6372 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6973) );
  INV_X1 U6373 ( .A(n9917), .ZN(n9970) );
  INV_X1 U6374 ( .A(n9924), .ZN(n9959) );
  AND2_X1 U6375 ( .A1(n7312), .A2(n7811), .ZN(n7933) );
  AND2_X1 U6376 ( .A1(n7907), .A2(n6518), .ZN(n9984) );
  NAND2_X1 U6377 ( .A1(n10090), .A2(n6239), .ZN(n6240) );
  AND3_X1 U6378 ( .A1(n6497), .A2(n5550), .A3(n5549), .ZN(n6592) );
  NOR2_X1 U6379 ( .A1(n10074), .A2(n5481), .ZN(n5586) );
  NAND2_X1 U6380 ( .A1(n7762), .A2(n7761), .ZN(n10054) );
  INV_X1 U6381 ( .A(n10061), .ZN(n10068) );
  AND2_X1 U6382 ( .A1(n5531), .A2(n5530), .ZN(n6268) );
  INV_X1 U6383 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6205) );
  OR2_X1 U6384 ( .A1(n6181), .A2(n6180), .ZN(n6182) );
  INV_X1 U6385 ( .A(n8594), .ZN(n9670) );
  OR2_X1 U6386 ( .A1(n9681), .A2(n8873), .ZN(n8960) );
  INV_X1 U6387 ( .A(n9691), .ZN(n8975) );
  INV_X1 U6388 ( .A(n9403), .ZN(n9750) );
  INV_X1 U6389 ( .A(n9415), .ZN(n9755) );
  INV_X1 U6390 ( .A(n9413), .ZN(n9754) );
  AND2_X1 U6391 ( .A1(n6188), .A2(n9544), .ZN(n6761) );
  INV_X1 U6392 ( .A(n9632), .ZN(n9850) );
  XNOR2_X1 U6393 ( .A(n4970), .B(SI_7_), .ZN(n5168) );
  XNOR2_X1 U6394 ( .A(n4967), .B(SI_6_), .ZN(n5152) );
  XNOR2_X1 U6395 ( .A(n4953), .B(SI_2_), .ZN(n5085) );
  AND2_X1 U6396 ( .A1(n6489), .A2(n6488), .ZN(n7724) );
  NAND2_X1 U6397 ( .A1(n5470), .A2(n5469), .ZN(n7967) );
  INV_X1 U6398 ( .A(n9914), .ZN(n9980) );
  OR2_X1 U6399 ( .A1(n6438), .A2(n9882), .ZN(n9965) );
  INV_X1 U6400 ( .A(n5583), .ZN(n8177) );
  NAND2_X1 U6401 ( .A1(n6596), .A2(n6595), .ZN(n8329) );
  NAND2_X1 U6402 ( .A1(n10092), .A2(n10073), .ZN(n8394) );
  INV_X1 U6403 ( .A(n10092), .ZN(n10090) );
  NOR2_X1 U6404 ( .A1(n5585), .A2(n5586), .ZN(n5587) );
  INV_X1 U6405 ( .A(n7547), .ZN(n8446) );
  AND2_X1 U6406 ( .A1(n5546), .A2(n5545), .ZN(n10076) );
  AND2_X1 U6407 ( .A1(n6496), .A2(n5538), .ZN(n6284) );
  INV_X1 U6408 ( .A(n7962), .ZN(n7761) );
  INV_X1 U6409 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6622) );
  INV_X1 U6410 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6275) );
  AND2_X1 U6411 ( .A1(n6216), .A2(n6215), .ZN(n9674) );
  AND2_X1 U6412 ( .A1(n6236), .A2(n9741), .ZN(n8594) );
  OR2_X1 U6413 ( .A1(n9681), .A2(n6300), .ZN(n9689) );
  AND2_X1 U6414 ( .A1(n7161), .A2(n7160), .ZN(n9837) );
  OR2_X1 U6415 ( .A1(n9758), .A2(n6781), .ZN(n9415) );
  INV_X1 U6416 ( .A(n9257), .ZN(n9514) );
  AND2_X1 U6417 ( .A1(n9837), .A2(n9836), .ZN(n9874) );
  INV_X1 U6418 ( .A(n9862), .ZN(n9860) );
  INV_X1 U6419 ( .A(n9763), .ZN(n9764) );
  AND2_X1 U6420 ( .A1(n8877), .A2(n6271), .ZN(n9763) );
  INV_X1 U6421 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6406) );
  INV_X1 U6422 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6250) );
  NOR2_X1 U6423 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  AND2_X1 U6424 ( .A1(n6424), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3893) );
  NAND2_X1 U6425 ( .A1(n5547), .A2(n4901), .ZN(P2_U3455) );
  NOR2_X1 U6426 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4913) );
  NOR2_X1 U6427 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4912) );
  NOR2_X1 U6428 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n4911) );
  NAND4_X1 U6429 ( .A1(n4913), .A2(n4912), .A3(n4911), .A4(n9111), .ZN(n4915)
         );
  NAND3_X1 U6430 ( .A1(n5034), .A2(n5036), .A3(n5032), .ZN(n4914) );
  NAND2_X1 U6431 ( .A1(n5509), .A2(n9109), .ZN(n4917) );
  INV_X1 U6432 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4918) );
  INV_X1 U6433 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4919) );
  INV_X1 U6434 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4922) );
  XNOR2_X2 U6435 ( .A(n4923), .B(n4922), .ZN(n8455) );
  INV_X1 U6436 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7273) );
  INV_X1 U6437 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n4930) );
  INV_X1 U6438 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4932) );
  INV_X1 U6439 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9097) );
  INV_X1 U6440 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4935) );
  NAND2_X1 U6441 ( .A1(n5049), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6442 ( .A1(n5328), .A2(n4937), .ZN(n8276) );
  NAND2_X1 U6443 ( .A1(n5069), .A2(n8276), .ZN(n4944) );
  NAND2_X2 U6444 ( .A1(n7603), .A2(n4938), .ZN(n5378) );
  INV_X1 U6445 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8375) );
  OR2_X1 U6446 ( .A1(n5378), .A2(n8375), .ZN(n4943) );
  INV_X1 U6447 ( .A(n7603), .ZN(n4939) );
  INV_X1 U6448 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n4940) );
  OR2_X1 U6449 ( .A1(n5078), .A2(n4940), .ZN(n4942) );
  INV_X1 U6450 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8432) );
  OR2_X1 U6451 ( .A1(n6844), .A2(n8432), .ZN(n4941) );
  INV_X1 U6452 ( .A(n5060), .ZN(n4949) );
  NAND2_X1 U6453 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4948) );
  AND2_X1 U6454 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4947) );
  NAND2_X1 U6455 ( .A1(n6249), .A2(n4947), .ZN(n5668) );
  OAI21_X1 U6456 ( .B1(n6249), .B2(n4948), .A(n5668), .ZN(n5059) );
  NAND2_X1 U6457 ( .A1(n4949), .A2(n5059), .ZN(n4952) );
  NAND2_X1 U6458 ( .A1(n4950), .A2(SI_1_), .ZN(n4951) );
  INV_X1 U6459 ( .A(n4953), .ZN(n4954) );
  NAND2_X1 U6460 ( .A1(n4954), .A2(SI_2_), .ZN(n4955) );
  MUX2_X1 U6461 ( .A(n6257), .B(n6252), .S(n6249), .Z(n4956) );
  INV_X1 U6462 ( .A(n4956), .ZN(n4957) );
  NAND2_X1 U6463 ( .A1(n4957), .A2(SI_3_), .ZN(n4958) );
  MUX2_X1 U6464 ( .A(n6255), .B(n9102), .S(n6249), .Z(n4959) );
  INV_X1 U6465 ( .A(n4959), .ZN(n4960) );
  NAND2_X1 U6466 ( .A1(n4960), .A2(SI_4_), .ZN(n4961) );
  MUX2_X1 U6467 ( .A(n6260), .B(n6258), .S(n6249), .Z(n4963) );
  INV_X1 U6468 ( .A(n4963), .ZN(n4964) );
  NAND2_X1 U6469 ( .A1(n4964), .A2(SI_5_), .ZN(n4965) );
  MUX2_X1 U6470 ( .A(n6264), .B(n6262), .S(n6249), .Z(n4967) );
  INV_X1 U6471 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6472 ( .A1(n4968), .A2(SI_6_), .ZN(n4969) );
  MUX2_X1 U6473 ( .A(n6265), .B(n6266), .S(n7747), .Z(n4970) );
  INV_X1 U6474 ( .A(n4970), .ZN(n4971) );
  NAND2_X1 U6475 ( .A1(n4971), .A2(SI_7_), .ZN(n4972) );
  MUX2_X1 U6476 ( .A(n6275), .B(n6276), .S(n7747), .Z(n4974) );
  INV_X1 U6477 ( .A(n4974), .ZN(n4975) );
  NAND2_X1 U6478 ( .A1(n4975), .A2(SI_8_), .ZN(n4976) );
  MUX2_X1 U6479 ( .A(n6289), .B(n6290), .S(n7747), .Z(n4979) );
  INV_X1 U6480 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6481 ( .A1(n4980), .A2(SI_9_), .ZN(n4981) );
  MUX2_X1 U6482 ( .A(n6295), .B(n6296), .S(n7747), .Z(n4984) );
  INV_X1 U6483 ( .A(n4984), .ZN(n4985) );
  MUX2_X1 U6484 ( .A(n9103), .B(n6376), .S(n7747), .Z(n4988) );
  INV_X1 U6485 ( .A(SI_11_), .ZN(n4987) );
  INV_X1 U6486 ( .A(n4988), .ZN(n4989) );
  NAND2_X1 U6487 ( .A1(n4989), .A2(SI_11_), .ZN(n4990) );
  MUX2_X1 U6488 ( .A(n6404), .B(n6406), .S(n7747), .Z(n4993) );
  INV_X1 U6489 ( .A(n4993), .ZN(n4994) );
  MUX2_X1 U6490 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7747), .Z(n4997) );
  NAND2_X1 U6491 ( .A1(n4997), .A2(SI_13_), .ZN(n4998) );
  INV_X1 U6492 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6620) );
  MUX2_X1 U6493 ( .A(n6622), .B(n6620), .S(n7747), .Z(n5000) );
  INV_X1 U6494 ( .A(SI_14_), .ZN(n4999) );
  INV_X1 U6495 ( .A(n5000), .ZN(n5001) );
  NAND2_X1 U6496 ( .A1(n5001), .A2(SI_14_), .ZN(n5002) );
  INV_X1 U6497 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6677) );
  INV_X1 U6498 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6701) );
  MUX2_X1 U6499 ( .A(n6677), .B(n6701), .S(n7747), .Z(n5004) );
  INV_X1 U6500 ( .A(n5004), .ZN(n5005) );
  NAND2_X1 U6501 ( .A1(n5005), .A2(SI_15_), .ZN(n5006) );
  MUX2_X1 U6502 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7747), .Z(n5009) );
  XNOR2_X1 U6503 ( .A(n5009), .B(SI_16_), .ZN(n5284) );
  NAND2_X1 U6504 ( .A1(n5009), .A2(SI_16_), .ZN(n5010) );
  INV_X1 U6505 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6751) );
  INV_X1 U6506 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6749) );
  MUX2_X1 U6507 ( .A(n6751), .B(n6749), .S(n7747), .Z(n5012) );
  INV_X1 U6508 ( .A(SI_17_), .ZN(n5011) );
  INV_X1 U6509 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6510 ( .A1(n5013), .A2(SI_17_), .ZN(n5014) );
  NAND2_X1 U6511 ( .A1(n5015), .A2(n5014), .ZN(n5302) );
  INV_X1 U6512 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6933) );
  INV_X1 U6513 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5016) );
  MUX2_X1 U6514 ( .A(n6933), .B(n5016), .S(n7747), .Z(n5017) );
  XNOR2_X1 U6515 ( .A(n5017), .B(SI_18_), .ZN(n5040) );
  INV_X1 U6516 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6517 ( .A1(n5018), .A2(SI_18_), .ZN(n5019) );
  INV_X1 U6518 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6949) );
  INV_X1 U6519 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6947) );
  MUX2_X1 U6520 ( .A(n6949), .B(n6947), .S(n7747), .Z(n5022) );
  INV_X1 U6521 ( .A(SI_19_), .ZN(n5021) );
  NAND2_X1 U6522 ( .A1(n5022), .A2(n5021), .ZN(n5317) );
  INV_X1 U6523 ( .A(n5022), .ZN(n5023) );
  NAND2_X1 U6524 ( .A1(n5023), .A2(SI_19_), .ZN(n5024) );
  NAND2_X1 U6525 ( .A1(n5317), .A2(n5024), .ZN(n5318) );
  XNOR2_X1 U6526 ( .A(n5319), .B(n5318), .ZN(n6946) );
  XNOR2_X2 U6527 ( .A(n5027), .B(n5026), .ZN(n6423) );
  XNOR2_X2 U6528 ( .A(n5030), .B(n5029), .ZN(n6449) );
  NAND2_X1 U6529 ( .A1(n6246), .A2(n5642), .ZN(n5086) );
  NAND2_X1 U6530 ( .A1(n6946), .A2(n7753), .ZN(n5039) );
  NAND2_X1 U6531 ( .A1(n6246), .A2(n7747), .ZN(n5058) );
  NOR2_X1 U6532 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n5033) );
  INV_X1 U6533 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5035) );
  NAND2_X1 U6534 ( .A1(n5042), .A2(n5035), .ZN(n5471) );
  NAND2_X1 U6535 ( .A1(n5471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5037) );
  INV_X1 U6536 ( .A(n6246), .ZN(n5088) );
  AOI22_X1 U6537 ( .A1(n7752), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7957), .B2(
        n5305), .ZN(n5038) );
  XNOR2_X1 U6538 ( .A(n5041), .B(n5040), .ZN(n6825) );
  NAND2_X1 U6539 ( .A1(n6825), .A2(n7753), .ZN(n5047) );
  INV_X1 U6540 ( .A(n5042), .ZN(n5043) );
  NAND2_X1 U6541 ( .A1(n5043), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5044) );
  MUX2_X1 U6542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5044), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5045) );
  NAND2_X1 U6543 ( .A1(n5045), .A2(n5471), .ZN(n8150) );
  INV_X1 U6544 ( .A(n8150), .ZN(n8124) );
  AOI22_X1 U6545 ( .A1(n7752), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5305), .B2(
        n8124), .ZN(n5046) );
  NAND2_X1 U6546 ( .A1(n6839), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5053) );
  INV_X1 U6547 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8436) );
  OR2_X1 U6548 ( .A1(n6844), .A2(n8436), .ZN(n5052) );
  NAND2_X1 U6549 ( .A1(n5310), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5048) );
  AND2_X1 U6550 ( .A1(n5049), .A2(n5048), .ZN(n8288) );
  OR2_X1 U6551 ( .A1(n8288), .A2(n5076), .ZN(n5051) );
  INV_X1 U6552 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8379) );
  OR2_X1 U6553 ( .A1(n5378), .A2(n8379), .ZN(n5050) );
  INV_X1 U6554 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U6555 ( .A1(n5065), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5056) );
  INV_X1 U6556 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6427) );
  OR2_X1 U6557 ( .A1(n5076), .A2(n6427), .ZN(n5054) );
  AND4_X2 U6558 ( .A1(n5057), .A2(n5056), .A3(n5055), .A4(n5054), .ZN(n5073)
         );
  INV_X1 U6559 ( .A(n5073), .ZN(n6492) );
  OR2_X1 U6560 ( .A1(n5058), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U6561 ( .A(n5060), .B(n5059), .ZN(n5641) );
  OR2_X1 U6562 ( .A1(n5086), .A2(n5641), .ZN(n5063) );
  NAND2_X1 U6563 ( .A1(n5088), .A2(n6435), .ZN(n5062) );
  NAND3_X1 U6564 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n5061) );
  NAND2_X1 U6565 ( .A1(n6492), .A2(n5061), .ZN(n7765) );
  AND3_X2 U6566 ( .A1(n5064), .A2(n5063), .A3(n5062), .ZN(n6794) );
  INV_X1 U6567 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9096) );
  INV_X1 U6568 ( .A(n5378), .ZN(n5065) );
  NAND2_X1 U6569 ( .A1(n5065), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5066) );
  OAI21_X1 U6570 ( .B1(n9096), .B2(n5078), .A(n5066), .ZN(n5067) );
  NOR2_X1 U6571 ( .A1(n5068), .A2(n5067), .ZN(n5071) );
  INV_X1 U6572 ( .A(n5076), .ZN(n5069) );
  NAND2_X1 U6573 ( .A1(n5069), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5070) );
  NAND2_X1 U6574 ( .A1(n5642), .A2(SI_0_), .ZN(n5072) );
  XNOR2_X1 U6575 ( .A(n5072), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8468) );
  MUX2_X1 U6576 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8468), .S(n6246), .Z(n6483) );
  NAND2_X1 U6577 ( .A1(n7989), .A2(n6483), .ZN(n6680) );
  NAND2_X1 U6578 ( .A1(n5486), .A2(n6680), .ZN(n5075) );
  NAND2_X1 U6579 ( .A1(n10006), .A2(n5061), .ZN(n5074) );
  NAND2_X1 U6580 ( .A1(n5075), .A2(n5074), .ZN(n10004) );
  NAND2_X1 U6581 ( .A1(n5343), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5083) );
  INV_X1 U6582 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6571) );
  OR2_X1 U6583 ( .A1(n5378), .A2(n6571), .ZN(n5081) );
  INV_X1 U6584 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10001) );
  OR2_X1 U6585 ( .A1(n5076), .A2(n10001), .ZN(n5080) );
  INV_X1 U6586 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5077) );
  OR2_X1 U6587 ( .A1(n7739), .A2(n6248), .ZN(n5091) );
  XNOR2_X1 U6588 ( .A(n5084), .B(n5085), .ZN(n6251) );
  OR2_X1 U6589 ( .A1(n5086), .A2(n6251), .ZN(n5090) );
  NAND2_X1 U6590 ( .A1(n5088), .A2(n4295), .ZN(n5089) );
  NAND2_X1 U6591 ( .A1(n10004), .A2(n7929), .ZN(n5094) );
  NAND2_X1 U6592 ( .A1(n6641), .A2(n10018), .ZN(n5093) );
  NAND2_X1 U6593 ( .A1(n6839), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U6594 ( .A1(n5343), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5096) );
  INV_X1 U6595 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6596 ( .A1(n5101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  OR2_X1 U6597 ( .A1(n7739), .A2(n6257), .ZN(n5106) );
  XNOR2_X1 U6598 ( .A(n5103), .B(n5104), .ZN(n6256) );
  NOR2_X1 U6599 ( .A1(n7988), .A2(n6726), .ZN(n5108) );
  NAND2_X1 U6600 ( .A1(n7988), .A2(n6726), .ZN(n5107) );
  OAI21_X2 U6601 ( .B1(n6719), .B2(n5108), .A(n5107), .ZN(n6914) );
  NAND2_X1 U6602 ( .A1(n6839), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6603 ( .A1(n5343), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6604 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5109) );
  AND2_X1 U6605 ( .A1(n5125), .A2(n5109), .ZN(n6715) );
  OR2_X1 U6606 ( .A1(n5076), .A2(n6715), .ZN(n5111) );
  INV_X1 U6607 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6579) );
  OR2_X1 U6608 ( .A1(n5378), .A2(n6579), .ZN(n5110) );
  NAND4_X1 U6609 ( .A1(n5113), .A2(n5112), .A3(n5111), .A4(n5110), .ZN(n7987)
         );
  XNOR2_X1 U6610 ( .A(n5114), .B(n5115), .ZN(n6254) );
  OR2_X1 U6611 ( .A1(n5169), .A2(n6254), .ZN(n5122) );
  NAND2_X1 U6612 ( .A1(n5117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5116) );
  MUX2_X1 U6613 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5116), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5119) );
  INV_X1 U6614 ( .A(n5133), .ZN(n5118) );
  NAND2_X1 U6615 ( .A1(n5305), .A2(n9915), .ZN(n5120) );
  NAND2_X1 U6616 ( .A1(n6840), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5130) );
  NAND2_X1 U6617 ( .A1(n5343), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5129) );
  INV_X1 U6618 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5124) );
  OR2_X1 U6619 ( .A1(n5078), .A2(n5124), .ZN(n5128) );
  NAND2_X1 U6620 ( .A1(n5125), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5126) );
  AND2_X1 U6621 ( .A1(n5142), .A2(n5126), .ZN(n6982) );
  OR2_X1 U6622 ( .A1(n5076), .A2(n6982), .ZN(n5127) );
  NAND4_X1 U6623 ( .A1(n5130), .A2(n5129), .A3(n5128), .A4(n5127), .ZN(n9983)
         );
  NOR2_X1 U6624 ( .A1(n5133), .A2(n8452), .ZN(n5131) );
  MUX2_X1 U6625 ( .A(n8452), .B(n5131), .S(P2_IR_REG_5__SCAN_IN), .Z(n5135) );
  NAND2_X1 U6626 ( .A1(n5133), .A2(n5132), .ZN(n5164) );
  INV_X1 U6627 ( .A(n5164), .ZN(n5134) );
  XNOR2_X1 U6628 ( .A(n5136), .B(n5137), .ZN(n6259) );
  OR2_X1 U6629 ( .A1(n5169), .A2(n6259), .ZN(n5139) );
  OR2_X1 U6630 ( .A1(n7739), .A2(n6260), .ZN(n5138) );
  OAI211_X1 U6631 ( .C1(n6246), .C2(n9928), .A(n5139), .B(n5138), .ZN(n6822)
         );
  NOR2_X1 U6632 ( .A1(n9983), .A2(n6822), .ZN(n5141) );
  INV_X1 U6633 ( .A(n9983), .ZN(n6829) );
  INV_X1 U6634 ( .A(n6822), .ZN(n10034) );
  NAND2_X1 U6635 ( .A1(n6840), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5148) );
  NAND2_X1 U6636 ( .A1(n6839), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6637 ( .A1(n5142), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5143) );
  AND2_X1 U6638 ( .A1(n5158), .A2(n5143), .ZN(n9992) );
  OR2_X1 U6639 ( .A1(n5076), .A2(n9992), .ZN(n5146) );
  INV_X1 U6640 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6641 ( .A1(n6844), .A2(n5144), .ZN(n5145) );
  NAND4_X1 U6642 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n7986)
         );
  NAND2_X1 U6643 ( .A1(n5164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5150) );
  XNOR2_X1 U6644 ( .A(n5150), .B(n5149), .ZN(n6900) );
  XNOR2_X1 U6645 ( .A(n5151), .B(n5152), .ZN(n6263) );
  OR2_X1 U6646 ( .A1(n5169), .A2(n6263), .ZN(n5154) );
  OR2_X1 U6647 ( .A1(n5460), .A2(n6264), .ZN(n5153) );
  OAI211_X1 U6648 ( .C1(n6246), .C2(n6900), .A(n5154), .B(n5153), .ZN(n10039)
         );
  AND2_X1 U6649 ( .A1(n7986), .A2(n10039), .ZN(n5156) );
  INV_X1 U6650 ( .A(n10039), .ZN(n6834) );
  NAND2_X1 U6651 ( .A1(n7119), .A2(n6834), .ZN(n5155) );
  OAI21_X2 U6652 ( .B1(n9981), .B2(n5156), .A(n5155), .ZN(n7118) );
  NAND2_X1 U6653 ( .A1(n5343), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5163) );
  INV_X1 U6654 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6655 ( .A1(n5378), .A2(n5157), .ZN(n5162) );
  INV_X1 U6656 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6890) );
  OR2_X1 U6657 ( .A1(n5078), .A2(n6890), .ZN(n5161) );
  NAND2_X1 U6658 ( .A1(n5158), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5159) );
  AND2_X1 U6659 ( .A1(n5174), .A2(n5159), .ZN(n7123) );
  OR2_X1 U6660 ( .A1(n5076), .A2(n7123), .ZN(n5160) );
  NAND2_X1 U6661 ( .A1(n5181), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6662 ( .A(n5166), .B(n5165), .ZN(n9942) );
  XNOR2_X1 U6663 ( .A(n5167), .B(n5168), .ZN(n6267) );
  OR2_X1 U6664 ( .A1(n5169), .A2(n6267), .ZN(n5171) );
  OR2_X1 U6665 ( .A1(n7739), .A2(n6265), .ZN(n5170) );
  OAI211_X1 U6666 ( .C1(n6246), .C2(n9942), .A(n5171), .B(n5170), .ZN(n7125)
         );
  NAND2_X1 U6667 ( .A1(n7129), .A2(n7125), .ZN(n7799) );
  INV_X1 U6668 ( .A(n7125), .ZN(n10043) );
  NAND2_X1 U6669 ( .A1(n9985), .A2(n10043), .ZN(n7045) );
  NAND2_X1 U6670 ( .A1(n7799), .A2(n7045), .ZN(n7804) );
  NAND2_X1 U6671 ( .A1(n7118), .A2(n7804), .ZN(n5173) );
  NAND2_X1 U6672 ( .A1(n7129), .A2(n10043), .ZN(n5172) );
  NAND2_X1 U6673 ( .A1(n6840), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6674 ( .A1(n6839), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6675 ( .A1(n5174), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5175) );
  AND2_X1 U6676 ( .A1(n5189), .A2(n5175), .ZN(n7047) );
  OR2_X1 U6677 ( .A1(n5076), .A2(n7047), .ZN(n5178) );
  INV_X1 U6678 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5176) );
  OR2_X1 U6679 ( .A1(n6844), .A2(n5176), .ZN(n5177) );
  OAI21_X1 U6680 ( .B1(n5181), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5182) );
  XNOR2_X1 U6681 ( .A(n5182), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7079) );
  AOI22_X1 U6682 ( .A1(n7752), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5305), .B2(
        n7079), .ZN(n5186) );
  XNOR2_X1 U6683 ( .A(n5183), .B(n5184), .ZN(n6274) );
  NAND2_X1 U6684 ( .A1(n6274), .A2(n7753), .ZN(n5185) );
  NOR2_X1 U6685 ( .A1(n7985), .A2(n7139), .ZN(n5188) );
  NAND2_X1 U6686 ( .A1(n7985), .A2(n7139), .ZN(n5187) );
  NAND2_X1 U6687 ( .A1(n6840), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U6688 ( .A1(n5343), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5193) );
  NAND2_X1 U6689 ( .A1(n5189), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5190) );
  AND2_X1 U6690 ( .A1(n5209), .A2(n5190), .ZN(n7183) );
  OR2_X1 U6691 ( .A1(n5076), .A2(n7183), .ZN(n5192) );
  INV_X1 U6692 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7094) );
  OR2_X1 U6693 ( .A1(n5078), .A2(n7094), .ZN(n5191) );
  NAND4_X1 U6694 ( .A1(n5194), .A2(n5193), .A3(n5192), .A4(n5191), .ZN(n7984)
         );
  XNOR2_X1 U6695 ( .A(n5196), .B(n5195), .ZN(n6288) );
  NAND2_X1 U6696 ( .A1(n6288), .A2(n7753), .ZN(n5202) );
  NOR2_X1 U6697 ( .A1(n5197), .A2(n8452), .ZN(n5198) );
  MUX2_X1 U6698 ( .A(n8452), .B(n5198), .S(P2_IR_REG_9__SCAN_IN), .Z(n5200) );
  OR2_X1 U6699 ( .A1(n5200), .A2(n5199), .ZN(n7082) );
  INV_X1 U6700 ( .A(n7082), .ZN(n7996) );
  AOI22_X1 U6701 ( .A1(n7752), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5305), .B2(
        n7996), .ZN(n5201) );
  NAND2_X1 U6702 ( .A1(n6294), .A2(n7753), .ZN(n5207) );
  OR2_X1 U6703 ( .A1(n5199), .A2(n8452), .ZN(n5205) );
  XNOR2_X1 U6704 ( .A(n5205), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7093) );
  AOI22_X1 U6705 ( .A1(n7752), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5305), .B2(
        n7093), .ZN(n5206) );
  NAND2_X1 U6706 ( .A1(n5207), .A2(n5206), .ZN(n7323) );
  INV_X1 U6707 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5208) );
  OR2_X1 U6708 ( .A1(n5378), .A2(n5208), .ZN(n5214) );
  NAND2_X1 U6709 ( .A1(n5343), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5213) );
  INV_X1 U6710 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7088) );
  OR2_X1 U6711 ( .A1(n5078), .A2(n7088), .ZN(n5212) );
  NAND2_X1 U6712 ( .A1(n5209), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5210) );
  AND2_X1 U6713 ( .A1(n5222), .A2(n5210), .ZN(n7321) );
  OR2_X1 U6714 ( .A1(n5076), .A2(n7321), .ZN(n5211) );
  NAND4_X1 U6715 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n7983)
         );
  NOR2_X1 U6716 ( .A1(n7323), .A2(n7983), .ZN(n5215) );
  INV_X1 U6717 ( .A(n7323), .ZN(n10055) );
  XNOR2_X1 U6718 ( .A(n5217), .B(n5216), .ZN(n6375) );
  NAND2_X1 U6719 ( .A1(n6375), .A2(n7753), .ZN(n5221) );
  NAND2_X1 U6720 ( .A1(n5218), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5219) );
  XNOR2_X1 U6721 ( .A(n5219), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7268) );
  AOI22_X1 U6722 ( .A1(n7752), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5305), .B2(
        n7268), .ZN(n5220) );
  NAND2_X1 U6723 ( .A1(n6840), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5227) );
  NAND2_X1 U6724 ( .A1(n5343), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5226) );
  INV_X1 U6725 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7433) );
  OR2_X1 U6726 ( .A1(n5078), .A2(n7433), .ZN(n5225) );
  NAND2_X1 U6727 ( .A1(n5222), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5223) );
  AND2_X1 U6728 ( .A1(n5235), .A2(n5223), .ZN(n7432) );
  OR2_X1 U6729 ( .A1(n5076), .A2(n7432), .ZN(n5224) );
  NAND4_X1 U6730 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n7982)
         );
  OR2_X1 U6731 ( .A1(n10065), .A2(n7982), .ZN(n5228) );
  NAND2_X1 U6732 ( .A1(n7428), .A2(n5228), .ZN(n7424) );
  NAND2_X1 U6733 ( .A1(n10065), .A2(n7982), .ZN(n7425) );
  NAND2_X1 U6734 ( .A1(n7424), .A2(n7425), .ZN(n7450) );
  XNOR2_X1 U6735 ( .A(n5230), .B(n5229), .ZN(n6403) );
  NAND2_X1 U6736 ( .A1(n6403), .A2(n7753), .ZN(n5234) );
  NAND2_X1 U6737 ( .A1(n5231), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5232) );
  XNOR2_X1 U6738 ( .A(n5232), .B(n4817), .ZN(n8023) );
  INV_X1 U6739 ( .A(n8023), .ZN(n7275) );
  AOI22_X1 U6740 ( .A1(n7752), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5305), .B2(
        n7275), .ZN(n5233) );
  NAND2_X1 U6741 ( .A1(n6839), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U6742 ( .A1(n5343), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6743 ( .A1(n5235), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5236) );
  AND2_X1 U6744 ( .A1(n5248), .A2(n5236), .ZN(n7452) );
  OR2_X1 U6745 ( .A1(n5076), .A2(n7452), .ZN(n5238) );
  INV_X1 U6746 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7254) );
  OR2_X1 U6747 ( .A1(n5378), .A2(n7254), .ZN(n5237) );
  NAND4_X1 U6748 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n7981)
         );
  AND2_X1 U6749 ( .A1(n10072), .A2(n7981), .ZN(n5241) );
  OR2_X1 U6750 ( .A1(n10072), .A2(n7981), .ZN(n5242) );
  XNOR2_X1 U6751 ( .A(n5244), .B(n5243), .ZN(n6510) );
  NAND2_X1 U6752 ( .A1(n6510), .A2(n7753), .ZN(n5247) );
  OR2_X1 U6753 ( .A1(n4399), .A2(n8452), .ZN(n5245) );
  XNOR2_X1 U6754 ( .A(n5245), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8019) );
  AOI22_X1 U6755 ( .A1(n7752), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5305), .B2(
        n8019), .ZN(n5246) );
  NAND2_X1 U6756 ( .A1(n6839), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6757 ( .A1(n5343), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5253) );
  NAND2_X1 U6758 ( .A1(n5248), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5249) );
  AND2_X1 U6759 ( .A1(n5264), .A2(n5249), .ZN(n7496) );
  OR2_X1 U6760 ( .A1(n5076), .A2(n7496), .ZN(n5252) );
  INV_X1 U6761 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5250) );
  OR2_X1 U6762 ( .A1(n5378), .A2(n5250), .ZN(n5251) );
  NAND4_X1 U6763 ( .A1(n5254), .A2(n5253), .A3(n5252), .A4(n5251), .ZN(n7980)
         );
  NOR2_X1 U6764 ( .A1(n9627), .A2(n7980), .ZN(n5255) );
  NAND2_X1 U6765 ( .A1(n6619), .A2(n7753), .ZN(n5262) );
  NAND2_X1 U6766 ( .A1(n5258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5287) );
  INV_X1 U6767 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U6768 ( .A1(n5287), .A2(n5259), .ZN(n5273) );
  OR2_X1 U6769 ( .A1(n5287), .A2(n5259), .ZN(n5260) );
  NAND2_X1 U6770 ( .A1(n5273), .A2(n5260), .ZN(n9979) );
  INV_X1 U6771 ( .A(n9979), .ZN(n8047) );
  AOI22_X1 U6772 ( .A1(n7752), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5305), .B2(
        n8047), .ZN(n5261) );
  NAND2_X1 U6773 ( .A1(n5343), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5269) );
  INV_X1 U6774 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8044) );
  OR2_X1 U6775 ( .A1(n5078), .A2(n8044), .ZN(n5268) );
  INV_X1 U6776 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5263) );
  OR2_X1 U6777 ( .A1(n5378), .A2(n5263), .ZN(n5267) );
  NAND2_X1 U6778 ( .A1(n5264), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5265) );
  AND2_X1 U6779 ( .A1(n5277), .A2(n5265), .ZN(n7539) );
  OR2_X1 U6780 ( .A1(n5076), .A2(n7539), .ZN(n5266) );
  NAND2_X1 U6781 ( .A1(n9619), .A2(n8326), .ZN(n7835) );
  NAND2_X1 U6782 ( .A1(n7836), .A2(n7835), .ZN(n7535) );
  INV_X1 U6783 ( .A(n8326), .ZN(n7979) );
  AND2_X1 U6784 ( .A1(n9619), .A2(n7979), .ZN(n5270) );
  XNOR2_X1 U6785 ( .A(n5272), .B(n5271), .ZN(n6676) );
  NAND2_X1 U6786 ( .A1(n6676), .A2(n7753), .ZN(n5276) );
  NAND2_X1 U6787 ( .A1(n5273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  XNOR2_X1 U6788 ( .A(n5274), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8078) );
  AOI22_X1 U6789 ( .A1(n7752), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5305), .B2(
        n8078), .ZN(n5275) );
  NAND2_X1 U6790 ( .A1(n5276), .A2(n5275), .ZN(n7525) );
  NAND2_X1 U6791 ( .A1(n5343), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5282) );
  INV_X1 U6792 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8392) );
  OR2_X1 U6793 ( .A1(n5378), .A2(n8392), .ZN(n5281) );
  OR2_X1 U6794 ( .A1(n5078), .A2(n8039), .ZN(n5280) );
  NAND2_X1 U6795 ( .A1(n5277), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5278) );
  AND2_X1 U6796 ( .A1(n5292), .A2(n5278), .ZN(n8330) );
  OR2_X1 U6797 ( .A1(n5076), .A2(n8330), .ZN(n5279) );
  NAND2_X1 U6798 ( .A1(n7525), .A2(n8308), .ZN(n5492) );
  NAND2_X1 U6799 ( .A1(n7839), .A2(n5492), .ZN(n8321) );
  INV_X1 U6800 ( .A(n7525), .ZN(n8451) );
  NAND2_X1 U6801 ( .A1(n8451), .A2(n8308), .ZN(n5283) );
  NAND2_X1 U6802 ( .A1(n6703), .A2(n7753), .ZN(n5291) );
  OAI21_X1 U6803 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U6804 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  OR2_X1 U6805 ( .A1(n5288), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6806 ( .A1(n5288), .A2(P2_IR_REG_16__SCAN_IN), .ZN(n5289) );
  NAND2_X1 U6807 ( .A1(n5303), .A2(n5289), .ZN(n8090) );
  INV_X1 U6808 ( .A(n8090), .ZN(n8096) );
  AOI22_X1 U6809 ( .A1(n7752), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5305), .B2(
        n8096), .ZN(n5290) );
  NAND2_X1 U6810 ( .A1(n5343), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5297) );
  INV_X1 U6811 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8316) );
  OR2_X1 U6812 ( .A1(n5078), .A2(n8316), .ZN(n5296) );
  NAND2_X1 U6813 ( .A1(n5292), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5293) );
  AND2_X1 U6814 ( .A1(n5308), .A2(n5293), .ZN(n8315) );
  OR2_X1 U6815 ( .A1(n5076), .A2(n8315), .ZN(n5295) );
  INV_X1 U6816 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8388) );
  OR2_X1 U6817 ( .A1(n5378), .A2(n8388), .ZN(n5294) );
  NAND2_X1 U6818 ( .A1(n7547), .A2(n8325), .ZN(n7849) );
  INV_X1 U6819 ( .A(n8325), .ZN(n5299) );
  NAND2_X1 U6820 ( .A1(n7547), .A2(n5299), .ZN(n5300) );
  XNOR2_X1 U6821 ( .A(n5301), .B(n5302), .ZN(n6748) );
  NAND2_X1 U6822 ( .A1(n6748), .A2(n7753), .ZN(n5307) );
  NAND2_X1 U6823 ( .A1(n5303), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5304) );
  XNOR2_X1 U6824 ( .A(n5304), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8130) );
  AOI22_X1 U6825 ( .A1(n7752), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5305), .B2(
        n8130), .ZN(n5306) );
  NAND2_X1 U6826 ( .A1(n5343), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5314) );
  INV_X1 U6827 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8383) );
  OR2_X1 U6828 ( .A1(n5378), .A2(n8383), .ZN(n5313) );
  INV_X1 U6829 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8301) );
  OR2_X1 U6830 ( .A1(n5078), .A2(n8301), .ZN(n5312) );
  NAND2_X1 U6831 ( .A1(n5308), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5309) );
  AND2_X1 U6832 ( .A1(n5310), .A2(n5309), .ZN(n8300) );
  OR2_X1 U6833 ( .A1(n5076), .A2(n8300), .ZN(n5311) );
  NAND2_X1 U6834 ( .A1(n8299), .A2(n8309), .ZN(n7854) );
  NAND2_X1 U6835 ( .A1(n7847), .A2(n7854), .ZN(n8297) );
  INV_X1 U6836 ( .A(n8309), .ZN(n7977) );
  NAND2_X1 U6837 ( .A1(n7644), .A2(n8283), .ZN(n7859) );
  INV_X1 U6838 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7013) );
  INV_X1 U6839 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7015) );
  MUX2_X1 U6840 ( .A(n7013), .B(n7015), .S(n7747), .Z(n5321) );
  INV_X1 U6841 ( .A(SI_20_), .ZN(n5320) );
  NAND2_X1 U6842 ( .A1(n5321), .A2(n5320), .ZN(n5336) );
  INV_X1 U6843 ( .A(n5321), .ZN(n5322) );
  NAND2_X1 U6844 ( .A1(n5322), .A2(SI_20_), .ZN(n5323) );
  NAND2_X1 U6845 ( .A1(n7012), .A2(n7753), .ZN(n5325) );
  OR2_X1 U6846 ( .A1(n7739), .A2(n7013), .ZN(n5324) );
  NAND2_X1 U6847 ( .A1(n6839), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6848 ( .A1(n6840), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5326) );
  AND2_X1 U6849 ( .A1(n5327), .A2(n5326), .ZN(n5332) );
  OR2_X2 U6850 ( .A1(n5328), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6851 ( .A1(n5328), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5329) );
  NAND2_X1 U6852 ( .A1(n5341), .A2(n5329), .ZN(n8264) );
  NAND2_X1 U6853 ( .A1(n8264), .A2(n5069), .ZN(n5331) );
  NAND2_X1 U6854 ( .A1(n5343), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5330) );
  NAND2_X1 U6855 ( .A1(n7692), .A2(n8271), .ZN(n8248) );
  NAND2_X1 U6856 ( .A1(n7863), .A2(n8248), .ZN(n8263) );
  INV_X1 U6857 ( .A(n8271), .ZN(n7974) );
  INV_X1 U6858 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7019) );
  INV_X1 U6859 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7040) );
  MUX2_X1 U6860 ( .A(n7019), .B(n7040), .S(n7747), .Z(n5349) );
  XNOR2_X1 U6861 ( .A(n5349), .B(SI_21_), .ZN(n5347) );
  XNOR2_X1 U6862 ( .A(n5348), .B(n5347), .ZN(n7018) );
  NAND2_X1 U6863 ( .A1(n7018), .A2(n7753), .ZN(n5338) );
  OR2_X1 U6864 ( .A1(n5460), .A2(n7019), .ZN(n5337) );
  INV_X1 U6865 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6866 ( .A1(n5341), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6867 ( .A1(n5359), .A2(n5342), .ZN(n8252) );
  NAND2_X1 U6868 ( .A1(n8252), .A2(n5069), .ZN(n5346) );
  AOI22_X1 U6869 ( .A1(n6840), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6839), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U6870 ( .A1(n5343), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6871 ( .A1(n7562), .A2(n8261), .ZN(n7868) );
  INV_X1 U6872 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6873 ( .A1(n5350), .A2(SI_21_), .ZN(n5351) );
  INV_X1 U6874 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7189) );
  INV_X1 U6875 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7604) );
  MUX2_X1 U6876 ( .A(n7189), .B(n7604), .S(n7747), .Z(n5354) );
  INV_X1 U6877 ( .A(SI_22_), .ZN(n5353) );
  NAND2_X1 U6878 ( .A1(n5354), .A2(n5353), .ZN(n5364) );
  INV_X1 U6879 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6880 ( .A1(n5355), .A2(SI_22_), .ZN(n5356) );
  NAND2_X1 U6881 ( .A1(n5364), .A2(n5356), .ZN(n5365) );
  NAND2_X1 U6882 ( .A1(n7188), .A2(n7753), .ZN(n5358) );
  OR2_X1 U6883 ( .A1(n5460), .A2(n7189), .ZN(n5357) );
  NAND2_X1 U6884 ( .A1(n5359), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5360) );
  NAND2_X1 U6885 ( .A1(n5376), .A2(n5360), .ZN(n8240) );
  NAND2_X1 U6886 ( .A1(n8240), .A2(n5069), .ZN(n5363) );
  AOI22_X1 U6887 ( .A1(n6840), .A2(P2_REG1_REG_22__SCAN_IN), .B1(n6839), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6888 ( .A1(n5343), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5361) );
  NAND2_X1 U6889 ( .A1(n7703), .A2(n8247), .ZN(n7874) );
  INV_X1 U6890 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7196) );
  INV_X1 U6891 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7192) );
  MUX2_X1 U6892 ( .A(n7196), .B(n7192), .S(n7747), .Z(n5368) );
  INV_X1 U6893 ( .A(SI_23_), .ZN(n5367) );
  NAND2_X1 U6894 ( .A1(n5368), .A2(n5367), .ZN(n5385) );
  INV_X1 U6895 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6896 ( .A1(n5369), .A2(SI_23_), .ZN(n5370) );
  OR2_X1 U6897 ( .A1(n5372), .A2(n5371), .ZN(n5373) );
  NAND2_X1 U6898 ( .A1(n7193), .A2(n7753), .ZN(n5375) );
  OR2_X1 U6899 ( .A1(n7739), .A2(n7196), .ZN(n5374) );
  NAND2_X1 U6900 ( .A1(n5376), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6901 ( .A1(n5396), .A2(n5377), .ZN(n8230) );
  NAND2_X1 U6902 ( .A1(n8230), .A2(n5069), .ZN(n5383) );
  INV_X1 U6903 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9035) );
  NAND2_X1 U6904 ( .A1(n6839), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5380) );
  INV_X1 U6905 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9095) );
  OR2_X1 U6906 ( .A1(n5378), .A2(n9095), .ZN(n5379) );
  OAI211_X1 U6907 ( .C1(n9035), .C2(n6844), .A(n5380), .B(n5379), .ZN(n5381)
         );
  INV_X1 U6908 ( .A(n5381), .ZN(n5382) );
  NOR2_X1 U6909 ( .A1(n7641), .A2(n7971), .ZN(n5384) );
  INV_X1 U6910 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7367) );
  INV_X1 U6911 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7368) );
  MUX2_X1 U6912 ( .A(n7367), .B(n7368), .S(n7747), .Z(n5388) );
  INV_X1 U6913 ( .A(SI_24_), .ZN(n5387) );
  NAND2_X1 U6914 ( .A1(n5388), .A2(n5387), .ZN(n5403) );
  INV_X1 U6915 ( .A(n5388), .ZN(n5389) );
  NAND2_X1 U6916 ( .A1(n5389), .A2(SI_24_), .ZN(n5390) );
  INV_X1 U6917 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6918 ( .A1(n5396), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6919 ( .A1(n5413), .A2(n5397), .ZN(n8220) );
  NAND2_X1 U6920 ( .A1(n8220), .A2(n5069), .ZN(n5402) );
  INV_X1 U6921 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U6922 ( .A1(n6840), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6923 ( .A1(n6839), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5398) );
  OAI211_X1 U6924 ( .C1(n9083), .C2(n6844), .A(n5399), .B(n5398), .ZN(n5400)
         );
  INV_X1 U6925 ( .A(n5400), .ZN(n5401) );
  INV_X1 U6926 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7417) );
  INV_X1 U6927 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7419) );
  MUX2_X1 U6928 ( .A(n7417), .B(n7419), .S(n7747), .Z(n5406) );
  INV_X1 U6929 ( .A(SI_25_), .ZN(n5405) );
  NAND2_X1 U6930 ( .A1(n5406), .A2(n5405), .ZN(n5422) );
  INV_X1 U6931 ( .A(n5406), .ZN(n5407) );
  NAND2_X1 U6932 ( .A1(n5407), .A2(SI_25_), .ZN(n5408) );
  NAND2_X1 U6933 ( .A1(n7416), .A2(n7753), .ZN(n5410) );
  OR2_X1 U6934 ( .A1(n7739), .A2(n7417), .ZN(n5409) );
  INV_X1 U6935 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6936 ( .A1(n5413), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6937 ( .A1(n5430), .A2(n5414), .ZN(n8211) );
  NAND2_X1 U6938 ( .A1(n8211), .A2(n5069), .ZN(n5419) );
  INV_X1 U6939 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U6940 ( .A1(n6840), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U6941 ( .A1(n6839), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U6942 ( .C1(n8410), .C2(n6844), .A(n5416), .B(n5415), .ZN(n5417)
         );
  INV_X1 U6943 ( .A(n5417), .ZN(n5418) );
  INV_X1 U6944 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7460) );
  INV_X1 U6945 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9560) );
  MUX2_X1 U6946 ( .A(n7460), .B(n9560), .S(n7747), .Z(n5425) );
  INV_X1 U6947 ( .A(SI_26_), .ZN(n5424) );
  NAND2_X1 U6948 ( .A1(n5425), .A2(n5424), .ZN(n5439) );
  INV_X1 U6949 ( .A(n5425), .ZN(n5426) );
  NAND2_X1 U6950 ( .A1(n5426), .A2(SI_26_), .ZN(n5427) );
  NAND2_X1 U6951 ( .A1(n7459), .A2(n7753), .ZN(n5429) );
  OR2_X1 U6952 ( .A1(n5460), .A2(n7460), .ZN(n5428) );
  NAND2_X1 U6953 ( .A1(n5430), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6954 ( .A1(n5449), .A2(n5431), .ZN(n8202) );
  NAND2_X1 U6955 ( .A1(n8202), .A2(n5069), .ZN(n5436) );
  INV_X1 U6956 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8406) );
  NAND2_X1 U6957 ( .A1(n6839), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U6958 ( .A1(n6840), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5432) );
  OAI211_X1 U6959 ( .C1(n6844), .C2(n8406), .A(n5433), .B(n5432), .ZN(n5434)
         );
  INV_X1 U6960 ( .A(n5434), .ZN(n5435) );
  INV_X1 U6961 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9104) );
  INV_X1 U6962 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U6963 ( .A(n9104), .B(n9556), .S(n7747), .Z(n5442) );
  INV_X1 U6964 ( .A(SI_27_), .ZN(n5441) );
  NAND2_X1 U6965 ( .A1(n5442), .A2(n5441), .ZN(n5459) );
  INV_X1 U6966 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U6967 ( .A1(n5443), .A2(SI_27_), .ZN(n5444) );
  AND2_X1 U6968 ( .A1(n5459), .A2(n5444), .ZN(n5457) );
  NAND2_X1 U6969 ( .A1(n8463), .A2(n7753), .ZN(n5446) );
  OR2_X1 U6970 ( .A1(n5460), .A2(n9104), .ZN(n5445) );
  INV_X1 U6971 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6972 ( .A1(n5449), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6973 ( .A1(n5463), .A2(n5450), .ZN(n8191) );
  NAND2_X1 U6974 ( .A1(n8191), .A2(n5069), .ZN(n5455) );
  INV_X1 U6975 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U6976 ( .A1(n6840), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5452) );
  NAND2_X1 U6977 ( .A1(n6839), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6978 ( .C1(n8402), .C2(n6844), .A(n5452), .B(n5451), .ZN(n5453)
         );
  INV_X1 U6979 ( .A(n5453), .ZN(n5454) );
  NOR2_X1 U6980 ( .A1(n8404), .A2(n8199), .ZN(n5456) );
  INV_X1 U6981 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8462) );
  INV_X1 U6982 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7612) );
  MUX2_X1 U6983 ( .A(n8462), .B(n7612), .S(n7747), .Z(n5565) );
  XNOR2_X1 U6984 ( .A(n5565), .B(SI_28_), .ZN(n5562) );
  NAND2_X1 U6985 ( .A1(n8459), .A2(n7753), .ZN(n5462) );
  OR2_X1 U6986 ( .A1(n5460), .A2(n8462), .ZN(n5461) );
  NAND2_X1 U6987 ( .A1(n5463), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5464) );
  NAND2_X1 U6988 ( .A1(n8164), .A2(n5464), .ZN(n8179) );
  NAND2_X1 U6989 ( .A1(n8179), .A2(n5069), .ZN(n5470) );
  INV_X1 U6990 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U6991 ( .A1(n6840), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6992 ( .A1(n6839), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5465) );
  OAI211_X1 U6993 ( .C1(n5467), .C2(n6844), .A(n5466), .B(n5465), .ZN(n5468)
         );
  INV_X1 U6994 ( .A(n5468), .ZN(n5469) );
  XNOR2_X1 U6995 ( .A(n5561), .B(n7950), .ZN(n5485) );
  INV_X1 U6996 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6997 ( .A1(n5474), .A2(n5472), .ZN(n5475) );
  XNOR2_X1 U6998 ( .A(n5473), .B(P2_IR_REG_21__SCAN_IN), .ZN(n5539) );
  NAND2_X1 U6999 ( .A1(n5476), .A2(n5475), .ZN(n7014) );
  INV_X1 U7000 ( .A(n7014), .ZN(n7918) );
  NAND2_X1 U7001 ( .A1(n5539), .A2(n7918), .ZN(n7756) );
  NAND2_X1 U7002 ( .A1(n4324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7003 ( .A1(n7957), .A2(n7962), .ZN(n5540) );
  INV_X1 U7004 ( .A(n8164), .ZN(n5478) );
  NAND2_X1 U7005 ( .A1(n5478), .A2(n5069), .ZN(n6842) );
  INV_X1 U7006 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U7007 ( .A1(n6839), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5480) );
  NAND2_X1 U7008 ( .A1(n6840), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5479) );
  OAI211_X1 U7009 ( .C1(n6844), .C2(n5481), .A(n5480), .B(n5479), .ZN(n5482)
         );
  INV_X1 U7010 ( .A(n5482), .ZN(n5483) );
  INV_X1 U7011 ( .A(n6423), .ZN(n7959) );
  XNOR2_X1 U7012 ( .A(n7959), .B(n8145), .ZN(n6518) );
  OAI22_X1 U7013 ( .A1(n7585), .A2(n10007), .B1(n8199), .B2(n8307), .ZN(n5484)
         );
  NAND2_X1 U7014 ( .A1(n6678), .A2(n5489), .ZN(n9999) );
  INV_X1 U7015 ( .A(n7929), .ZN(n10005) );
  NAND2_X1 U7016 ( .A1(n9999), .A2(n10005), .ZN(n10000) );
  INV_X1 U7017 ( .A(n10018), .ZN(n6530) );
  NAND2_X1 U7018 ( .A1(n6641), .A2(n6530), .ZN(n7775) );
  NAND2_X1 U7019 ( .A1(n10000), .A2(n7775), .ZN(n6721) );
  NAND2_X1 U7020 ( .A1(n10008), .A2(n6726), .ZN(n7790) );
  INV_X1 U7021 ( .A(n6726), .ZN(n10024) );
  NAND2_X1 U7022 ( .A1(n7988), .A2(n10024), .ZN(n7782) );
  NAND2_X1 U7023 ( .A1(n7987), .A2(n10030), .ZN(n7792) );
  NAND2_X1 U7024 ( .A1(n5123), .A2(n4856), .ZN(n7784) );
  NOR2_X1 U7025 ( .A1(n9983), .A2(n10034), .ZN(n7783) );
  NAND2_X1 U7026 ( .A1(n9983), .A2(n10034), .ZN(n9988) );
  NAND2_X1 U7027 ( .A1(n7986), .A2(n6834), .ZN(n7927) );
  AND2_X1 U7028 ( .A1(n9988), .A2(n7927), .ZN(n7793) );
  NAND2_X1 U7029 ( .A1(n7119), .A2(n10039), .ZN(n7928) );
  INV_X1 U7030 ( .A(n7139), .ZN(n7049) );
  NAND2_X1 U7031 ( .A1(n7985), .A2(n7049), .ZN(n7808) );
  AND2_X1 U7032 ( .A1(n7045), .A2(n7808), .ZN(n7802) );
  NOR2_X1 U7033 ( .A1(n7985), .A2(n7049), .ZN(n7806) );
  NAND2_X1 U7034 ( .A1(n10049), .A2(n7984), .ZN(n7312) );
  INV_X1 U7035 ( .A(n10049), .ZN(n7185) );
  NAND2_X1 U7036 ( .A1(n7316), .A2(n7185), .ZN(n7811) );
  NAND2_X1 U7037 ( .A1(n7177), .A2(n7933), .ZN(n7313) );
  OR2_X1 U7038 ( .A1(n7323), .A2(n7431), .ZN(n7820) );
  AND2_X1 U7039 ( .A1(n7820), .A2(n7312), .ZN(n7813) );
  NAND2_X1 U7040 ( .A1(n7323), .A2(n7431), .ZN(n7816) );
  XNOR2_X1 U7041 ( .A(n10065), .B(n7982), .ZN(n7422) );
  INV_X1 U7042 ( .A(n7982), .ZN(n7817) );
  NAND2_X1 U7043 ( .A1(n10065), .A2(n7817), .ZN(n7822) );
  XNOR2_X1 U7044 ( .A(n10072), .B(n7826), .ZN(n7938) );
  OR2_X1 U7045 ( .A1(n10072), .A2(n7826), .ZN(n7828) );
  INV_X1 U7046 ( .A(n7980), .ZN(n7538) );
  NAND2_X1 U7047 ( .A1(n9627), .A2(n7538), .ZN(n7831) );
  OR2_X1 U7048 ( .A1(n9627), .A2(n7538), .ZN(n7832) );
  INV_X1 U7049 ( .A(n5492), .ZN(n7840) );
  NAND2_X1 U7050 ( .A1(n7722), .A2(n8296), .ZN(n7853) );
  NAND2_X1 U7051 ( .A1(n7856), .A2(n7853), .ZN(n8286) );
  INV_X1 U7052 ( .A(n7857), .ZN(n5494) );
  NAND2_X1 U7053 ( .A1(n8262), .A2(n7863), .ZN(n8249) );
  AND2_X1 U7054 ( .A1(n7868), .A2(n8248), .ZN(n7864) );
  NAND2_X1 U7055 ( .A1(n8249), .A2(n7864), .ZN(n5495) );
  NAND2_X1 U7056 ( .A1(n5495), .A2(n7869), .ZN(n8238) );
  NAND2_X1 U7057 ( .A1(n7641), .A2(n8237), .ZN(n7878) );
  INV_X1 U7058 ( .A(n7879), .ZN(n5496) );
  INV_X1 U7059 ( .A(n7885), .ZN(n5498) );
  NAND2_X1 U7060 ( .A1(n5499), .A2(n8199), .ZN(n7888) );
  INV_X1 U7061 ( .A(n5573), .ZN(n5502) );
  AOI21_X1 U7062 ( .B1(n7950), .B2(n5501), .A(n5502), .ZN(n8178) );
  INV_X1 U7063 ( .A(n6514), .ZN(n5505) );
  AND2_X1 U7064 ( .A1(n8154), .A2(n7962), .ZN(n5551) );
  INV_X1 U7065 ( .A(n5551), .ZN(n5503) );
  NAND2_X1 U7066 ( .A1(n5505), .A2(n5503), .ZN(n5504) );
  AND2_X1 U7067 ( .A1(n10054), .A2(n5504), .ZN(n5506) );
  AND2_X1 U7068 ( .A1(n7014), .A2(n7957), .ZN(n6722) );
  NAND2_X1 U7069 ( .A1(n8185), .A2(n5507), .ZN(n5557) );
  NAND2_X1 U7070 ( .A1(n5508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7071 ( .A1(n5511), .A2(n9109), .ZN(n5513) );
  NAND2_X1 U7072 ( .A1(n5513), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5510) );
  XNOR2_X1 U7073 ( .A(n5510), .B(n5509), .ZN(n7418) );
  OR2_X1 U7074 ( .A1(n5511), .A2(n9109), .ZN(n5512) );
  XNOR2_X1 U7075 ( .A(n7366), .B(P2_B_REG_SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7076 ( .A1(n7418), .A2(n5514), .ZN(n5516) );
  NAND2_X1 U7077 ( .A1(n4367), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5515) );
  INV_X1 U7078 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n5517) );
  INV_X1 U7079 ( .A(n6286), .ZN(n7461) );
  NAND2_X1 U7080 ( .A1(n7461), .A2(n7366), .ZN(n5518) );
  NOR2_X1 U7081 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .ZN(
        n9124) );
  NOR4_X1 U7082 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5522) );
  NOR4_X1 U7083 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5521) );
  NOR4_X1 U7084 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n5520) );
  NAND4_X1 U7085 ( .A1(n9124), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n5528)
         );
  NOR4_X1 U7086 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5526) );
  NOR4_X1 U7087 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n5525) );
  NOR4_X1 U7088 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n5524) );
  NOR4_X1 U7089 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n5523) );
  NAND4_X1 U7090 ( .A1(n5526), .A2(n5525), .A3(n5524), .A4(n5523), .ZN(n5527)
         );
  NOR2_X1 U7091 ( .A1(n5528), .A2(n5527), .ZN(n5529) );
  OR2_X1 U7092 ( .A1(n6283), .A2(n5529), .ZN(n5548) );
  INV_X1 U7093 ( .A(n5548), .ZN(n5543) );
  NOR2_X1 U7094 ( .A1(n6594), .A2(n5543), .ZN(n5532) );
  OR2_X1 U7095 ( .A1(n6283), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7096 ( .A1(n7418), .A2(n7461), .ZN(n5530) );
  INV_X1 U7097 ( .A(n6268), .ZN(n6590) );
  AND2_X1 U7098 ( .A1(n5532), .A2(n6590), .ZN(n6502) );
  INV_X1 U7099 ( .A(n7366), .ZN(n6285) );
  NAND2_X1 U7100 ( .A1(n6286), .A2(n6285), .ZN(n5533) );
  INV_X1 U7101 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7102 ( .A1(n5535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5537) );
  XNOR2_X1 U7103 ( .A(n5537), .B(n5536), .ZN(n6495) );
  AND2_X1 U7104 ( .A1(n6495), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5538) );
  AND2_X1 U7105 ( .A1(n6502), .A2(n6284), .ZN(n6490) );
  INV_X1 U7106 ( .A(n5540), .ZN(n5541) );
  NAND2_X1 U7107 ( .A1(n4326), .A2(n5541), .ZN(n6500) );
  AND2_X1 U7108 ( .A1(n7903), .A2(n10054), .ZN(n5542) );
  NAND2_X1 U7109 ( .A1(n6500), .A2(n5542), .ZN(n6484) );
  NAND2_X1 U7110 ( .A1(n6484), .A2(n10003), .ZN(n6494) );
  NAND2_X1 U7111 ( .A1(n6490), .A2(n6494), .ZN(n5546) );
  NAND2_X1 U7112 ( .A1(n6594), .A2(n6268), .ZN(n5549) );
  OR2_X1 U7113 ( .A1(n5549), .A2(n5543), .ZN(n6493) );
  NOR2_X1 U7114 ( .A1(n6493), .A2(n6503), .ZN(n6486) );
  NAND2_X1 U7115 ( .A1(n6500), .A2(n6504), .ZN(n5544) );
  NAND2_X1 U7116 ( .A1(n6486), .A2(n5544), .ZN(n5545) );
  OR2_X1 U7117 ( .A1(n7903), .A2(n6514), .ZN(n6497) );
  AND2_X1 U7118 ( .A1(n6284), .A2(n5548), .ZN(n5550) );
  NAND2_X1 U7119 ( .A1(n7918), .A2(n5551), .ZN(n5552) );
  INV_X1 U7120 ( .A(n6593), .ZN(n5553) );
  NAND2_X1 U7121 ( .A1(n5553), .A2(n6590), .ZN(n5556) );
  NAND2_X1 U7122 ( .A1(n10046), .A2(n7762), .ZN(n6481) );
  NAND2_X1 U7123 ( .A1(n6481), .A2(n6594), .ZN(n5554) );
  NAND2_X1 U7124 ( .A1(n5554), .A2(n6593), .ZN(n5555) );
  NAND2_X1 U7125 ( .A1(n5557), .A2(n10092), .ZN(n5559) );
  NAND2_X1 U7126 ( .A1(n10090), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5558) );
  INV_X1 U7127 ( .A(n10054), .ZN(n10073) );
  NAND2_X1 U7128 ( .A1(n4905), .A2(n4899), .ZN(P2_U3487) );
  NOR2_X1 U7129 ( .A1(n7589), .A2(n7967), .ZN(n5560) );
  OAI22_X1 U7130 ( .A1(n5561), .A2(n5560), .B1(n8188), .B2(n8181), .ZN(n5571)
         );
  INV_X1 U7131 ( .A(SI_28_), .ZN(n5564) );
  NAND2_X1 U7132 ( .A1(n5565), .A2(n5564), .ZN(n5566) );
  INV_X1 U7133 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5568) );
  INV_X1 U7134 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8721) );
  MUX2_X1 U7135 ( .A(n5568), .B(n8721), .S(n7747), .Z(n7592) );
  NAND2_X1 U7136 ( .A1(n8720), .A2(n7753), .ZN(n5570) );
  OR2_X1 U7137 ( .A1(n7739), .A2(n5568), .ZN(n5569) );
  NAND2_X1 U7138 ( .A1(n5584), .A2(n7585), .ZN(n7742) );
  XNOR2_X1 U7139 ( .A(n5571), .B(n7897), .ZN(n5582) );
  NAND2_X1 U7140 ( .A1(n7589), .A2(n8188), .ZN(n5572) );
  INV_X1 U7141 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7142 ( .A1(n6840), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7143 ( .A1(n6839), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n5574) );
  OAI211_X1 U7144 ( .C1(n5576), .C2(n6844), .A(n5575), .B(n5574), .ZN(n5577)
         );
  INV_X1 U7145 ( .A(n5577), .ZN(n5578) );
  AND2_X1 U7146 ( .A1(n6842), .A2(n5578), .ZN(n7902) );
  NAND2_X1 U7147 ( .A1(n6246), .A2(P2_B_REG_SCAN_IN), .ZN(n5579) );
  NAND2_X1 U7148 ( .A1(n9984), .A2(n5579), .ZN(n8162) );
  OAI22_X1 U7149 ( .A1(n8188), .A2(n8307), .B1(n7902), .B2(n8162), .ZN(n5580)
         );
  INV_X1 U7150 ( .A(n10046), .ZN(n10056) );
  NAND2_X1 U7151 ( .A1(n6241), .A2(n10074), .ZN(n5588) );
  NOR2_X1 U7152 ( .A1(n8171), .A2(n8450), .ZN(n5585) );
  NAND2_X1 U7153 ( .A1(n5588), .A2(n5587), .ZN(P2_U3456) );
  NOR2_X1 U7154 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5597) );
  NOR2_X1 U7155 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5596) );
  INV_X1 U7156 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U7157 ( .A1(n5601), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5603) );
  INV_X1 U7158 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5602) );
  INV_X1 U7159 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6306) );
  OR2_X1 U7160 ( .A1(n8615), .A2(n6306), .ZN(n5610) );
  NAND2_X1 U7161 ( .A1(n8616), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5609) );
  NAND2_X4 U7162 ( .A1(n5606), .A2(n5605), .ZN(n6542) );
  INV_X1 U7163 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9020) );
  OR2_X1 U7164 ( .A1(n8620), .A2(n9020), .ZN(n5607) );
  NAND4_X2 U7165 ( .A1(n5610), .A2(n5609), .A3(n5608), .A4(n5607), .ZN(n6752)
         );
  MUX2_X1 U7166 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5611), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5612) );
  NAND2_X1 U7167 ( .A1(n5612), .A2(n5634), .ZN(n9563) );
  NAND2_X1 U7168 ( .A1(n5613), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5614) );
  MUX2_X1 U7169 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5614), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5616) );
  NAND2_X1 U7170 ( .A1(n5616), .A2(n5615), .ZN(n7421) );
  INV_X1 U7171 ( .A(n5617), .ZN(n5618) );
  NAND2_X1 U7172 ( .A1(n5618), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5619) );
  MUX2_X1 U7173 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5619), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5620) );
  NAND2_X1 U7174 ( .A1(n5620), .A2(n5613), .ZN(n7370) );
  NOR2_X1 U7175 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5622) );
  INV_X1 U7176 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7177 ( .A1(n5643), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  INV_X1 U7178 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5624) );
  XNOR2_X2 U7179 ( .A(n5625), .B(n5624), .ZN(n8737) );
  INV_X1 U7181 ( .A(n5626), .ZN(n5627) );
  NAND2_X1 U7182 ( .A1(n5627), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5628) );
  MUX2_X1 U7183 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5628), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5629) );
  NAND2_X1 U7184 ( .A1(n5629), .A2(n5643), .ZN(n7017) );
  AND2_X1 U7185 ( .A1(n8786), .A2(n7017), .ZN(n5630) );
  NAND2_X1 U7186 ( .A1(n6752), .A2(n5655), .ZN(n5653) );
  XNOR2_X2 U7187 ( .A(n5633), .B(n5632), .ZN(n7611) );
  XNOR2_X2 U7188 ( .A(n5636), .B(n5635), .ZN(n9677) );
  NAND2_X1 U7189 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5637) );
  MUX2_X1 U7190 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5637), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5640) );
  INV_X1 U7191 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7192 ( .A1(n5640), .A2(n5639), .ZN(n6305) );
  NAND2_X2 U7193 ( .A1(n4310), .A2(n7747), .ZN(n5797) );
  INV_X1 U7194 ( .A(n5641), .ZN(n6261) );
  INV_X1 U7195 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6202) );
  INV_X1 U7196 ( .A(n5644), .ZN(n5645) );
  INV_X1 U7197 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U7198 ( .A1(n6002), .A2(n9119), .ZN(n5646) );
  XNOR2_X2 U7199 ( .A(n5648), .B(n5647), .ZN(n8866) );
  NAND2_X1 U7200 ( .A1(n7017), .A2(n8866), .ZN(n6231) );
  INV_X2 U7201 ( .A(n6231), .ZN(n8834) );
  NAND2_X1 U7202 ( .A1(n8868), .A2(n8834), .ZN(n5649) );
  INV_X2 U7203 ( .A(n8866), .ZN(n8980) );
  AND2_X1 U7204 ( .A1(n7017), .A2(n8980), .ZN(n8835) );
  NAND2_X1 U7205 ( .A1(n8835), .A2(n8786), .ZN(n6872) );
  AND2_X1 U7206 ( .A1(n6872), .A2(n5649), .ZN(n5650) );
  NAND2_X1 U7207 ( .A1(n6243), .A2(n5650), .ZN(n6138) );
  NAND2_X1 U7208 ( .A1(n8737), .A2(n8980), .ZN(n5651) );
  NAND2_X1 U7209 ( .A1(n8786), .A2(n8853), .ZN(n8870) );
  XNOR2_X1 U7210 ( .A(n5654), .B(n6173), .ZN(n5658) );
  INV_X2 U7211 ( .A(n6138), .ZN(n7615) );
  AND2_X1 U7212 ( .A1(n6874), .A2(n7620), .ZN(n5656) );
  AOI21_X1 U7213 ( .B1(n6752), .B2(n7615), .A(n5656), .ZN(n5657) );
  NAND2_X1 U7214 ( .A1(n5658), .A2(n5657), .ZN(n6668) );
  NAND2_X1 U7215 ( .A1(n4306), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5665) );
  INV_X1 U7216 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5660) );
  OR2_X1 U7217 ( .A1(n4309), .A2(n5660), .ZN(n5664) );
  INV_X1 U7218 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9676) );
  OR2_X1 U7219 ( .A1(n8615), .A2(n9676), .ZN(n5663) );
  INV_X1 U7220 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5661) );
  NAND2_X1 U7221 ( .A1(n7747), .A2(SI_0_), .ZN(n5667) );
  INV_X1 U7222 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7223 ( .A1(n5667), .A2(n5666), .ZN(n5669) );
  AND2_X1 U7224 ( .A1(n5669), .A2(n5668), .ZN(n9564) );
  MUX2_X1 U7225 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9564), .S(n4310), .Z(n6770) );
  AND2_X1 U7226 ( .A1(n6770), .A2(n5687), .ZN(n5670) );
  INV_X1 U7227 ( .A(n6243), .ZN(n5672) );
  NAND2_X1 U7228 ( .A1(n5672), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5671) );
  NAND2_X1 U7229 ( .A1(n5675), .A2(n5671), .ZN(n6477) );
  NAND2_X1 U7230 ( .A1(n6771), .A2(n7615), .ZN(n5674) );
  INV_X2 U7231 ( .A(n6139), .ZN(n6035) );
  AOI22_X1 U7232 ( .A1(n6770), .A2(n6035), .B1(n5672), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7233 ( .A1(n5674), .A2(n5673), .ZN(n6476) );
  NAND2_X1 U7234 ( .A1(n6477), .A2(n6476), .ZN(n5677) );
  INV_X4 U7235 ( .A(n7618), .ZN(n6173) );
  NAND2_X1 U7236 ( .A1(n5675), .A2(n6173), .ZN(n5676) );
  NAND2_X1 U7237 ( .A1(n5677), .A2(n5676), .ZN(n6624) );
  INV_X1 U7238 ( .A(n6624), .ZN(n5678) );
  NAND2_X1 U7239 ( .A1(n4307), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5683) );
  INV_X1 U7240 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6307) );
  OR2_X1 U7241 ( .A1(n8615), .A2(n6307), .ZN(n5682) );
  INV_X1 U7242 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5679) );
  OR2_X1 U7243 ( .A1(n4309), .A2(n5679), .ZN(n5681) );
  INV_X1 U7244 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9740) );
  OR2_X1 U7245 ( .A1(n6542), .A2(n9740), .ZN(n5680) );
  NAND2_X1 U7246 ( .A1(n8898), .A2(n6035), .ZN(n5689) );
  OR2_X1 U7247 ( .A1(n5704), .A2(n6250), .ZN(n5685) );
  NAND2_X1 U7248 ( .A1(n6767), .A2(n5687), .ZN(n5688) );
  NAND2_X1 U7249 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  XNOR2_X1 U7250 ( .A(n5690), .B(n6173), .ZN(n5692) );
  AND2_X1 U7251 ( .A1(n6767), .A2(n7620), .ZN(n5691) );
  AOI21_X1 U7252 ( .B1(n8898), .B2(n7615), .A(n5691), .ZN(n5693) );
  NAND2_X1 U7253 ( .A1(n5692), .A2(n5693), .ZN(n5697) );
  INV_X1 U7254 ( .A(n5692), .ZN(n5695) );
  INV_X1 U7255 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7256 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  AND2_X1 U7257 ( .A1(n5697), .A2(n5696), .ZN(n6669) );
  NAND2_X1 U7258 ( .A1(n6670), .A2(n5697), .ZN(n8493) );
  NAND2_X1 U7259 ( .A1(n4306), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5701) );
  INV_X1 U7260 ( .A(n4308), .ZN(n6145) );
  NAND2_X1 U7261 ( .A1(n6145), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5700) );
  OR2_X1 U7262 ( .A1(n6542), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5699) );
  INV_X1 U7263 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6321) );
  OR2_X1 U7264 ( .A1(n8615), .A2(n6321), .ZN(n5698) );
  NAND4_X1 U7265 ( .A1(n5701), .A2(n5700), .A3(n5699), .A4(n5698), .ZN(n8897)
         );
  NAND2_X1 U7266 ( .A1(n8897), .A2(n6035), .ZN(n5708) );
  OR2_X1 U7267 ( .A1(n5702), .A2(n5838), .ZN(n5703) );
  XNOR2_X1 U7268 ( .A(n5703), .B(n5716), .ZN(n6329) );
  OR2_X1 U7269 ( .A1(n5797), .A2(n6256), .ZN(n5706) );
  OR2_X1 U7270 ( .A1(n8729), .A2(n6252), .ZN(n5705) );
  NAND2_X1 U7271 ( .A1(n8497), .A2(n5687), .ZN(n5707) );
  NAND2_X1 U7272 ( .A1(n5708), .A2(n5707), .ZN(n5709) );
  XNOR2_X1 U7273 ( .A(n5709), .B(n7618), .ZN(n5727) );
  AND2_X1 U7274 ( .A1(n8497), .A2(n7620), .ZN(n5710) );
  AOI21_X1 U7275 ( .B1(n8897), .B2(n7615), .A(n5710), .ZN(n5728) );
  XNOR2_X1 U7276 ( .A(n5727), .B(n5728), .ZN(n8494) );
  NAND2_X1 U7277 ( .A1(n6145), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7278 ( .A1(n6218), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5714) );
  XNOR2_X1 U7279 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9673) );
  OR2_X1 U7280 ( .A1(n6542), .A2(n9673), .ZN(n5713) );
  INV_X1 U7281 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5711) );
  OR2_X1 U7282 ( .A1(n5736), .A2(n5711), .ZN(n5712) );
  NAND2_X1 U7283 ( .A1(n8896), .A2(n6035), .ZN(n5724) );
  NAND2_X1 U7284 ( .A1(n5702), .A2(n5716), .ZN(n5717) );
  INV_X1 U7285 ( .A(n5763), .ZN(n5720) );
  NAND2_X1 U7286 ( .A1(n5717), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5718) );
  MUX2_X1 U7287 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5718), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5719) );
  NAND2_X1 U7288 ( .A1(n5720), .A2(n5719), .ZN(n6689) );
  OR2_X1 U7289 ( .A1(n8729), .A2(n9102), .ZN(n5722) );
  OR2_X1 U7290 ( .A1(n5797), .A2(n6254), .ZN(n5721) );
  OAI211_X1 U7291 ( .C1(n4311), .C2(n6689), .A(n5722), .B(n5721), .ZN(n9671)
         );
  NAND2_X1 U7292 ( .A1(n9671), .A2(n4294), .ZN(n5723) );
  NAND2_X1 U7293 ( .A1(n5724), .A2(n5723), .ZN(n5725) );
  XNOR2_X1 U7294 ( .A(n5725), .B(n7618), .ZN(n5733) );
  AND2_X1 U7295 ( .A1(n9671), .A2(n7620), .ZN(n5726) );
  AOI21_X1 U7296 ( .B1(n8896), .B2(n7615), .A(n5726), .ZN(n5731) );
  XNOR2_X1 U7297 ( .A(n5733), .B(n5731), .ZN(n9662) );
  INV_X1 U7298 ( .A(n5727), .ZN(n5729) );
  NAND2_X1 U7299 ( .A1(n5729), .A2(n5728), .ZN(n9663) );
  AND2_X1 U7300 ( .A1(n9662), .A2(n9663), .ZN(n5730) );
  INV_X1 U7301 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7302 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  INV_X1 U7303 ( .A(n6542), .ZN(n6144) );
  AOI21_X1 U7304 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5735) );
  NOR2_X1 U7305 ( .A1(n5735), .A2(n5755), .ZN(n6929) );
  NAND2_X1 U7306 ( .A1(n6144), .A2(n6929), .ZN(n5742) );
  INV_X1 U7307 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5737) );
  OR2_X1 U7308 ( .A1(n5736), .A2(n5737), .ZN(n5741) );
  INV_X1 U7309 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6318) );
  OR2_X1 U7310 ( .A1(n8615), .A2(n6318), .ZN(n5740) );
  INV_X1 U7311 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5738) );
  OR2_X1 U7312 ( .A1(n4308), .A2(n5738), .ZN(n5739) );
  NAND4_X1 U7313 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n8895)
         );
  NAND2_X1 U7314 ( .A1(n8895), .A2(n6035), .ZN(n5747) );
  OR2_X1 U7315 ( .A1(n5763), .A2(n5838), .ZN(n5743) );
  XNOR2_X1 U7316 ( .A(n5743), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6333) );
  INV_X1 U7317 ( .A(n6333), .ZN(n6398) );
  OR2_X1 U7318 ( .A1(n5797), .A2(n6259), .ZN(n5745) );
  OR2_X1 U7319 ( .A1(n8729), .A2(n6258), .ZN(n5744) );
  OAI211_X1 U7320 ( .C1(n6281), .C2(n6398), .A(n5745), .B(n5744), .ZN(n6859)
         );
  NAND2_X1 U7321 ( .A1(n6859), .A2(n4294), .ZN(n5746) );
  NAND2_X1 U7322 ( .A1(n5747), .A2(n5746), .ZN(n5748) );
  XNOR2_X1 U7323 ( .A(n5748), .B(n7618), .ZN(n5751) );
  NAND2_X1 U7324 ( .A1(n8895), .A2(n7615), .ZN(n5750) );
  NAND2_X1 U7325 ( .A1(n6859), .A2(n6035), .ZN(n5749) );
  NAND2_X1 U7326 ( .A1(n5750), .A2(n5749), .ZN(n6925) );
  NAND2_X1 U7327 ( .A1(n6922), .A2(n6925), .ZN(n5753) );
  NAND2_X1 U7328 ( .A1(n5752), .A2(n5751), .ZN(n6923) );
  NAND2_X1 U7329 ( .A1(n5753), .A2(n6923), .ZN(n6934) );
  NAND2_X1 U7330 ( .A1(n6218), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5761) );
  INV_X1 U7331 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5754) );
  OR2_X1 U7332 ( .A1(n5736), .A2(n5754), .ZN(n5760) );
  INV_X1 U7333 ( .A(n5778), .ZN(n5780) );
  INV_X1 U7334 ( .A(n5755), .ZN(n5756) );
  INV_X1 U7335 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7336 ( .A1(n5756), .A2(n6328), .ZN(n5757) );
  NAND2_X1 U7337 ( .A1(n5780), .A2(n5757), .ZN(n9725) );
  OR2_X1 U7338 ( .A1(n6542), .A2(n9725), .ZN(n5759) );
  INV_X1 U7339 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6334) );
  OR2_X1 U7340 ( .A1(n4309), .A2(n6334), .ZN(n5758) );
  NAND4_X1 U7341 ( .A1(n5761), .A2(n5760), .A3(n5759), .A4(n5758), .ZN(n8894)
         );
  NAND2_X1 U7342 ( .A1(n8894), .A2(n6035), .ZN(n5769) );
  NAND2_X1 U7343 ( .A1(n5763), .A2(n5762), .ZN(n5786) );
  NAND2_X1 U7344 ( .A1(n5786), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5765) );
  XNOR2_X1 U7345 ( .A(n5765), .B(n5764), .ZN(n6347) );
  OR2_X1 U7346 ( .A1(n5797), .A2(n6263), .ZN(n5767) );
  OR2_X1 U7347 ( .A1(n8729), .A2(n6262), .ZN(n5766) );
  OAI211_X1 U7348 ( .C1(n6281), .C2(n6347), .A(n5767), .B(n5766), .ZN(n6995)
         );
  NAND2_X1 U7349 ( .A1(n6995), .A2(n4294), .ZN(n5768) );
  NAND2_X1 U7350 ( .A1(n5769), .A2(n5768), .ZN(n5770) );
  XNOR2_X1 U7351 ( .A(n5770), .B(n7618), .ZN(n5773) );
  NAND2_X1 U7352 ( .A1(n8894), .A2(n7615), .ZN(n5772) );
  NAND2_X1 U7353 ( .A1(n6995), .A2(n6035), .ZN(n5771) );
  NAND2_X1 U7354 ( .A1(n5772), .A2(n5771), .ZN(n5774) );
  AND2_X1 U7355 ( .A1(n5773), .A2(n5774), .ZN(n6936) );
  INV_X1 U7356 ( .A(n5773), .ZN(n5776) );
  INV_X1 U7357 ( .A(n5774), .ZN(n5775) );
  NAND2_X1 U7358 ( .A1(n5776), .A2(n5775), .ZN(n6935) );
  NAND2_X1 U7359 ( .A1(n4306), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7360 ( .A1(n5778), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5814) );
  INV_X1 U7361 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7362 ( .A1(n5780), .A2(n5779), .ZN(n5781) );
  NAND2_X1 U7363 ( .A1(n5814), .A2(n5781), .ZN(n9658) );
  OR2_X1 U7364 ( .A1(n6542), .A2(n9658), .ZN(n5784) );
  INV_X1 U7365 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7005) );
  OR2_X1 U7366 ( .A1(n4309), .A2(n7005), .ZN(n5783) );
  INV_X1 U7367 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6343) );
  OR2_X1 U7368 ( .A1(n8615), .A2(n6343), .ZN(n5782) );
  NAND4_X1 U7369 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n8893)
         );
  NAND2_X1 U7370 ( .A1(n8893), .A2(n6035), .ZN(n5791) );
  OAI21_X1 U7371 ( .B1(n5786), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5787) );
  XNOR2_X1 U7372 ( .A(n5787), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6350) );
  INV_X1 U7373 ( .A(n6350), .ZN(n6372) );
  OR2_X1 U7374 ( .A1(n8729), .A2(n6266), .ZN(n5788) );
  NAND2_X1 U7375 ( .A1(n9656), .A2(n4293), .ZN(n5790) );
  NAND2_X1 U7376 ( .A1(n5791), .A2(n5790), .ZN(n5792) );
  XNOR2_X1 U7377 ( .A(n5792), .B(n7618), .ZN(n5795) );
  AOI22_X1 U7378 ( .A1(n8893), .A2(n7615), .B1(n7620), .B2(n9656), .ZN(n5793)
         );
  XNOR2_X1 U7379 ( .A(n5795), .B(n5793), .ZN(n9651) );
  INV_X1 U7380 ( .A(n5793), .ZN(n5794) );
  NAND2_X1 U7381 ( .A1(n5795), .A2(n5794), .ZN(n5796) );
  NAND2_X1 U7382 ( .A1(n6288), .A2(n8730), .ZN(n5802) );
  INV_X1 U7383 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U7384 ( .A1(n4299), .A2(n5799), .ZN(n5837) );
  NAND2_X1 U7385 ( .A1(n5837), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5800) );
  XNOR2_X1 U7386 ( .A(n5800), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6411) );
  AOI22_X1 U7387 ( .A1(n6021), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6020), .B2(
        n6411), .ZN(n5801) );
  NAND2_X1 U7388 ( .A1(n7339), .A2(n4294), .ZN(n5812) );
  NAND2_X1 U7389 ( .A1(n4307), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5810) );
  INV_X1 U7390 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5803) );
  OR2_X1 U7391 ( .A1(n8615), .A2(n5803), .ZN(n5809) );
  INV_X1 U7392 ( .A(n5814), .ZN(n5804) );
  NAND2_X1 U7393 ( .A1(n5804), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5816) );
  INV_X1 U7394 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5805) );
  NAND2_X1 U7395 ( .A1(n5816), .A2(n5805), .ZN(n5806) );
  NAND2_X1 U7396 ( .A1(n5842), .A2(n5806), .ZN(n7337) );
  OR2_X1 U7397 ( .A1(n6542), .A2(n7337), .ZN(n5808) );
  INV_X1 U7398 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7034) );
  OR2_X1 U7399 ( .A1(n4309), .A2(n7034), .ZN(n5807) );
  NAND4_X1 U7400 ( .A1(n5810), .A2(n5809), .A3(n5808), .A4(n5807), .ZN(n8891)
         );
  NAND2_X1 U7401 ( .A1(n8891), .A2(n6097), .ZN(n5811) );
  NAND2_X1 U7402 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  XNOR2_X1 U7403 ( .A(n5813), .B(n6173), .ZN(n5833) );
  AOI22_X1 U7404 ( .A1(n7339), .A2(n6035), .B1(n7615), .B2(n8891), .ZN(n5832)
         );
  OR2_X1 U7405 ( .A1(n5833), .A2(n5832), .ZN(n7329) );
  NAND2_X1 U7406 ( .A1(n4307), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5821) );
  INV_X1 U7407 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6342) );
  OR2_X1 U7408 ( .A1(n8615), .A2(n6342), .ZN(n5820) );
  INV_X1 U7409 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7289) );
  NAND2_X1 U7410 ( .A1(n5814), .A2(n7289), .ZN(n5815) );
  NAND2_X1 U7411 ( .A1(n5816), .A2(n5815), .ZN(n9710) );
  OR2_X1 U7412 ( .A1(n6542), .A2(n9710), .ZN(n5819) );
  INV_X1 U7413 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5817) );
  OR2_X1 U7414 ( .A1(n4309), .A2(n5817), .ZN(n5818) );
  NAND4_X1 U7415 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n8892)
         );
  NAND2_X1 U7416 ( .A1(n8892), .A2(n6097), .ZN(n5826) );
  NAND2_X1 U7417 ( .A1(n6274), .A2(n8730), .ZN(n5824) );
  OR2_X1 U7418 ( .A1(n4299), .A2(n5838), .ZN(n5822) );
  XNOR2_X1 U7419 ( .A(n5822), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6352) );
  AOI22_X1 U7420 ( .A1(n6021), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6020), .B2(
        n6352), .ZN(n5823) );
  NAND2_X1 U7421 ( .A1(n5824), .A2(n5823), .ZN(n7031) );
  NAND2_X1 U7422 ( .A1(n7031), .A2(n4294), .ZN(n5825) );
  NAND2_X1 U7423 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  XNOR2_X1 U7424 ( .A(n5827), .B(n6173), .ZN(n7283) );
  INV_X1 U7425 ( .A(n7283), .ZN(n7327) );
  NAND2_X1 U7426 ( .A1(n8892), .A2(n7615), .ZN(n5829) );
  NAND2_X1 U7427 ( .A1(n7031), .A2(n6097), .ZN(n5828) );
  INV_X1 U7428 ( .A(n7285), .ZN(n5830) );
  NAND2_X1 U7429 ( .A1(n7327), .A2(n5830), .ZN(n5831) );
  NAND2_X1 U7430 ( .A1(n7329), .A2(n5831), .ZN(n5836) );
  NAND3_X1 U7431 ( .A1(n7329), .A2(n7285), .A3(n7283), .ZN(n5834) );
  NAND2_X1 U7432 ( .A1(n5833), .A2(n5832), .ZN(n7328) );
  AND2_X1 U7433 ( .A1(n5834), .A2(n7328), .ZN(n5835) );
  NAND2_X1 U7434 ( .A1(n6294), .A2(n8730), .ZN(n5840) );
  NOR2_X1 U7435 ( .A1(n5837), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5874) );
  OR2_X1 U7436 ( .A1(n5874), .A2(n5838), .ZN(n5855) );
  XNOR2_X1 U7437 ( .A(n5855), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7438 ( .A1(n6021), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6020), .B2(
        n6606), .ZN(n5839) );
  NAND2_X1 U7439 ( .A1(n7154), .A2(n4293), .ZN(n5849) );
  NAND2_X1 U7440 ( .A1(n4306), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5847) );
  INV_X1 U7441 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7062) );
  OR2_X1 U7442 ( .A1(n4308), .A2(n7062), .ZN(n5846) );
  INV_X1 U7443 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7444 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  NAND2_X1 U7445 ( .A1(n5881), .A2(n5843), .ZN(n7359) );
  OR2_X1 U7446 ( .A1(n6542), .A2(n7359), .ZN(n5845) );
  INV_X1 U7447 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6414) );
  OR2_X1 U7448 ( .A1(n8615), .A2(n6414), .ZN(n5844) );
  NAND4_X1 U7449 ( .A1(n5847), .A2(n5846), .A3(n5845), .A4(n5844), .ZN(n8890)
         );
  NAND2_X1 U7450 ( .A1(n8890), .A2(n6097), .ZN(n5848) );
  NAND2_X1 U7451 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  XNOR2_X1 U7452 ( .A(n5850), .B(n6173), .ZN(n5851) );
  NAND2_X1 U7453 ( .A1(n5852), .A2(n5851), .ZN(n7437) );
  AND2_X1 U7454 ( .A1(n8890), .A2(n7615), .ZN(n5853) );
  AOI21_X1 U7455 ( .B1(n7154), .B2(n6035), .A(n5853), .ZN(n7357) );
  NAND2_X1 U7456 ( .A1(n6375), .A2(n8730), .ZN(n5859) );
  INV_X1 U7457 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5854) );
  NAND2_X1 U7458 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  NAND2_X1 U7459 ( .A1(n5856), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5857) );
  XNOR2_X1 U7460 ( .A(n5857), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6733) );
  AOI22_X1 U7461 ( .A1(n6021), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6020), .B2(
        n6733), .ZN(n5858) );
  NAND2_X1 U7462 ( .A1(n7305), .A2(n4293), .ZN(n5865) );
  NAND2_X1 U7463 ( .A1(n4306), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5863) );
  INV_X1 U7464 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7163) );
  OR2_X1 U7465 ( .A1(n4308), .A2(n7163), .ZN(n5862) );
  INV_X1 U7466 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5880) );
  XNOR2_X1 U7467 ( .A(n5881), .B(n5880), .ZN(n7444) );
  OR2_X1 U7468 ( .A1(n6542), .A2(n7444), .ZN(n5861) );
  INV_X1 U7469 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6612) );
  OR2_X1 U7470 ( .A1(n8615), .A2(n6612), .ZN(n5860) );
  NAND4_X1 U7471 ( .A1(n5863), .A2(n5862), .A3(n5861), .A4(n5860), .ZN(n8889)
         );
  NAND2_X1 U7472 ( .A1(n8889), .A2(n6097), .ZN(n5864) );
  NAND2_X1 U7473 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  XNOR2_X1 U7474 ( .A(n5866), .B(n6173), .ZN(n5868) );
  AND2_X1 U7475 ( .A1(n8889), .A2(n7615), .ZN(n5867) );
  AOI21_X1 U7476 ( .B1(n7305), .B2(n6035), .A(n5867), .ZN(n5869) );
  NAND2_X1 U7477 ( .A1(n5868), .A2(n5869), .ZN(n7505) );
  INV_X1 U7478 ( .A(n5868), .ZN(n5871) );
  INV_X1 U7479 ( .A(n5869), .ZN(n5870) );
  NAND2_X1 U7480 ( .A1(n5871), .A2(n5870), .ZN(n5872) );
  AND2_X1 U7481 ( .A1(n7505), .A2(n5872), .ZN(n7438) );
  NAND2_X1 U7482 ( .A1(n6403), .A2(n8730), .ZN(n5877) );
  NOR2_X1 U7483 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5873) );
  NAND2_X1 U7484 ( .A1(n5874), .A2(n5873), .ZN(n5899) );
  NAND2_X1 U7485 ( .A1(n5899), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5875) );
  XNOR2_X1 U7486 ( .A(n5875), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6738) );
  AOI22_X1 U7487 ( .A1(n6021), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6020), .B2(
        n6738), .ZN(n5876) );
  NAND2_X1 U7488 ( .A1(n7510), .A2(n4293), .ZN(n5889) );
  NAND2_X1 U7489 ( .A1(n4307), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5887) );
  INV_X1 U7490 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7304) );
  OR2_X1 U7491 ( .A1(n4308), .A2(n7304), .ZN(n5886) );
  NAND2_X1 U7492 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n5878) );
  INV_X1 U7493 ( .A(n5903), .ZN(n5905) );
  INV_X1 U7494 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5879) );
  OAI21_X1 U7495 ( .B1(n5881), .B2(n5880), .A(n5879), .ZN(n5882) );
  NAND2_X1 U7496 ( .A1(n5905), .A2(n5882), .ZN(n7502) );
  OR2_X1 U7497 ( .A1(n6542), .A2(n7502), .ZN(n5885) );
  INV_X1 U7498 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5883) );
  OR2_X1 U7499 ( .A1(n8615), .A2(n5883), .ZN(n5884) );
  NAND4_X1 U7500 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n8888)
         );
  NAND2_X1 U7501 ( .A1(n8888), .A2(n6097), .ZN(n5888) );
  NAND2_X1 U7502 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  XNOR2_X1 U7503 ( .A(n5890), .B(n6173), .ZN(n5892) );
  AND2_X1 U7504 ( .A1(n8888), .A2(n7615), .ZN(n5891) );
  AOI21_X1 U7505 ( .B1(n7510), .B2(n6035), .A(n5891), .ZN(n5893) );
  NAND2_X1 U7506 ( .A1(n5892), .A2(n5893), .ZN(n5898) );
  INV_X1 U7507 ( .A(n5892), .ZN(n5895) );
  INV_X1 U7508 ( .A(n5893), .ZN(n5894) );
  NAND2_X1 U7509 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  AND2_X1 U7510 ( .A1(n5898), .A2(n5896), .ZN(n7503) );
  NAND2_X1 U7511 ( .A1(n5897), .A2(n7503), .ZN(n7507) );
  NAND2_X1 U7512 ( .A1(n7507), .A2(n5898), .ZN(n7513) );
  NAND2_X1 U7513 ( .A1(n6510), .A2(n8730), .ZN(n5902) );
  NAND2_X1 U7514 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X1 U7515 ( .A(n5900), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6958) );
  AOI22_X1 U7516 ( .A1(n6021), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6020), .B2(
        n6958), .ZN(n5901) );
  NAND2_X2 U7517 ( .A1(n5902), .A2(n5901), .ZN(n7400) );
  NAND2_X1 U7518 ( .A1(n7400), .A2(n4294), .ZN(n5913) );
  NAND2_X1 U7519 ( .A1(n4306), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5911) );
  INV_X1 U7520 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7394) );
  OR2_X1 U7521 ( .A1(n4309), .A2(n7394), .ZN(n5910) );
  NAND2_X1 U7522 ( .A1(n5903), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5945) );
  INV_X1 U7523 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7524 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  NAND2_X1 U7525 ( .A1(n5945), .A2(n5906), .ZN(n7516) );
  OR2_X1 U7526 ( .A1(n6542), .A2(n7516), .ZN(n5909) );
  INV_X1 U7527 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5907) );
  OR2_X1 U7528 ( .A1(n8615), .A2(n5907), .ZN(n5908) );
  NAND4_X1 U7529 ( .A1(n5911), .A2(n5910), .A3(n5909), .A4(n5908), .ZN(n8887)
         );
  NAND2_X1 U7530 ( .A1(n8887), .A2(n6097), .ZN(n5912) );
  NAND2_X1 U7531 ( .A1(n5913), .A2(n5912), .ZN(n5914) );
  XNOR2_X1 U7532 ( .A(n5914), .B(n7618), .ZN(n5916) );
  AND2_X1 U7533 ( .A1(n8887), .A2(n7615), .ZN(n5915) );
  AOI21_X1 U7534 ( .B1(n7400), .B2(n6035), .A(n5915), .ZN(n5917) );
  XNOR2_X1 U7535 ( .A(n5916), .B(n5917), .ZN(n7514) );
  INV_X1 U7536 ( .A(n5916), .ZN(n5918) );
  NAND2_X1 U7537 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  NAND2_X1 U7538 ( .A1(n6619), .A2(n8730), .ZN(n5923) );
  OR2_X1 U7539 ( .A1(n5920), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7540 ( .A1(n5921), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5937) );
  XNOR2_X1 U7541 ( .A(n5937), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7143) );
  AOI22_X1 U7542 ( .A1(n6021), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6020), .B2(
        n7143), .ZN(n5922) );
  NAND2_X2 U7543 ( .A1(n5923), .A2(n5922), .ZN(n8476) );
  NAND2_X1 U7544 ( .A1(n8476), .A2(n4293), .ZN(n5929) );
  NAND2_X1 U7545 ( .A1(n4307), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5927) );
  INV_X1 U7546 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5943) );
  XNOR2_X1 U7547 ( .A(n5945), .B(n5943), .ZN(n8474) );
  OR2_X1 U7548 ( .A1(n6542), .A2(n8474), .ZN(n5926) );
  INV_X1 U7549 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7385) );
  OR2_X1 U7550 ( .A1(n4308), .A2(n7385), .ZN(n5925) );
  INV_X1 U7551 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6952) );
  OR2_X1 U7552 ( .A1(n8615), .A2(n6952), .ZN(n5924) );
  NAND4_X1 U7553 ( .A1(n5927), .A2(n5926), .A3(n5925), .A4(n5924), .ZN(n8886)
         );
  NAND2_X1 U7554 ( .A1(n8886), .A2(n6097), .ZN(n5928) );
  NAND2_X1 U7555 ( .A1(n5929), .A2(n5928), .ZN(n5930) );
  XNOR2_X1 U7556 ( .A(n5930), .B(n6173), .ZN(n5932) );
  INV_X1 U7557 ( .A(n5932), .ZN(n5931) );
  NAND2_X1 U7558 ( .A1(n8476), .A2(n6097), .ZN(n5935) );
  NAND2_X1 U7559 ( .A1(n8886), .A2(n7615), .ZN(n5934) );
  NAND2_X1 U7560 ( .A1(n5935), .A2(n5934), .ZN(n8470) );
  NAND2_X1 U7561 ( .A1(n6676), .A2(n8730), .ZN(n5941) );
  INV_X1 U7562 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7563 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7564 ( .A1(n5938), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5939) );
  XNOR2_X1 U7565 ( .A(n5939), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8912) );
  AOI22_X1 U7566 ( .A1(n6021), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6020), .B2(
        n8912), .ZN(n5940) );
  NAND2_X1 U7567 ( .A1(n9139), .A2(n4293), .ZN(n5953) );
  NAND2_X1 U7568 ( .A1(n4307), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5951) );
  INV_X1 U7569 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7469) );
  OR2_X1 U7570 ( .A1(n4308), .A2(n7469), .ZN(n5950) );
  INV_X1 U7571 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5942) );
  OAI21_X1 U7572 ( .B1(n5945), .B2(n5943), .A(n5942), .ZN(n5946) );
  NAND2_X1 U7573 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n5944) );
  NAND2_X1 U7574 ( .A1(n5946), .A2(n5964), .ZN(n8603) );
  OR2_X1 U7575 ( .A1(n6542), .A2(n8603), .ZN(n5949) );
  INV_X1 U7576 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5947) );
  OR2_X1 U7577 ( .A1(n8615), .A2(n5947), .ZN(n5948) );
  NAND4_X1 U7578 ( .A1(n5951), .A2(n5950), .A3(n5949), .A4(n5948), .ZN(n8885)
         );
  NAND2_X1 U7579 ( .A1(n8885), .A2(n6097), .ZN(n5952) );
  NAND2_X1 U7580 ( .A1(n5953), .A2(n5952), .ZN(n5954) );
  XNOR2_X1 U7581 ( .A(n5954), .B(n6173), .ZN(n5955) );
  NAND2_X1 U7582 ( .A1(n9139), .A2(n6097), .ZN(n5958) );
  NAND2_X1 U7583 ( .A1(n8885), .A2(n7615), .ZN(n5957) );
  NAND2_X1 U7584 ( .A1(n5958), .A2(n5957), .ZN(n8597) );
  NAND2_X1 U7585 ( .A1(n5961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7586 ( .A(n5962), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8934) );
  AOI22_X1 U7587 ( .A1(n6021), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6020), .B2(
        n8934), .ZN(n5963) );
  NAND2_X1 U7588 ( .A1(n4457), .A2(n4294), .ZN(n5972) );
  NAND2_X1 U7589 ( .A1(n4306), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5970) );
  INV_X1 U7590 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8915) );
  OR2_X1 U7591 ( .A1(n8615), .A2(n8915), .ZN(n5969) );
  INV_X1 U7592 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8927) );
  INV_X1 U7593 ( .A(n5986), .ZN(n5988) );
  NAND2_X1 U7594 ( .A1(n5964), .A2(n8927), .ZN(n5965) );
  NAND2_X1 U7595 ( .A1(n5988), .A2(n5965), .ZN(n9408) );
  OR2_X1 U7596 ( .A1(n6542), .A2(n9408), .ZN(n5968) );
  INV_X1 U7597 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5966) );
  OR2_X1 U7598 ( .A1(n4309), .A2(n5966), .ZN(n5967) );
  NAND4_X1 U7599 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n9141)
         );
  NAND2_X1 U7600 ( .A1(n9141), .A2(n6097), .ZN(n5971) );
  NAND2_X1 U7601 ( .A1(n5972), .A2(n5971), .ZN(n5973) );
  XNOR2_X1 U7602 ( .A(n5973), .B(n6173), .ZN(n5975) );
  AND2_X1 U7603 ( .A1(n9141), .A2(n7615), .ZN(n5974) );
  AOI21_X1 U7604 ( .B1(n4457), .B2(n7620), .A(n5974), .ZN(n5976) );
  NAND2_X1 U7605 ( .A1(n5975), .A2(n5976), .ZN(n5980) );
  INV_X1 U7606 ( .A(n5975), .ZN(n5978) );
  INV_X1 U7607 ( .A(n5976), .ZN(n5977) );
  NAND2_X1 U7608 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  AND2_X1 U7609 ( .A1(n5980), .A2(n5979), .ZN(n8530) );
  NAND2_X1 U7610 ( .A1(n6748), .A2(n8730), .ZN(n5984) );
  NAND2_X1 U7611 ( .A1(n5981), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5982) );
  XNOR2_X1 U7612 ( .A(n5982), .B(P1_IR_REG_17__SCAN_IN), .ZN(n8957) );
  AOI22_X1 U7613 ( .A1(n6021), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6020), .B2(
        n8957), .ZN(n5983) );
  NAND2_X1 U7614 ( .A1(n9392), .A2(n4294), .ZN(n5995) );
  NAND2_X1 U7615 ( .A1(n4306), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5993) );
  INV_X1 U7616 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5985) );
  OR2_X1 U7617 ( .A1(n4309), .A2(n5985), .ZN(n5992) );
  INV_X1 U7618 ( .A(n6005), .ZN(n6006) );
  INV_X1 U7619 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7620 ( .A1(n5988), .A2(n5987), .ZN(n5989) );
  NAND2_X1 U7621 ( .A1(n6006), .A2(n5989), .ZN(n9393) );
  OR2_X1 U7622 ( .A1(n6542), .A2(n9393), .ZN(n5991) );
  INV_X1 U7623 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n8938) );
  OR2_X1 U7624 ( .A1(n8615), .A2(n8938), .ZN(n5990) );
  NAND4_X1 U7625 ( .A1(n5993), .A2(n5992), .A3(n5991), .A4(n5990), .ZN(n9144)
         );
  NAND2_X1 U7626 ( .A1(n9144), .A2(n6097), .ZN(n5994) );
  NAND2_X1 U7627 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  XNOR2_X1 U7628 ( .A(n5996), .B(n7618), .ZN(n5998) );
  AND2_X1 U7629 ( .A1(n9144), .A2(n7615), .ZN(n5997) );
  AOI21_X1 U7630 ( .B1(n9392), .B2(n6035), .A(n5997), .ZN(n5999) );
  XNOR2_X1 U7631 ( .A(n5998), .B(n5999), .ZN(n8538) );
  INV_X1 U7632 ( .A(n5998), .ZN(n6000) );
  NAND2_X1 U7633 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  NAND2_X1 U7634 ( .A1(n6825), .A2(n8730), .ZN(n6004) );
  XNOR2_X1 U7635 ( .A(n6002), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8971) );
  AOI22_X1 U7636 ( .A1(n6021), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6020), .B2(
        n8971), .ZN(n6003) );
  NAND2_X1 U7637 ( .A1(n9377), .A2(n4294), .ZN(n6013) );
  NAND2_X1 U7638 ( .A1(n6218), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6011) );
  INV_X1 U7639 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9536) );
  OR2_X1 U7640 ( .A1(n5736), .A2(n9536), .ZN(n6010) );
  NAND2_X1 U7641 ( .A1(n6005), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6025) );
  INV_X1 U7642 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U7643 ( .A1(n6006), .A2(n8955), .ZN(n6007) );
  NAND2_X1 U7644 ( .A1(n6025), .A2(n6007), .ZN(n9378) );
  OR2_X1 U7645 ( .A1(n6542), .A2(n9378), .ZN(n6009) );
  INV_X1 U7646 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9379) );
  OR2_X1 U7647 ( .A1(n4308), .A2(n9379), .ZN(n6008) );
  NAND4_X1 U7648 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n9147)
         );
  NAND2_X1 U7649 ( .A1(n9147), .A2(n6097), .ZN(n6012) );
  NAND2_X1 U7650 ( .A1(n6013), .A2(n6012), .ZN(n6014) );
  XNOR2_X1 U7651 ( .A(n6014), .B(n6173), .ZN(n6017) );
  INV_X1 U7652 ( .A(n6017), .ZN(n6015) );
  AND2_X1 U7653 ( .A1(n9147), .A2(n7615), .ZN(n6016) );
  AOI21_X1 U7654 ( .B1(n9377), .B2(n7620), .A(n6016), .ZN(n8575) );
  NAND2_X1 U7655 ( .A1(n8574), .A2(n8575), .ZN(n6019) );
  NAND2_X1 U7656 ( .A1(n6018), .A2(n6017), .ZN(n8573) );
  NAND2_X1 U7657 ( .A1(n6946), .A2(n8730), .ZN(n6023) );
  AOI22_X1 U7658 ( .A1(n6021), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n8980), .B2(
        n6020), .ZN(n6022) );
  NAND2_X1 U7659 ( .A1(n9356), .A2(n4293), .ZN(n6032) );
  NAND2_X1 U7660 ( .A1(n4307), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6030) );
  INV_X1 U7661 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9478) );
  OR2_X1 U7662 ( .A1(n8615), .A2(n9478), .ZN(n6029) );
  INV_X1 U7663 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7664 ( .A1(n6025), .A2(n6024), .ZN(n6026) );
  NAND2_X1 U7665 ( .A1(n6044), .A2(n6026), .ZN(n9357) );
  OR2_X1 U7666 ( .A1(n6542), .A2(n9357), .ZN(n6028) );
  INV_X1 U7667 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9358) );
  OR2_X1 U7668 ( .A1(n4309), .A2(n9358), .ZN(n6027) );
  NAND4_X1 U7669 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n9150)
         );
  NAND2_X1 U7670 ( .A1(n9150), .A2(n6097), .ZN(n6031) );
  NAND2_X1 U7671 ( .A1(n6032), .A2(n6031), .ZN(n6033) );
  XNOR2_X1 U7672 ( .A(n6033), .B(n6173), .ZN(n6036) );
  AND2_X1 U7673 ( .A1(n9150), .A2(n7615), .ZN(n6034) );
  AOI21_X1 U7674 ( .B1(n9356), .B2(n6035), .A(n6034), .ZN(n6037) );
  INV_X1 U7675 ( .A(n6036), .ZN(n6039) );
  INV_X1 U7676 ( .A(n6037), .ZN(n6038) );
  NAND2_X1 U7677 ( .A1(n6039), .A2(n6038), .ZN(n8503) );
  NAND2_X1 U7678 ( .A1(n7012), .A2(n8730), .ZN(n6041) );
  OR2_X1 U7679 ( .A1(n8729), .A2(n7015), .ZN(n6040) );
  NAND2_X1 U7680 ( .A1(n9471), .A2(n4293), .ZN(n6052) );
  NAND2_X1 U7681 ( .A1(n6218), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n6050) );
  INV_X1 U7682 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7683 ( .A1(n5736), .A2(n6042), .ZN(n6049) );
  INV_X1 U7684 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6043) );
  INV_X1 U7685 ( .A(n6060), .ZN(n6061) );
  NAND2_X1 U7686 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NAND2_X1 U7687 ( .A1(n6061), .A2(n6045), .ZN(n9334) );
  OR2_X1 U7688 ( .A1(n6542), .A2(n9334), .ZN(n6048) );
  INV_X1 U7689 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7690 ( .A1(n4309), .A2(n6046), .ZN(n6047) );
  NAND4_X1 U7691 ( .A1(n6050), .A2(n6049), .A3(n6048), .A4(n6047), .ZN(n9153)
         );
  NAND2_X1 U7692 ( .A1(n9153), .A2(n6097), .ZN(n6051) );
  NAND2_X1 U7693 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  XNOR2_X1 U7694 ( .A(n6053), .B(n6173), .ZN(n6056) );
  AND2_X1 U7695 ( .A1(n9153), .A2(n7615), .ZN(n6054) );
  AOI21_X1 U7696 ( .B1(n9471), .B2(n7620), .A(n6054), .ZN(n6055) );
  XNOR2_X1 U7697 ( .A(n6056), .B(n6055), .ZN(n8557) );
  NAND2_X1 U7698 ( .A1(n6056), .A2(n6055), .ZN(n6057) );
  NAND2_X1 U7699 ( .A1(n7018), .A2(n8730), .ZN(n6059) );
  OR2_X1 U7700 ( .A1(n8729), .A2(n7040), .ZN(n6058) );
  NAND2_X1 U7701 ( .A1(n9323), .A2(n4294), .ZN(n6069) );
  INV_X1 U7702 ( .A(n6077), .ZN(n6087) );
  INV_X1 U7703 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U7704 ( .A1(n6061), .A2(n8513), .ZN(n6062) );
  AND2_X1 U7705 ( .A1(n6087), .A2(n6062), .ZN(n9324) );
  NAND2_X1 U7706 ( .A1(n6144), .A2(n9324), .ZN(n6067) );
  NAND2_X1 U7707 ( .A1(n4306), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6066) );
  INV_X1 U7708 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9468) );
  OR2_X1 U7709 ( .A1(n8615), .A2(n9468), .ZN(n6065) );
  INV_X1 U7710 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6063) );
  OR2_X1 U7711 ( .A1(n4308), .A2(n6063), .ZN(n6064) );
  NAND4_X1 U7712 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n9155)
         );
  NAND2_X1 U7713 ( .A1(n9155), .A2(n6097), .ZN(n6068) );
  NAND2_X1 U7714 ( .A1(n6069), .A2(n6068), .ZN(n6070) );
  XNOR2_X1 U7715 ( .A(n6070), .B(n7618), .ZN(n6072) );
  AND2_X1 U7716 ( .A1(n9155), .A2(n7615), .ZN(n6071) );
  AOI21_X1 U7717 ( .B1(n9323), .B2(n7620), .A(n6071), .ZN(n6073) );
  XNOR2_X1 U7718 ( .A(n6072), .B(n6073), .ZN(n8512) );
  INV_X1 U7719 ( .A(n6072), .ZN(n6074) );
  NAND2_X1 U7720 ( .A1(n7193), .A2(n8730), .ZN(n6076) );
  OR2_X1 U7721 ( .A1(n8729), .A2(n7192), .ZN(n6075) );
  NAND2_X1 U7722 ( .A1(n9291), .A2(n4293), .ZN(n6082) );
  INV_X1 U7723 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9292) );
  NAND2_X1 U7724 ( .A1(n6077), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6089) );
  INV_X1 U7725 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8488) );
  NAND2_X1 U7726 ( .A1(n6089), .A2(n8488), .ZN(n6078) );
  NAND2_X1 U7727 ( .A1(n6111), .A2(n6078), .ZN(n9282) );
  OR2_X1 U7728 ( .A1(n9282), .A2(n6542), .ZN(n6080) );
  AOI22_X1 U7729 ( .A1(n4307), .A2(P1_REG0_REG_23__SCAN_IN), .B1(n6218), .B2(
        P1_REG1_REG_23__SCAN_IN), .ZN(n6079) );
  OAI211_X1 U7730 ( .C1(n4309), .C2(n9292), .A(n6080), .B(n6079), .ZN(n9160)
         );
  NAND2_X1 U7731 ( .A1(n9160), .A2(n6097), .ZN(n6081) );
  NAND2_X1 U7732 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  XNOR2_X1 U7733 ( .A(n6083), .B(n7618), .ZN(n8481) );
  INV_X1 U7734 ( .A(n9160), .ZN(n8695) );
  OAI22_X1 U7735 ( .A1(n9522), .A2(n6139), .B1(n8695), .B2(n6138), .ZN(n8480)
         );
  NAND2_X1 U7736 ( .A1(n8481), .A2(n8480), .ZN(n8479) );
  INV_X1 U7737 ( .A(n8479), .ZN(n6101) );
  NAND2_X1 U7738 ( .A1(n7188), .A2(n8730), .ZN(n6085) );
  OR2_X1 U7739 ( .A1(n8729), .A2(n7604), .ZN(n6084) );
  NAND2_X1 U7740 ( .A1(n9307), .A2(n4293), .ZN(n6095) );
  INV_X1 U7741 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9463) );
  INV_X1 U7742 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7743 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7744 ( .A1(n6089), .A2(n6088), .ZN(n9308) );
  OR2_X1 U7745 ( .A1(n9308), .A2(n6542), .ZN(n6093) );
  INV_X1 U7746 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9524) );
  OR2_X1 U7747 ( .A1(n5736), .A2(n9524), .ZN(n6091) );
  OR2_X1 U7748 ( .A1(n4308), .A2(n9026), .ZN(n6090) );
  AND2_X1 U7749 ( .A1(n6091), .A2(n6090), .ZN(n6092) );
  OAI211_X1 U7750 ( .C1(n8615), .C2(n9463), .A(n6093), .B(n6092), .ZN(n9157)
         );
  NAND2_X1 U7751 ( .A1(n9157), .A2(n6097), .ZN(n6094) );
  NAND2_X1 U7752 ( .A1(n6095), .A2(n6094), .ZN(n6096) );
  NAND2_X1 U7753 ( .A1(n9307), .A2(n6097), .ZN(n6099) );
  NAND2_X1 U7754 ( .A1(n9157), .A2(n7615), .ZN(n6098) );
  NAND2_X1 U7755 ( .A1(n8482), .A2(n6102), .ZN(n6108) );
  INV_X1 U7756 ( .A(n8480), .ZN(n6104) );
  AOI21_X1 U7757 ( .B1(n8484), .B2(n8483), .A(n6104), .ZN(n6103) );
  NAND3_X1 U7758 ( .A1(n6104), .A2(n8483), .A3(n8484), .ZN(n6105) );
  NAND2_X1 U7759 ( .A1(n6108), .A2(n6107), .ZN(n8546) );
  NAND2_X1 U7760 ( .A1(n7365), .A2(n8730), .ZN(n6110) );
  OR2_X1 U7761 ( .A1(n8729), .A2(n7368), .ZN(n6109) );
  NAND2_X2 U7762 ( .A1(n6110), .A2(n6109), .ZN(n9275) );
  NAND2_X1 U7763 ( .A1(n9275), .A2(n4294), .ZN(n6119) );
  INV_X1 U7764 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U7765 ( .A1(n6111), .A2(n8550), .ZN(n6112) );
  AND2_X1 U7766 ( .A1(n6129), .A2(n6112), .ZN(n9276) );
  NAND2_X1 U7767 ( .A1(n9276), .A2(n6144), .ZN(n6117) );
  INV_X1 U7768 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9516) );
  NAND2_X1 U7769 ( .A1(n6218), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7770 ( .A1(n6145), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6113) );
  OAI211_X1 U7771 ( .C1(n5736), .C2(n9516), .A(n6114), .B(n6113), .ZN(n6115)
         );
  INV_X1 U7772 ( .A(n6115), .ZN(n6116) );
  NAND2_X1 U7773 ( .A1(n6117), .A2(n6116), .ZN(n9162) );
  NAND2_X1 U7774 ( .A1(n9162), .A2(n6097), .ZN(n6118) );
  NAND2_X1 U7775 ( .A1(n6119), .A2(n6118), .ZN(n6120) );
  XNOR2_X1 U7776 ( .A(n6120), .B(n7618), .ZN(n6124) );
  NAND2_X1 U7777 ( .A1(n9275), .A2(n6097), .ZN(n6122) );
  NAND2_X1 U7778 ( .A1(n9162), .A2(n7615), .ZN(n6121) );
  NAND2_X1 U7779 ( .A1(n6122), .A2(n6121), .ZN(n6123) );
  AOI21_X1 U7780 ( .B1(n6124), .B2(n6123), .A(n6125), .ZN(n8547) );
  INV_X1 U7781 ( .A(n6125), .ZN(n6126) );
  NAND2_X1 U7782 ( .A1(n7416), .A2(n8730), .ZN(n6128) );
  OR2_X1 U7783 ( .A1(n8729), .A2(n7419), .ZN(n6127) );
  NAND2_X1 U7784 ( .A1(n9257), .A2(n4294), .ZN(n6136) );
  INV_X1 U7785 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8524) );
  AND2_X1 U7786 ( .A1(n6129), .A2(n8524), .ZN(n6130) );
  NOR2_X1 U7787 ( .A1(n6129), .A2(n8524), .ZN(n6142) );
  OR2_X1 U7788 ( .A1(n6130), .A2(n6142), .ZN(n8522) );
  INV_X1 U7789 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U7790 ( .A1(n6145), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7791 ( .A1(n6218), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6131) );
  OAI211_X1 U7792 ( .C1(n5736), .C2(n9511), .A(n6132), .B(n6131), .ZN(n6133)
         );
  INV_X1 U7793 ( .A(n6133), .ZN(n6134) );
  OAI21_X1 U7794 ( .B1(n8522), .B2(n6542), .A(n6134), .ZN(n9165) );
  NAND2_X1 U7795 ( .A1(n9165), .A2(n6097), .ZN(n6135) );
  NAND2_X1 U7796 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  XNOR2_X1 U7797 ( .A(n6137), .B(n6173), .ZN(n6155) );
  INV_X1 U7798 ( .A(n9165), .ZN(n8702) );
  OAI22_X1 U7799 ( .A1(n9514), .A2(n6139), .B1(n8702), .B2(n6138), .ZN(n6156)
         );
  XNOR2_X1 U7800 ( .A(n6155), .B(n6156), .ZN(n8519) );
  NAND2_X1 U7801 ( .A1(n7459), .A2(n8730), .ZN(n6141) );
  OR2_X1 U7802 ( .A1(n8729), .A2(n9560), .ZN(n6140) );
  NAND2_X1 U7803 ( .A1(n9241), .A2(n4293), .ZN(n6152) );
  OR2_X1 U7804 ( .A1(n6142), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6143) );
  NAND2_X1 U7805 ( .A1(n6142), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6165) );
  AND2_X1 U7806 ( .A1(n6143), .A2(n6165), .ZN(n9242) );
  NAND2_X1 U7807 ( .A1(n9242), .A2(n6144), .ZN(n6150) );
  INV_X1 U7808 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9509) );
  NAND2_X1 U7809 ( .A1(n6145), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7810 ( .A1(n6218), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6146) );
  OAI211_X1 U7811 ( .C1(n5736), .C2(n9509), .A(n6147), .B(n6146), .ZN(n6148)
         );
  INV_X1 U7812 ( .A(n6148), .ZN(n6149) );
  NAND2_X1 U7813 ( .A1(n6150), .A2(n6149), .ZN(n8884) );
  NAND2_X1 U7814 ( .A1(n8884), .A2(n6097), .ZN(n6151) );
  NAND2_X1 U7815 ( .A1(n6152), .A2(n6151), .ZN(n6153) );
  XNOR2_X1 U7816 ( .A(n6153), .B(n6173), .ZN(n6159) );
  AND2_X1 U7817 ( .A1(n8884), .A2(n7615), .ZN(n6154) );
  AOI21_X1 U7818 ( .B1(n9241), .B2(n7620), .A(n6154), .ZN(n6160) );
  XNOR2_X1 U7819 ( .A(n6159), .B(n6160), .ZN(n8584) );
  INV_X1 U7820 ( .A(n6155), .ZN(n6157) );
  NOR2_X1 U7821 ( .A1(n6157), .A2(n6156), .ZN(n8585) );
  INV_X1 U7822 ( .A(n6183), .ZN(n8587) );
  INV_X1 U7823 ( .A(n6159), .ZN(n6162) );
  INV_X1 U7824 ( .A(n6160), .ZN(n6161) );
  INV_X1 U7825 ( .A(n6180), .ZN(n6179) );
  NAND2_X1 U7826 ( .A1(n8463), .A2(n8730), .ZN(n6164) );
  OR2_X1 U7827 ( .A1(n8729), .A2(n9556), .ZN(n6163) );
  NAND2_X1 U7828 ( .A1(n9228), .A2(n4294), .ZN(n6172) );
  NAND2_X1 U7829 ( .A1(n6218), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6170) );
  INV_X1 U7830 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9505) );
  OR2_X1 U7831 ( .A1(n5736), .A2(n9505), .ZN(n6169) );
  INV_X1 U7832 ( .A(n6165), .ZN(n6220) );
  XNOR2_X1 U7833 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6220), .ZN(n6217) );
  OR2_X1 U7834 ( .A1(n6542), .A2(n6217), .ZN(n6168) );
  INV_X1 U7835 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7836 ( .A1(n4308), .A2(n6166), .ZN(n6167) );
  NAND4_X1 U7837 ( .A1(n6170), .A2(n6169), .A3(n6168), .A4(n6167), .ZN(n9169)
         );
  NAND2_X1 U7838 ( .A1(n9169), .A2(n6097), .ZN(n6171) );
  NAND2_X1 U7839 ( .A1(n6172), .A2(n6171), .ZN(n6174) );
  XNOR2_X1 U7840 ( .A(n6174), .B(n6173), .ZN(n6177) );
  AND2_X1 U7841 ( .A1(n9169), .A2(n7615), .ZN(n6175) );
  AOI21_X1 U7842 ( .B1(n9228), .B2(n7620), .A(n6175), .ZN(n6176) );
  NAND2_X1 U7843 ( .A1(n6177), .A2(n6176), .ZN(n7627) );
  OAI21_X1 U7844 ( .B1(n6177), .B2(n6176), .A(n7627), .ZN(n6181) );
  INV_X1 U7845 ( .A(n6181), .ZN(n6178) );
  AOI21_X1 U7846 ( .B1(n8587), .B2(n6179), .A(n6178), .ZN(n6210) );
  NOR2_X2 U7847 ( .A1(n6183), .A2(n6182), .ZN(n7634) );
  NAND2_X1 U7848 ( .A1(n7421), .A2(P1_B_REG_SCAN_IN), .ZN(n6184) );
  MUX2_X1 U7849 ( .A(P1_B_REG_SCAN_IN), .B(n6184), .S(n7370), .Z(n6186) );
  NAND2_X1 U7850 ( .A1(n6186), .A2(n6185), .ZN(n6271) );
  INV_X1 U7851 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7852 ( .A1(n6201), .A2(n6187), .ZN(n6188) );
  NAND2_X1 U7853 ( .A1(n9563), .A2(n7370), .ZN(n9544) );
  INV_X1 U7854 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7855 ( .A1(n9563), .A2(n7421), .ZN(n6272) );
  INV_X1 U7856 ( .A(n6272), .ZN(n6189) );
  AOI21_X1 U7857 ( .B1(n6201), .B2(n6190), .A(n6189), .ZN(n6762) );
  NOR4_X1 U7858 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6199) );
  NOR4_X1 U7859 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n6198) );
  INV_X1 U7860 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9761) );
  INV_X1 U7861 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n9759) );
  INV_X1 U7862 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9760) );
  INV_X1 U7863 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9762) );
  NAND4_X1 U7864 ( .A1(n9761), .A2(n9759), .A3(n9760), .A4(n9762), .ZN(n6196)
         );
  NOR4_X1 U7865 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6194) );
  NOR4_X1 U7866 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6193) );
  NOR4_X1 U7867 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6192) );
  NOR4_X1 U7868 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n6191) );
  NAND4_X1 U7869 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n6195)
         );
  NOR4_X1 U7870 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n6196), .A4(n6195), .ZN(n6197) );
  NAND3_X1 U7871 ( .A1(n6199), .A2(n6198), .A3(n6197), .ZN(n6200) );
  NAND2_X1 U7872 ( .A1(n6201), .A2(n6200), .ZN(n6473) );
  NAND3_X1 U7873 ( .A1(n6761), .A2(n6762), .A3(n6473), .ZN(n6214) );
  INV_X1 U7874 ( .A(n6214), .ZN(n6207) );
  NAND2_X1 U7875 ( .A1(n6203), .A2(n6202), .ZN(n6204) );
  NAND2_X1 U7876 ( .A1(n6204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6206) );
  XNOR2_X1 U7877 ( .A(n6206), .B(n6205), .ZN(n6279) );
  AND2_X1 U7878 ( .A1(n6207), .A2(n8877), .ZN(n6230) );
  NAND2_X1 U7879 ( .A1(n6784), .A2(n6231), .ZN(n9853) );
  INV_X1 U7880 ( .A(n8868), .ZN(n6208) );
  INV_X1 U7881 ( .A(n6465), .ZN(n8854) );
  AND2_X1 U7882 ( .A1(n9853), .A2(n8854), .ZN(n6209) );
  OAI21_X1 U7883 ( .B1(n6210), .B2(n7634), .A(n9649), .ZN(n6238) );
  NAND2_X1 U7884 ( .A1(n6214), .A2(n9853), .ZN(n6212) );
  NAND2_X1 U7885 ( .A1(n6465), .A2(n6231), .ZN(n6211) );
  AND3_X1 U7886 ( .A1(n6243), .A2(n6211), .A3(n6279), .ZN(n6472) );
  NAND2_X1 U7887 ( .A1(n6212), .A2(n6472), .ZN(n6213) );
  NAND2_X1 U7888 ( .A1(n6213), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6216) );
  AND2_X1 U7889 ( .A1(n6784), .A2(n8853), .ZN(n6234) );
  NAND3_X1 U7890 ( .A1(n6214), .A2(P1_STATE_REG_SCAN_IN), .A3(n6234), .ZN(
        n6215) );
  INV_X1 U7891 ( .A(n9674), .ZN(n8591) );
  INV_X1 U7892 ( .A(n6217), .ZN(n9229) );
  INV_X1 U7893 ( .A(n7611), .ZN(n6300) );
  AND2_X2 U7894 ( .A1(n6300), .A2(n6465), .ZN(n9199) );
  NAND2_X1 U7895 ( .A1(n6218), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6228) );
  INV_X1 U7896 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n6219) );
  OR2_X1 U7897 ( .A1(n5736), .A2(n6219), .ZN(n6227) );
  AND2_X1 U7898 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6220), .ZN(n6221) );
  NAND2_X1 U7899 ( .A1(n6221), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9175) );
  INV_X1 U7900 ( .A(n6221), .ZN(n6223) );
  INV_X1 U7901 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6222) );
  NAND2_X1 U7902 ( .A1(n6223), .A2(n6222), .ZN(n6224) );
  NAND2_X1 U7903 ( .A1(n9175), .A2(n6224), .ZN(n9211) );
  OR2_X1 U7904 ( .A1(n6542), .A2(n9211), .ZN(n6226) );
  INV_X1 U7905 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9215) );
  OR2_X1 U7906 ( .A1(n4309), .A2(n9215), .ZN(n6225) );
  NAND4_X1 U7907 ( .A1(n6228), .A2(n6227), .A3(n6226), .A4(n6225), .ZN(n9200)
         );
  AND2_X1 U7908 ( .A1(n7611), .A2(n6465), .ZN(n8577) );
  INV_X1 U7909 ( .A(n8577), .ZN(n6939) );
  AND2_X1 U7910 ( .A1(n9200), .A2(n8988), .ZN(n6229) );
  AOI21_X1 U7911 ( .B1(n8884), .B2(n9199), .A(n6229), .ZN(n9224) );
  INV_X1 U7912 ( .A(n6230), .ZN(n6235) );
  INV_X1 U7913 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n6232) );
  OAI22_X1 U7914 ( .A1(n9224), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6232), .ZN(n6233) );
  AOI21_X1 U7915 ( .B1(n8591), .B2(n9229), .A(n6233), .ZN(n6237) );
  INV_X1 U7916 ( .A(n6234), .ZN(n6765) );
  OR2_X1 U7917 ( .A1(n6235), .A2(n6765), .ZN(n6236) );
  NOR2_X1 U7918 ( .A1(n9767), .A2(n8786), .ZN(n6471) );
  NAND3_X1 U7919 ( .A1(n6238), .A2(n6237), .A3(n4898), .ZN(P1_U3214) );
  INV_X1 U7920 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7921 ( .A1(n6242), .A2(n4900), .ZN(P2_U3488) );
  NOR2_X1 U7922 ( .A1(n6243), .A2(P1_U3086), .ZN(n6244) );
  NAND2_X1 U7923 ( .A1(n7903), .A2(n6496), .ZN(n6245) );
  NAND2_X1 U7924 ( .A1(n6245), .A2(n6495), .ZN(n6429) );
  NAND2_X1 U7925 ( .A1(n6429), .A2(n6246), .ZN(n6247) );
  NAND2_X1 U7926 ( .A1(n6247), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U7927 ( .A(n6495), .ZN(n7194) );
  NOR2_X1 U7928 ( .A1(n6496), .A2(n7194), .ZN(n6424) );
  XNOR2_X1 U7929 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AND2_X1 U7930 ( .A1(n6249), .A2(P2_U3151), .ZN(n8465) );
  OR2_X1 U7931 ( .A1(n6249), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8467) );
  INV_X1 U7932 ( .A(n4295), .ZN(n6561) );
  OAI222_X1 U7933 ( .A1(n8456), .A2(n6248), .B1(n8467), .B2(n6251), .C1(
        P2_U3151), .C2(n6561), .ZN(P2_U3293) );
  NAND2_X1 U7934 ( .A1(n7747), .A2(P1_U3086), .ZN(n9551) );
  OR2_X1 U7935 ( .A1(n7747), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9554) );
  OAI222_X1 U7936 ( .A1(n6657), .A2(P1_U3086), .B1(n9551), .B2(n6251), .C1(
        n6250), .C2(n9554), .ZN(P1_U3353) );
  OAI222_X1 U7937 ( .A1(n6329), .A2(P1_U3086), .B1(n9551), .B2(n6256), .C1(
        n6252), .C2(n9554), .ZN(P1_U3352) );
  INV_X1 U7938 ( .A(n9554), .ZN(n6826) );
  INV_X1 U7939 ( .A(n6826), .ZN(n9559) );
  OAI222_X1 U7940 ( .A1(n9559), .A2(n9102), .B1(n9551), .B2(n6254), .C1(n6689), 
        .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U7941 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6253) );
  OAI222_X1 U7942 ( .A1(n8456), .A2(n6253), .B1(n8467), .B2(n6261), .C1(
        P2_U3151), .C2(n6435), .ZN(P2_U3294) );
  INV_X1 U7943 ( .A(n8467), .ZN(n8458) );
  INV_X1 U7944 ( .A(n8458), .ZN(n8457) );
  OAI222_X1 U7945 ( .A1(n8456), .A2(n6255), .B1(n8457), .B2(n6254), .C1(
        P2_U3151), .C2(n6577), .ZN(P2_U3291) );
  OAI222_X1 U7946 ( .A1(n8456), .A2(n6257), .B1(n8457), .B2(n6256), .C1(
        P2_U3151), .C2(n9888), .ZN(P2_U3292) );
  OAI222_X1 U7947 ( .A1(n6398), .A2(P1_U3086), .B1(n9551), .B2(n6259), .C1(
        n6258), .C2(n9554), .ZN(P1_U3350) );
  OAI222_X1 U7948 ( .A1(n8456), .A2(n6260), .B1(n8467), .B2(n6259), .C1(
        P2_U3151), .C2(n9928), .ZN(P2_U3290) );
  INV_X1 U7949 ( .A(n9551), .ZN(n7190) );
  INV_X1 U7950 ( .A(n7190), .ZN(n9562) );
  OAI222_X1 U7951 ( .A1(n6305), .A2(P1_U3086), .B1(n9562), .B2(n6261), .C1(
        n4461), .C2(n9554), .ZN(P1_U3354) );
  OAI222_X1 U7952 ( .A1(n6347), .A2(P1_U3086), .B1(n9551), .B2(n6263), .C1(
        n6262), .C2(n9554), .ZN(P1_U3349) );
  OAI222_X1 U7953 ( .A1(n8456), .A2(n6264), .B1(n8457), .B2(n6263), .C1(
        P2_U3151), .C2(n6900), .ZN(P2_U3289) );
  OAI222_X1 U7954 ( .A1(n8456), .A2(n6265), .B1(n8467), .B2(n6267), .C1(
        P2_U3151), .C2(n9942), .ZN(P2_U3288) );
  OAI222_X1 U7955 ( .A1(n6372), .A2(P1_U3086), .B1(n9551), .B2(n6267), .C1(
        n6266), .C2(n9554), .ZN(P1_U3348) );
  INV_X1 U7956 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7957 ( .A1(n6268), .A2(n6284), .ZN(n6269) );
  OAI21_X1 U7958 ( .B1(n6284), .B2(n6270), .A(n6269), .ZN(P2_U3377) );
  NAND2_X1 U7959 ( .A1(n9763), .A2(n6272), .ZN(n6273) );
  OAI21_X1 U7960 ( .B1(n9763), .B2(n6190), .A(n6273), .ZN(P1_U3440) );
  INV_X1 U7961 ( .A(n6274), .ZN(n6277) );
  INV_X1 U7962 ( .A(n7079), .ZN(n6909) );
  OAI222_X1 U7963 ( .A1(n8456), .A2(n6275), .B1(n8457), .B2(n6277), .C1(
        P2_U3151), .C2(n6909), .ZN(P2_U3287) );
  INV_X1 U7964 ( .A(n6352), .ZN(n6387) );
  OAI222_X1 U7965 ( .A1(n6387), .A2(P1_U3086), .B1(n9551), .B2(n6277), .C1(
        n6276), .C2(n9554), .ZN(P1_U3347) );
  INV_X1 U7966 ( .A(n8877), .ZN(n6278) );
  OR2_X1 U7967 ( .A1(n6279), .A2(P1_U3086), .ZN(n8882) );
  NAND2_X1 U7968 ( .A1(n6278), .A2(n8882), .ZN(n6299) );
  NAND2_X1 U7969 ( .A1(n6465), .A2(n6279), .ZN(n6280) );
  AND2_X1 U7970 ( .A1(n6281), .A2(n6280), .ZN(n6298) );
  INV_X1 U7971 ( .A(n6298), .ZN(n6282) );
  AND2_X1 U7972 ( .A1(n6299), .A2(n6282), .ZN(n9679) );
  NOR2_X1 U7973 ( .A1(n9679), .A2(P1_U3973), .ZN(P1_U3085) );
  NAND2_X1 U7974 ( .A1(n6284), .A2(n6283), .ZN(n6292) );
  NOR4_X1 U7975 ( .A1(n6286), .A2(n6285), .A3(n7194), .A4(P2_U3151), .ZN(n6287) );
  AOI21_X1 U7976 ( .B1(n6292), .B2(n5517), .A(n6287), .ZN(P2_U3376) );
  AND2_X1 U7977 ( .A1(n6292), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7978 ( .A1(n6292), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7979 ( .A1(n6292), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7980 ( .A1(n6292), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7981 ( .A1(n6292), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7982 ( .A1(n6292), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7983 ( .A1(n6292), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7984 ( .A1(n6292), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7985 ( .A1(n6292), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7986 ( .A1(n6292), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7987 ( .A1(n6292), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7988 ( .A1(n6292), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7989 ( .A1(n6292), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7990 ( .A1(n6292), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7991 ( .A1(n6292), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7992 ( .A1(n6292), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U7993 ( .A1(n6292), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7994 ( .A1(n6292), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7995 ( .A1(n6292), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7996 ( .A1(n6292), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7997 ( .A1(n6292), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7998 ( .A1(n6292), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7999 ( .A1(n6292), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8000 ( .A1(n6292), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8001 ( .A1(n6292), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8002 ( .A1(n6292), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8003 ( .A(n6288), .ZN(n6291) );
  OAI222_X1 U8004 ( .A1(n8457), .A2(n6291), .B1(n7082), .B2(P2_U3151), .C1(
        n6289), .C2(n8456), .ZN(P2_U3286) );
  INV_X1 U8005 ( .A(n6411), .ZN(n6341) );
  OAI222_X1 U8006 ( .A1(P1_U3086), .A2(n6341), .B1(n9551), .B2(n6291), .C1(
        n6290), .C2(n9554), .ZN(P1_U3346) );
  INV_X1 U8007 ( .A(n6292), .ZN(n6293) );
  INV_X1 U8008 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n9037) );
  NOR2_X1 U8009 ( .A1(n6293), .A2(n9037), .ZN(P2_U3262) );
  INV_X1 U8010 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n9010) );
  NOR2_X1 U8011 ( .A1(n6293), .A2(n9010), .ZN(P2_U3236) );
  INV_X1 U8012 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n9009) );
  NOR2_X1 U8013 ( .A1(n6293), .A2(n9009), .ZN(P2_U3256) );
  INV_X1 U8014 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n9044) );
  NOR2_X1 U8015 ( .A1(n6293), .A2(n9044), .ZN(P2_U3246) );
  INV_X1 U8016 ( .A(n6294), .ZN(n6297) );
  INV_X1 U8017 ( .A(n7093), .ZN(n7234) );
  OAI222_X1 U8018 ( .A1(n8457), .A2(n6297), .B1(n7234), .B2(P2_U3151), .C1(
        n6295), .C2(n8456), .ZN(P2_U3285) );
  INV_X1 U8019 ( .A(n6606), .ZN(n6611) );
  OAI222_X1 U8020 ( .A1(P1_U3086), .A2(n6611), .B1(n9551), .B2(n6297), .C1(
        n6296), .C2(n9554), .ZN(P1_U3345) );
  NAND2_X1 U8021 ( .A1(n6299), .A2(n6298), .ZN(n9681) );
  INV_X1 U8022 ( .A(n6657), .ZN(n6656) );
  XNOR2_X1 U8023 ( .A(n6305), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n8901) );
  AND2_X1 U8024 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n8900) );
  NAND2_X1 U8025 ( .A1(n8901), .A2(n8900), .ZN(n8899) );
  INV_X1 U8026 ( .A(n6305), .ZN(n8905) );
  NAND2_X1 U8027 ( .A1(n8905), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U8028 ( .A1(n8899), .A2(n6301), .ZN(n6654) );
  INV_X1 U8029 ( .A(n6653), .ZN(n6302) );
  AOI21_X1 U8030 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6656), .A(n6302), .ZN(
        n6304) );
  INV_X1 U8031 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6766) );
  XNOR2_X1 U8032 ( .A(n6329), .B(n6766), .ZN(n6303) );
  NOR2_X1 U8033 ( .A1(n6304), .A2(n6303), .ZN(n6330) );
  OR2_X1 U8034 ( .A1(n7611), .A2(n9677), .ZN(n8873) );
  AOI211_X1 U8035 ( .C1(n6304), .C2(n6303), .A(n6330), .B(n8960), .ZN(n6314)
         );
  INV_X1 U8036 ( .A(n9677), .ZN(n6648) );
  OR2_X1 U8037 ( .A1(n9681), .A2(n6648), .ZN(n9691) );
  MUX2_X1 U8038 ( .A(n6306), .B(P1_REG1_REG_1__SCAN_IN), .S(n6305), .Z(n8903)
         );
  AND2_X1 U8039 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n8904) );
  NAND2_X1 U8040 ( .A1(n8903), .A2(n8904), .ZN(n8902) );
  NAND2_X1 U8041 ( .A1(n8905), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6659) );
  NAND2_X1 U8042 ( .A1(n8902), .A2(n6659), .ZN(n6309) );
  MUX2_X1 U8043 ( .A(n6307), .B(P1_REG1_REG_2__SCAN_IN), .S(n6657), .Z(n6308)
         );
  NAND2_X1 U8044 ( .A1(n6309), .A2(n6308), .ZN(n6661) );
  NAND2_X1 U8045 ( .A1(n6656), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6310) );
  MUX2_X1 U8046 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6321), .S(n6329), .Z(n6311)
         );
  AOI21_X1 U8047 ( .B1(n6661), .B2(n6310), .A(n6311), .ZN(n6319) );
  AND3_X1 U8048 ( .A1(n6661), .A2(n6311), .A3(n6310), .ZN(n6312) );
  NOR3_X1 U8049 ( .A1(n9691), .A2(n6319), .A3(n6312), .ZN(n6313) );
  NOR2_X1 U8050 ( .A1(n6314), .A2(n6313), .ZN(n6317) );
  AND2_X1 U8051 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6315) );
  AOI21_X1 U8052 ( .B1(n9679), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6315), .ZN(
        n6316) );
  OAI211_X1 U8053 ( .C1(n6329), .C2(n9689), .A(n6317), .B(n6316), .ZN(P1_U3246) );
  NAND2_X1 U8054 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6333), .ZN(n6324) );
  MUX2_X1 U8055 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6318), .S(n6333), .Z(n6393)
         );
  INV_X1 U8056 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6323) );
  MUX2_X1 U8057 ( .A(n6323), .B(P1_REG1_REG_4__SCAN_IN), .S(n6689), .Z(n6694)
         );
  INV_X1 U8058 ( .A(n6319), .ZN(n6320) );
  OAI21_X1 U8059 ( .B1(n6321), .B2(n6329), .A(n6320), .ZN(n6693) );
  NAND2_X1 U8060 ( .A1(n6694), .A2(n6693), .ZN(n6322) );
  OAI21_X1 U8061 ( .B1(n6689), .B2(n6323), .A(n6322), .ZN(n6394) );
  NAND2_X1 U8062 ( .A1(n6393), .A2(n6394), .ZN(n6392) );
  AND2_X1 U8063 ( .A1(n6324), .A2(n6392), .ZN(n6326) );
  INV_X1 U8064 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9868) );
  MUX2_X1 U8065 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9868), .S(n6347), .Z(n6325)
         );
  NOR2_X1 U8066 ( .A1(n6326), .A2(n6325), .ZN(n6366) );
  AOI211_X1 U8067 ( .C1(n6326), .C2(n6325), .A(n6366), .B(n9691), .ZN(n6327)
         );
  INV_X1 U8068 ( .A(n6327), .ZN(n6340) );
  NOR2_X1 U8069 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6328), .ZN(n6338) );
  INV_X1 U8070 ( .A(n6689), .ZN(n6331) );
  INV_X1 U8071 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6808) );
  XNOR2_X1 U8072 ( .A(n6689), .B(n6808), .ZN(n6691) );
  NAND2_X1 U8073 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6333), .ZN(n6332) );
  OAI21_X1 U8074 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6333), .A(n6332), .ZN(
        n6390) );
  AOI21_X1 U8075 ( .B1(n6333), .B2(P1_REG2_REG_5__SCAN_IN), .A(n4350), .ZN(
        n6336) );
  MUX2_X1 U8076 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6334), .S(n6347), .Z(n6335)
         );
  NOR2_X1 U8077 ( .A1(n6336), .A2(n6335), .ZN(n6348) );
  AOI211_X1 U8078 ( .C1(n6336), .C2(n6335), .A(n6348), .B(n8960), .ZN(n6337)
         );
  AOI211_X1 U8079 ( .C1(n9679), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n6338), .B(
        n6337), .ZN(n6339) );
  OAI211_X1 U8080 ( .C1(n9689), .C2(n6347), .A(n6340), .B(n6339), .ZN(P1_U3249) );
  AOI22_X1 U8081 ( .A1(n6411), .A2(n5803), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n6341), .ZN(n6345) );
  MUX2_X1 U8082 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6342), .S(n6352), .Z(n6382)
         );
  NOR2_X1 U8083 ( .A1(n6347), .A2(n9868), .ZN(n6365) );
  MUX2_X1 U8084 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6343), .S(n6350), .Z(n6364)
         );
  OAI21_X1 U8085 ( .B1(n6366), .B2(n6365), .A(n6364), .ZN(n6368) );
  OAI21_X1 U8086 ( .B1(n6343), .B2(n6372), .A(n6368), .ZN(n6383) );
  NAND2_X1 U8087 ( .A1(n6382), .A2(n6383), .ZN(n6381) );
  OAI21_X1 U8088 ( .B1(n6387), .B2(n6342), .A(n6381), .ZN(n6344) );
  NOR2_X1 U8089 ( .A1(n6345), .A2(n6344), .ZN(n6413) );
  AOI21_X1 U8090 ( .B1(n6345), .B2(n6344), .A(n6413), .ZN(n6360) );
  NOR2_X1 U8091 ( .A1(n6411), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6346) );
  AOI21_X1 U8092 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n6411), .A(n6346), .ZN(
        n6354) );
  INV_X1 U8093 ( .A(n6347), .ZN(n6349) );
  AOI21_X1 U8094 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6349), .A(n6348), .ZN(
        n6363) );
  AOI22_X1 U8095 ( .A1(n6350), .A2(n7005), .B1(P1_REG2_REG_7__SCAN_IN), .B2(
        n6372), .ZN(n6362) );
  NOR2_X1 U8096 ( .A1(n6363), .A2(n6362), .ZN(n6361) );
  NAND2_X1 U8097 ( .A1(P1_REG2_REG_8__SCAN_IN), .A2(n6352), .ZN(n6351) );
  OAI21_X1 U8098 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n6352), .A(n6351), .ZN(
        n6379) );
  OAI21_X1 U8099 ( .B1(n6354), .B2(n6353), .A(n6408), .ZN(n6355) );
  INV_X1 U8100 ( .A(n8960), .ZN(n9695) );
  NAND2_X1 U8101 ( .A1(n6355), .A2(n9695), .ZN(n6359) );
  INV_X1 U8102 ( .A(n9689), .ZN(n8906) );
  INV_X1 U8103 ( .A(n9679), .ZN(n9699) );
  INV_X1 U8104 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8105 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7335) );
  OAI21_X1 U8106 ( .B1(n9699), .B2(n6356), .A(n7335), .ZN(n6357) );
  AOI21_X1 U8107 ( .B1(n6411), .B2(n8906), .A(n6357), .ZN(n6358) );
  OAI211_X1 U8108 ( .C1(n6360), .C2(n9691), .A(n6359), .B(n6358), .ZN(P1_U3252) );
  AOI211_X1 U8109 ( .C1(n6363), .C2(n6362), .A(n6361), .B(n8960), .ZN(n6374)
         );
  OR3_X1 U8110 ( .A1(n6366), .A2(n6365), .A3(n6364), .ZN(n6367) );
  NAND3_X1 U8111 ( .A1(n8975), .A2(n6368), .A3(n6367), .ZN(n6371) );
  NOR2_X1 U8112 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5779), .ZN(n6369) );
  AOI21_X1 U8113 ( .B1(n9679), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6369), .ZN(
        n6370) );
  OAI211_X1 U8114 ( .C1(n9689), .C2(n6372), .A(n6371), .B(n6370), .ZN(n6373)
         );
  OR2_X1 U8115 ( .A1(n6374), .A2(n6373), .ZN(P1_U3250) );
  INV_X1 U8116 ( .A(n6375), .ZN(n6377) );
  OAI222_X1 U8117 ( .A1(n8456), .A2(n9103), .B1(n8467), .B2(n6377), .C1(
        P2_U3151), .C2(n4511), .ZN(P2_U3284) );
  INV_X1 U8118 ( .A(n6733), .ZN(n6737) );
  OAI222_X1 U8119 ( .A1(n6737), .A2(P1_U3086), .B1(n9551), .B2(n6377), .C1(
        n6376), .C2(n9554), .ZN(P1_U3344) );
  AOI211_X1 U8120 ( .C1(n6380), .C2(n6379), .A(n6378), .B(n8960), .ZN(n6389)
         );
  OAI211_X1 U8121 ( .C1(n6383), .C2(n6382), .A(n8975), .B(n6381), .ZN(n6386)
         );
  NOR2_X1 U8122 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7289), .ZN(n6384) );
  AOI21_X1 U8123 ( .B1(n9679), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n6384), .ZN(
        n6385) );
  OAI211_X1 U8124 ( .C1(n9689), .C2(n6387), .A(n6386), .B(n6385), .ZN(n6388)
         );
  OR2_X1 U8125 ( .A1(n6389), .A2(n6388), .ZN(P1_U3251) );
  AOI211_X1 U8126 ( .C1(n6391), .C2(n6390), .A(n4350), .B(n8960), .ZN(n6400)
         );
  OAI211_X1 U8127 ( .C1(n6394), .C2(n6393), .A(n8975), .B(n6392), .ZN(n6397)
         );
  AND2_X1 U8128 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6395) );
  AOI21_X1 U8129 ( .B1(n9679), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6395), .ZN(
        n6396) );
  OAI211_X1 U8130 ( .C1(n9689), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6399)
         );
  OR2_X1 U8131 ( .A1(n6400), .A2(n6399), .ZN(P1_U3248) );
  INV_X1 U8132 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U8133 ( .A1(n6771), .A2(P1_U3973), .ZN(n6401) );
  OAI21_X1 U8134 ( .B1(P1_U3973), .B2(n6402), .A(n6401), .ZN(P1_U3554) );
  INV_X1 U8135 ( .A(n6403), .ZN(n6405) );
  OAI222_X1 U8136 ( .A1(n8457), .A2(n6405), .B1(n8023), .B2(P2_U3151), .C1(
        n6404), .C2(n8456), .ZN(P2_U3283) );
  INV_X1 U8137 ( .A(n6738), .ZN(n9690) );
  OAI222_X1 U8138 ( .A1(n9559), .A2(n6406), .B1(n9562), .B2(n6405), .C1(
        P1_U3086), .C2(n9690), .ZN(P1_U3343) );
  NAND2_X1 U8139 ( .A1(n6606), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6407) );
  OAI21_X1 U8140 ( .B1(n6606), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6407), .ZN(
        n6410) );
  OAI21_X1 U8141 ( .B1(n6411), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6408), .ZN(
        n6409) );
  NOR2_X1 U8142 ( .A1(n6410), .A2(n6409), .ZN(n6605) );
  AOI211_X1 U8143 ( .C1(n6410), .C2(n6409), .A(n6605), .B(n8960), .ZN(n6420)
         );
  NOR2_X1 U8144 ( .A1(n6411), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6412) );
  NOR2_X1 U8145 ( .A1(n6413), .A2(n6412), .ZN(n6416) );
  MUX2_X1 U8146 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6414), .S(n6606), .Z(n6415)
         );
  NAND2_X1 U8147 ( .A1(n6415), .A2(n6416), .ZN(n6610) );
  OAI211_X1 U8148 ( .C1(n6416), .C2(n6415), .A(n6610), .B(n8975), .ZN(n6418)
         );
  AND2_X1 U8149 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n7361) );
  AOI21_X1 U8150 ( .B1(n9679), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7361), .ZN(
        n6417) );
  OAI211_X1 U8151 ( .C1(n9689), .C2(n6611), .A(n6418), .B(n6417), .ZN(n6419)
         );
  OR2_X1 U8152 ( .A1(n6420), .A2(n6419), .ZN(P1_U3253) );
  NAND2_X1 U8153 ( .A1(P2_U3893), .A2(n6423), .ZN(n9917) );
  MUX2_X1 U8154 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6449), .Z(n6445) );
  XNOR2_X1 U8155 ( .A(n6445), .B(n6435), .ZN(n6448) );
  INV_X1 U8156 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9881) );
  MUX2_X1 U8157 ( .A(n9096), .B(n9881), .S(n6449), .Z(n6421) );
  AND2_X1 U8158 ( .A1(n6421), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n9884) );
  XNOR2_X1 U8159 ( .A(n6448), .B(n9884), .ZN(n6444) );
  OR2_X1 U8160 ( .A1(P2_U3150), .A2(n6424), .ZN(n9924) );
  INV_X4 U8161 ( .A(n8145), .ZN(n9882) );
  NOR2_X1 U8162 ( .A1(n9882), .A2(P2_U3151), .ZN(n8464) );
  AND2_X1 U8163 ( .A1(n8464), .A2(n6423), .ZN(n6422) );
  NAND2_X1 U8164 ( .A1(n6429), .A2(n6422), .ZN(n6426) );
  OR2_X1 U8165 ( .A1(n6423), .A2(P2_U3151), .ZN(n8460) );
  INV_X1 U8166 ( .A(n8460), .ZN(n6428) );
  NAND2_X1 U8167 ( .A1(n6428), .A2(n6424), .ZN(n6425) );
  NAND2_X1 U8168 ( .A1(n6426), .A2(n6425), .ZN(n9914) );
  OAI22_X1 U8169 ( .A1(n9980), .A2(n6435), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6427), .ZN(n6442) );
  AND2_X1 U8170 ( .A1(n6429), .A2(n6428), .ZN(n9885) );
  INV_X1 U8171 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U8172 ( .A1(n6430), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U8173 ( .A1(n6431), .A2(n6454), .ZN(n6433) );
  OR2_X1 U8174 ( .A1(n6433), .A2(n6682), .ZN(n6455) );
  INV_X1 U8175 ( .A(n6455), .ZN(n6432) );
  AOI21_X1 U8176 ( .B1(n6682), .B2(n6433), .A(n6432), .ZN(n6440) );
  NOR2_X1 U8177 ( .A1(n9096), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6434) );
  NAND2_X1 U8178 ( .A1(n6430), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6450) );
  INV_X1 U8179 ( .A(n6451), .ZN(n6436) );
  AOI21_X1 U8180 ( .B1(n6793), .B2(n6437), .A(n6436), .ZN(n6439) );
  INV_X1 U8181 ( .A(n9885), .ZN(n6438) );
  OAI22_X1 U8182 ( .A1(n9974), .A2(n6440), .B1(n6439), .B2(n9965), .ZN(n6441)
         );
  AOI211_X1 U8183 ( .C1(n9959), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6442), .B(
        n6441), .ZN(n6443) );
  OAI21_X1 U8184 ( .B1(n9917), .B2(n6444), .A(n6443), .ZN(P2_U3183) );
  INV_X1 U8185 ( .A(n6445), .ZN(n6446) );
  OAI22_X1 U8186 ( .A1(n6448), .A2(n9884), .B1(n6447), .B2(n6446), .ZN(n6556)
         );
  MUX2_X1 U8187 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6449), .Z(n6554) );
  XNOR2_X1 U8188 ( .A(n6554), .B(n4295), .ZN(n6555) );
  XNOR2_X1 U8189 ( .A(n6556), .B(n6555), .ZN(n6463) );
  INV_X1 U8190 ( .A(n9965), .ZN(n6584) );
  NAND2_X1 U8191 ( .A1(n6451), .A2(n6450), .ZN(n6452) );
  OAI21_X1 U8192 ( .B1(n6453), .B2(n6452), .A(n6563), .ZN(n6458) );
  NAND2_X1 U8193 ( .A1(n6455), .A2(n6454), .ZN(n6456) );
  AOI22_X1 U8194 ( .A1(n6584), .A2(n6458), .B1(n9951), .B2(n6457), .ZN(n6460)
         );
  AOI22_X1 U8195 ( .A1(n9914), .A2(n4295), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n6459) );
  NAND2_X1 U8196 ( .A1(n6460), .A2(n6459), .ZN(n6461) );
  AOI21_X1 U8197 ( .B1(n9959), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n6461), .ZN(
        n6462) );
  OAI21_X1 U8198 ( .B1(n9917), .B2(n6463), .A(n6462), .ZN(P2_U3184) );
  NAND2_X1 U8199 ( .A1(n6752), .A2(n8988), .ZN(n6786) );
  INV_X1 U8200 ( .A(n6786), .ZN(n6470) );
  OR2_X1 U8201 ( .A1(n8868), .A2(n8866), .ZN(n6464) );
  NAND2_X1 U8202 ( .A1(n6464), .A2(n8870), .ZN(n9738) );
  NOR2_X1 U8203 ( .A1(n8868), .A2(n8980), .ZN(n6466) );
  NAND2_X1 U8204 ( .A1(n6465), .A2(n8834), .ZN(n8872) );
  OAI211_X1 U8205 ( .C1(n6466), .C2(n8834), .A(n6785), .B(n8872), .ZN(n7004)
         );
  INV_X1 U8206 ( .A(n6771), .ZN(n6467) );
  NAND2_X1 U8207 ( .A1(n6467), .A2(n6770), .ZN(n6867) );
  INV_X1 U8208 ( .A(n6770), .ZN(n6873) );
  NAND2_X1 U8209 ( .A1(n6771), .A2(n6873), .ZN(n8787) );
  NAND2_X1 U8210 ( .A1(n6867), .A2(n8787), .ZN(n8747) );
  INV_X1 U8211 ( .A(n8747), .ZN(n6468) );
  AOI21_X1 U8212 ( .B1(n9706), .B2(n9632), .A(n6468), .ZN(n6469) );
  AOI211_X1 U8213 ( .C1(n6770), .C2(n6784), .A(n6470), .B(n6469), .ZN(n9766)
         );
  OR2_X1 U8214 ( .A1(n6762), .A2(n6471), .ZN(n6474) );
  NAND3_X1 U8215 ( .A1(n6473), .A2(n6472), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n6760) );
  AND2_X2 U8216 ( .A1(n9491), .A2(n6761), .ZN(n9879) );
  NAND2_X1 U8217 ( .A1(n9877), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6475) );
  OAI21_X1 U8218 ( .B1(n9766), .B2(n9877), .A(n6475), .ZN(P1_U3522) );
  XOR2_X1 U8219 ( .A(n6477), .B(n6476), .Z(n6649) );
  AND2_X1 U8220 ( .A1(n9674), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6675) );
  NOR2_X1 U8221 ( .A1(n6675), .A2(n5661), .ZN(n6479) );
  OAI22_X1 U8222 ( .A1(n8594), .A2(n6873), .B1(n6786), .B2(n9660), .ZN(n6478)
         );
  AOI211_X1 U8223 ( .C1(n6649), .C2(n9649), .A(n6479), .B(n6478), .ZN(n6480)
         );
  INV_X1 U8224 ( .A(n6480), .ZN(P1_U3232) );
  NAND2_X1 U8225 ( .A1(n6486), .A2(n10073), .ZN(n6482) );
  NAND2_X1 U8226 ( .A1(n6482), .A2(n10002), .ZN(n7721) );
  INV_X1 U8227 ( .A(n7721), .ZN(n7737) );
  INV_X1 U8228 ( .A(n6483), .ZN(n6604) );
  NAND2_X1 U8229 ( .A1(n7989), .A2(n6604), .ZN(n7768) );
  AND2_X1 U8230 ( .A1(n7763), .A2(n7768), .ZN(n7924) );
  INV_X1 U8231 ( .A(n7924), .ZN(n6536) );
  INV_X1 U8232 ( .A(n6484), .ZN(n6485) );
  NAND2_X1 U8233 ( .A1(n6486), .A2(n6485), .ZN(n6489) );
  INV_X1 U8234 ( .A(n6500), .ZN(n6487) );
  NAND2_X1 U8235 ( .A1(n6490), .A2(n6487), .ZN(n6488) );
  INV_X1 U8236 ( .A(n6504), .ZN(n6597) );
  NAND2_X1 U8237 ( .A1(n6490), .A2(n6597), .ZN(n6519) );
  INV_X1 U8238 ( .A(n6518), .ZN(n6491) );
  INV_X1 U8239 ( .A(n7731), .ZN(n7717) );
  AOI22_X1 U8240 ( .A1(n6536), .A2(n7727), .B1(n7717), .B2(n6492), .ZN(n6509)
         );
  NAND2_X1 U8241 ( .A1(n6494), .A2(n6493), .ZN(n6499) );
  AND3_X1 U8242 ( .A1(n6497), .A2(n6496), .A3(n6495), .ZN(n6498) );
  OAI211_X1 U8243 ( .C1(n6502), .C2(n6500), .A(n6499), .B(n6498), .ZN(n6501)
         );
  NAND2_X1 U8244 ( .A1(n6501), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6507) );
  INV_X1 U8245 ( .A(n6502), .ZN(n6505) );
  NOR2_X1 U8246 ( .A1(n6504), .A2(n6503), .ZN(n7960) );
  NAND2_X1 U8247 ( .A1(n6505), .A2(n7960), .ZN(n6506) );
  INV_X1 U8248 ( .A(n7734), .ZN(n7719) );
  NAND2_X1 U8249 ( .A1(n7719), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6533) );
  NAND2_X1 U8250 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(n6533), .ZN(n6508) );
  OAI211_X1 U8251 ( .C1(n7737), .C2(n6604), .A(n6509), .B(n6508), .ZN(P2_U3172) );
  INV_X1 U8252 ( .A(n6958), .ZN(n6951) );
  INV_X1 U8253 ( .A(n6510), .ZN(n6512) );
  INV_X1 U8254 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6511) );
  OAI222_X1 U8255 ( .A1(n6951), .A2(P1_U3086), .B1(n9562), .B2(n6512), .C1(
        n6511), .C2(n9554), .ZN(P1_U3342) );
  INV_X1 U8256 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6513) );
  INV_X1 U8257 ( .A(n8019), .ZN(n8050) );
  OAI222_X1 U8258 ( .A1(n8456), .A2(n6513), .B1(n8467), .B2(n6512), .C1(
        P2_U3151), .C2(n8050), .ZN(P2_U3282) );
  NAND2_X1 U8259 ( .A1(n4326), .A2(n6594), .ZN(n6516) );
  NAND2_X1 U8260 ( .A1(n7571), .A2(n6604), .ZN(n6517) );
  XNOR2_X1 U8261 ( .A(n6526), .B(n10006), .ZN(n6525) );
  XOR2_X1 U8262 ( .A(n6524), .B(n6525), .Z(n6523) );
  INV_X1 U8263 ( .A(n7730), .ZN(n7708) );
  AOI22_X1 U8264 ( .A1(n7708), .A2(n7989), .B1(n6794), .B2(n7721), .ZN(n6520)
         );
  OAI21_X1 U8265 ( .B1(n6641), .B2(n7731), .A(n6520), .ZN(n6521) );
  AOI21_X1 U8266 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6533), .A(n6521), .ZN(
        n6522) );
  OAI21_X1 U8267 ( .B1(n7724), .B2(n6523), .A(n6522), .ZN(P2_U3162) );
  INV_X2 U8268 ( .A(n7571), .ZN(n7210) );
  XNOR2_X1 U8269 ( .A(n10018), .B(n7210), .ZN(n6632) );
  XNOR2_X1 U8270 ( .A(n6632), .B(n6641), .ZN(n6630) );
  NAND2_X1 U8271 ( .A1(n6525), .A2(n6524), .ZN(n6529) );
  INV_X1 U8272 ( .A(n6526), .ZN(n6527) );
  NAND2_X1 U8273 ( .A1(n6527), .A2(n10006), .ZN(n6528) );
  NAND2_X1 U8274 ( .A1(n6529), .A2(n6528), .ZN(n6631) );
  XOR2_X1 U8275 ( .A(n6630), .B(n6631), .Z(n6535) );
  AOI22_X1 U8276 ( .A1(n7708), .A2(n6492), .B1(n6530), .B2(n7721), .ZN(n6531)
         );
  OAI21_X1 U8277 ( .B1(n10008), .B2(n7731), .A(n6531), .ZN(n6532) );
  AOI21_X1 U8278 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6533), .A(n6532), .ZN(
        n6534) );
  OAI21_X1 U8279 ( .B1(n6535), .B2(n7724), .A(n6534), .ZN(P2_U3177) );
  INV_X1 U8280 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6540) );
  OAI21_X1 U8281 ( .B1(n10068), .B2(n9987), .A(n6536), .ZN(n6538) );
  NOR2_X1 U8282 ( .A1(n10006), .A2(n10007), .ZN(n6598) );
  INV_X1 U8283 ( .A(n6598), .ZN(n6537) );
  OAI211_X1 U8284 ( .C1(n6604), .C2(n10054), .A(n6538), .B(n6537), .ZN(n6549)
         );
  NAND2_X1 U8285 ( .A1(n6549), .A2(n10074), .ZN(n6539) );
  OAI21_X1 U8286 ( .B1(n6540), .B2(n10074), .A(n6539), .ZN(P2_U3390) );
  NAND2_X1 U8287 ( .A1(n4306), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6547) );
  INV_X1 U8288 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6541) );
  OR2_X1 U8289 ( .A1(n8615), .A2(n6541), .ZN(n6546) );
  OR2_X1 U8290 ( .A1(n6542), .A2(n9175), .ZN(n6545) );
  INV_X1 U8291 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6543) );
  OR2_X1 U8292 ( .A1(n4308), .A2(n6543), .ZN(n6544) );
  NAND4_X1 U8293 ( .A1(n6547), .A2(n6546), .A3(n6545), .A4(n6544), .ZN(n8724)
         );
  NAND2_X1 U8294 ( .A1(n8724), .A2(P1_U3973), .ZN(n6548) );
  OAI21_X1 U8295 ( .B1(n5568), .B2(P1_U3973), .A(n6548), .ZN(P1_U3583) );
  NAND2_X1 U8296 ( .A1(n6549), .A2(n10092), .ZN(n6550) );
  OAI21_X1 U8297 ( .B1(n10092), .B2(n9881), .A(n6550), .ZN(P2_U3459) );
  MUX2_X1 U8298 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9882), .Z(n6893) );
  XNOR2_X1 U8299 ( .A(n6893), .B(n6900), .ZN(n6894) );
  MUX2_X1 U8300 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9882), .Z(n6558) );
  INV_X1 U8301 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6551) );
  OR2_X1 U8302 ( .A1(n6449), .A2(n6551), .ZN(n6553) );
  NAND2_X1 U8303 ( .A1(n9882), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8304 ( .A1(n6553), .A2(n6552), .ZN(n6557) );
  AOI22_X1 U8305 ( .A1(n6556), .A2(n6555), .B1(n6554), .B2(n6561), .ZN(n9899)
         );
  XOR2_X1 U8306 ( .A(n9888), .B(n6557), .Z(n9900) );
  NAND2_X1 U8307 ( .A1(n9899), .A2(n9900), .ZN(n9898) );
  OAI21_X1 U8308 ( .B1(n6557), .B2(n9888), .A(n9898), .ZN(n9918) );
  XNOR2_X1 U8309 ( .A(n6558), .B(n6577), .ZN(n9919) );
  NOR2_X1 U8310 ( .A1(n9918), .A2(n9919), .ZN(n9916) );
  AOI21_X1 U8311 ( .B1(n6558), .B2(n6577), .A(n9916), .ZN(n9931) );
  MUX2_X1 U8312 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9882), .Z(n6559) );
  XNOR2_X1 U8313 ( .A(n6559), .B(n9928), .ZN(n9932) );
  INV_X1 U8314 ( .A(n6559), .ZN(n6560) );
  OAI22_X1 U8315 ( .A1(n9931), .A2(n9932), .B1(n6565), .B2(n6560), .ZN(n6895)
         );
  XOR2_X1 U8316 ( .A(n6894), .B(n6895), .Z(n6589) );
  INV_X1 U8317 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9998) );
  MUX2_X1 U8318 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n9998), .S(n6900), .Z(n6569)
         );
  NAND2_X1 U8319 ( .A1(n6561), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6562) );
  OR2_X1 U8320 ( .A1(n6567), .A2(n9925), .ZN(n6568) );
  NAND2_X1 U8321 ( .A1(n6568), .A2(n6569), .ZN(n6882) );
  OAI21_X1 U8322 ( .B1(n6569), .B2(n6568), .A(n6882), .ZN(n6583) );
  INV_X1 U8323 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10082) );
  MUX2_X1 U8324 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10082), .S(n6900), .Z(n6581)
         );
  OAI21_X1 U8325 ( .B1(n4295), .B2(n6571), .A(n6570), .ZN(n6573) );
  NAND2_X1 U8326 ( .A1(n6573), .A2(n9888), .ZN(n6574) );
  OAI21_X1 U8327 ( .B1(n6573), .B2(n9888), .A(n6574), .ZN(n9890) );
  NOR2_X1 U8328 ( .A1(n9890), .A2(n5097), .ZN(n9889) );
  INV_X1 U8329 ( .A(n6574), .ZN(n6575) );
  NAND2_X1 U8330 ( .A1(P2_REG1_REG_4__SCAN_IN), .A2(n6577), .ZN(n6576) );
  OAI21_X1 U8331 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6577), .A(n6576), .ZN(
        n9906) );
  INV_X1 U8332 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10080) );
  NAND2_X1 U8333 ( .A1(n6580), .A2(n6581), .ZN(n6902) );
  OAI21_X1 U8334 ( .B1(n6581), .B2(n6580), .A(n6902), .ZN(n6582) );
  AOI22_X1 U8335 ( .A1(n6584), .A2(n6583), .B1(n9951), .B2(n6582), .ZN(n6586)
         );
  AND2_X1 U8336 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6836) );
  INV_X1 U8337 ( .A(n6836), .ZN(n6585) );
  OAI211_X1 U8338 ( .C1(n9980), .C2(n6900), .A(n6586), .B(n6585), .ZN(n6587)
         );
  AOI21_X1 U8339 ( .B1(n9959), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n6587), .ZN(
        n6588) );
  OAI21_X1 U8340 ( .B1(n6589), .B2(n9917), .A(n6588), .ZN(P2_U3188) );
  NAND2_X1 U8341 ( .A1(n6593), .A2(n6590), .ZN(n6591) );
  OAI211_X1 U8342 ( .C1(n6594), .C2(n6593), .A(n6592), .B(n6591), .ZN(n6600)
         );
  INV_X1 U8343 ( .A(n6600), .ZN(n6596) );
  INV_X1 U8344 ( .A(n10003), .ZN(n6595) );
  NOR3_X1 U8345 ( .A1(n7924), .A2(n10073), .A3(n6597), .ZN(n6599) );
  NOR2_X1 U8346 ( .A1(n6599), .A2(n6598), .ZN(n6601) );
  NAND2_X2 U8347 ( .A1(n6600), .A2(n10002), .ZN(n10016) );
  MUX2_X1 U8348 ( .A(n9096), .B(n6601), .S(n10016), .Z(n6603) );
  NAND2_X1 U8349 ( .A1(n9994), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6602) );
  OAI211_X1 U8350 ( .C1(n8329), .C2(n6604), .A(n6603), .B(n6602), .ZN(P2_U3233) );
  NAND2_X1 U8351 ( .A1(n6733), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U8352 ( .B1(n6733), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6607), .ZN(
        n6608) );
  AOI211_X1 U8353 ( .C1(n6609), .C2(n6608), .A(n6732), .B(n8960), .ZN(n6618)
         );
  OAI21_X1 U8354 ( .B1(n6611), .B2(n6414), .A(n6610), .ZN(n6614) );
  MUX2_X1 U8355 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n6612), .S(n6733), .Z(n6613)
         );
  NAND2_X1 U8356 ( .A1(n6613), .A2(n6614), .ZN(n6736) );
  OAI211_X1 U8357 ( .C1(n6614), .C2(n6613), .A(n8975), .B(n6736), .ZN(n6616)
         );
  AND2_X1 U8358 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7446) );
  AOI21_X1 U8359 ( .B1(n9679), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n7446), .ZN(
        n6615) );
  OAI211_X1 U8360 ( .C1(n9689), .C2(n6737), .A(n6616), .B(n6615), .ZN(n6617)
         );
  OR2_X1 U8361 ( .A1(n6618), .A2(n6617), .ZN(P1_U3254) );
  INV_X1 U8362 ( .A(n7143), .ZN(n7146) );
  INV_X1 U8363 ( .A(n6619), .ZN(n6621) );
  OAI222_X1 U8364 ( .A1(n7146), .A2(P1_U3086), .B1(n9562), .B2(n6621), .C1(
        n6620), .C2(n9559), .ZN(P1_U3341) );
  OAI222_X1 U8365 ( .A1(n8456), .A2(n6622), .B1(n8467), .B2(n6621), .C1(
        P2_U3151), .C2(n9979), .ZN(P2_U3281) );
  AOI21_X1 U8366 ( .B1(n6624), .B2(n6623), .A(n4325), .ZN(n6629) );
  AOI22_X1 U8367 ( .A1(n9199), .A2(n6771), .B1(n8898), .B2(n8577), .ZN(n6870)
         );
  INV_X1 U8368 ( .A(n6870), .ZN(n6625) );
  AOI22_X1 U8369 ( .A1(n6625), .A2(n8599), .B1(n6874), .B2(n9670), .ZN(n6628)
         );
  INV_X1 U8370 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6626) );
  OR2_X1 U8371 ( .A1(n6675), .A2(n6626), .ZN(n6627) );
  OAI211_X1 U8372 ( .C1(n6629), .C2(n9665), .A(n6628), .B(n6627), .ZN(P1_U3222) );
  NAND2_X1 U8373 ( .A1(n6631), .A2(n6630), .ZN(n6635) );
  INV_X1 U8374 ( .A(n6632), .ZN(n6633) );
  NAND2_X1 U8375 ( .A1(n6633), .A2(n6641), .ZN(n6634) );
  NAND2_X1 U8376 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  XNOR2_X1 U8377 ( .A(n7210), .B(n6726), .ZN(n6707) );
  XNOR2_X1 U8378 ( .A(n6707), .B(n10008), .ZN(n6637) );
  AOI21_X1 U8379 ( .B1(n6636), .B2(n6637), .A(n7724), .ZN(n6640) );
  INV_X1 U8380 ( .A(n6636), .ZN(n6639) );
  INV_X1 U8381 ( .A(n6637), .ZN(n6638) );
  NAND2_X1 U8382 ( .A1(n6640), .A2(n6710), .ZN(n6644) );
  INV_X1 U8383 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6725) );
  NOR2_X1 U8384 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6725), .ZN(n9896) );
  OAI22_X1 U8385 ( .A1(n6641), .A2(n7730), .B1(n7731), .B2(n5123), .ZN(n6642)
         );
  AOI211_X1 U8386 ( .C1(n6726), .C2(n7721), .A(n9896), .B(n6642), .ZN(n6643)
         );
  OAI211_X1 U8387 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7719), .A(n6644), .B(
        n6643), .ZN(P2_U3158) );
  INV_X1 U8388 ( .A(n8873), .ZN(n6652) );
  NOR2_X1 U8389 ( .A1(n9677), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6645) );
  OR2_X1 U8390 ( .A1(n6645), .A2(n7611), .ZN(n9675) );
  INV_X1 U8391 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8392 ( .A1(n9675), .A2(n6646), .ZN(n6647) );
  NAND2_X1 U8393 ( .A1(P1_U3973), .A2(n6647), .ZN(n6651) );
  NOR3_X1 U8394 ( .A1(n6649), .A2(n6648), .A3(n7611), .ZN(n6650) );
  AOI211_X1 U8395 ( .C1(n6652), .C2(n8900), .A(n6651), .B(n6650), .ZN(n6700)
         );
  OAI211_X1 U8396 ( .C1(n6655), .C2(n6654), .A(n9695), .B(n6653), .ZN(n6665)
         );
  AOI22_X1 U8397 ( .A1(n9679), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6664) );
  NAND2_X1 U8398 ( .A1(n8906), .A2(n6656), .ZN(n6663) );
  MUX2_X1 U8399 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6307), .S(n6657), .Z(n6658)
         );
  NAND3_X1 U8400 ( .A1(n8902), .A2(n6659), .A3(n6658), .ZN(n6660) );
  NAND3_X1 U8401 ( .A1(n8975), .A2(n6661), .A3(n6660), .ZN(n6662) );
  NAND4_X1 U8402 ( .A1(n6665), .A2(n6664), .A3(n6663), .A4(n6662), .ZN(n6666)
         );
  OR2_X1 U8403 ( .A1(n6700), .A2(n6666), .ZN(P1_U3245) );
  NAND2_X1 U8404 ( .A1(n8122), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n6667) );
  OAI21_X1 U8405 ( .B1(n8218), .B2(n8122), .A(n6667), .ZN(P2_U3516) );
  NOR3_X1 U8406 ( .A1(n4325), .A2(n4564), .A3(n6669), .ZN(n6672) );
  INV_X1 U8407 ( .A(n6670), .ZN(n6671) );
  OAI21_X1 U8408 ( .B1(n6672), .B2(n6671), .A(n9649), .ZN(n6674) );
  INV_X1 U8409 ( .A(n8897), .ZN(n6799) );
  INV_X1 U8410 ( .A(n9199), .ZN(n6940) );
  OAI22_X1 U8411 ( .A1(n6799), .A2(n6939), .B1(n6773), .B2(n6940), .ZN(n9737)
         );
  AOI22_X1 U8412 ( .A1(n9737), .A2(n8599), .B1(n6767), .B2(n9670), .ZN(n6673)
         );
  OAI211_X1 U8413 ( .C1(n6675), .C2(n9740), .A(n6674), .B(n6673), .ZN(P1_U3237) );
  INV_X1 U8414 ( .A(n6676), .ZN(n6702) );
  INV_X1 U8415 ( .A(n8078), .ZN(n8069) );
  OAI222_X1 U8416 ( .A1(n8457), .A2(n6702), .B1(n8069), .B2(P2_U3151), .C1(
        n6677), .C2(n8456), .ZN(P2_U3280) );
  INV_X1 U8417 ( .A(n6678), .ZN(n6679) );
  AOI21_X1 U8418 ( .B1(n7763), .B2(n5486), .A(n6679), .ZN(n6797) );
  XNOR2_X1 U8419 ( .A(n5486), .B(n6680), .ZN(n6681) );
  INV_X1 U8420 ( .A(n8307), .ZN(n9982) );
  AOI222_X1 U8421 ( .A1(n9987), .A2(n6681), .B1(n7989), .B2(n9982), .C1(n5092), 
        .C2(n9984), .ZN(n6792) );
  OAI21_X1 U8422 ( .B1(n10061), .B2(n6797), .A(n6792), .ZN(n6687) );
  OAI22_X1 U8423 ( .A1(n8394), .A2(n5061), .B1(n10092), .B2(n6682), .ZN(n6683)
         );
  AOI21_X1 U8424 ( .B1(n6687), .B2(n10092), .A(n6683), .ZN(n6684) );
  INV_X1 U8425 ( .A(n6684), .ZN(P2_U3460) );
  INV_X1 U8426 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6685) );
  OAI22_X1 U8427 ( .A1(n5061), .A2(n8450), .B1(n10074), .B2(n6685), .ZN(n6686)
         );
  AOI21_X1 U8428 ( .B1(n6687), .B2(n10074), .A(n6686), .ZN(n6688) );
  INV_X1 U8429 ( .A(n6688), .ZN(P2_U3393) );
  NOR2_X1 U8430 ( .A1(n9689), .A2(n6689), .ZN(n6699) );
  AOI211_X1 U8431 ( .C1(n6692), .C2(n6691), .A(n6690), .B(n8960), .ZN(n6698)
         );
  INV_X1 U8432 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9572) );
  XOR2_X1 U8433 ( .A(n6694), .B(n6693), .Z(n6695) );
  NAND2_X1 U8434 ( .A1(n8975), .A2(n6695), .ZN(n6696) );
  NAND2_X1 U8435 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9659) );
  OAI211_X1 U8436 ( .C1(n9572), .C2(n9699), .A(n6696), .B(n9659), .ZN(n6697)
         );
  OR4_X1 U8437 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(P1_U3247)
         );
  INV_X1 U8438 ( .A(n8912), .ZN(n8919) );
  OAI222_X1 U8439 ( .A1(P1_U3086), .A2(n8919), .B1(n9562), .B2(n6702), .C1(
        n6701), .C2(n9559), .ZN(P1_U3340) );
  INV_X1 U8440 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6704) );
  INV_X1 U8441 ( .A(n6703), .ZN(n6705) );
  OAI222_X1 U8442 ( .A1(n8456), .A2(n6704), .B1(n8467), .B2(n6705), .C1(
        P2_U3151), .C2(n8090), .ZN(P2_U3279) );
  INV_X1 U8443 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6706) );
  INV_X1 U8444 ( .A(n8934), .ZN(n8941) );
  OAI222_X1 U8445 ( .A1(n9559), .A2(n6706), .B1(n9562), .B2(n6705), .C1(n8941), 
        .C2(P1_U3086), .ZN(P1_U3339) );
  XNOR2_X1 U8446 ( .A(n10030), .B(n7210), .ZN(n6816) );
  XNOR2_X1 U8447 ( .A(n6816), .B(n7987), .ZN(n6713) );
  INV_X1 U8448 ( .A(n6707), .ZN(n6708) );
  NAND2_X1 U8449 ( .A1(n6708), .A2(n7988), .ZN(n6709) );
  INV_X1 U8450 ( .A(n6819), .ZN(n6711) );
  AOI21_X1 U8451 ( .B1(n6713), .B2(n6712), .A(n6711), .ZN(n6718) );
  AND2_X1 U8452 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9913) );
  OAI22_X1 U8453 ( .A1(n6829), .A2(n7731), .B1(n7730), .B2(n10008), .ZN(n6714)
         );
  AOI211_X1 U8454 ( .C1(n4856), .C2(n7721), .A(n9913), .B(n6714), .ZN(n6717)
         );
  INV_X1 U8455 ( .A(n6715), .ZN(n6919) );
  NAND2_X1 U8456 ( .A1(n7734), .A2(n6919), .ZN(n6716) );
  OAI211_X1 U8457 ( .C1(n6718), .C2(n7724), .A(n6717), .B(n6716), .ZN(P2_U3170) );
  XOR2_X1 U8458 ( .A(n6719), .B(n7926), .Z(n6720) );
  AOI222_X1 U8459 ( .A1(n9987), .A2(n6720), .B1(n7987), .B2(n9984), .C1(n5092), 
        .C2(n9982), .ZN(n10023) );
  XNOR2_X1 U8460 ( .A(n6721), .B(n7926), .ZN(n10026) );
  INV_X1 U8461 ( .A(n10010), .ZN(n7182) );
  AND2_X1 U8462 ( .A1(n5539), .A2(n6722), .ZN(n10015) );
  INV_X1 U8463 ( .A(n10015), .ZN(n6723) );
  NAND2_X1 U8464 ( .A1(n7182), .A2(n6723), .ZN(n6724) );
  AOI22_X1 U8465 ( .A1(n9993), .A2(n6726), .B1(n6725), .B2(n9994), .ZN(n6727)
         );
  OAI21_X1 U8466 ( .B1(n6551), .B2(n10016), .A(n6727), .ZN(n6728) );
  AOI21_X1 U8467 ( .B1(n10026), .B2(n9996), .A(n6728), .ZN(n6729) );
  OAI21_X1 U8468 ( .B1(n10023), .B2(n8334), .A(n6729), .ZN(P2_U3230) );
  NAND2_X1 U8469 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n6958), .ZN(n6730) );
  OAI21_X1 U8470 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6958), .A(n6730), .ZN(
        n6735) );
  NOR2_X1 U8471 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6738), .ZN(n6731) );
  AOI21_X1 U8472 ( .B1(n6738), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6731), .ZN(
        n9685) );
  OAI21_X1 U8473 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n6738), .A(n9683), .ZN(
        n6734) );
  NOR2_X1 U8474 ( .A1(n6735), .A2(n6734), .ZN(n6957) );
  AOI211_X1 U8475 ( .C1(n6735), .C2(n6734), .A(n6957), .B(n8960), .ZN(n6747)
         );
  OAI21_X1 U8476 ( .B1(n6612), .B2(n6737), .A(n6736), .ZN(n9688) );
  AOI22_X1 U8477 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(n9690), .B1(n6738), .B2(
        n5883), .ZN(n9687) );
  NOR2_X1 U8478 ( .A1(n9688), .A2(n9687), .ZN(n9686) );
  NOR2_X1 U8479 ( .A1(n6738), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U8480 ( .A1(n9686), .A2(n6739), .ZN(n6743) );
  OR2_X1 U8481 ( .A1(n6958), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6741) );
  NAND2_X1 U8482 ( .A1(n6958), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6740) );
  AND2_X1 U8483 ( .A1(n6741), .A2(n6740), .ZN(n6742) );
  NAND2_X1 U8484 ( .A1(n6742), .A2(n6743), .ZN(n6950) );
  OAI211_X1 U8485 ( .C1(n6743), .C2(n6742), .A(n6950), .B(n8975), .ZN(n6745)
         );
  AND2_X1 U8486 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7518) );
  AOI21_X1 U8487 ( .B1(n9679), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n7518), .ZN(
        n6744) );
  OAI211_X1 U8488 ( .C1(n9689), .C2(n6951), .A(n6745), .B(n6744), .ZN(n6746)
         );
  OR2_X1 U8489 ( .A1(n6747), .A2(n6746), .ZN(P1_U3256) );
  INV_X1 U8490 ( .A(n8957), .ZN(n8949) );
  INV_X1 U8491 ( .A(n6748), .ZN(n6750) );
  OAI222_X1 U8492 ( .A1(n8949), .A2(P1_U3086), .B1(n9562), .B2(n6750), .C1(
        n6749), .C2(n9559), .ZN(P1_U3338) );
  INV_X1 U8493 ( .A(n8130), .ZN(n8116) );
  OAI222_X1 U8494 ( .A1(n8456), .A2(n6751), .B1(n8467), .B2(n6750), .C1(
        P2_U3151), .C2(n8116), .ZN(P2_U3278) );
  OR2_X1 U8495 ( .A1(n6772), .A2(n6867), .ZN(n6865) );
  NAND2_X1 U8496 ( .A1(n6865), .A2(n6753), .ZN(n9736) );
  INV_X2 U8497 ( .A(n6767), .ZN(n9775) );
  NAND2_X1 U8498 ( .A1(n8898), .A2(n9775), .ZN(n8791) );
  INV_X1 U8499 ( .A(n6754), .ZN(n6756) );
  NAND2_X1 U8500 ( .A1(n6799), .A2(n8497), .ZN(n6802) );
  NAND2_X1 U8501 ( .A1(n8897), .A2(n9783), .ZN(n8788) );
  INV_X1 U8502 ( .A(n8746), .ZN(n6755) );
  OR2_X2 U8503 ( .A1(n6754), .A2(n8746), .ZN(n6803) );
  OAI21_X1 U8504 ( .B1(n6756), .B2(n6755), .A(n6803), .ZN(n6759) );
  NAND2_X1 U8505 ( .A1(n8896), .A2(n8577), .ZN(n6758) );
  NAND2_X1 U8506 ( .A1(n8898), .A2(n9199), .ZN(n6757) );
  NAND2_X1 U8507 ( .A1(n6758), .A2(n6757), .ZN(n8496) );
  AOI21_X1 U8508 ( .B1(n6759), .B2(n9738), .A(n8496), .ZN(n9782) );
  INV_X1 U8509 ( .A(n6760), .ZN(n6763) );
  INV_X1 U8510 ( .A(n6761), .ZN(n9490) );
  NAND3_X1 U8511 ( .A1(n6763), .A2(n9490), .A3(n6762), .ZN(n6764) );
  OAI22_X1 U8512 ( .A1(n9394), .A2(n6766), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9741), .ZN(n6769) );
  OR2_X1 U8513 ( .A1(n6874), .A2(n6770), .ZN(n9748) );
  NOR2_X1 U8514 ( .A1(n9748), .A2(n6767), .ZN(n9749) );
  NAND2_X1 U8515 ( .A1(n6784), .A2(n7017), .ZN(n9403) );
  OAI211_X1 U8516 ( .C1(n9749), .C2(n9783), .A(n9750), .B(n6809), .ZN(n9781)
         );
  NOR2_X1 U8517 ( .A1(n9781), .A2(n9413), .ZN(n6768) );
  AOI211_X1 U8518 ( .C1(n9410), .C2(n8497), .A(n6769), .B(n6768), .ZN(n6783)
         );
  NAND2_X1 U8519 ( .A1(n6771), .A2(n6770), .ZN(n6868) );
  NAND2_X1 U8520 ( .A1(n6772), .A2(n6868), .ZN(n6775) );
  NAND2_X1 U8521 ( .A1(n6773), .A2(n9769), .ZN(n6774) );
  NAND2_X1 U8522 ( .A1(n6775), .A2(n6774), .ZN(n9746) );
  INV_X1 U8523 ( .A(n6776), .ZN(n6777) );
  NAND2_X1 U8524 ( .A1(n9747), .A2(n9746), .ZN(n6780) );
  INV_X1 U8525 ( .A(n8898), .ZN(n6778) );
  NAND2_X1 U8526 ( .A1(n6778), .A2(n9775), .ZN(n6779) );
  NAND2_X1 U8527 ( .A1(n6780), .A2(n6779), .ZN(n6798) );
  XNOR2_X1 U8528 ( .A(n6798), .B(n8746), .ZN(n9785) );
  AND2_X1 U8529 ( .A1(n7004), .A2(n6872), .ZN(n6781) );
  NAND2_X1 U8530 ( .A1(n9785), .A2(n9755), .ZN(n6782) );
  OAI211_X1 U8531 ( .C1(n9782), .C2(n9758), .A(n6783), .B(n6782), .ZN(P1_U3290) );
  AOI21_X1 U8532 ( .B1(n9754), .B2(n6784), .A(n9410), .ZN(n6791) );
  NAND3_X1 U8533 ( .A1(n8747), .A2(n6785), .A3(n8872), .ZN(n6787) );
  OAI211_X1 U8534 ( .C1(n5661), .C2(n9741), .A(n6787), .B(n6786), .ZN(n6789)
         );
  NOR2_X1 U8535 ( .A1(n9394), .A2(n5660), .ZN(n6788) );
  AOI21_X1 U8536 ( .B1(n6789), .B2(n9394), .A(n6788), .ZN(n6790) );
  OAI21_X1 U8537 ( .B1(n6791), .B2(n6873), .A(n6790), .ZN(P1_U3293) );
  INV_X1 U8538 ( .A(n9996), .ZN(n7543) );
  MUX2_X1 U8539 ( .A(n6793), .B(n6792), .S(n10016), .Z(n6796) );
  AOI22_X1 U8540 ( .A1(n9993), .A2(n6794), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9994), .ZN(n6795) );
  OAI211_X1 U8541 ( .C1(n6797), .C2(n7543), .A(n6796), .B(n6795), .ZN(P2_U3232) );
  NAND2_X1 U8542 ( .A1(n6799), .A2(n9783), .ZN(n6800) );
  NAND2_X1 U8543 ( .A1(n8896), .A2(n9789), .ZN(n8790) );
  NAND2_X1 U8544 ( .A1(n4351), .A2(n8790), .ZN(n8745) );
  XNOR2_X1 U8545 ( .A(n4303), .B(n8745), .ZN(n9792) );
  INV_X1 U8546 ( .A(n9792), .ZN(n6815) );
  XNOR2_X1 U8547 ( .A(n6847), .B(n8745), .ZN(n6804) );
  NOR2_X1 U8548 ( .A1(n6804), .A2(n9706), .ZN(n9790) );
  NAND2_X1 U8549 ( .A1(n8897), .A2(n9199), .ZN(n6806) );
  NAND2_X1 U8550 ( .A1(n8895), .A2(n8988), .ZN(n6805) );
  AND2_X1 U8551 ( .A1(n6806), .A2(n6805), .ZN(n9787) );
  INV_X1 U8552 ( .A(n9787), .ZN(n6807) );
  OAI21_X1 U8553 ( .B1(n9790), .B2(n6807), .A(n9394), .ZN(n6814) );
  OAI22_X1 U8554 ( .A1(n9394), .A2(n6808), .B1(n9673), .B2(n9741), .ZN(n6812)
         );
  AOI21_X1 U8555 ( .B1(n6809), .B2(n9671), .A(n9403), .ZN(n6810) );
  NAND2_X1 U8556 ( .A1(n6810), .A2(n6857), .ZN(n9788) );
  NOR2_X1 U8557 ( .A1(n9788), .A2(n9413), .ZN(n6811) );
  AOI211_X1 U8558 ( .C1(n9410), .C2(n9671), .A(n6812), .B(n6811), .ZN(n6813)
         );
  OAI211_X1 U8559 ( .C1(n6815), .C2(n9415), .A(n6814), .B(n6813), .ZN(P1_U3289) );
  INV_X1 U8560 ( .A(n6816), .ZN(n6817) );
  NAND2_X1 U8561 ( .A1(n6817), .A2(n5123), .ZN(n6818) );
  NAND2_X1 U8562 ( .A1(n6819), .A2(n6818), .ZN(n6831) );
  XNOR2_X1 U8563 ( .A(n7583), .B(n6822), .ZN(n6828) );
  XNOR2_X1 U8564 ( .A(n6828), .B(n9983), .ZN(n6830) );
  XNOR2_X1 U8565 ( .A(n6831), .B(n6830), .ZN(n6820) );
  NAND2_X1 U8566 ( .A1(n6820), .A2(n7727), .ZN(n6824) );
  NOR2_X1 U8567 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9081), .ZN(n9930) );
  OAI22_X1 U8568 ( .A1(n5123), .A2(n7730), .B1(n7731), .B2(n7119), .ZN(n6821)
         );
  AOI211_X1 U8569 ( .C1(n6822), .C2(n7721), .A(n9930), .B(n6821), .ZN(n6823)
         );
  OAI211_X1 U8570 ( .C1(n6982), .C2(n7719), .A(n6824), .B(n6823), .ZN(P2_U3167) );
  INV_X1 U8571 ( .A(n6825), .ZN(n6932) );
  AOI22_X1 U8572 ( .A1(n8971), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n6826), .ZN(n6827) );
  OAI21_X1 U8573 ( .B1(n6932), .B2(n9551), .A(n6827), .ZN(P1_U3337) );
  XNOR2_X1 U8574 ( .A(n7583), .B(n10039), .ZN(n6965) );
  XNOR2_X1 U8575 ( .A(n6965), .B(n7986), .ZN(n6832) );
  OAI211_X1 U8576 ( .C1(n6833), .C2(n6832), .A(n6968), .B(n7727), .ZN(n6838)
         );
  OAI22_X1 U8577 ( .A1(n7737), .A2(n6834), .B1(n7731), .B2(n7129), .ZN(n6835)
         );
  AOI211_X1 U8578 ( .C1(n7708), .C2(n9983), .A(n6836), .B(n6835), .ZN(n6837)
         );
  OAI211_X1 U8579 ( .C1(n9992), .C2(n7719), .A(n6838), .B(n6837), .ZN(P2_U3179) );
  INV_X1 U8580 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6846) );
  INV_X1 U8581 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6843) );
  AOI22_X1 U8582 ( .A1(n6840), .A2(P2_REG1_REG_31__SCAN_IN), .B1(n6839), .B2(
        P2_REG2_REG_31__SCAN_IN), .ZN(n6841) );
  OAI211_X1 U8583 ( .C1(n6844), .C2(n6843), .A(n6842), .B(n6841), .ZN(n7760)
         );
  NAND2_X1 U8584 ( .A1(n7760), .A2(P2_U3893), .ZN(n6845) );
  OAI21_X1 U8585 ( .B1(P2_U3893), .B2(n6846), .A(n6845), .ZN(P2_U3522) );
  INV_X1 U8586 ( .A(n8895), .ZN(n6992) );
  NAND2_X1 U8587 ( .A1(n6992), .A2(n6859), .ZN(n6998) );
  INV_X1 U8588 ( .A(n6859), .ZN(n9794) );
  NAND2_X1 U8589 ( .A1(n8895), .A2(n9794), .ZN(n8792) );
  NAND2_X1 U8590 ( .A1(n6998), .A2(n8792), .ZN(n6990) );
  INV_X1 U8591 ( .A(n6990), .ZN(n8749) );
  XNOR2_X1 U8592 ( .A(n6999), .B(n8749), .ZN(n6851) );
  NAND2_X1 U8593 ( .A1(n8896), .A2(n9199), .ZN(n6849) );
  NAND2_X1 U8594 ( .A1(n8894), .A2(n8577), .ZN(n6848) );
  NAND2_X1 U8595 ( .A1(n6849), .A2(n6848), .ZN(n6926) );
  INV_X1 U8596 ( .A(n6926), .ZN(n6850) );
  OAI21_X1 U8597 ( .B1(n6851), .B2(n9706), .A(n6850), .ZN(n9795) );
  INV_X1 U8598 ( .A(n9795), .ZN(n6864) );
  NAND2_X1 U8599 ( .A1(n6852), .A2(n8745), .ZN(n6855) );
  INV_X1 U8600 ( .A(n8896), .ZN(n6853) );
  NAND2_X1 U8601 ( .A1(n6853), .A2(n9789), .ZN(n6854) );
  XNOR2_X1 U8602 ( .A(n4302), .B(n6990), .ZN(n9797) );
  NAND2_X1 U8603 ( .A1(n6857), .A2(n6859), .ZN(n6856) );
  NAND2_X1 U8604 ( .A1(n6856), .A2(n9750), .ZN(n6858) );
  OR2_X1 U8605 ( .A1(n6858), .A2(n9732), .ZN(n9793) );
  INV_X1 U8606 ( .A(n9741), .ZN(n9335) );
  AOI22_X1 U8607 ( .A1(n9758), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n6929), .B2(
        n9335), .ZN(n6861) );
  NAND2_X1 U8608 ( .A1(n9410), .A2(n6859), .ZN(n6860) );
  OAI211_X1 U8609 ( .C1(n9793), .C2(n9413), .A(n6861), .B(n6860), .ZN(n6862)
         );
  AOI21_X1 U8610 ( .B1(n9797), .B2(n9755), .A(n6862), .ZN(n6863) );
  OAI21_X1 U8611 ( .B1(n6864), .B2(n9758), .A(n6863), .ZN(P1_U3288) );
  INV_X1 U8612 ( .A(n6865), .ZN(n6866) );
  AOI21_X1 U8613 ( .B1(n6772), .B2(n6867), .A(n6866), .ZN(n6871) );
  XNOR2_X1 U8614 ( .A(n6772), .B(n6868), .ZN(n9772) );
  INV_X1 U8615 ( .A(n7004), .ZN(n9709) );
  NAND2_X1 U8616 ( .A1(n9772), .A2(n9709), .ZN(n6869) );
  OAI211_X1 U8617 ( .C1(n6871), .C2(n9706), .A(n6870), .B(n6869), .ZN(n9770)
         );
  INV_X1 U8618 ( .A(n9770), .ZN(n6879) );
  NOR2_X1 U8619 ( .A1(n9758), .A2(n6872), .ZN(n9719) );
  OAI211_X1 U8620 ( .C1(n9769), .C2(n6873), .A(n9750), .B(n9748), .ZN(n9768)
         );
  NAND2_X1 U8621 ( .A1(n9410), .A2(n6874), .ZN(n6876) );
  AOI22_X1 U8622 ( .A1(n9758), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9335), .ZN(n6875) );
  OAI211_X1 U8623 ( .C1(n9768), .C2(n9413), .A(n6876), .B(n6875), .ZN(n6877)
         );
  AOI21_X1 U8624 ( .B1(n9772), .B2(n9719), .A(n6877), .ZN(n6878) );
  OAI21_X1 U8625 ( .B1(n6879), .B2(n9758), .A(n6878), .ZN(P1_U3292) );
  INV_X1 U8626 ( .A(n7585), .ZN(n6880) );
  NAND2_X1 U8627 ( .A1(n6880), .A2(P2_U3893), .ZN(n6881) );
  OAI21_X1 U8628 ( .B1(P2_U3893), .B2(n8721), .A(n6881), .ZN(P2_U3520) );
  INV_X1 U8629 ( .A(n9942), .ZN(n6883) );
  NAND2_X1 U8630 ( .A1(n6884), .A2(n6883), .ZN(n6885) );
  AOI22_X1 U8631 ( .A1(n7079), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7070), .B2(
        n6909), .ZN(n6887) );
  AOI21_X1 U8632 ( .B1(n6888), .B2(n6887), .A(n7072), .ZN(n6912) );
  MUX2_X1 U8633 ( .A(P2_REG1_REG_8__SCAN_IN), .B(P2_REG2_REG_8__SCAN_IN), .S(
        n8145), .Z(n6889) );
  NOR2_X1 U8634 ( .A1(n6909), .A2(n6889), .ZN(n7098) );
  AOI21_X1 U8635 ( .B1(n6909), .B2(n6889), .A(n7098), .ZN(n6898) );
  OR2_X1 U8636 ( .A1(n9882), .A2(n6890), .ZN(n6892) );
  NAND2_X1 U8637 ( .A1(n9882), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8638 ( .A1(n6892), .A2(n6891), .ZN(n6896) );
  OAI22_X1 U8639 ( .A1(n6895), .A2(n6894), .B1(n6893), .B2(n6900), .ZN(n9946)
         );
  XOR2_X1 U8640 ( .A(n9942), .B(n6896), .Z(n9947) );
  NAND2_X1 U8641 ( .A1(n9946), .A2(n9947), .ZN(n9945) );
  OAI21_X1 U8642 ( .B1(n6896), .B2(n9942), .A(n9945), .ZN(n6897) );
  AND2_X1 U8643 ( .A1(n6898), .A2(n6897), .ZN(n7097) );
  NOR2_X1 U8644 ( .A1(n6898), .A2(n6897), .ZN(n6899) );
  OAI21_X1 U8645 ( .B1(n7097), .B2(n6899), .A(n9970), .ZN(n6908) );
  NAND2_X1 U8646 ( .A1(n6900), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8647 ( .A1(n6902), .A2(n6901), .ZN(n6903) );
  XNOR2_X1 U8648 ( .A(n6903), .B(n9942), .ZN(n9949) );
  NOR2_X1 U8649 ( .A1(n9949), .A2(n5157), .ZN(n9953) );
  INV_X1 U8650 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7078) );
  MUX2_X1 U8651 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n7078), .S(n7079), .Z(n6904)
         );
  AOI21_X1 U8652 ( .B1(n6905), .B2(n6904), .A(n7080), .ZN(n6906) );
  OR2_X1 U8653 ( .A1(n6906), .A2(n9974), .ZN(n6907) );
  OAI211_X1 U8654 ( .C1(n9980), .C2(n6909), .A(n6908), .B(n6907), .ZN(n6910)
         );
  AND2_X1 U8655 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7133) );
  AOI211_X1 U8656 ( .C1(n9959), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6910), .B(
        n7133), .ZN(n6911) );
  OAI21_X1 U8657 ( .B1(n6912), .B2(n9965), .A(n6911), .ZN(P2_U3190) );
  NAND2_X1 U8658 ( .A1(n7784), .A2(n7792), .ZN(n7779) );
  XNOR2_X1 U8659 ( .A(n6913), .B(n7779), .ZN(n10028) );
  INV_X1 U8660 ( .A(n7779), .ZN(n7925) );
  XNOR2_X1 U8661 ( .A(n6914), .B(n7925), .ZN(n6915) );
  NAND2_X1 U8662 ( .A1(n6915), .A2(n9987), .ZN(n6917) );
  AOI22_X1 U8663 ( .A1(n9984), .A2(n9983), .B1(n7988), .B2(n9982), .ZN(n6916)
         );
  AND2_X1 U8664 ( .A1(n6917), .A2(n6916), .ZN(n10029) );
  INV_X1 U8665 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6918) );
  MUX2_X1 U8666 ( .A(n10029), .B(n6918), .S(n8334), .Z(n6921) );
  AOI22_X1 U8667 ( .A1(n9993), .A2(n4856), .B1(n9994), .B2(n6919), .ZN(n6920)
         );
  OAI211_X1 U8668 ( .C1(n7543), .C2(n10028), .A(n6921), .B(n6920), .ZN(
        P2_U3229) );
  NAND2_X1 U8669 ( .A1(n6922), .A2(n6923), .ZN(n6924) );
  XOR2_X1 U8670 ( .A(n6925), .B(n6924), .Z(n6931) );
  AOI22_X1 U8671 ( .A1(n6926), .A2(n8599), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        P1_U3086), .ZN(n6927) );
  OAI21_X1 U8672 ( .B1(n9794), .B2(n8594), .A(n6927), .ZN(n6928) );
  AOI21_X1 U8673 ( .B1(n6929), .B2(n8591), .A(n6928), .ZN(n6930) );
  OAI21_X1 U8674 ( .B1(n6931), .B2(n9665), .A(n6930), .ZN(P1_U3227) );
  OAI222_X1 U8675 ( .A1(n8456), .A2(n6933), .B1(n8150), .B2(P2_U3151), .C1(
        n8457), .C2(n6932), .ZN(P2_U3277) );
  INV_X1 U8676 ( .A(n6935), .ZN(n6937) );
  NOR2_X1 U8677 ( .A1(n6937), .A2(n6936), .ZN(n6938) );
  XNOR2_X1 U8678 ( .A(n6934), .B(n6938), .ZN(n6945) );
  INV_X1 U8679 ( .A(n9725), .ZN(n6943) );
  INV_X1 U8680 ( .A(n8893), .ZN(n7027) );
  OAI22_X1 U8681 ( .A1(n6992), .A2(n6940), .B1(n7027), .B2(n6939), .ZN(n9723)
         );
  AOI22_X1 U8682 ( .A1(n9723), .A2(n8599), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n6941) );
  OAI21_X1 U8683 ( .B1(n9799), .B2(n8594), .A(n6941), .ZN(n6942) );
  AOI21_X1 U8684 ( .B1(n6943), .B2(n8591), .A(n6942), .ZN(n6944) );
  OAI21_X1 U8685 ( .B1(n6945), .B2(n9665), .A(n6944), .ZN(P1_U3239) );
  INV_X1 U8686 ( .A(n6946), .ZN(n6948) );
  OAI222_X1 U8687 ( .A1(n8866), .A2(P1_U3086), .B1(n9562), .B2(n6948), .C1(
        n6947), .C2(n9559), .ZN(P1_U3336) );
  OAI222_X1 U8688 ( .A1(n8456), .A2(n6949), .B1(n8467), .B2(n6948), .C1(n8154), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U8689 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n6956) );
  OAI21_X1 U8690 ( .B1(n6951), .B2(n5907), .A(n6950), .ZN(n6954) );
  MUX2_X1 U8691 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n6952), .S(n7143), .Z(n6953)
         );
  NAND2_X1 U8692 ( .A1(n6953), .A2(n6954), .ZN(n7145) );
  OAI211_X1 U8693 ( .C1(n6954), .C2(n6953), .A(n8975), .B(n7145), .ZN(n6955)
         );
  NAND2_X1 U8694 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8472) );
  OAI211_X1 U8695 ( .C1(n9699), .C2(n6956), .A(n6955), .B(n8472), .ZN(n6963)
         );
  NAND2_X1 U8696 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n7143), .ZN(n6959) );
  OAI21_X1 U8697 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7143), .A(n6959), .ZN(
        n6960) );
  AOI211_X1 U8698 ( .C1(n6961), .C2(n6960), .A(n7142), .B(n8960), .ZN(n6962)
         );
  AOI211_X1 U8699 ( .C1(n8906), .C2(n7143), .A(n6963), .B(n6962), .ZN(n6964)
         );
  INV_X1 U8700 ( .A(n6964), .ZN(P1_U3257) );
  XNOR2_X1 U8701 ( .A(n7583), .B(n7125), .ZN(n7130) );
  XNOR2_X1 U8702 ( .A(n7130), .B(n7129), .ZN(n6972) );
  INV_X1 U8703 ( .A(n6965), .ZN(n6966) );
  NAND2_X1 U8704 ( .A1(n6966), .A2(n7986), .ZN(n6967) );
  INV_X1 U8705 ( .A(n6972), .ZN(n6970) );
  INV_X1 U8706 ( .A(n7132), .ZN(n6971) );
  AOI21_X1 U8707 ( .B1(n6972), .B2(n6969), .A(n6971), .ZN(n6979) );
  INV_X1 U8708 ( .A(n7123), .ZN(n6977) );
  NOR2_X1 U8709 ( .A1(n7737), .A2(n10043), .ZN(n6976) );
  NAND2_X1 U8710 ( .A1(n7717), .A2(n7985), .ZN(n6974) );
  OR2_X1 U8711 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6973), .ZN(n9956) );
  OAI211_X1 U8712 ( .C1(n7119), .C2(n7730), .A(n6974), .B(n9956), .ZN(n6975)
         );
  AOI211_X1 U8713 ( .C1(n6977), .C2(n7734), .A(n6976), .B(n6975), .ZN(n6978)
         );
  OAI21_X1 U8714 ( .B1(n6979), .B2(n7724), .A(n6978), .ZN(P2_U3153) );
  INV_X1 U8715 ( .A(n9988), .ZN(n6980) );
  OR2_X1 U8716 ( .A1(n6980), .A2(n7783), .ZN(n7930) );
  XOR2_X1 U8717 ( .A(n6981), .B(n7930), .Z(n10037) );
  OAI22_X1 U8718 ( .A1(n8329), .A2(n10034), .B1(n6982), .B2(n10002), .ZN(n6988) );
  XNOR2_X1 U8719 ( .A(n6983), .B(n7930), .ZN(n6984) );
  NAND2_X1 U8720 ( .A1(n6984), .A2(n9987), .ZN(n6986) );
  AOI22_X1 U8721 ( .A1(n9982), .A2(n7987), .B1(n7986), .B2(n9984), .ZN(n6985)
         );
  NAND2_X1 U8722 ( .A1(n6986), .A2(n6985), .ZN(n10035) );
  MUX2_X1 U8723 ( .A(n10035), .B(P2_REG2_REG_5__SCAN_IN), .S(n8334), .Z(n6987)
         );
  AOI211_X1 U8724 ( .C1(n9996), .C2(n10037), .A(n6988), .B(n6987), .ZN(n6989)
         );
  INV_X1 U8725 ( .A(n6989), .ZN(P2_U3228) );
  NAND2_X1 U8726 ( .A1(n6991), .A2(n6990), .ZN(n6994) );
  NAND2_X1 U8727 ( .A1(n6992), .A2(n9794), .ZN(n6993) );
  NAND2_X1 U8728 ( .A1(n6994), .A2(n6993), .ZN(n9729) );
  INV_X1 U8729 ( .A(n8894), .ZN(n6996) );
  NAND2_X1 U8730 ( .A1(n6996), .A2(n6995), .ZN(n8623) );
  NAND2_X1 U8731 ( .A1(n8894), .A2(n9799), .ZN(n8622) );
  NAND2_X1 U8732 ( .A1(n8623), .A2(n8622), .ZN(n9730) );
  NAND2_X1 U8733 ( .A1(n6996), .A2(n9799), .ZN(n6997) );
  NAND2_X1 U8734 ( .A1(n7027), .A2(n9656), .ZN(n9701) );
  NAND2_X1 U8735 ( .A1(n8893), .A2(n9808), .ZN(n7055) );
  INV_X1 U8736 ( .A(n7025), .ZN(n8627) );
  XNOR2_X1 U8737 ( .A(n7026), .B(n8627), .ZN(n9804) );
  INV_X1 U8738 ( .A(n9719), .ZN(n7011) );
  NAND2_X1 U8739 ( .A1(n7053), .A2(n8622), .ZN(n8625) );
  XNOR2_X1 U8740 ( .A(n8625), .B(n7025), .ZN(n7000) );
  NAND2_X1 U8741 ( .A1(n7000), .A2(n9738), .ZN(n7003) );
  NAND2_X1 U8742 ( .A1(n8892), .A2(n8988), .ZN(n7002) );
  NAND2_X1 U8743 ( .A1(n8894), .A2(n9199), .ZN(n7001) );
  AND2_X1 U8744 ( .A1(n7002), .A2(n7001), .ZN(n9648) );
  OAI211_X1 U8745 ( .C1(n9804), .C2(n7004), .A(n7003), .B(n9648), .ZN(n9810)
         );
  NAND2_X1 U8746 ( .A1(n9810), .A2(n9394), .ZN(n7010) );
  OAI22_X1 U8747 ( .A1(n9394), .A2(n7005), .B1(n9658), .B2(n9741), .ZN(n7008)
         );
  AOI21_X1 U8748 ( .B1(n9731), .B2(n9656), .A(n9403), .ZN(n7006) );
  NAND2_X1 U8749 ( .A1(n7006), .A2(n9714), .ZN(n9806) );
  NOR2_X1 U8750 ( .A1(n9806), .A2(n9413), .ZN(n7007) );
  AOI211_X1 U8751 ( .C1(n9410), .C2(n9656), .A(n7008), .B(n7007), .ZN(n7009)
         );
  OAI211_X1 U8752 ( .C1(n9804), .C2(n7011), .A(n7010), .B(n7009), .ZN(P1_U3286) );
  INV_X1 U8753 ( .A(n7012), .ZN(n7016) );
  OAI222_X1 U8754 ( .A1(n8457), .A2(n7016), .B1(P2_U3151), .B2(n7014), .C1(
        n7013), .C2(n8456), .ZN(P2_U3275) );
  OAI222_X1 U8755 ( .A1(P1_U3086), .A2(n7017), .B1(n9562), .B2(n7016), .C1(
        n7015), .C2(n9559), .ZN(P1_U3335) );
  INV_X1 U8756 ( .A(n7018), .ZN(n7041) );
  OAI222_X1 U8757 ( .A1(n8457), .A2(n7041), .B1(P2_U3151), .B2(n7762), .C1(
        n7019), .C2(n8456), .ZN(P2_U3274) );
  OR2_X1 U8758 ( .A1(n8625), .A2(n7025), .ZN(n9702) );
  INV_X1 U8759 ( .A(n8892), .ZN(n7028) );
  NAND2_X1 U8760 ( .A1(n7028), .A2(n7031), .ZN(n8632) );
  NAND2_X1 U8761 ( .A1(n9701), .A2(n8632), .ZN(n7054) );
  INV_X1 U8762 ( .A(n7054), .ZN(n8629) );
  NAND2_X1 U8763 ( .A1(n9702), .A2(n8629), .ZN(n7020) );
  NAND2_X1 U8764 ( .A1(n9813), .A2(n8892), .ZN(n7056) );
  NAND2_X1 U8765 ( .A1(n7020), .A2(n7056), .ZN(n7022) );
  INV_X1 U8766 ( .A(n8891), .ZN(n7021) );
  OR2_X1 U8767 ( .A1(n7021), .A2(n7339), .ZN(n8648) );
  NAND2_X1 U8768 ( .A1(n7339), .A2(n7021), .ZN(n8638) );
  NAND2_X1 U8769 ( .A1(n8648), .A2(n8638), .ZN(n8753) );
  XNOR2_X1 U8770 ( .A(n7022), .B(n8753), .ZN(n7023) );
  NAND2_X1 U8771 ( .A1(n7023), .A2(n9738), .ZN(n7024) );
  NAND2_X1 U8772 ( .A1(n8892), .A2(n9199), .ZN(n7332) );
  NAND2_X1 U8773 ( .A1(n7024), .A2(n7332), .ZN(n9824) );
  INV_X1 U8774 ( .A(n9824), .ZN(n7039) );
  NAND2_X1 U8775 ( .A1(n8632), .A2(n7056), .ZN(n9703) );
  NAND2_X1 U8776 ( .A1(n9700), .A2(n9703), .ZN(n7030) );
  NAND2_X1 U8777 ( .A1(n7028), .A2(n9813), .ZN(n7029) );
  NAND2_X1 U8778 ( .A1(n7030), .A2(n7029), .ZN(n7066) );
  XNOR2_X1 U8779 ( .A(n7066), .B(n8753), .ZN(n9819) );
  XNOR2_X1 U8780 ( .A(n9715), .B(n7339), .ZN(n7033) );
  NAND2_X1 U8781 ( .A1(n8890), .A2(n8577), .ZN(n7333) );
  INV_X1 U8782 ( .A(n7333), .ZN(n7032) );
  AOI21_X1 U8783 ( .B1(n7033), .B2(n9750), .A(n7032), .ZN(n9820) );
  OAI22_X1 U8784 ( .A1(n9394), .A2(n7034), .B1(n7337), .B2(n9741), .ZN(n7035)
         );
  AOI21_X1 U8785 ( .B1(n9410), .B2(n7339), .A(n7035), .ZN(n7036) );
  OAI21_X1 U8786 ( .B1(n9820), .B2(n9413), .A(n7036), .ZN(n7037) );
  AOI21_X1 U8787 ( .B1(n9819), .B2(n9755), .A(n7037), .ZN(n7038) );
  OAI21_X1 U8788 ( .B1(n7039), .B2(n9758), .A(n7038), .ZN(P1_U3284) );
  OAI222_X1 U8789 ( .A1(P1_U3086), .A2(n8737), .B1(n9562), .B2(n7041), .C1(
        n7040), .C2(n9559), .ZN(P1_U3334) );
  INV_X1 U8790 ( .A(n7808), .ZN(n7043) );
  NOR2_X1 U8791 ( .A1(n7806), .A2(n7043), .ZN(n7932) );
  XNOR2_X1 U8792 ( .A(n7042), .B(n7932), .ZN(n7044) );
  OAI222_X1 U8793 ( .A1(n8307), .A2(n7129), .B1(n10007), .B2(n7316), .C1(
        n10013), .C2(n7044), .ZN(n7110) );
  INV_X1 U8794 ( .A(n7110), .ZN(n7052) );
  NAND2_X1 U8795 ( .A1(n7115), .A2(n7045), .ZN(n7046) );
  XOR2_X1 U8796 ( .A(n7046), .B(n7932), .Z(n7111) );
  INV_X1 U8797 ( .A(n7047), .ZN(n7134) );
  AOI22_X1 U8798 ( .A1(n8334), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n9994), .B2(
        n7134), .ZN(n7048) );
  OAI21_X1 U8799 ( .B1(n7049), .B2(n8329), .A(n7048), .ZN(n7050) );
  AOI21_X1 U8800 ( .B1(n7111), .B2(n9996), .A(n7050), .ZN(n7051) );
  OAI21_X1 U8801 ( .B1(n7052), .B2(n8334), .A(n7051), .ZN(P2_U3225) );
  AND2_X1 U8802 ( .A1(n8648), .A2(n7056), .ZN(n8634) );
  NAND2_X1 U8803 ( .A1(n8634), .A2(n7054), .ZN(n8754) );
  AND2_X1 U8804 ( .A1(n7056), .A2(n7055), .ZN(n8755) );
  NAND3_X1 U8805 ( .A1(n8755), .A2(n8648), .A3(n8622), .ZN(n7057) );
  NAND2_X1 U8806 ( .A1(n4357), .A2(n7057), .ZN(n8794) );
  INV_X1 U8807 ( .A(n8890), .ZN(n7058) );
  NAND2_X1 U8808 ( .A1(n7154), .A2(n7058), .ZN(n8650) );
  OAI21_X1 U8809 ( .B1(n4406), .B2(n4636), .A(n7294), .ZN(n7061) );
  NAND2_X1 U8810 ( .A1(n8889), .A2(n8577), .ZN(n7060) );
  NAND2_X1 U8811 ( .A1(n8891), .A2(n9199), .ZN(n7059) );
  NAND2_X1 U8812 ( .A1(n7060), .A2(n7059), .ZN(n7362) );
  AOI21_X1 U8813 ( .B1(n7061), .B2(n9738), .A(n7362), .ZN(n9827) );
  OAI22_X1 U8814 ( .A1(n9394), .A2(n7062), .B1(n7359), .B2(n9741), .ZN(n7065)
         );
  INV_X1 U8815 ( .A(n7339), .ZN(n9821) );
  INV_X1 U8816 ( .A(n7154), .ZN(n9828) );
  OAI211_X1 U8817 ( .C1(n7063), .C2(n9828), .A(n9750), .B(n4405), .ZN(n9826)
         );
  NOR2_X1 U8818 ( .A1(n9826), .A2(n9413), .ZN(n7064) );
  AOI211_X1 U8819 ( .C1(n9410), .C2(n7154), .A(n7065), .B(n7064), .ZN(n7069)
         );
  OR2_X1 U8820 ( .A1(n7339), .A2(n8891), .ZN(n7067) );
  XNOR2_X1 U8821 ( .A(n7153), .B(n8758), .ZN(n9830) );
  NAND2_X1 U8822 ( .A1(n9830), .A2(n9755), .ZN(n7068) );
  OAI211_X1 U8823 ( .C1(n9827), .C2(n9758), .A(n7069), .B(n7068), .ZN(P1_U3283) );
  INV_X1 U8824 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U8825 ( .A1(n7079), .A2(n7070), .ZN(n7071) );
  INV_X1 U8826 ( .A(n7073), .ZN(n7075) );
  OAI21_X1 U8827 ( .B1(n7074), .B2(n7082), .A(n7073), .ZN(n7991) );
  NOR2_X1 U8828 ( .A1(n7094), .A2(n7991), .ZN(n7990) );
  AOI22_X1 U8829 ( .A1(n7093), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7088), .B2(
        n7234), .ZN(n7076) );
  AOI21_X1 U8830 ( .B1(n7077), .B2(n7076), .A(n7231), .ZN(n7109) );
  OR2_X1 U8831 ( .A1(n7079), .A2(n7078), .ZN(n7081) );
  INV_X1 U8832 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U8833 ( .A1(n7093), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n5208), .B2(
        n7234), .ZN(n7084) );
  AOI21_X1 U8834 ( .B1(n7085), .B2(n7084), .A(n7233), .ZN(n7086) );
  NOR2_X1 U8835 ( .A1(n7086), .A2(n9974), .ZN(n7107) );
  INV_X1 U8836 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7087) );
  NOR2_X1 U8837 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7087), .ZN(n7222) );
  INV_X1 U8838 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9588) );
  OAI22_X1 U8839 ( .A1(n9980), .A2(n7234), .B1(n9924), .B2(n9588), .ZN(n7106)
         );
  OR2_X1 U8840 ( .A1(n9882), .A2(n7088), .ZN(n7090) );
  NAND2_X1 U8841 ( .A1(n9882), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7089) );
  AND2_X1 U8842 ( .A1(n7090), .A2(n7089), .ZN(n7092) );
  AND2_X1 U8843 ( .A1(n7092), .A2(n7093), .ZN(n7242) );
  INV_X1 U8844 ( .A(n7242), .ZN(n7091) );
  OAI21_X1 U8845 ( .B1(n7093), .B2(n7092), .A(n7091), .ZN(n7103) );
  OR2_X1 U8846 ( .A1(n9882), .A2(n7094), .ZN(n7096) );
  NAND2_X1 U8847 ( .A1(n9882), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7095) );
  AND2_X1 U8848 ( .A1(n7096), .A2(n7095), .ZN(n7100) );
  AND2_X1 U8849 ( .A1(n7100), .A2(n7996), .ZN(n7101) );
  NOR2_X1 U8850 ( .A1(n7098), .A2(n7097), .ZN(n7994) );
  INV_X1 U8851 ( .A(n7101), .ZN(n7099) );
  OAI21_X1 U8852 ( .B1(n7996), .B2(n7100), .A(n7099), .ZN(n7995) );
  NOR2_X1 U8853 ( .A1(n7994), .A2(n7995), .ZN(n7993) );
  NOR2_X1 U8854 ( .A1(n7101), .A2(n7993), .ZN(n7102) );
  NOR2_X1 U8855 ( .A1(n7102), .A2(n7103), .ZN(n7241) );
  AOI21_X1 U8856 ( .B1(n7103), .B2(n7102), .A(n7241), .ZN(n7104) );
  NOR2_X1 U8857 ( .A1(n7104), .A2(n9917), .ZN(n7105) );
  NOR4_X1 U8858 ( .A1(n7107), .A2(n7222), .A3(n7106), .A4(n7105), .ZN(n7108)
         );
  OAI21_X1 U8859 ( .B1(n7109), .B2(n9965), .A(n7108), .ZN(P2_U3192) );
  AOI21_X1 U8860 ( .B1(n10068), .B2(n7111), .A(n7110), .ZN(n7114) );
  INV_X1 U8861 ( .A(n8450), .ZN(n8398) );
  AOI22_X1 U8862 ( .A1(n8398), .A2(n7139), .B1(n10076), .B2(
        P2_REG0_REG_8__SCAN_IN), .ZN(n7112) );
  OAI21_X1 U8863 ( .B1(n7114), .B2(n10076), .A(n7112), .ZN(P2_U3414) );
  INV_X1 U8864 ( .A(n8394), .ZN(n8338) );
  AOI22_X1 U8865 ( .A1(n8338), .A2(n7139), .B1(n10090), .B2(
        P2_REG1_REG_8__SCAN_IN), .ZN(n7113) );
  OAI21_X1 U8866 ( .B1(n7114), .B2(n10090), .A(n7113), .ZN(P2_U3467) );
  INV_X1 U8867 ( .A(n7115), .ZN(n7116) );
  AOI21_X1 U8868 ( .B1(n7117), .B2(n7804), .A(n7116), .ZN(n10047) );
  INV_X1 U8869 ( .A(n10047), .ZN(n7128) );
  NAND2_X1 U8870 ( .A1(n10016), .A2(n10015), .ZN(n8176) );
  XNOR2_X1 U8871 ( .A(n7118), .B(n5491), .ZN(n7122) );
  INV_X1 U8872 ( .A(n7985), .ZN(n7198) );
  OAI22_X1 U8873 ( .A1(n7198), .A2(n10007), .B1(n7119), .B2(n8307), .ZN(n7120)
         );
  AOI21_X1 U8874 ( .B1(n10047), .B2(n10010), .A(n7120), .ZN(n7121) );
  OAI21_X1 U8875 ( .B1(n10013), .B2(n7122), .A(n7121), .ZN(n10044) );
  NAND2_X1 U8876 ( .A1(n10044), .A2(n10016), .ZN(n7127) );
  OAI22_X1 U8877 ( .A1(n10016), .A2(n6890), .B1(n7123), .B2(n10002), .ZN(n7124) );
  AOI21_X1 U8878 ( .B1(n9993), .B2(n7125), .A(n7124), .ZN(n7126) );
  OAI211_X1 U8879 ( .C1(n7128), .C2(n8176), .A(n7127), .B(n7126), .ZN(P2_U3226) );
  NAND2_X1 U8880 ( .A1(n7130), .A2(n7129), .ZN(n7131) );
  XNOR2_X1 U8881 ( .A(n7571), .B(n7139), .ZN(n7197) );
  XNOR2_X1 U8882 ( .A(n7206), .B(n7197), .ZN(n7168) );
  XNOR2_X1 U8883 ( .A(n7168), .B(n7985), .ZN(n7141) );
  AOI21_X1 U8884 ( .B1(n7708), .B2(n9985), .A(n7133), .ZN(n7137) );
  NAND2_X1 U8885 ( .A1(n7734), .A2(n7134), .ZN(n7136) );
  NAND2_X1 U8886 ( .A1(n7717), .A2(n7984), .ZN(n7135) );
  NAND3_X1 U8887 ( .A1(n7137), .A2(n7136), .A3(n7135), .ZN(n7138) );
  AOI21_X1 U8888 ( .B1(n7139), .B2(n7721), .A(n7138), .ZN(n7140) );
  OAI21_X1 U8889 ( .B1(n7141), .B2(n7724), .A(n7140), .ZN(P2_U3161) );
  AOI211_X1 U8890 ( .C1(n7469), .C2(n7144), .A(n8921), .B(n8960), .ZN(n7152)
         );
  OAI21_X1 U8891 ( .B1(n7146), .B2(n6952), .A(n7145), .ZN(n8911) );
  XNOR2_X1 U8892 ( .A(n8919), .B(n8911), .ZN(n7147) );
  NAND2_X1 U8893 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7147), .ZN(n8913) );
  OAI211_X1 U8894 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7147), .A(n8975), .B(
        n8913), .ZN(n7150) );
  NAND2_X1 U8895 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8601) );
  INV_X1 U8896 ( .A(n8601), .ZN(n7148) );
  AOI21_X1 U8897 ( .B1(n9679), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n7148), .ZN(
        n7149) );
  OAI211_X1 U8898 ( .C1(n9689), .C2(n8919), .A(n7150), .B(n7149), .ZN(n7151)
         );
  OR2_X1 U8899 ( .A1(n7152), .A2(n7151), .ZN(P1_U3258) );
  INV_X1 U8900 ( .A(n8889), .ZN(n7155) );
  OR2_X1 U8901 ( .A1(n7305), .A2(n7155), .ZN(n8652) );
  NAND2_X1 U8902 ( .A1(n7305), .A2(n7155), .ZN(n8655) );
  NAND2_X1 U8903 ( .A1(n8652), .A2(n8655), .ZN(n7300) );
  XNOR2_X1 U8904 ( .A(n4298), .B(n7300), .ZN(n9835) );
  NAND2_X1 U8905 ( .A1(n9835), .A2(n9709), .ZN(n7161) );
  NAND2_X1 U8906 ( .A1(n7294), .A2(n8650), .ZN(n7156) );
  INV_X1 U8907 ( .A(n7300), .ZN(n8761) );
  XNOR2_X1 U8908 ( .A(n7156), .B(n8761), .ZN(n7159) );
  NAND2_X1 U8909 ( .A1(n8888), .A2(n8577), .ZN(n7158) );
  NAND2_X1 U8910 ( .A1(n8890), .A2(n9199), .ZN(n7157) );
  NAND2_X1 U8911 ( .A1(n7158), .A2(n7157), .ZN(n7447) );
  AOI21_X1 U8912 ( .B1(n7159), .B2(n9738), .A(n7447), .ZN(n7160) );
  INV_X1 U8913 ( .A(n7305), .ZN(n9833) );
  XNOR2_X1 U8914 ( .A(n4405), .B(n9833), .ZN(n7162) );
  NAND2_X1 U8915 ( .A1(n7162), .A2(n9750), .ZN(n9832) );
  OAI22_X1 U8916 ( .A1(n9394), .A2(n7163), .B1(n7444), .B2(n9741), .ZN(n7164)
         );
  AOI21_X1 U8917 ( .B1(n7305), .B2(n9410), .A(n7164), .ZN(n7165) );
  OAI21_X1 U8918 ( .B1(n9832), .B2(n9413), .A(n7165), .ZN(n7166) );
  AOI21_X1 U8919 ( .B1(n9835), .B2(n9719), .A(n7166), .ZN(n7167) );
  OAI21_X1 U8920 ( .B1(n9837), .B2(n9758), .A(n7167), .ZN(P1_U3282) );
  INV_X1 U8921 ( .A(n7197), .ZN(n7199) );
  AOI22_X1 U8922 ( .A1(n7168), .A2(n7198), .B1(n7206), .B2(n7199), .ZN(n7170)
         );
  XNOR2_X1 U8923 ( .A(n10049), .B(n7571), .ZN(n7200) );
  XNOR2_X1 U8924 ( .A(n7200), .B(n7984), .ZN(n7169) );
  XNOR2_X1 U8925 ( .A(n7170), .B(n7169), .ZN(n7176) );
  INV_X1 U8926 ( .A(n7183), .ZN(n7174) );
  NOR2_X1 U8927 ( .A1(n7737), .A2(n10049), .ZN(n7173) );
  NAND2_X1 U8928 ( .A1(n7708), .A2(n7985), .ZN(n7171) );
  NAND2_X1 U8929 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7997) );
  OAI211_X1 U8930 ( .C1(n7431), .C2(n7731), .A(n7171), .B(n7997), .ZN(n7172)
         );
  AOI211_X1 U8931 ( .C1(n7174), .C2(n7734), .A(n7173), .B(n7172), .ZN(n7175)
         );
  OAI21_X1 U8932 ( .B1(n7176), .B2(n7724), .A(n7175), .ZN(P2_U3171) );
  OAI21_X1 U8933 ( .B1(n7177), .B2(n7933), .A(n7313), .ZN(n10050) );
  XNOR2_X1 U8934 ( .A(n7178), .B(n7933), .ZN(n7179) );
  NAND2_X1 U8935 ( .A1(n7179), .A2(n9987), .ZN(n7181) );
  AOI22_X1 U8936 ( .A1(n9982), .A2(n7985), .B1(n7983), .B2(n9984), .ZN(n7180)
         );
  OAI211_X1 U8937 ( .C1(n7182), .C2(n10050), .A(n7181), .B(n7180), .ZN(n10052)
         );
  NAND2_X1 U8938 ( .A1(n10052), .A2(n10016), .ZN(n7187) );
  OAI22_X1 U8939 ( .A1(n10016), .A2(n7094), .B1(n7183), .B2(n10002), .ZN(n7184) );
  AOI21_X1 U8940 ( .B1(n9993), .B2(n7185), .A(n7184), .ZN(n7186) );
  OAI211_X1 U8941 ( .C1(n10050), .C2(n8176), .A(n7187), .B(n7186), .ZN(
        P2_U3224) );
  INV_X1 U8942 ( .A(n7188), .ZN(n7605) );
  OAI222_X1 U8943 ( .A1(n8456), .A2(n7189), .B1(n8467), .B2(n7605), .C1(n7761), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  NAND2_X1 U8944 ( .A1(n7193), .A2(n7190), .ZN(n7191) );
  OAI211_X1 U8945 ( .C1(n7192), .C2(n9554), .A(n7191), .B(n8882), .ZN(P1_U3332) );
  NAND2_X1 U8946 ( .A1(n7193), .A2(n8458), .ZN(n7195) );
  NAND2_X1 U8947 ( .A1(n7194), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7964) );
  OAI211_X1 U8948 ( .C1(n7196), .C2(n8456), .A(n7195), .B(n7964), .ZN(P2_U3272) );
  INV_X1 U8949 ( .A(n10065), .ZN(n7217) );
  NAND2_X1 U8950 ( .A1(n7200), .A2(n7316), .ZN(n7203) );
  OAI21_X1 U8951 ( .B1(n7197), .B2(n7985), .A(n7203), .ZN(n7205) );
  NOR2_X1 U8952 ( .A1(n7199), .A2(n7198), .ZN(n7202) );
  INV_X1 U8953 ( .A(n7200), .ZN(n7201) );
  AOI22_X1 U8954 ( .A1(n7203), .A2(n7202), .B1(n7201), .B2(n7984), .ZN(n7204)
         );
  INV_X1 U8955 ( .A(n7208), .ZN(n7207) );
  NAND2_X1 U8956 ( .A1(n7207), .A2(n7431), .ZN(n7218) );
  XNOR2_X1 U8957 ( .A(n7323), .B(n7571), .ZN(n7220) );
  NAND2_X1 U8958 ( .A1(n7218), .A2(n7220), .ZN(n7209) );
  NAND2_X1 U8959 ( .A1(n7208), .A2(n7983), .ZN(n7219) );
  NAND2_X1 U8960 ( .A1(n7209), .A2(n7219), .ZN(n7211) );
  XNOR2_X1 U8961 ( .A(n7422), .B(n7583), .ZN(n7342) );
  OAI211_X1 U8962 ( .C1(n7211), .C2(n7342), .A(n7345), .B(n7727), .ZN(n7216)
         );
  INV_X1 U8963 ( .A(n7432), .ZN(n7214) );
  AND2_X1 U8964 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7248) );
  AOI21_X1 U8965 ( .B1(n7708), .B2(n7983), .A(n7248), .ZN(n7212) );
  OAI21_X1 U8966 ( .B1(n7826), .B2(n7731), .A(n7212), .ZN(n7213) );
  AOI21_X1 U8967 ( .B1(n7214), .B2(n7734), .A(n7213), .ZN(n7215) );
  OAI211_X1 U8968 ( .C1(n7217), .C2(n7737), .A(n7216), .B(n7215), .ZN(P2_U3176) );
  NAND2_X1 U8969 ( .A1(n7218), .A2(n7219), .ZN(n7221) );
  XNOR2_X1 U8970 ( .A(n7221), .B(n7220), .ZN(n7229) );
  AOI21_X1 U8971 ( .B1(n7708), .B2(n7984), .A(n7222), .ZN(n7227) );
  NAND2_X1 U8972 ( .A1(n7323), .A2(n7721), .ZN(n7226) );
  INV_X1 U8973 ( .A(n7321), .ZN(n7223) );
  NAND2_X1 U8974 ( .A1(n7734), .A2(n7223), .ZN(n7225) );
  NAND2_X1 U8975 ( .A1(n7717), .A2(n7982), .ZN(n7224) );
  NAND4_X1 U8976 ( .A1(n7227), .A2(n7226), .A3(n7225), .A4(n7224), .ZN(n7228)
         );
  AOI21_X1 U8977 ( .B1(n7229), .B2(n7727), .A(n7228), .ZN(n7230) );
  INV_X1 U8978 ( .A(n7230), .ZN(P2_U3157) );
  AOI21_X1 U8979 ( .B1(n7433), .B2(n7232), .A(n7261), .ZN(n7251) );
  INV_X1 U8980 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10088) );
  AOI21_X1 U8981 ( .B1(n10088), .B2(n7235), .A(n7269), .ZN(n7236) );
  NOR2_X1 U8982 ( .A1(n7236), .A2(n9974), .ZN(n7249) );
  INV_X1 U8983 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n9592) );
  OAI22_X1 U8984 ( .A1(n9980), .A2(n4511), .B1(n9924), .B2(n9592), .ZN(n7247)
         );
  OR2_X1 U8985 ( .A1(n9882), .A2(n7433), .ZN(n7238) );
  NAND2_X1 U8986 ( .A1(n9882), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7237) );
  AND2_X1 U8987 ( .A1(n7238), .A2(n7237), .ZN(n7240) );
  AND2_X1 U8988 ( .A1(n7240), .A2(n7268), .ZN(n7253) );
  INV_X1 U8989 ( .A(n7253), .ZN(n7239) );
  OAI21_X1 U8990 ( .B1(n7268), .B2(n7240), .A(n7239), .ZN(n7244) );
  NOR2_X1 U8991 ( .A1(n7242), .A2(n7241), .ZN(n7243) );
  NOR2_X1 U8992 ( .A1(n7243), .A2(n7244), .ZN(n7252) );
  AOI21_X1 U8993 ( .B1(n7244), .B2(n7243), .A(n7252), .ZN(n7245) );
  NOR2_X1 U8994 ( .A1(n7245), .A2(n9917), .ZN(n7246) );
  NOR4_X1 U8995 ( .A1(n7249), .A2(n7248), .A3(n7247), .A4(n7246), .ZN(n7250)
         );
  OAI21_X1 U8996 ( .B1(n7251), .B2(n9965), .A(n7250), .ZN(P2_U3193) );
  NOR2_X1 U8997 ( .A1(n7253), .A2(n7252), .ZN(n8010) );
  OR2_X1 U8998 ( .A1(n9882), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U8999 ( .A1(n9882), .A2(n7254), .ZN(n7255) );
  AND3_X1 U9000 ( .A1(n7256), .A2(n7255), .A3(n8023), .ZN(n8008) );
  INV_X1 U9001 ( .A(n8008), .ZN(n7258) );
  INV_X1 U9002 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7453) );
  AOI21_X1 U9003 ( .B1(n9882), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8023), .ZN(
        n7257) );
  OAI21_X1 U9004 ( .B1(n9882), .B2(n7453), .A(n7257), .ZN(n8009) );
  NAND2_X1 U9005 ( .A1(n7258), .A2(n8009), .ZN(n7259) );
  XNOR2_X1 U9006 ( .A(n8010), .B(n7259), .ZN(n7280) );
  NOR2_X1 U9007 ( .A1(n7268), .A2(n7260), .ZN(n7262) );
  NAND2_X1 U9008 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8023), .ZN(n7263) );
  OAI21_X1 U9009 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8023), .A(n7263), .ZN(
        n7264) );
  AOI21_X1 U9010 ( .B1(n7265), .B2(n7264), .A(n8025), .ZN(n7266) );
  NOR2_X1 U9011 ( .A1(n7266), .A2(n9965), .ZN(n7279) );
  NAND2_X1 U9012 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8023), .ZN(n7270) );
  OAI21_X1 U9013 ( .B1(n8023), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7270), .ZN(
        n7271) );
  NOR2_X1 U9014 ( .A1(n7272), .A2(n7271), .ZN(n8013) );
  AOI21_X1 U9015 ( .B1(n7272), .B2(n7271), .A(n8013), .ZN(n7277) );
  NOR2_X1 U9016 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7273), .ZN(n7348) );
  INV_X1 U9017 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9596) );
  NOR2_X1 U9018 ( .A1(n9924), .A2(n9596), .ZN(n7274) );
  AOI211_X1 U9019 ( .C1(n7275), .C2(n9914), .A(n7348), .B(n7274), .ZN(n7276)
         );
  OAI21_X1 U9020 ( .B1(n7277), .B2(n9974), .A(n7276), .ZN(n7278) );
  AOI211_X1 U9021 ( .C1(n7280), .C2(n9970), .A(n7279), .B(n7278), .ZN(n7281)
         );
  INV_X1 U9022 ( .A(n7281), .ZN(P2_U3194) );
  XNOR2_X1 U9023 ( .A(n7282), .B(n7283), .ZN(n7284) );
  NAND2_X1 U9024 ( .A1(n7284), .A2(n7285), .ZN(n7326) );
  OAI21_X1 U9025 ( .B1(n7285), .B2(n7284), .A(n7326), .ZN(n7286) );
  NAND2_X1 U9026 ( .A1(n7286), .A2(n9649), .ZN(n7293) );
  INV_X1 U9027 ( .A(n9710), .ZN(n7291) );
  NAND2_X1 U9028 ( .A1(n8891), .A2(n8988), .ZN(n7288) );
  NAND2_X1 U9029 ( .A1(n8893), .A2(n9199), .ZN(n7287) );
  AND2_X1 U9030 ( .A1(n7288), .A2(n7287), .ZN(n9705) );
  OAI22_X1 U9031 ( .A1(n9705), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7289), .ZN(n7290) );
  AOI21_X1 U9032 ( .B1(n7291), .B2(n8591), .A(n7290), .ZN(n7292) );
  OAI211_X1 U9033 ( .C1(n9813), .C2(n8594), .A(n7293), .B(n7292), .ZN(P1_U3221) );
  AND2_X1 U9034 ( .A1(n8655), .A2(n8650), .ZN(n8639) );
  NAND2_X1 U9035 ( .A1(n7294), .A2(n8639), .ZN(n7295) );
  INV_X1 U9036 ( .A(n8888), .ZN(n7296) );
  NAND2_X1 U9037 ( .A1(n7510), .A2(n7296), .ZN(n8656) );
  XNOR2_X1 U9038 ( .A(n7378), .B(n7371), .ZN(n7299) );
  NAND2_X1 U9039 ( .A1(n8887), .A2(n8577), .ZN(n7298) );
  NAND2_X1 U9040 ( .A1(n8889), .A2(n9199), .ZN(n7297) );
  NAND2_X1 U9041 ( .A1(n7298), .A2(n7297), .ZN(n7500) );
  AOI21_X1 U9042 ( .B1(n7299), .B2(n9738), .A(n7500), .ZN(n9840) );
  NAND2_X1 U9043 ( .A1(n7301), .A2(n7300), .ZN(n7303) );
  OR2_X1 U9044 ( .A1(n7305), .A2(n8889), .ZN(n7302) );
  NAND2_X1 U9045 ( .A1(n7303), .A2(n7302), .ZN(n7372) );
  XNOR2_X1 U9046 ( .A(n7372), .B(n7371), .ZN(n9843) );
  NAND2_X1 U9047 ( .A1(n9843), .A2(n9755), .ZN(n7311) );
  OAI22_X1 U9048 ( .A1(n9394), .A2(n7304), .B1(n7502), .B2(n9741), .ZN(n7309)
         );
  INV_X1 U9049 ( .A(n7510), .ZN(n9841) );
  INV_X1 U9050 ( .A(n7397), .ZN(n7307) );
  OAI211_X1 U9051 ( .C1(n9841), .C2(n4646), .A(n7307), .B(n9750), .ZN(n9839)
         );
  NOR2_X1 U9052 ( .A1(n9839), .A2(n9413), .ZN(n7308) );
  AOI211_X1 U9053 ( .C1(n9410), .C2(n7510), .A(n7309), .B(n7308), .ZN(n7310)
         );
  OAI211_X1 U9054 ( .C1(n9758), .C2(n9840), .A(n7311), .B(n7310), .ZN(P1_U3281) );
  NAND2_X1 U9055 ( .A1(n7313), .A2(n7312), .ZN(n7314) );
  NAND2_X1 U9056 ( .A1(n7820), .A2(n7816), .ZN(n7935) );
  XNOR2_X1 U9057 ( .A(n7314), .B(n7935), .ZN(n7318) );
  INV_X1 U9058 ( .A(n7318), .ZN(n10057) );
  XOR2_X1 U9059 ( .A(n7935), .B(n7315), .Z(n7320) );
  OAI22_X1 U9060 ( .A1(n7316), .A2(n8307), .B1(n7817), .B2(n10007), .ZN(n7317)
         );
  AOI21_X1 U9061 ( .B1(n7318), .B2(n10010), .A(n7317), .ZN(n7319) );
  OAI21_X1 U9062 ( .B1(n7320), .B2(n10013), .A(n7319), .ZN(n10059) );
  NAND2_X1 U9063 ( .A1(n10059), .A2(n10016), .ZN(n7325) );
  OAI22_X1 U9064 ( .A1(n10016), .A2(n7088), .B1(n7321), .B2(n10002), .ZN(n7322) );
  AOI21_X1 U9065 ( .B1(n9993), .B2(n7323), .A(n7322), .ZN(n7324) );
  OAI211_X1 U9066 ( .C1(n10057), .C2(n8176), .A(n7325), .B(n7324), .ZN(
        P2_U3223) );
  OAI21_X1 U9067 ( .B1(n7327), .B2(n7282), .A(n7326), .ZN(n7331) );
  NAND2_X1 U9068 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  XNOR2_X1 U9069 ( .A(n7331), .B(n7330), .ZN(n7341) );
  NAND2_X1 U9070 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  NAND2_X1 U9071 ( .A1(n7334), .A2(n8599), .ZN(n7336) );
  OAI211_X1 U9072 ( .C1(n9674), .C2(n7337), .A(n7336), .B(n7335), .ZN(n7338)
         );
  AOI21_X1 U9073 ( .B1(n7339), .B2(n9670), .A(n7338), .ZN(n7340) );
  OAI21_X1 U9074 ( .B1(n7341), .B2(n9665), .A(n7340), .ZN(P1_U3231) );
  INV_X1 U9075 ( .A(n10072), .ZN(n7354) );
  INV_X1 U9076 ( .A(n7342), .ZN(n7343) );
  NAND2_X1 U9077 ( .A1(n7343), .A2(n7982), .ZN(n7344) );
  NAND2_X1 U9078 ( .A1(n7345), .A2(n7344), .ZN(n7347) );
  XNOR2_X1 U9079 ( .A(n10072), .B(n7583), .ZN(n7405) );
  XNOR2_X1 U9080 ( .A(n7405), .B(n7981), .ZN(n7346) );
  OAI211_X1 U9081 ( .C1(n7347), .C2(n7346), .A(n7408), .B(n7727), .ZN(n7353)
         );
  INV_X1 U9082 ( .A(n7452), .ZN(n7351) );
  AOI21_X1 U9083 ( .B1(n7708), .B2(n7982), .A(n7348), .ZN(n7349) );
  OAI21_X1 U9084 ( .B1(n7538), .B2(n7731), .A(n7349), .ZN(n7350) );
  AOI21_X1 U9085 ( .B1(n7351), .B2(n7734), .A(n7350), .ZN(n7352) );
  OAI211_X1 U9086 ( .C1(n7354), .C2(n7737), .A(n7353), .B(n7352), .ZN(P2_U3164) );
  OAI21_X1 U9087 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(n7358) );
  NAND2_X1 U9088 ( .A1(n7358), .A2(n9649), .ZN(n7364) );
  NOR2_X1 U9089 ( .A1(n9674), .A2(n7359), .ZN(n7360) );
  AOI211_X1 U9090 ( .C1(n8599), .C2(n7362), .A(n7361), .B(n7360), .ZN(n7363)
         );
  OAI211_X1 U9091 ( .C1(n9828), .C2(n8594), .A(n7364), .B(n7363), .ZN(P1_U3217) );
  INV_X1 U9092 ( .A(n7365), .ZN(n7369) );
  OAI222_X1 U9093 ( .A1(n8456), .A2(n7367), .B1(n8467), .B2(n7369), .C1(n7366), 
        .C2(P2_U3151), .ZN(P2_U3271) );
  OAI222_X1 U9094 ( .A1(n7370), .A2(P1_U3086), .B1(n9562), .B2(n7369), .C1(
        n7368), .C2(n9559), .ZN(P1_U3331) );
  OR2_X1 U9095 ( .A1(n7510), .A2(n8888), .ZN(n7373) );
  INV_X1 U9096 ( .A(n8887), .ZN(n7375) );
  OR2_X1 U9097 ( .A1(n7400), .A2(n7375), .ZN(n8661) );
  NAND2_X1 U9098 ( .A1(n7400), .A2(n7375), .ZN(n8799) );
  NAND2_X1 U9099 ( .A1(n8661), .A2(n8799), .ZN(n7402) );
  OR2_X1 U9100 ( .A1(n7400), .A2(n8887), .ZN(n7376) );
  INV_X1 U9101 ( .A(n8886), .ZN(n7377) );
  NAND2_X1 U9102 ( .A1(n8476), .A2(n7377), .ZN(n8662) );
  XNOR2_X1 U9103 ( .A(n7474), .B(n8763), .ZN(n9857) );
  NAND2_X1 U9104 ( .A1(n7378), .A2(n8762), .ZN(n7379) );
  XNOR2_X1 U9105 ( .A(n7462), .B(n8763), .ZN(n7383) );
  NAND2_X1 U9106 ( .A1(n8885), .A2(n8577), .ZN(n7381) );
  NAND2_X1 U9107 ( .A1(n8887), .A2(n9199), .ZN(n7380) );
  NAND2_X1 U9108 ( .A1(n7381), .A2(n7380), .ZN(n8471) );
  INV_X1 U9109 ( .A(n8471), .ZN(n7382) );
  OAI21_X1 U9110 ( .B1(n7383), .B2(n9706), .A(n7382), .ZN(n7384) );
  AOI21_X1 U9111 ( .B1(n9857), .B2(n9709), .A(n7384), .ZN(n9859) );
  INV_X1 U9112 ( .A(n7400), .ZN(n9847) );
  INV_X1 U9113 ( .A(n8476), .ZN(n9854) );
  OAI211_X1 U9114 ( .C1(n7395), .C2(n9854), .A(n9750), .B(n7470), .ZN(n9852)
         );
  OAI22_X1 U9115 ( .A1(n9394), .A2(n7385), .B1(n8474), .B2(n9741), .ZN(n7386)
         );
  AOI21_X1 U9116 ( .B1(n8476), .B2(n9410), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9117 ( .B1(n9852), .B2(n9413), .A(n7387), .ZN(n7388) );
  AOI21_X1 U9118 ( .B1(n9857), .B2(n9719), .A(n7388), .ZN(n7389) );
  OAI21_X1 U9119 ( .B1(n9859), .B2(n9758), .A(n7389), .ZN(P1_U3279) );
  OAI21_X1 U9120 ( .B1(n4394), .B2(n4635), .A(n7390), .ZN(n7393) );
  NAND2_X1 U9121 ( .A1(n8886), .A2(n8577), .ZN(n7392) );
  NAND2_X1 U9122 ( .A1(n8888), .A2(n9199), .ZN(n7391) );
  NAND2_X1 U9123 ( .A1(n7392), .A2(n7391), .ZN(n7519) );
  AOI21_X1 U9124 ( .B1(n7393), .B2(n9738), .A(n7519), .ZN(n9846) );
  OAI22_X1 U9125 ( .A1(n9394), .A2(n7394), .B1(n7516), .B2(n9741), .ZN(n7399)
         );
  INV_X1 U9126 ( .A(n7395), .ZN(n7396) );
  OAI211_X1 U9127 ( .C1(n9847), .C2(n7397), .A(n7396), .B(n9750), .ZN(n9845)
         );
  NOR2_X1 U9128 ( .A1(n9845), .A2(n9413), .ZN(n7398) );
  AOI211_X1 U9129 ( .C1(n9410), .C2(n7400), .A(n7399), .B(n7398), .ZN(n7404)
         );
  XNOR2_X1 U9130 ( .A(n7401), .B(n7402), .ZN(n9849) );
  NAND2_X1 U9131 ( .A1(n9849), .A2(n9755), .ZN(n7403) );
  OAI211_X1 U9132 ( .C1(n9846), .C2(n9758), .A(n7404), .B(n7403), .ZN(P1_U3280) );
  INV_X1 U9133 ( .A(n9627), .ZN(n7415) );
  INV_X1 U9134 ( .A(n7405), .ZN(n7406) );
  NAND2_X1 U9135 ( .A1(n7406), .A2(n7981), .ZN(n7407) );
  NAND2_X1 U9136 ( .A1(n7408), .A2(n7407), .ZN(n7410) );
  XNOR2_X1 U9137 ( .A(n9627), .B(n7210), .ZN(n7479) );
  XNOR2_X1 U9138 ( .A(n7479), .B(n7980), .ZN(n7409) );
  NAND2_X1 U9139 ( .A1(n7410), .A2(n7409), .ZN(n7482) );
  OAI211_X1 U9140 ( .C1(n7410), .C2(n7409), .A(n7482), .B(n7727), .ZN(n7414)
         );
  NAND2_X1 U9141 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3151), .ZN(n8017) );
  OAI21_X1 U9142 ( .B1(n7730), .B2(n7826), .A(n8017), .ZN(n7412) );
  NOR2_X1 U9143 ( .A1(n7719), .A2(n7496), .ZN(n7411) );
  AOI211_X1 U9144 ( .C1(n7717), .C2(n7979), .A(n7412), .B(n7411), .ZN(n7413)
         );
  OAI211_X1 U9145 ( .C1(n7415), .C2(n7737), .A(n7414), .B(n7413), .ZN(P2_U3174) );
  INV_X1 U9146 ( .A(n7416), .ZN(n7420) );
  OAI222_X1 U9147 ( .A1(n8457), .A2(n7420), .B1(P2_U3151), .B2(n7418), .C1(
        n7417), .C2(n8456), .ZN(P2_U3270) );
  OAI222_X1 U9148 ( .A1(P1_U3086), .A2(n7421), .B1(n9562), .B2(n7420), .C1(
        n7419), .C2(n9559), .ZN(P1_U3330) );
  INV_X1 U9149 ( .A(n7422), .ZN(n7936) );
  XNOR2_X1 U9150 ( .A(n7423), .B(n7936), .ZN(n10062) );
  INV_X1 U9151 ( .A(n7424), .ZN(n7426) );
  NAND2_X1 U9152 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  OAI211_X1 U9153 ( .C1(n7936), .C2(n7428), .A(n7427), .B(n9987), .ZN(n7430)
         );
  NAND2_X1 U9154 ( .A1(n7981), .A2(n9984), .ZN(n7429) );
  OAI211_X1 U9155 ( .C1(n7431), .C2(n8307), .A(n7430), .B(n7429), .ZN(n10063)
         );
  NAND2_X1 U9156 ( .A1(n10063), .A2(n10016), .ZN(n7436) );
  OAI22_X1 U9157 ( .A1(n10016), .A2(n7433), .B1(n7432), .B2(n10002), .ZN(n7434) );
  AOI21_X1 U9158 ( .B1(n10065), .B2(n9993), .A(n7434), .ZN(n7435) );
  OAI211_X1 U9159 ( .C1(n10062), .C2(n7543), .A(n7436), .B(n7435), .ZN(
        P2_U3222) );
  INV_X1 U9160 ( .A(n7355), .ZN(n7440) );
  INV_X1 U9161 ( .A(n7437), .ZN(n7439) );
  NOR3_X1 U9162 ( .A1(n7440), .A2(n7439), .A3(n7438), .ZN(n7443) );
  INV_X1 U9163 ( .A(n7441), .ZN(n7442) );
  OAI21_X1 U9164 ( .B1(n7443), .B2(n7442), .A(n9649), .ZN(n7449) );
  NOR2_X1 U9165 ( .A1(n9674), .A2(n7444), .ZN(n7445) );
  AOI211_X1 U9166 ( .C1(n8599), .C2(n7447), .A(n7446), .B(n7445), .ZN(n7448)
         );
  OAI211_X1 U9167 ( .C1(n9833), .C2(n8594), .A(n7449), .B(n7448), .ZN(P1_U3236) );
  XNOR2_X1 U9168 ( .A(n7450), .B(n7938), .ZN(n7451) );
  OAI222_X1 U9169 ( .A1(n10007), .A2(n7538), .B1(n8307), .B2(n7817), .C1(
        n10013), .C2(n7451), .ZN(n10070) );
  INV_X1 U9170 ( .A(n10070), .ZN(n7458) );
  OAI22_X1 U9171 ( .A1(n10016), .A2(n7453), .B1(n7452), .B2(n10002), .ZN(n7454) );
  AOI21_X1 U9172 ( .B1(n10072), .B2(n9993), .A(n7454), .ZN(n7457) );
  NAND2_X1 U9173 ( .A1(n7455), .A2(n7938), .ZN(n10067) );
  NAND3_X1 U9174 ( .A1(n10069), .A2(n10067), .A3(n9996), .ZN(n7456) );
  OAI211_X1 U9175 ( .C1(n7458), .C2(n8334), .A(n7457), .B(n7456), .ZN(P2_U3221) );
  INV_X1 U9176 ( .A(n7459), .ZN(n9561) );
  OAI222_X1 U9177 ( .A1(n8457), .A2(n9561), .B1(P2_U3151), .B2(n7461), .C1(
        n7460), .C2(n8456), .ZN(P2_U3269) );
  INV_X1 U9178 ( .A(n7464), .ZN(n7465) );
  INV_X1 U9179 ( .A(n8885), .ZN(n9137) );
  OR2_X1 U9180 ( .A1(n9139), .A2(n9137), .ZN(n8665) );
  NAND2_X1 U9181 ( .A1(n9139), .A2(n9137), .ZN(n8836) );
  NAND2_X1 U9182 ( .A1(n8665), .A2(n8836), .ZN(n7463) );
  INV_X1 U9183 ( .A(n7463), .ZN(n8766) );
  OAI21_X1 U9184 ( .B1(n7465), .B2(n8766), .A(n8837), .ZN(n7468) );
  NAND2_X1 U9185 ( .A1(n9141), .A2(n8577), .ZN(n7467) );
  NAND2_X1 U9186 ( .A1(n8886), .A2(n9199), .ZN(n7466) );
  NAND2_X1 U9187 ( .A1(n7467), .A2(n7466), .ZN(n8600) );
  AOI21_X1 U9188 ( .B1(n7468), .B2(n9738), .A(n8600), .ZN(n9640) );
  OAI22_X1 U9189 ( .A1(n9394), .A2(n7469), .B1(n8603), .B2(n9741), .ZN(n7473)
         );
  INV_X1 U9190 ( .A(n7470), .ZN(n7471) );
  INV_X1 U9191 ( .A(n9139), .ZN(n9641) );
  OAI211_X1 U9192 ( .C1(n7471), .C2(n9641), .A(n9750), .B(n9404), .ZN(n9639)
         );
  NOR2_X1 U9193 ( .A1(n9639), .A2(n9413), .ZN(n7472) );
  AOI211_X1 U9194 ( .C1(n9410), .C2(n9139), .A(n7473), .B(n7472), .ZN(n7478)
         );
  NAND2_X1 U9195 ( .A1(n8476), .A2(n8886), .ZN(n7475) );
  XNOR2_X1 U9196 ( .A(n9138), .B(n8766), .ZN(n9643) );
  NAND2_X1 U9197 ( .A1(n9643), .A2(n9755), .ZN(n7477) );
  OAI211_X1 U9198 ( .C1(n9640), .C2(n9758), .A(n7478), .B(n7477), .ZN(P1_U3278) );
  XNOR2_X1 U9199 ( .A(n9619), .B(n7583), .ZN(n7522) );
  XNOR2_X1 U9200 ( .A(n7522), .B(n8326), .ZN(n7487) );
  INV_X1 U9201 ( .A(n7479), .ZN(n7480) );
  NAND2_X1 U9202 ( .A1(n7480), .A2(n7980), .ZN(n7481) );
  NAND2_X1 U9203 ( .A1(n7482), .A2(n7481), .ZN(n7486) );
  INV_X1 U9204 ( .A(n7486), .ZN(n7484) );
  INV_X1 U9205 ( .A(n7487), .ZN(n7483) );
  INV_X1 U9206 ( .A(n7524), .ZN(n7485) );
  AOI21_X1 U9207 ( .B1(n7487), .B2(n7486), .A(n7485), .ZN(n7492) );
  AOI22_X1 U9208 ( .A1(n7708), .A2(n7980), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n7489) );
  INV_X1 U9209 ( .A(n8308), .ZN(n7978) );
  NAND2_X1 U9210 ( .A1(n7717), .A2(n7978), .ZN(n7488) );
  OAI211_X1 U9211 ( .C1(n7719), .C2(n7539), .A(n7489), .B(n7488), .ZN(n7490)
         );
  AOI21_X1 U9212 ( .B1(n9619), .B2(n7721), .A(n7490), .ZN(n7491) );
  OAI21_X1 U9213 ( .B1(n7492), .B2(n7724), .A(n7491), .ZN(P2_U3155) );
  XNOR2_X1 U9214 ( .A(n7493), .B(n7923), .ZN(n9624) );
  XNOR2_X1 U9215 ( .A(n7494), .B(n7923), .ZN(n7495) );
  OAI222_X1 U9216 ( .A1(n10007), .A2(n8326), .B1(n8307), .B2(n7826), .C1(
        n10013), .C2(n7495), .ZN(n9625) );
  NAND2_X1 U9217 ( .A1(n9625), .A2(n10016), .ZN(n7499) );
  INV_X1 U9218 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8027) );
  OAI22_X1 U9219 ( .A1(n10016), .A2(n8027), .B1(n7496), .B2(n10002), .ZN(n7497) );
  AOI21_X1 U9220 ( .B1(n9627), .B2(n9993), .A(n7497), .ZN(n7498) );
  OAI211_X1 U9221 ( .C1(n9624), .C2(n7543), .A(n7499), .B(n7498), .ZN(P2_U3220) );
  NAND2_X1 U9222 ( .A1(n7500), .A2(n8599), .ZN(n7501) );
  NAND2_X1 U9223 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9696) );
  OAI211_X1 U9224 ( .C1(n9674), .C2(n7502), .A(n7501), .B(n9696), .ZN(n7509)
         );
  INV_X1 U9225 ( .A(n7503), .ZN(n7504) );
  NAND3_X1 U9226 ( .A1(n7441), .A2(n7505), .A3(n7504), .ZN(n7506) );
  AOI21_X1 U9227 ( .B1(n7507), .B2(n7506), .A(n9665), .ZN(n7508) );
  AOI211_X1 U9228 ( .C1(n7510), .C2(n9670), .A(n7509), .B(n7508), .ZN(n7511)
         );
  INV_X1 U9229 ( .A(n7511), .ZN(P1_U3224) );
  OAI21_X1 U9230 ( .B1(n7514), .B2(n7513), .A(n7512), .ZN(n7515) );
  NAND2_X1 U9231 ( .A1(n7515), .A2(n9649), .ZN(n7521) );
  NOR2_X1 U9232 ( .A1(n9674), .A2(n7516), .ZN(n7517) );
  AOI211_X1 U9233 ( .C1(n8599), .C2(n7519), .A(n7518), .B(n7517), .ZN(n7520)
         );
  OAI211_X1 U9234 ( .C1(n9847), .C2(n8594), .A(n7521), .B(n7520), .ZN(P1_U3234) );
  NAND2_X1 U9235 ( .A1(n7522), .A2(n8326), .ZN(n7523) );
  XNOR2_X1 U9236 ( .A(n7525), .B(n7210), .ZN(n7544) );
  XNOR2_X1 U9237 ( .A(n7544), .B(n8308), .ZN(n7527) );
  AOI21_X1 U9238 ( .B1(n7526), .B2(n7527), .A(n7724), .ZN(n7529) );
  INV_X1 U9239 ( .A(n7527), .ZN(n7528) );
  NAND2_X1 U9240 ( .A1(n7529), .A2(n7546), .ZN(n7533) );
  NAND2_X1 U9241 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8056) );
  OAI21_X1 U9242 ( .B1(n7730), .B2(n8326), .A(n8056), .ZN(n7531) );
  NOR2_X1 U9243 ( .A1(n7719), .A2(n8330), .ZN(n7530) );
  AOI211_X1 U9244 ( .C1(n7717), .C2(n5299), .A(n7531), .B(n7530), .ZN(n7532)
         );
  OAI211_X1 U9245 ( .C1(n8451), .C2(n7737), .A(n7533), .B(n7532), .ZN(P2_U3181) );
  INV_X1 U9246 ( .A(n7535), .ZN(n7942) );
  XNOR2_X1 U9247 ( .A(n7534), .B(n7942), .ZN(n9621) );
  XNOR2_X1 U9248 ( .A(n7536), .B(n7535), .ZN(n7537) );
  OAI222_X1 U9249 ( .A1(n10007), .A2(n8308), .B1(n8307), .B2(n7538), .C1(n7537), .C2(n10013), .ZN(n9623) );
  NAND2_X1 U9250 ( .A1(n9623), .A2(n10016), .ZN(n7542) );
  OAI22_X1 U9251 ( .A1(n10016), .A2(n8044), .B1(n7539), .B2(n10002), .ZN(n7540) );
  AOI21_X1 U9252 ( .B1(n9619), .B2(n9993), .A(n7540), .ZN(n7541) );
  OAI211_X1 U9253 ( .C1(n9621), .C2(n7543), .A(n7542), .B(n7541), .ZN(P2_U3219) );
  INV_X1 U9254 ( .A(n7544), .ZN(n7545) );
  XNOR2_X1 U9255 ( .A(n7547), .B(n7571), .ZN(n7548) );
  XNOR2_X1 U9256 ( .A(n7548), .B(n8325), .ZN(n7670) );
  NAND2_X1 U9257 ( .A1(n7548), .A2(n5299), .ZN(n7549) );
  NAND2_X1 U9258 ( .A1(n7669), .A2(n7549), .ZN(n7678) );
  XNOR2_X1 U9259 ( .A(n8299), .B(n7583), .ZN(n7676) );
  NAND2_X1 U9260 ( .A1(n7676), .A2(n8309), .ZN(n7550) );
  NAND2_X1 U9261 ( .A1(n7678), .A2(n7550), .ZN(n7553) );
  INV_X1 U9262 ( .A(n7676), .ZN(n7551) );
  NAND2_X1 U9263 ( .A1(n7551), .A2(n7977), .ZN(n7552) );
  NAND2_X1 U9264 ( .A1(n7553), .A2(n7552), .ZN(n7714) );
  XNOR2_X1 U9265 ( .A(n8438), .B(n7210), .ZN(n7554) );
  XNOR2_X1 U9266 ( .A(n7554), .B(n7976), .ZN(n7715) );
  INV_X1 U9267 ( .A(n7554), .ZN(n7555) );
  XNOR2_X1 U9268 ( .A(n7644), .B(n7583), .ZN(n7559) );
  XNOR2_X1 U9269 ( .A(n7559), .B(n7975), .ZN(n7645) );
  XNOR2_X1 U9270 ( .A(n7692), .B(n7210), .ZN(n7556) );
  NAND2_X1 U9271 ( .A1(n7556), .A2(n8271), .ZN(n7650) );
  INV_X1 U9272 ( .A(n7556), .ZN(n7557) );
  NAND2_X1 U9273 ( .A1(n7557), .A2(n7974), .ZN(n7558) );
  NAND2_X1 U9274 ( .A1(n7650), .A2(n7558), .ZN(n7694) );
  INV_X1 U9275 ( .A(n7559), .ZN(n7560) );
  AND2_X1 U9276 ( .A1(n7560), .A2(n7975), .ZN(n7693) );
  NOR2_X1 U9277 ( .A1(n7694), .A2(n7693), .ZN(n7561) );
  XNOR2_X1 U9278 ( .A(n7562), .B(n7571), .ZN(n7563) );
  XNOR2_X1 U9279 ( .A(n7563), .B(n8261), .ZN(n7651) );
  INV_X1 U9280 ( .A(n7563), .ZN(n7564) );
  NAND2_X1 U9281 ( .A1(n7564), .A2(n8261), .ZN(n7565) );
  XNOR2_X1 U9282 ( .A(n7703), .B(n7583), .ZN(n7566) );
  XNOR2_X1 U9283 ( .A(n7566), .B(n8247), .ZN(n7704) );
  INV_X1 U9284 ( .A(n7566), .ZN(n7567) );
  NAND2_X1 U9285 ( .A1(n7567), .A2(n7972), .ZN(n7568) );
  INV_X1 U9286 ( .A(n7569), .ZN(n7570) );
  NAND2_X1 U9287 ( .A1(n7572), .A2(n8227), .ZN(n7660) );
  INV_X1 U9288 ( .A(n7572), .ZN(n7573) );
  NAND2_X1 U9289 ( .A1(n7573), .A2(n7970), .ZN(n7574) );
  XNOR2_X1 U9290 ( .A(n7575), .B(n7583), .ZN(n7576) );
  XNOR2_X1 U9291 ( .A(n7576), .B(n8218), .ZN(n7661) );
  XNOR2_X1 U9292 ( .A(n7578), .B(n7210), .ZN(n7580) );
  XNOR2_X1 U9293 ( .A(n7579), .B(n7580), .ZN(n7726) );
  INV_X1 U9294 ( .A(n7580), .ZN(n7581) );
  XNOR2_X1 U9295 ( .A(n8404), .B(n7583), .ZN(n7584) );
  NOR2_X1 U9296 ( .A1(n7585), .A2(n7731), .ZN(n7588) );
  AOI22_X1 U9297 ( .A1(n8179), .A2(n7734), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7586) );
  OAI21_X1 U9298 ( .B1(n8199), .B2(n7730), .A(n7586), .ZN(n7587) );
  AOI211_X1 U9299 ( .C1(n7589), .C2(n7721), .A(n7588), .B(n7587), .ZN(n7590)
         );
  OAI21_X1 U9300 ( .B1(n7591), .B2(n7724), .A(n7590), .ZN(P2_U3160) );
  INV_X1 U9301 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7738) );
  INV_X1 U9302 ( .A(SI_29_), .ZN(n9118) );
  INV_X1 U9303 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8608) );
  MUX2_X1 U9304 ( .A(n7738), .B(n8608), .S(n7747), .Z(n7597) );
  INV_X1 U9305 ( .A(SI_30_), .ZN(n7596) );
  NAND2_X1 U9306 ( .A1(n7597), .A2(n7596), .ZN(n7745) );
  INV_X1 U9307 ( .A(n7597), .ZN(n7598) );
  NAND2_X1 U9308 ( .A1(n7598), .A2(SI_30_), .ZN(n7599) );
  NAND2_X1 U9309 ( .A1(n7745), .A2(n7599), .ZN(n7600) );
  NAND2_X1 U9310 ( .A1(n7601), .A2(n7600), .ZN(n7602) );
  INV_X1 U9311 ( .A(n8607), .ZN(n7636) );
  OAI222_X1 U9312 ( .A1(n8456), .A2(n7738), .B1(n8467), .B2(n7636), .C1(
        P2_U3151), .C2(n7603), .ZN(P2_U3265) );
  OAI222_X1 U9313 ( .A1(n8868), .A2(P1_U3086), .B1(n9562), .B2(n7605), .C1(
        n7604), .C2(n9554), .ZN(P1_U3333) );
  AOI22_X1 U9314 ( .A1(n8191), .A2(n7734), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7606) );
  OAI21_X1 U9315 ( .B1(n8208), .B2(n7730), .A(n7606), .ZN(n7607) );
  AOI21_X1 U9316 ( .B1(n7717), .B2(n7967), .A(n7607), .ZN(n7608) );
  OAI211_X1 U9317 ( .C1(n8404), .C2(n7737), .A(n7609), .B(n7608), .ZN(P2_U3154) );
  INV_X1 U9318 ( .A(n8459), .ZN(n7610) );
  OAI222_X1 U9319 ( .A1(P1_U3086), .A2(n7611), .B1(n9562), .B2(n7610), .C1(
        n7612), .C2(n9554), .ZN(P1_U3327) );
  NAND2_X1 U9320 ( .A1(n8459), .A2(n8730), .ZN(n7614) );
  OR2_X1 U9321 ( .A1(n8729), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U9322 ( .A1(n9212), .A2(n6097), .ZN(n7617) );
  NAND2_X1 U9323 ( .A1(n9200), .A2(n7615), .ZN(n7616) );
  NAND2_X1 U9324 ( .A1(n7617), .A2(n7616), .ZN(n7619) );
  XNOR2_X1 U9325 ( .A(n7619), .B(n7618), .ZN(n7622) );
  AOI22_X1 U9326 ( .A1(n9212), .A2(n4293), .B1(n7620), .B2(n9200), .ZN(n7621)
         );
  XNOR2_X1 U9327 ( .A(n7622), .B(n7621), .ZN(n7623) );
  INV_X1 U9328 ( .A(n7623), .ZN(n7628) );
  NAND3_X1 U9329 ( .A1(n7628), .A2(n9649), .A3(n7627), .ZN(n7633) );
  NAND3_X1 U9330 ( .A1(n7634), .A2(n9649), .A3(n7623), .ZN(n7632) );
  NAND2_X1 U9331 ( .A1(n8724), .A2(n8577), .ZN(n7625) );
  NAND2_X1 U9332 ( .A1(n9169), .A2(n9199), .ZN(n7624) );
  NAND2_X1 U9333 ( .A1(n7625), .A2(n7624), .ZN(n9209) );
  AOI22_X1 U9334 ( .A1(n9209), .A2(n8599), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n7626) );
  OAI21_X1 U9335 ( .B1(n9674), .B2(n9211), .A(n7626), .ZN(n7630) );
  NOR3_X1 U9336 ( .A1(n7628), .A2(n9665), .A3(n7627), .ZN(n7629) );
  AOI211_X1 U9337 ( .C1(n9670), .C2(n9212), .A(n7630), .B(n7629), .ZN(n7631)
         );
  OAI211_X1 U9338 ( .C1(n7634), .C2(n7633), .A(n7632), .B(n7631), .ZN(P1_U3220) );
  OAI222_X1 U9339 ( .A1(n9559), .A2(n8608), .B1(n9551), .B2(n7636), .C1(
        P1_U3086), .C2(n7635), .ZN(P1_U3325) );
  AOI21_X1 U9340 ( .B1(n7971), .B2(n7637), .A(n4314), .ZN(n7643) );
  AOI22_X1 U9341 ( .A1(n7970), .A2(n7717), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7639) );
  NAND2_X1 U9342 ( .A1(n7734), .A2(n8230), .ZN(n7638) );
  OAI211_X1 U9343 ( .C1(n8247), .C2(n7730), .A(n7639), .B(n7638), .ZN(n7640)
         );
  AOI21_X1 U9344 ( .B1(n7641), .B2(n7721), .A(n7640), .ZN(n7642) );
  OAI21_X1 U9345 ( .B1(n7643), .B2(n7724), .A(n7642), .ZN(P2_U3156) );
  INV_X1 U9346 ( .A(n7644), .ZN(n8434) );
  OAI211_X1 U9347 ( .C1(n4356), .C2(n7645), .A(n7697), .B(n7727), .ZN(n7649)
         );
  NAND2_X1 U9348 ( .A1(n7708), .A2(n7976), .ZN(n7646) );
  NAND2_X1 U9349 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8153) );
  OAI211_X1 U9350 ( .C1(n8271), .C2(n7731), .A(n7646), .B(n8153), .ZN(n7647)
         );
  AOI21_X1 U9351 ( .B1(n8276), .B2(n7734), .A(n7647), .ZN(n7648) );
  OAI211_X1 U9352 ( .C1(n8434), .C2(n7737), .A(n7649), .B(n7648), .ZN(P2_U3159) );
  NOR3_X1 U9353 ( .A1(n4328), .A2(n4483), .A3(n7651), .ZN(n7654) );
  INV_X1 U9354 ( .A(n7652), .ZN(n7653) );
  OAI21_X1 U9355 ( .B1(n7654), .B2(n7653), .A(n7727), .ZN(n7658) );
  AOI22_X1 U9356 ( .A1(n7972), .A2(n7717), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7655) );
  OAI21_X1 U9357 ( .B1(n8271), .B2(n7730), .A(n7655), .ZN(n7656) );
  AOI21_X1 U9358 ( .B1(n8252), .B2(n7734), .A(n7656), .ZN(n7657) );
  OAI211_X1 U9359 ( .C1(n8426), .C2(n7737), .A(n7658), .B(n7657), .ZN(P2_U3163) );
  AND3_X1 U9360 ( .A1(n7659), .A2(n7661), .A3(n7660), .ZN(n7662) );
  OAI21_X1 U9361 ( .B1(n7663), .B2(n7662), .A(n7727), .ZN(n7668) );
  INV_X1 U9362 ( .A(n8211), .ZN(n7665) );
  AOI22_X1 U9363 ( .A1(n7970), .A2(n7708), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7664) );
  OAI21_X1 U9364 ( .B1(n7665), .B2(n7719), .A(n7664), .ZN(n7666) );
  AOI21_X1 U9365 ( .B1(n7717), .B2(n7969), .A(n7666), .ZN(n7667) );
  OAI211_X1 U9366 ( .C1(n8412), .C2(n7737), .A(n7668), .B(n7667), .ZN(P2_U3165) );
  OAI211_X1 U9367 ( .C1(n7671), .C2(n7670), .A(n7669), .B(n7727), .ZN(n7675)
         );
  NAND2_X1 U9368 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8075) );
  OAI21_X1 U9369 ( .B1(n7731), .B2(n8309), .A(n8075), .ZN(n7673) );
  NOR2_X1 U9370 ( .A1(n7719), .A2(n8315), .ZN(n7672) );
  AOI211_X1 U9371 ( .C1(n7708), .C2(n7978), .A(n7673), .B(n7672), .ZN(n7674)
         );
  OAI211_X1 U9372 ( .C1(n8446), .C2(n7737), .A(n7675), .B(n7674), .ZN(P2_U3166) );
  XNOR2_X1 U9373 ( .A(n7676), .B(n7977), .ZN(n7677) );
  XNOR2_X1 U9374 ( .A(n7678), .B(n7677), .ZN(n7683) );
  AND2_X1 U9375 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8102) );
  NOR2_X1 U9376 ( .A1(n7730), .A2(n8325), .ZN(n7679) );
  AOI211_X1 U9377 ( .C1(n7717), .C2(n7976), .A(n8102), .B(n7679), .ZN(n7680)
         );
  OAI21_X1 U9378 ( .B1(n8300), .B2(n7719), .A(n7680), .ZN(n7681) );
  AOI21_X1 U9379 ( .B1(n8299), .B2(n7721), .A(n7681), .ZN(n7682) );
  OAI21_X1 U9380 ( .B1(n7683), .B2(n7724), .A(n7682), .ZN(P2_U3168) );
  INV_X1 U9381 ( .A(n7659), .ZN(n7687) );
  NOR3_X1 U9382 ( .A1(n4314), .A2(n7685), .A3(n7684), .ZN(n7686) );
  OAI21_X1 U9383 ( .B1(n7687), .B2(n7686), .A(n7727), .ZN(n7691) );
  AOI22_X1 U9384 ( .A1(n7971), .A2(n7708), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7688) );
  OAI21_X1 U9385 ( .B1(n8218), .B2(n7731), .A(n7688), .ZN(n7689) );
  AOI21_X1 U9386 ( .B1(n8220), .B2(n7734), .A(n7689), .ZN(n7690) );
  OAI211_X1 U9387 ( .C1(n8415), .C2(n7737), .A(n7691), .B(n7690), .ZN(P2_U3169) );
  INV_X1 U9388 ( .A(n7692), .ZN(n8430) );
  INV_X1 U9389 ( .A(n7693), .ZN(n7696) );
  INV_X1 U9390 ( .A(n7694), .ZN(n7695) );
  AOI21_X1 U9391 ( .B1(n7697), .B2(n7696), .A(n7695), .ZN(n7698) );
  OAI21_X1 U9392 ( .B1(n4328), .B2(n7698), .A(n7727), .ZN(n7702) );
  INV_X1 U9393 ( .A(n8261), .ZN(n7973) );
  AOI22_X1 U9394 ( .A1(n7973), .A2(n7717), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7699) );
  OAI21_X1 U9395 ( .B1(n8283), .B2(n7730), .A(n7699), .ZN(n7700) );
  AOI21_X1 U9396 ( .B1(n8264), .B2(n7734), .A(n7700), .ZN(n7701) );
  OAI211_X1 U9397 ( .C1(n8430), .C2(n7737), .A(n7702), .B(n7701), .ZN(P2_U3173) );
  INV_X1 U9398 ( .A(n7703), .ZN(n8422) );
  AOI21_X1 U9399 ( .B1(n7705), .B2(n7704), .A(n7724), .ZN(n7707) );
  NAND2_X1 U9400 ( .A1(n7707), .A2(n7706), .ZN(n7712) );
  AOI22_X1 U9401 ( .A1(n7973), .A2(n7708), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7709) );
  OAI21_X1 U9402 ( .B1(n8237), .B2(n7731), .A(n7709), .ZN(n7710) );
  AOI21_X1 U9403 ( .B1(n8240), .B2(n7734), .A(n7710), .ZN(n7711) );
  OAI211_X1 U9404 ( .C1(n8422), .C2(n7737), .A(n7712), .B(n7711), .ZN(P2_U3175) );
  AOI21_X1 U9405 ( .B1(n7715), .B2(n7714), .A(n7713), .ZN(n7725) );
  AND2_X1 U9406 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8128) );
  NOR2_X1 U9407 ( .A1(n7730), .A2(n8309), .ZN(n7716) );
  AOI211_X1 U9408 ( .C1(n7717), .C2(n7975), .A(n8128), .B(n7716), .ZN(n7718)
         );
  OAI21_X1 U9409 ( .B1(n8288), .B2(n7719), .A(n7718), .ZN(n7720) );
  AOI21_X1 U9410 ( .B1(n7722), .B2(n7721), .A(n7720), .ZN(n7723) );
  OAI21_X1 U9411 ( .B1(n7725), .B2(n7724), .A(n7723), .ZN(P2_U3178) );
  OAI21_X1 U9412 ( .B1(n8208), .B2(n7726), .A(n4449), .ZN(n7728) );
  NAND2_X1 U9413 ( .A1(n7728), .A2(n7727), .ZN(n7736) );
  INV_X1 U9414 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n7729) );
  OAI22_X1 U9415 ( .A1(n8218), .A2(n7730), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7729), .ZN(n7733) );
  NOR2_X1 U9416 ( .A1(n8199), .A2(n7731), .ZN(n7732) );
  AOI211_X1 U9417 ( .C1(n8202), .C2(n7734), .A(n7733), .B(n7732), .ZN(n7735)
         );
  OAI211_X1 U9418 ( .C1(n8408), .C2(n7737), .A(n7736), .B(n7735), .ZN(P2_U3180) );
  NAND2_X1 U9419 ( .A1(n8607), .A2(n7753), .ZN(n7741) );
  OR2_X1 U9420 ( .A1(n7739), .A2(n7738), .ZN(n7740) );
  NAND2_X1 U9421 ( .A1(n7951), .A2(n7742), .ZN(n7906) );
  INV_X1 U9422 ( .A(n7952), .ZN(n7754) );
  MUX2_X1 U9423 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7747), .Z(n7749) );
  INV_X1 U9424 ( .A(SI_31_), .ZN(n7748) );
  XNOR2_X1 U9425 ( .A(n7749), .B(n7748), .ZN(n7750) );
  INV_X1 U9426 ( .A(n7744), .ZN(n8169) );
  INV_X1 U9427 ( .A(n7760), .ZN(n8163) );
  NAND3_X1 U9428 ( .A1(n7755), .A2(n8169), .A3(n8163), .ZN(n7757) );
  AOI21_X1 U9429 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7759) );
  INV_X1 U9430 ( .A(n7759), .ZN(n7956) );
  NOR2_X1 U9431 ( .A1(n8166), .A2(n7760), .ZN(n7910) );
  INV_X1 U9432 ( .A(n7910), .ZN(n7917) );
  MUX2_X1 U9433 ( .A(n8188), .B(n8181), .S(n7903), .Z(n7899) );
  MUX2_X1 U9434 ( .A(n7888), .B(n7889), .S(n7903), .Z(n7896) );
  NAND2_X1 U9435 ( .A1(n7768), .A2(n7761), .ZN(n7764) );
  INV_X1 U9436 ( .A(n7765), .ZN(n7766) );
  OAI21_X1 U9437 ( .B1(n7770), .B2(n7766), .A(n5489), .ZN(n7767) );
  MUX2_X1 U9438 ( .A(n7767), .B(n5489), .S(n7907), .Z(n7773) );
  INV_X1 U9439 ( .A(n7768), .ZN(n7769) );
  NOR2_X1 U9440 ( .A1(n5486), .A2(n7769), .ZN(n7771) );
  AOI21_X1 U9441 ( .B1(n7771), .B2(n7770), .A(n7929), .ZN(n7772) );
  NAND2_X1 U9442 ( .A1(n7773), .A2(n7772), .ZN(n7781) );
  NAND2_X1 U9443 ( .A1(n5092), .A2(n10018), .ZN(n7774) );
  NAND2_X1 U9444 ( .A1(n7782), .A2(n7774), .ZN(n7777) );
  NAND2_X1 U9445 ( .A1(n7790), .A2(n7775), .ZN(n7776) );
  MUX2_X1 U9446 ( .A(n7777), .B(n7776), .S(n7903), .Z(n7778) );
  INV_X1 U9447 ( .A(n7778), .ZN(n7780) );
  AOI21_X1 U9448 ( .B1(n7781), .B2(n7780), .A(n7779), .ZN(n7791) );
  NAND2_X1 U9449 ( .A1(n7791), .A2(n7782), .ZN(n7789) );
  NAND2_X1 U9450 ( .A1(n5490), .A2(n7928), .ZN(n7794) );
  INV_X1 U9451 ( .A(n7784), .ZN(n7785) );
  NOR2_X1 U9452 ( .A1(n7794), .A2(n7785), .ZN(n7788) );
  INV_X1 U9453 ( .A(n7928), .ZN(n7786) );
  NOR2_X1 U9454 ( .A1(n7786), .A2(n7793), .ZN(n7787) );
  AOI21_X1 U9455 ( .B1(n7789), .B2(n7788), .A(n7787), .ZN(n7798) );
  NAND2_X1 U9456 ( .A1(n7791), .A2(n7790), .ZN(n7796) );
  AND2_X1 U9457 ( .A1(n7793), .A2(n7792), .ZN(n7795) );
  AOI22_X1 U9458 ( .A1(n7796), .A2(n7795), .B1(n7927), .B2(n7794), .ZN(n7797)
         );
  MUX2_X1 U9459 ( .A(n7798), .B(n7797), .S(n7907), .Z(n7805) );
  INV_X1 U9460 ( .A(n7799), .ZN(n7800) );
  NOR2_X1 U9461 ( .A1(n7800), .A2(n7806), .ZN(n7801) );
  MUX2_X1 U9462 ( .A(n7802), .B(n7801), .S(n7907), .Z(n7803) );
  OAI21_X1 U9463 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7810) );
  INV_X1 U9464 ( .A(n7806), .ZN(n7807) );
  MUX2_X1 U9465 ( .A(n7808), .B(n7807), .S(n7903), .Z(n7809) );
  NAND3_X1 U9466 ( .A1(n7810), .A2(n7933), .A3(n7809), .ZN(n7815) );
  AND2_X1 U9467 ( .A1(n7816), .A2(n7811), .ZN(n7812) );
  MUX2_X1 U9468 ( .A(n7813), .B(n7812), .S(n7907), .Z(n7814) );
  NAND2_X1 U9469 ( .A1(n7815), .A2(n7814), .ZN(n7821) );
  NAND3_X1 U9470 ( .A1(n7821), .A2(n7816), .A3(n7822), .ZN(n7818) );
  OR2_X1 U9471 ( .A1(n10065), .A2(n7817), .ZN(n7819) );
  NAND2_X1 U9472 ( .A1(n7818), .A2(n7819), .ZN(n7825) );
  NAND3_X1 U9473 ( .A1(n7821), .A2(n7820), .A3(n7819), .ZN(n7823) );
  NAND2_X1 U9474 ( .A1(n7823), .A2(n7822), .ZN(n7824) );
  MUX2_X1 U9475 ( .A(n7825), .B(n7824), .S(n7907), .Z(n7830) );
  NAND2_X1 U9476 ( .A1(n10072), .A2(n7826), .ZN(n7827) );
  MUX2_X1 U9477 ( .A(n7828), .B(n7827), .S(n7903), .Z(n7829) );
  OAI211_X1 U9478 ( .C1(n7830), .C2(n7938), .A(n7923), .B(n7829), .ZN(n7834)
         );
  MUX2_X1 U9479 ( .A(n7832), .B(n7831), .S(n7907), .Z(n7833) );
  NAND3_X1 U9480 ( .A1(n7834), .A2(n7942), .A3(n7833), .ZN(n7838) );
  INV_X1 U9481 ( .A(n8321), .ZN(n8327) );
  MUX2_X1 U9482 ( .A(n7836), .B(n7835), .S(n7903), .Z(n7837) );
  NAND3_X1 U9483 ( .A1(n7838), .A2(n8327), .A3(n7837), .ZN(n7845) );
  NAND2_X1 U9484 ( .A1(n7846), .A2(n7839), .ZN(n7841) );
  INV_X1 U9485 ( .A(n7849), .ZN(n7842) );
  AOI21_X1 U9486 ( .B1(n7845), .B2(n7844), .A(n8297), .ZN(n7850) );
  NAND2_X1 U9487 ( .A1(n7850), .A2(n7846), .ZN(n7851) );
  NAND2_X1 U9488 ( .A1(n7856), .A2(n7847), .ZN(n7848) );
  NAND2_X1 U9489 ( .A1(n7859), .A2(n7853), .ZN(n7852) );
  OAI211_X1 U9490 ( .C1(n7855), .C2(n7852), .A(n7863), .B(n7857), .ZN(n7862)
         );
  NAND3_X1 U9491 ( .A1(n7855), .A2(n7854), .A3(n7853), .ZN(n7858) );
  NAND3_X1 U9492 ( .A1(n7858), .A2(n7857), .A3(n7856), .ZN(n7860) );
  NAND2_X1 U9493 ( .A1(n7860), .A2(n7859), .ZN(n7861) );
  INV_X1 U9494 ( .A(n8248), .ZN(n7867) );
  AND2_X1 U9495 ( .A1(n7869), .A2(n7863), .ZN(n7865) );
  MUX2_X1 U9496 ( .A(n7865), .B(n7864), .S(n7903), .Z(n7866) );
  MUX2_X1 U9497 ( .A(n7869), .B(n7868), .S(n7907), .Z(n7870) );
  NAND3_X1 U9498 ( .A1(n7871), .A2(n7922), .A3(n7870), .ZN(n7877) );
  INV_X1 U9499 ( .A(n7872), .ZN(n7873) );
  NOR2_X1 U9500 ( .A1(n7921), .A2(n7873), .ZN(n7875) );
  MUX2_X1 U9501 ( .A(n7875), .B(n7874), .S(n7903), .Z(n7876) );
  INV_X1 U9502 ( .A(n7878), .ZN(n7920) );
  OAI21_X1 U9503 ( .B1(n7879), .B2(n7920), .A(n7880), .ZN(n7882) );
  OAI21_X1 U9504 ( .B1(n4296), .B2(n7921), .A(n5496), .ZN(n7881) );
  MUX2_X1 U9505 ( .A(n7882), .B(n7881), .S(n7903), .Z(n7883) );
  INV_X1 U9506 ( .A(n7884), .ZN(n7890) );
  MUX2_X1 U9507 ( .A(n7886), .B(n7885), .S(n7903), .Z(n7887) );
  NAND2_X1 U9508 ( .A1(n8200), .A2(n7887), .ZN(n7893) );
  MUX2_X1 U9509 ( .A(n7891), .B(n7890), .S(n7903), .Z(n7892) );
  OAI211_X1 U9510 ( .C1(n7894), .C2(n7893), .A(n7919), .B(n7892), .ZN(n7895)
         );
  NAND2_X1 U9511 ( .A1(n7952), .A2(n7898), .ZN(n7901) );
  AOI211_X1 U9512 ( .C1(n8181), .C2(n7909), .A(n7901), .B(n7908), .ZN(n7915)
         );
  INV_X1 U9513 ( .A(n7902), .ZN(n7966) );
  AOI21_X1 U9514 ( .B1(n7907), .B2(n7966), .A(n8169), .ZN(n7905) );
  NOR3_X1 U9515 ( .A1(n7908), .A2(n7907), .A3(n7906), .ZN(n7912) );
  NAND2_X1 U9516 ( .A1(n7909), .A2(n8188), .ZN(n7911) );
  INV_X1 U9517 ( .A(n7922), .ZN(n8239) );
  INV_X1 U9518 ( .A(n7923), .ZN(n7940) );
  NAND4_X1 U9519 ( .A1(n5487), .A2(n7926), .A3(n7925), .A4(n7924), .ZN(n7931)
         );
  NAND2_X1 U9520 ( .A1(n7928), .A2(n7927), .ZN(n9990) );
  NOR4_X1 U9521 ( .A1(n7931), .A2(n7930), .A3(n9990), .A4(n7929), .ZN(n7934)
         );
  NAND4_X1 U9522 ( .A1(n7934), .A2(n5491), .A3(n7933), .A4(n7932), .ZN(n7937)
         );
  OR3_X1 U9523 ( .A1(n7937), .A2(n7936), .A3(n7935), .ZN(n7939) );
  NOR3_X1 U9524 ( .A1(n7940), .A2(n7939), .A3(n7938), .ZN(n7941) );
  NAND4_X1 U9525 ( .A1(n8314), .A2(n8327), .A3(n7942), .A4(n7941), .ZN(n7943)
         );
  NOR2_X1 U9526 ( .A1(n7943), .A2(n8297), .ZN(n7944) );
  NAND3_X1 U9527 ( .A1(n8274), .A2(n4763), .A3(n7944), .ZN(n7945) );
  OR3_X1 U9528 ( .A1(n8251), .A2(n8263), .A3(n7945), .ZN(n7946) );
  NOR3_X1 U9529 ( .A1(n8228), .A2(n8239), .A3(n7946), .ZN(n7947) );
  NAND2_X1 U9530 ( .A1(n8221), .A2(n7947), .ZN(n7948) );
  OR4_X1 U9531 ( .A1(n8196), .A2(n8190), .A3(n7948), .A4(n8209), .ZN(n7949) );
  NAND4_X1 U9532 ( .A1(n4342), .A2(n7954), .A3(n7953), .A4(n7952), .ZN(n7955)
         );
  NAND3_X1 U9533 ( .A1(n7960), .A2(n7959), .A3(n9882), .ZN(n7961) );
  OAI211_X1 U9534 ( .C1(n7962), .C2(n7964), .A(n7961), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7963) );
  OAI21_X1 U9535 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(P2_U3296) );
  MUX2_X1 U9536 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n7966), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9537 ( .A(n7967), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8122), .Z(
        P2_U3519) );
  MUX2_X1 U9538 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n7968), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9539 ( .A(n7969), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8122), .Z(
        P2_U3517) );
  MUX2_X1 U9540 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n7970), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9541 ( .A(n7971), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8122), .Z(
        P2_U3514) );
  MUX2_X1 U9542 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n7972), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9543 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n7973), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9544 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n7974), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9545 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n7975), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9546 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n7976), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9547 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n7977), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9548 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n5299), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9549 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n7978), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9550 ( .A(n7979), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8122), .Z(
        P2_U3505) );
  MUX2_X1 U9551 ( .A(n7980), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8122), .Z(
        P2_U3504) );
  MUX2_X1 U9552 ( .A(n7981), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8122), .Z(
        P2_U3503) );
  MUX2_X1 U9553 ( .A(n7982), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8122), .Z(
        P2_U3502) );
  MUX2_X1 U9554 ( .A(n7983), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8122), .Z(
        P2_U3501) );
  MUX2_X1 U9555 ( .A(n7984), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8122), .Z(
        P2_U3500) );
  MUX2_X1 U9556 ( .A(n7985), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8122), .Z(
        P2_U3499) );
  MUX2_X1 U9557 ( .A(n9985), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8122), .Z(
        P2_U3498) );
  MUX2_X1 U9558 ( .A(n7986), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8122), .Z(
        P2_U3497) );
  MUX2_X1 U9559 ( .A(n9983), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8122), .Z(
        P2_U3496) );
  MUX2_X1 U9560 ( .A(n7987), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8122), .Z(
        P2_U3495) );
  MUX2_X1 U9561 ( .A(n7988), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8122), .Z(
        P2_U3494) );
  MUX2_X1 U9562 ( .A(n5092), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8122), .Z(
        P2_U3493) );
  MUX2_X1 U9563 ( .A(n6492), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8122), .Z(
        P2_U3492) );
  MUX2_X1 U9564 ( .A(n7989), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8122), .Z(
        P2_U3491) );
  AOI21_X1 U9565 ( .B1(n7991), .B2(n7094), .A(n7990), .ZN(n7992) );
  OR2_X1 U9566 ( .A1(n7992), .A2(n9965), .ZN(n8007) );
  AOI21_X1 U9567 ( .B1(n7995), .B2(n7994), .A(n7993), .ZN(n7999) );
  NAND2_X1 U9568 ( .A1(n9914), .A2(n7996), .ZN(n7998) );
  OAI211_X1 U9569 ( .C1(n7999), .C2(n9917), .A(n7998), .B(n7997), .ZN(n8000)
         );
  INV_X1 U9570 ( .A(n8000), .ZN(n8006) );
  INV_X1 U9571 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9585) );
  OR2_X1 U9572 ( .A1(n9924), .A2(n9585), .ZN(n8005) );
  AND2_X1 U9573 ( .A1(n8001), .A2(n10085), .ZN(n8002) );
  OAI21_X1 U9574 ( .B1(n8003), .B2(n8002), .A(n9951), .ZN(n8004) );
  NAND4_X1 U9575 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(
        P2_U3191) );
  AOI21_X1 U9576 ( .B1(n8010), .B2(n8009), .A(n8008), .ZN(n8012) );
  MUX2_X1 U9577 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9882), .Z(n8049) );
  XNOR2_X1 U9578 ( .A(n8049), .B(n8019), .ZN(n8011) );
  NAND2_X1 U9579 ( .A1(n8012), .A2(n8011), .ZN(n8051) );
  OAI21_X1 U9580 ( .B1(n8012), .B2(n8011), .A(n8051), .ZN(n8032) );
  INV_X1 U9581 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8022) );
  AND2_X1 U9582 ( .A1(n8015), .A2(n5250), .ZN(n8016) );
  OAI21_X1 U9583 ( .B1(n4401), .B2(n8016), .A(n9951), .ZN(n8021) );
  INV_X1 U9584 ( .A(n8017), .ZN(n8018) );
  AOI21_X1 U9585 ( .B1(n9914), .B2(n8019), .A(n8018), .ZN(n8020) );
  OAI211_X1 U9586 ( .C1(n8022), .C2(n9924), .A(n8021), .B(n8020), .ZN(n8031)
         );
  AND2_X1 U9587 ( .A1(n8023), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8024) );
  AOI21_X1 U9588 ( .B1(n8028), .B2(n8027), .A(n8035), .ZN(n8029) );
  NOR2_X1 U9589 ( .A1(n8029), .A2(n9965), .ZN(n8030) );
  AOI211_X1 U9590 ( .C1(n8032), .C2(n9970), .A(n8031), .B(n8030), .ZN(n8033)
         );
  INV_X1 U9591 ( .A(n8033), .ZN(P2_U3195) );
  INV_X1 U9592 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8039) );
  INV_X1 U9593 ( .A(n8034), .ZN(n8036) );
  NAND2_X1 U9594 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n9979), .ZN(n8037) );
  OAI21_X1 U9595 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n9979), .A(n8037), .ZN(
        n9963) );
  AOI21_X1 U9596 ( .B1(n8039), .B2(n8038), .A(n8064), .ZN(n8062) );
  NAND2_X1 U9597 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n9979), .ZN(n8040) );
  OAI21_X1 U9598 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9979), .A(n8040), .ZN(
        n9961) );
  NOR2_X1 U9599 ( .A1(n4346), .A2(n9961), .ZN(n9960) );
  AOI21_X1 U9600 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n9979), .A(n9960), .ZN(
        n8077) );
  INV_X1 U9601 ( .A(n8042), .ZN(n8041) );
  NOR2_X1 U9602 ( .A1(n8041), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8043) );
  OAI21_X1 U9603 ( .B1(n8043), .B2(n8079), .A(n9951), .ZN(n8061) );
  MUX2_X1 U9604 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9882), .Z(n8068) );
  XNOR2_X1 U9605 ( .A(n8068), .B(n8078), .ZN(n8055) );
  OR2_X1 U9606 ( .A1(n9882), .A2(n8044), .ZN(n8046) );
  NAND2_X1 U9607 ( .A1(n9882), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8045) );
  NAND2_X1 U9608 ( .A1(n8046), .A2(n8045), .ZN(n8048) );
  OR2_X1 U9609 ( .A1(n9979), .A2(n8048), .ZN(n8053) );
  XNOR2_X1 U9610 ( .A(n8048), .B(n8047), .ZN(n9969) );
  OR2_X1 U9611 ( .A1(n8050), .A2(n8049), .ZN(n8052) );
  NAND2_X1 U9612 ( .A1(n8052), .A2(n8051), .ZN(n9968) );
  NAND2_X1 U9613 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  NAND2_X1 U9614 ( .A1(n8053), .A2(n9967), .ZN(n8054) );
  NAND2_X1 U9615 ( .A1(n8055), .A2(n8054), .ZN(n8070) );
  OAI21_X1 U9616 ( .B1(n8055), .B2(n8054), .A(n8070), .ZN(n8059) );
  INV_X1 U9617 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9603) );
  NOR2_X1 U9618 ( .A1(n9924), .A2(n9603), .ZN(n8058) );
  OAI21_X1 U9619 ( .B1(n9980), .B2(n8069), .A(n8056), .ZN(n8057) );
  AOI211_X1 U9620 ( .C1(n9970), .C2(n8059), .A(n8058), .B(n8057), .ZN(n8060)
         );
  OAI211_X1 U9621 ( .C1(n8062), .C2(n9965), .A(n8061), .B(n8060), .ZN(P2_U3197) );
  NAND2_X1 U9622 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8090), .ZN(n8065) );
  OAI21_X1 U9623 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8090), .A(n8065), .ZN(
        n8066) );
  AOI21_X1 U9624 ( .B1(n8067), .B2(n8066), .A(n8087), .ZN(n8086) );
  MUX2_X1 U9625 ( .A(n8316), .B(n8388), .S(n9882), .Z(n8095) );
  XNOR2_X1 U9626 ( .A(n8095), .B(n8090), .ZN(n8073) );
  OR2_X1 U9627 ( .A1(n8069), .A2(n8068), .ZN(n8071) );
  NAND2_X1 U9628 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  NAND2_X1 U9629 ( .A1(n8073), .A2(n8072), .ZN(n8097) );
  OAI21_X1 U9630 ( .B1(n8073), .B2(n8072), .A(n8097), .ZN(n8074) );
  NAND2_X1 U9631 ( .A1(n8074), .A2(n9970), .ZN(n8076) );
  OAI211_X1 U9632 ( .C1(n9980), .C2(n8090), .A(n8076), .B(n8075), .ZN(n8084)
         );
  NOR2_X1 U9633 ( .A1(n8078), .A2(n8077), .ZN(n8080) );
  XNOR2_X1 U9634 ( .A(n8090), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8081) );
  AOI21_X1 U9635 ( .B1(n4358), .B2(n8081), .A(n8089), .ZN(n8082) );
  NOR2_X1 U9636 ( .A1(n8082), .A2(n9974), .ZN(n8083) );
  AOI211_X1 U9637 ( .C1(n9959), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8084), .B(
        n8083), .ZN(n8085) );
  OAI21_X1 U9638 ( .B1(n8086), .B2(n9965), .A(n8085), .ZN(P2_U3198) );
  AOI21_X1 U9639 ( .B1(n8301), .B2(n8088), .A(n8109), .ZN(n8107) );
  INV_X1 U9640 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9611) );
  AOI21_X1 U9641 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n8090), .A(n8089), .ZN(
        n8129) );
  NAND2_X1 U9642 ( .A1(n8091), .A2(n8383), .ZN(n8092) );
  OR2_X1 U9643 ( .A1(n9882), .A2(n8301), .ZN(n8094) );
  NAND2_X1 U9644 ( .A1(n9882), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U9645 ( .A1(n8094), .A2(n8093), .ZN(n8117) );
  XNOR2_X1 U9646 ( .A(n8117), .B(n8130), .ZN(n8100) );
  NAND2_X1 U9647 ( .A1(n8096), .A2(n8095), .ZN(n8098) );
  NAND2_X1 U9648 ( .A1(n8098), .A2(n8097), .ZN(n8099) );
  NAND2_X1 U9649 ( .A1(n8100), .A2(n8099), .ZN(n8115) );
  OAI21_X1 U9650 ( .B1(n8100), .B2(n8099), .A(n8115), .ZN(n8101) );
  AOI21_X1 U9651 ( .B1(n9914), .B2(n8130), .A(n8102), .ZN(n8103) );
  OAI211_X1 U9652 ( .C1(n9611), .C2(n9924), .A(n8104), .B(n8103), .ZN(n8105)
         );
  INV_X1 U9653 ( .A(n8105), .ZN(n8106) );
  OAI21_X1 U9654 ( .B1(n8107), .B2(n9965), .A(n8106), .ZN(P2_U3199) );
  NOR2_X1 U9655 ( .A1(n8130), .A2(n8108), .ZN(n8110) );
  NAND2_X1 U9656 ( .A1(n8150), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8137) );
  OAI21_X1 U9657 ( .B1(n8150), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8137), .ZN(
        n8112) );
  INV_X1 U9658 ( .A(n8138), .ZN(n8111) );
  AOI21_X1 U9659 ( .B1(n8113), .B2(n8112), .A(n8111), .ZN(n8136) );
  INV_X1 U9660 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8289) );
  NOR2_X1 U9661 ( .A1(n9882), .A2(n8289), .ZN(n8114) );
  AOI21_X1 U9662 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n9882), .A(n8114), .ZN(
        n8119) );
  OAI21_X1 U9663 ( .B1(n8117), .B2(n8116), .A(n8115), .ZN(n8118) );
  NOR2_X1 U9664 ( .A1(n8119), .A2(n8118), .ZN(n8148) );
  INV_X1 U9665 ( .A(n8148), .ZN(n8120) );
  NAND2_X1 U9666 ( .A1(n8119), .A2(n8118), .ZN(n8149) );
  NAND2_X1 U9667 ( .A1(n8120), .A2(n8149), .ZN(n8123) );
  INV_X1 U9668 ( .A(n8123), .ZN(n8121) );
  NOR2_X1 U9669 ( .A1(n8121), .A2(n9917), .ZN(n8126) );
  OAI21_X1 U9670 ( .B1(n8123), .B2(n8122), .A(n9980), .ZN(n8125) );
  MUX2_X1 U9671 ( .A(n8126), .B(n8125), .S(n8124), .Z(n8127) );
  NOR2_X1 U9672 ( .A1(n8130), .A2(n8129), .ZN(n8131) );
  NAND2_X1 U9673 ( .A1(n8150), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8140) );
  OAI21_X1 U9674 ( .B1(n8150), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8140), .ZN(
        n8132) );
  AND2_X1 U9675 ( .A1(n4379), .A2(n8132), .ZN(n8133) );
  OAI21_X1 U9676 ( .B1(n8142), .B2(n8133), .A(n9951), .ZN(n8134) );
  OAI211_X1 U9677 ( .C1(n8136), .C2(n9965), .A(n8135), .B(n8134), .ZN(P2_U3200) );
  MUX2_X1 U9678 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n4940), .S(n8154), .Z(n8146)
         );
  INV_X1 U9679 ( .A(n8146), .ZN(n8139) );
  INV_X1 U9680 ( .A(n8140), .ZN(n8141) );
  NOR2_X1 U9681 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  XNOR2_X1 U9682 ( .A(n8154), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8144) );
  XNOR2_X1 U9683 ( .A(n8143), .B(n8144), .ZN(n8159) );
  INV_X1 U9684 ( .A(n8144), .ZN(n8147) );
  MUX2_X1 U9685 ( .A(n8147), .B(n8146), .S(n8145), .Z(n8152) );
  AOI21_X1 U9686 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8151) );
  XOR2_X1 U9687 ( .A(n8152), .B(n8151), .Z(n8157) );
  OAI21_X1 U9688 ( .B1(n9980), .B2(n8154), .A(n8153), .ZN(n8155) );
  AOI21_X1 U9689 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n9959), .A(n8155), .ZN(
        n8156) );
  OAI21_X1 U9690 ( .B1(n8157), .B2(n9917), .A(n8156), .ZN(n8158) );
  AOI21_X1 U9691 ( .B1(n8159), .B2(n9951), .A(n8158), .ZN(n8160) );
  OAI21_X1 U9692 ( .B1(n8161), .B2(n9965), .A(n8160), .ZN(P2_U3201) );
  NOR2_X1 U9693 ( .A1(n8163), .A2(n8162), .ZN(n8396) );
  NOR2_X1 U9694 ( .A1(n8164), .A2(n10002), .ZN(n8173) );
  AOI21_X1 U9695 ( .B1(n8396), .B2(n10016), .A(n8173), .ZN(n8168) );
  NAND2_X1 U9696 ( .A1(n8334), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8165) );
  OAI211_X1 U9697 ( .C1(n8166), .C2(n8329), .A(n8168), .B(n8165), .ZN(P2_U3202) );
  NAND2_X1 U9698 ( .A1(n8334), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8167) );
  OAI211_X1 U9699 ( .C1(n8169), .C2(n8329), .A(n8168), .B(n8167), .ZN(P2_U3203) );
  NAND2_X1 U9700 ( .A1(n8170), .A2(n10016), .ZN(n8175) );
  NOR2_X1 U9701 ( .A1(n8171), .A2(n8329), .ZN(n8172) );
  AOI211_X1 U9702 ( .C1(n8334), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8173), .B(
        n8172), .ZN(n8174) );
  OAI211_X1 U9703 ( .C1(n8177), .C2(n8176), .A(n8175), .B(n8174), .ZN(P2_U3204) );
  INV_X1 U9704 ( .A(n8178), .ZN(n8183) );
  AOI22_X1 U9705 ( .A1(n8179), .A2(n9994), .B1(n8334), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8180) );
  OAI21_X1 U9706 ( .B1(n8181), .B2(n8329), .A(n8180), .ZN(n8182) );
  AOI21_X1 U9707 ( .B1(n8183), .B2(n9996), .A(n8182), .ZN(n8184) );
  OAI21_X1 U9708 ( .B1(n8185), .B2(n8334), .A(n8184), .ZN(P2_U3205) );
  XNOR2_X1 U9709 ( .A(n8186), .B(n8190), .ZN(n8187) );
  OAI222_X1 U9710 ( .A1(n8307), .A2(n8208), .B1(n10007), .B2(n8188), .C1(n8187), .C2(n10013), .ZN(n8342) );
  INV_X1 U9711 ( .A(n8342), .ZN(n8195) );
  XNOR2_X1 U9712 ( .A(n8189), .B(n8190), .ZN(n8343) );
  AOI22_X1 U9713 ( .A1(n8191), .A2(n9994), .B1(n8334), .B2(
        P2_REG2_REG_27__SCAN_IN), .ZN(n8192) );
  OAI21_X1 U9714 ( .B1(n8404), .B2(n8329), .A(n8192), .ZN(n8193) );
  AOI21_X1 U9715 ( .B1(n8343), .B2(n9996), .A(n8193), .ZN(n8194) );
  OAI21_X1 U9716 ( .B1(n8195), .B2(n8334), .A(n8194), .ZN(P2_U3206) );
  XNOR2_X1 U9717 ( .A(n8197), .B(n8196), .ZN(n8198) );
  OAI222_X1 U9718 ( .A1(n10007), .A2(n8199), .B1(n8307), .B2(n8218), .C1(
        n10013), .C2(n8198), .ZN(n8346) );
  INV_X1 U9719 ( .A(n8346), .ZN(n8206) );
  XNOR2_X1 U9720 ( .A(n8201), .B(n8200), .ZN(n8347) );
  AOI22_X1 U9721 ( .A1(n8202), .A2(n9994), .B1(n8334), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8203) );
  OAI21_X1 U9722 ( .B1(n8408), .B2(n8329), .A(n8203), .ZN(n8204) );
  AOI21_X1 U9723 ( .B1(n8347), .B2(n9996), .A(n8204), .ZN(n8205) );
  OAI21_X1 U9724 ( .B1(n8206), .B2(n8334), .A(n8205), .ZN(P2_U3207) );
  OAI222_X1 U9725 ( .A1(n10007), .A2(n8208), .B1(n8307), .B2(n8227), .C1(
        n10013), .C2(n8207), .ZN(n8350) );
  INV_X1 U9726 ( .A(n8350), .ZN(n8215) );
  XNOR2_X1 U9727 ( .A(n8210), .B(n8209), .ZN(n8351) );
  AOI22_X1 U9728 ( .A1(n8211), .A2(n9994), .B1(n8334), .B2(
        P2_REG2_REG_25__SCAN_IN), .ZN(n8212) );
  OAI21_X1 U9729 ( .B1(n8412), .B2(n8329), .A(n8212), .ZN(n8213) );
  AOI21_X1 U9730 ( .B1(n8351), .B2(n9996), .A(n8213), .ZN(n8214) );
  OAI21_X1 U9731 ( .B1(n8215), .B2(n8334), .A(n8214), .ZN(P2_U3208) );
  NOR2_X1 U9732 ( .A1(n8415), .A2(n10003), .ZN(n8219) );
  XOR2_X1 U9733 ( .A(n8221), .B(n8216), .Z(n8217) );
  OAI222_X1 U9734 ( .A1(n8307), .A2(n8237), .B1(n10007), .B2(n8218), .C1(n8217), .C2(n10013), .ZN(n8354) );
  AOI211_X1 U9735 ( .C1(n9994), .C2(n8220), .A(n8219), .B(n8354), .ZN(n8224)
         );
  XNOR2_X1 U9736 ( .A(n8222), .B(n8221), .ZN(n8355) );
  AOI22_X1 U9737 ( .A1(n8355), .A2(n9996), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8334), .ZN(n8223) );
  OAI21_X1 U9738 ( .B1(n8224), .B2(n8334), .A(n8223), .ZN(P2_U3209) );
  XOR2_X1 U9739 ( .A(n8228), .B(n8225), .Z(n8226) );
  OAI222_X1 U9740 ( .A1(n10007), .A2(n8227), .B1(n8307), .B2(n8247), .C1(
        n10013), .C2(n8226), .ZN(n8358) );
  INV_X1 U9741 ( .A(n8358), .ZN(n8234) );
  XNOR2_X1 U9742 ( .A(n8229), .B(n8228), .ZN(n8359) );
  AOI22_X1 U9743 ( .A1(n8334), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8230), .B2(
        n9994), .ZN(n8231) );
  OAI21_X1 U9744 ( .B1(n8418), .B2(n8329), .A(n8231), .ZN(n8232) );
  AOI21_X1 U9745 ( .B1(n8359), .B2(n9996), .A(n8232), .ZN(n8233) );
  OAI21_X1 U9746 ( .B1(n8234), .B2(n8334), .A(n8233), .ZN(P2_U3210) );
  XNOR2_X1 U9747 ( .A(n8235), .B(n8239), .ZN(n8236) );
  OAI222_X1 U9748 ( .A1(n8307), .A2(n8261), .B1(n10007), .B2(n8237), .C1(
        n10013), .C2(n8236), .ZN(n8361) );
  INV_X1 U9749 ( .A(n8361), .ZN(n8244) );
  XNOR2_X1 U9750 ( .A(n8238), .B(n8239), .ZN(n8362) );
  AOI22_X1 U9751 ( .A1(n8334), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9994), .B2(
        n8240), .ZN(n8241) );
  OAI21_X1 U9752 ( .B1(n8422), .B2(n8329), .A(n8241), .ZN(n8242) );
  AOI21_X1 U9753 ( .B1(n8362), .B2(n9996), .A(n8242), .ZN(n8243) );
  OAI21_X1 U9754 ( .B1(n8244), .B2(n8334), .A(n8243), .ZN(P2_U3211) );
  XOR2_X1 U9755 ( .A(n8245), .B(n8251), .Z(n8246) );
  OAI222_X1 U9756 ( .A1(n10007), .A2(n8247), .B1(n8307), .B2(n8271), .C1(
        n10013), .C2(n8246), .ZN(n8365) );
  INV_X1 U9757 ( .A(n8365), .ZN(n8256) );
  NAND2_X1 U9758 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  XOR2_X1 U9759 ( .A(n8251), .B(n8250), .Z(n8366) );
  AOI22_X1 U9760 ( .A1(n8334), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9994), .B2(
        n8252), .ZN(n8253) );
  OAI21_X1 U9761 ( .B1(n8426), .B2(n8329), .A(n8253), .ZN(n8254) );
  AOI21_X1 U9762 ( .B1(n8366), .B2(n9996), .A(n8254), .ZN(n8255) );
  OAI21_X1 U9763 ( .B1(n8256), .B2(n8334), .A(n8255), .ZN(P2_U3212) );
  OAI21_X1 U9764 ( .B1(n8258), .B2(n8263), .A(n8257), .ZN(n8259) );
  INV_X1 U9765 ( .A(n8259), .ZN(n8260) );
  OAI222_X1 U9766 ( .A1(n10007), .A2(n8261), .B1(n8307), .B2(n8283), .C1(
        n10013), .C2(n8260), .ZN(n8369) );
  INV_X1 U9767 ( .A(n8369), .ZN(n8268) );
  XOR2_X1 U9768 ( .A(n8262), .B(n8263), .Z(n8370) );
  AOI22_X1 U9769 ( .A1(n8334), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9994), .B2(
        n8264), .ZN(n8265) );
  OAI21_X1 U9770 ( .B1(n8430), .B2(n8329), .A(n8265), .ZN(n8266) );
  AOI21_X1 U9771 ( .B1(n8370), .B2(n9996), .A(n8266), .ZN(n8267) );
  OAI21_X1 U9772 ( .B1(n8268), .B2(n8334), .A(n8267), .ZN(P2_U3213) );
  AOI211_X1 U9773 ( .C1(n8274), .C2(n8269), .A(n10013), .B(n8270), .ZN(n8273)
         );
  OAI22_X1 U9774 ( .A1(n8271), .A2(n10007), .B1(n8296), .B2(n8307), .ZN(n8272)
         );
  OR2_X1 U9775 ( .A1(n8273), .A2(n8272), .ZN(n8373) );
  INV_X1 U9776 ( .A(n8373), .ZN(n8280) );
  XOR2_X1 U9777 ( .A(n8275), .B(n8274), .Z(n8374) );
  AOI22_X1 U9778 ( .A1(n8334), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n9994), .B2(
        n8276), .ZN(n8277) );
  OAI21_X1 U9779 ( .B1(n8434), .B2(n8329), .A(n8277), .ZN(n8278) );
  AOI21_X1 U9780 ( .B1(n8374), .B2(n9996), .A(n8278), .ZN(n8279) );
  OAI21_X1 U9781 ( .B1(n8280), .B2(n8334), .A(n8279), .ZN(P2_U3214) );
  XNOR2_X1 U9782 ( .A(n8281), .B(n4763), .ZN(n8282) );
  OAI222_X1 U9783 ( .A1(n10007), .A2(n8283), .B1(n8307), .B2(n8309), .C1(n8282), .C2(n10013), .ZN(n8377) );
  INV_X1 U9784 ( .A(n8377), .ZN(n8293) );
  INV_X1 U9785 ( .A(n8284), .ZN(n8285) );
  AOI21_X1 U9786 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8378) );
  NOR2_X1 U9787 ( .A1(n8438), .A2(n8329), .ZN(n8291) );
  OAI22_X1 U9788 ( .A1(n10016), .A2(n8289), .B1(n8288), .B2(n10002), .ZN(n8290) );
  AOI211_X1 U9789 ( .C1(n8378), .C2(n9996), .A(n8291), .B(n8290), .ZN(n8292)
         );
  OAI21_X1 U9790 ( .B1(n8293), .B2(n8334), .A(n8292), .ZN(P2_U3215) );
  XNOR2_X1 U9791 ( .A(n8294), .B(n8297), .ZN(n8295) );
  OAI222_X1 U9792 ( .A1(n10007), .A2(n8296), .B1(n8307), .B2(n8325), .C1(n8295), .C2(n10013), .ZN(n8381) );
  INV_X1 U9793 ( .A(n8381), .ZN(n8305) );
  XNOR2_X1 U9794 ( .A(n8298), .B(n8297), .ZN(n8382) );
  INV_X1 U9795 ( .A(n8299), .ZN(n8442) );
  NOR2_X1 U9796 ( .A1(n8442), .A2(n8329), .ZN(n8303) );
  OAI22_X1 U9797 ( .A1(n10016), .A2(n8301), .B1(n8300), .B2(n10002), .ZN(n8302) );
  AOI211_X1 U9798 ( .C1(n8382), .C2(n9996), .A(n8303), .B(n8302), .ZN(n8304)
         );
  OAI21_X1 U9799 ( .B1(n8305), .B2(n8334), .A(n8304), .ZN(P2_U3216) );
  AOI21_X1 U9800 ( .B1(n8306), .B2(n8314), .A(n10013), .ZN(n8312) );
  OAI22_X1 U9801 ( .A1(n8309), .A2(n10007), .B1(n8308), .B2(n8307), .ZN(n8310)
         );
  AOI21_X1 U9802 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(n8387) );
  XNOR2_X1 U9803 ( .A(n8313), .B(n5298), .ZN(n8385) );
  NOR2_X1 U9804 ( .A1(n8446), .A2(n8329), .ZN(n8318) );
  OAI22_X1 U9805 ( .A1(n10016), .A2(n8316), .B1(n8315), .B2(n10002), .ZN(n8317) );
  AOI211_X1 U9806 ( .C1(n8385), .C2(n9996), .A(n8318), .B(n8317), .ZN(n8319)
         );
  OAI21_X1 U9807 ( .B1(n8387), .B2(n8334), .A(n8319), .ZN(P2_U3217) );
  OAI21_X1 U9808 ( .B1(n8322), .B2(n8321), .A(n8320), .ZN(n8323) );
  INV_X1 U9809 ( .A(n8323), .ZN(n8324) );
  OAI222_X1 U9810 ( .A1(n8307), .A2(n8326), .B1(n10007), .B2(n8325), .C1(
        n10013), .C2(n8324), .ZN(n8390) );
  INV_X1 U9811 ( .A(n8390), .ZN(n8335) );
  XNOR2_X1 U9812 ( .A(n8328), .B(n8327), .ZN(n8391) );
  NOR2_X1 U9813 ( .A1(n8451), .A2(n8329), .ZN(n8332) );
  OAI22_X1 U9814 ( .A1(n10016), .A2(n8039), .B1(n8330), .B2(n10002), .ZN(n8331) );
  AOI211_X1 U9815 ( .C1(n8391), .C2(n9996), .A(n8332), .B(n8331), .ZN(n8333)
         );
  OAI21_X1 U9816 ( .B1(n8335), .B2(n8334), .A(n8333), .ZN(P2_U3218) );
  INV_X1 U9817 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U9818 ( .A1(n8395), .A2(n8338), .ZN(n8336) );
  NAND2_X1 U9819 ( .A1(n8396), .A2(n10092), .ZN(n8339) );
  OAI211_X1 U9820 ( .C1(n10092), .C2(n8337), .A(n8336), .B(n8339), .ZN(
        P2_U3490) );
  INV_X1 U9821 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8341) );
  NAND2_X1 U9822 ( .A1(n7744), .A2(n8338), .ZN(n8340) );
  OAI211_X1 U9823 ( .C1(n10092), .C2(n8341), .A(n8340), .B(n8339), .ZN(
        P2_U3489) );
  INV_X1 U9824 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8344) );
  AOI21_X1 U9825 ( .B1(n10068), .B2(n8343), .A(n8342), .ZN(n8401) );
  MUX2_X1 U9826 ( .A(n8344), .B(n8401), .S(n10092), .Z(n8345) );
  OAI21_X1 U9827 ( .B1(n8404), .B2(n8394), .A(n8345), .ZN(P2_U3486) );
  INV_X1 U9828 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8348) );
  AOI21_X1 U9829 ( .B1(n8347), .B2(n10068), .A(n8346), .ZN(n8405) );
  MUX2_X1 U9830 ( .A(n8348), .B(n8405), .S(n10092), .Z(n8349) );
  OAI21_X1 U9831 ( .B1(n8408), .B2(n8394), .A(n8349), .ZN(P2_U3485) );
  INV_X1 U9832 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8352) );
  AOI21_X1 U9833 ( .B1(n10068), .B2(n8351), .A(n8350), .ZN(n8409) );
  MUX2_X1 U9834 ( .A(n8352), .B(n8409), .S(n10092), .Z(n8353) );
  INV_X1 U9835 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8356) );
  AOI21_X1 U9836 ( .B1(n8355), .B2(n10068), .A(n8354), .ZN(n8413) );
  MUX2_X1 U9837 ( .A(n8356), .B(n8413), .S(n10092), .Z(n8357) );
  OAI21_X1 U9838 ( .B1(n8415), .B2(n8394), .A(n8357), .ZN(P2_U3483) );
  AOI21_X1 U9839 ( .B1(n10068), .B2(n8359), .A(n8358), .ZN(n8416) );
  MUX2_X1 U9840 ( .A(n9095), .B(n8416), .S(n10092), .Z(n8360) );
  OAI21_X1 U9841 ( .B1(n8418), .B2(n8394), .A(n8360), .ZN(P2_U3482) );
  INV_X1 U9842 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8363) );
  AOI21_X1 U9843 ( .B1(n10068), .B2(n8362), .A(n8361), .ZN(n8419) );
  MUX2_X1 U9844 ( .A(n8363), .B(n8419), .S(n10092), .Z(n8364) );
  OAI21_X1 U9845 ( .B1(n8422), .B2(n8394), .A(n8364), .ZN(P2_U3481) );
  INV_X1 U9846 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8367) );
  AOI21_X1 U9847 ( .B1(n8366), .B2(n10068), .A(n8365), .ZN(n8423) );
  MUX2_X1 U9848 ( .A(n8367), .B(n8423), .S(n10092), .Z(n8368) );
  OAI21_X1 U9849 ( .B1(n8426), .B2(n8394), .A(n8368), .ZN(P2_U3480) );
  INV_X1 U9850 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8371) );
  AOI21_X1 U9851 ( .B1(n8370), .B2(n10068), .A(n8369), .ZN(n8427) );
  MUX2_X1 U9852 ( .A(n8371), .B(n8427), .S(n10092), .Z(n8372) );
  OAI21_X1 U9853 ( .B1(n8430), .B2(n8394), .A(n8372), .ZN(P2_U3479) );
  AOI21_X1 U9854 ( .B1(n10068), .B2(n8374), .A(n8373), .ZN(n8431) );
  MUX2_X1 U9855 ( .A(n8375), .B(n8431), .S(n10092), .Z(n8376) );
  OAI21_X1 U9856 ( .B1(n8434), .B2(n8394), .A(n8376), .ZN(P2_U3478) );
  AOI21_X1 U9857 ( .B1(n8378), .B2(n10068), .A(n8377), .ZN(n8435) );
  MUX2_X1 U9858 ( .A(n8379), .B(n8435), .S(n10092), .Z(n8380) );
  OAI21_X1 U9859 ( .B1(n8438), .B2(n8394), .A(n8380), .ZN(P2_U3477) );
  AOI21_X1 U9860 ( .B1(n10068), .B2(n8382), .A(n8381), .ZN(n8439) );
  MUX2_X1 U9861 ( .A(n8383), .B(n8439), .S(n10092), .Z(n8384) );
  OAI21_X1 U9862 ( .B1(n8442), .B2(n8394), .A(n8384), .ZN(P2_U3476) );
  NAND2_X1 U9863 ( .A1(n8385), .A2(n10068), .ZN(n8386) );
  AND2_X1 U9864 ( .A1(n8387), .A2(n8386), .ZN(n8443) );
  MUX2_X1 U9865 ( .A(n8388), .B(n8443), .S(n10092), .Z(n8389) );
  OAI21_X1 U9866 ( .B1(n8446), .B2(n8394), .A(n8389), .ZN(P2_U3475) );
  AOI21_X1 U9867 ( .B1(n8391), .B2(n10068), .A(n8390), .ZN(n8447) );
  MUX2_X1 U9868 ( .A(n8392), .B(n8447), .S(n10092), .Z(n8393) );
  OAI21_X1 U9869 ( .B1(n8451), .B2(n8394), .A(n8393), .ZN(P2_U3474) );
  NAND2_X1 U9870 ( .A1(n8395), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U9871 ( .A1(n8396), .A2(n10074), .ZN(n8399) );
  OAI211_X1 U9872 ( .C1(n6843), .C2(n10074), .A(n8397), .B(n8399), .ZN(
        P2_U3458) );
  NAND2_X1 U9873 ( .A1(n7744), .A2(n8398), .ZN(n8400) );
  OAI211_X1 U9874 ( .C1(n5576), .C2(n10074), .A(n8400), .B(n8399), .ZN(
        P2_U3457) );
  MUX2_X1 U9875 ( .A(n8402), .B(n8401), .S(n10074), .Z(n8403) );
  OAI21_X1 U9876 ( .B1(n8404), .B2(n8450), .A(n8403), .ZN(P2_U3454) );
  MUX2_X1 U9877 ( .A(n8406), .B(n8405), .S(n10074), .Z(n8407) );
  OAI21_X1 U9878 ( .B1(n8408), .B2(n8450), .A(n8407), .ZN(P2_U3453) );
  MUX2_X1 U9879 ( .A(n8410), .B(n8409), .S(n10074), .Z(n8411) );
  OAI21_X1 U9880 ( .B1(n8412), .B2(n8450), .A(n8411), .ZN(P2_U3452) );
  MUX2_X1 U9881 ( .A(n9083), .B(n8413), .S(n10074), .Z(n8414) );
  OAI21_X1 U9882 ( .B1(n8415), .B2(n8450), .A(n8414), .ZN(P2_U3451) );
  MUX2_X1 U9883 ( .A(n9035), .B(n8416), .S(n10074), .Z(n8417) );
  OAI21_X1 U9884 ( .B1(n8418), .B2(n8450), .A(n8417), .ZN(P2_U3450) );
  INV_X1 U9885 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8420) );
  MUX2_X1 U9886 ( .A(n8420), .B(n8419), .S(n10074), .Z(n8421) );
  OAI21_X1 U9887 ( .B1(n8422), .B2(n8450), .A(n8421), .ZN(P2_U3449) );
  INV_X1 U9888 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8424) );
  MUX2_X1 U9889 ( .A(n8424), .B(n8423), .S(n10074), .Z(n8425) );
  OAI21_X1 U9890 ( .B1(n8426), .B2(n8450), .A(n8425), .ZN(P2_U3448) );
  INV_X1 U9891 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8428) );
  MUX2_X1 U9892 ( .A(n8428), .B(n8427), .S(n10074), .Z(n8429) );
  OAI21_X1 U9893 ( .B1(n8430), .B2(n8450), .A(n8429), .ZN(P2_U3447) );
  MUX2_X1 U9894 ( .A(n8432), .B(n8431), .S(n10074), .Z(n8433) );
  OAI21_X1 U9895 ( .B1(n8434), .B2(n8450), .A(n8433), .ZN(P2_U3446) );
  MUX2_X1 U9896 ( .A(n8436), .B(n8435), .S(n10074), .Z(n8437) );
  OAI21_X1 U9897 ( .B1(n8438), .B2(n8450), .A(n8437), .ZN(P2_U3444) );
  INV_X1 U9898 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8440) );
  MUX2_X1 U9899 ( .A(n8440), .B(n8439), .S(n10074), .Z(n8441) );
  OAI21_X1 U9900 ( .B1(n8442), .B2(n8450), .A(n8441), .ZN(P2_U3441) );
  INV_X1 U9901 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8444) );
  MUX2_X1 U9902 ( .A(n8444), .B(n8443), .S(n10074), .Z(n8445) );
  OAI21_X1 U9903 ( .B1(n8446), .B2(n8450), .A(n8445), .ZN(P2_U3438) );
  INV_X1 U9904 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8448) );
  MUX2_X1 U9905 ( .A(n8448), .B(n8447), .S(n10074), .Z(n8449) );
  OAI21_X1 U9906 ( .B1(n8451), .B2(n8450), .A(n8449), .ZN(P2_U3435) );
  INV_X1 U9907 ( .A(n8731), .ZN(n9552) );
  NOR4_X1 U9908 ( .A1(n4862), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n8452), .ZN(n8453) );
  AOI21_X1 U9909 ( .B1(n8465), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8453), .ZN(
        n8454) );
  OAI21_X1 U9910 ( .B1(n9552), .B2(n8467), .A(n8454), .ZN(P2_U3264) );
  INV_X1 U9911 ( .A(n8720), .ZN(n9553) );
  OAI222_X1 U9912 ( .A1(n8457), .A2(n9553), .B1(n8456), .B2(n5568), .C1(
        P2_U3151), .C2(n8455), .ZN(P2_U3266) );
  NAND2_X1 U9913 ( .A1(n8459), .A2(n8458), .ZN(n8461) );
  OAI211_X1 U9914 ( .C1(n8462), .C2(n8456), .A(n8461), .B(n8460), .ZN(P2_U3267) );
  INV_X1 U9915 ( .A(n8463), .ZN(n9557) );
  AOI21_X1 U9916 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(n8465), .A(n8464), .ZN(
        n8466) );
  OAI21_X1 U9917 ( .B1(n9557), .B2(n8467), .A(n8466), .ZN(P2_U3268) );
  MUX2_X1 U9918 ( .A(n8468), .B(P2_IR_REG_0__SCAN_IN), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  AOI21_X1 U9919 ( .B1(n8470), .B2(n8469), .A(n4396), .ZN(n8478) );
  NAND2_X1 U9920 ( .A1(n8471), .A2(n8599), .ZN(n8473) );
  OAI211_X1 U9921 ( .C1(n9674), .C2(n8474), .A(n8473), .B(n8472), .ZN(n8475)
         );
  AOI21_X1 U9922 ( .B1(n8476), .B2(n9670), .A(n8475), .ZN(n8477) );
  OAI21_X1 U9923 ( .B1(n8478), .B2(n9665), .A(n8477), .ZN(P1_U3215) );
  OAI21_X1 U9924 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8486) );
  INV_X1 U9925 ( .A(n8483), .ZN(n8565) );
  XOR2_X1 U9926 ( .A(n8486), .B(n8485), .Z(n8492) );
  NOR2_X1 U9927 ( .A1(n9674), .A2(n9282), .ZN(n8490) );
  AND2_X1 U9928 ( .A1(n9157), .A2(n9199), .ZN(n8487) );
  AOI21_X1 U9929 ( .B1(n9162), .B2(n8988), .A(n8487), .ZN(n9286) );
  OAI22_X1 U9930 ( .A1(n9286), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8488), .ZN(n8489) );
  AOI211_X1 U9931 ( .C1(n9291), .C2(n9670), .A(n8490), .B(n8489), .ZN(n8491)
         );
  OAI21_X1 U9932 ( .B1(n8492), .B2(n9665), .A(n8491), .ZN(P1_U3216) );
  OAI21_X1 U9933 ( .B1(n8494), .B2(n8493), .A(n9664), .ZN(n8495) );
  NAND2_X1 U9934 ( .A1(n8495), .A2(n9649), .ZN(n8500) );
  AOI22_X1 U9935 ( .A1(n9670), .A2(n8497), .B1(n8496), .B2(n8599), .ZN(n8499)
         );
  MUX2_X1 U9936 ( .A(n9674), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n8498) );
  NAND3_X1 U9937 ( .A1(n8500), .A2(n8499), .A3(n8498), .ZN(P1_U3218) );
  NAND2_X1 U9938 ( .A1(n4588), .A2(n8503), .ZN(n8504) );
  XNOR2_X1 U9939 ( .A(n8501), .B(n8504), .ZN(n8510) );
  NAND2_X1 U9940 ( .A1(n9147), .A2(n9199), .ZN(n8506) );
  NAND2_X1 U9941 ( .A1(n9153), .A2(n8988), .ZN(n8505) );
  NAND2_X1 U9942 ( .A1(n8506), .A2(n8505), .ZN(n9349) );
  AOI22_X1 U9943 ( .A1(n9349), .A2(n8599), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n8507) );
  OAI21_X1 U9944 ( .B1(n9674), .B2(n9357), .A(n8507), .ZN(n8508) );
  AOI21_X1 U9945 ( .B1(n9356), .B2(n9670), .A(n8508), .ZN(n8509) );
  OAI21_X1 U9946 ( .B1(n8510), .B2(n9665), .A(n8509), .ZN(P1_U3219) );
  XOR2_X1 U9947 ( .A(n8512), .B(n8511), .Z(n8517) );
  AOI22_X1 U9948 ( .A1(n9157), .A2(n8988), .B1(n9153), .B2(n9199), .ZN(n9319)
         );
  OAI22_X1 U9949 ( .A1(n9319), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8513), .ZN(n8514) );
  AOI21_X1 U9950 ( .B1(n9324), .B2(n8591), .A(n8514), .ZN(n8516) );
  NAND2_X1 U9951 ( .A1(n9323), .A2(n9670), .ZN(n8515) );
  OAI211_X1 U9952 ( .C1(n8517), .C2(n9665), .A(n8516), .B(n8515), .ZN(P1_U3223) );
  NOR2_X1 U9953 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  OAI21_X1 U9954 ( .B1(n8518), .B2(n8521), .A(n9649), .ZN(n8527) );
  INV_X1 U9955 ( .A(n8522), .ZN(n9258) );
  AND2_X1 U9956 ( .A1(n9162), .A2(n9199), .ZN(n8523) );
  AOI21_X1 U9957 ( .B1(n8884), .B2(n8988), .A(n8523), .ZN(n9253) );
  OAI22_X1 U9958 ( .A1(n9253), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8524), .ZN(n8525) );
  AOI21_X1 U9959 ( .B1(n9258), .B2(n8591), .A(n8525), .ZN(n8526) );
  OAI211_X1 U9960 ( .C1(n8594), .C2(n9514), .A(n8527), .B(n8526), .ZN(P1_U3225) );
  OAI21_X1 U9961 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8531) );
  NAND2_X1 U9962 ( .A1(n8531), .A2(n9649), .ZN(n8535) );
  INV_X1 U9963 ( .A(n9408), .ZN(n8533) );
  AOI22_X1 U9964 ( .A1(n9199), .A2(n8885), .B1(n9144), .B2(n8577), .ZN(n9401)
         );
  OAI22_X1 U9965 ( .A1(n9401), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8927), .ZN(n8532) );
  AOI21_X1 U9966 ( .B1(n8533), .B2(n8591), .A(n8532), .ZN(n8534) );
  OAI211_X1 U9967 ( .C1(n4652), .C2(n8594), .A(n8535), .B(n8534), .ZN(P1_U3226) );
  INV_X1 U9968 ( .A(n9392), .ZN(n9543) );
  OAI21_X1 U9969 ( .B1(n8538), .B2(n8537), .A(n8536), .ZN(n8539) );
  NAND2_X1 U9970 ( .A1(n8539), .A2(n9649), .ZN(n8544) );
  NAND2_X1 U9971 ( .A1(n9147), .A2(n8577), .ZN(n8541) );
  NAND2_X1 U9972 ( .A1(n9141), .A2(n9199), .ZN(n8540) );
  NAND2_X1 U9973 ( .A1(n8541), .A2(n8540), .ZN(n9388) );
  AND2_X1 U9974 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8946) );
  NOR2_X1 U9975 ( .A1(n9674), .A2(n9393), .ZN(n8542) );
  AOI211_X1 U9976 ( .C1(n8599), .C2(n9388), .A(n8946), .B(n8542), .ZN(n8543)
         );
  OAI211_X1 U9977 ( .C1(n9543), .C2(n8594), .A(n8544), .B(n8543), .ZN(P1_U3228) );
  OAI21_X1 U9978 ( .B1(n8547), .B2(n8546), .A(n8545), .ZN(n8548) );
  NAND2_X1 U9979 ( .A1(n8548), .A2(n9649), .ZN(n8553) );
  AND2_X1 U9980 ( .A1(n9160), .A2(n9199), .ZN(n8549) );
  AOI21_X1 U9981 ( .B1(n9165), .B2(n8988), .A(n8549), .ZN(n9270) );
  OAI22_X1 U9982 ( .A1(n9270), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8550), .ZN(n8551) );
  AOI21_X1 U9983 ( .B1(n9276), .B2(n8591), .A(n8551), .ZN(n8552) );
  OAI211_X1 U9984 ( .C1(n8594), .C2(n9518), .A(n8553), .B(n8552), .ZN(P1_U3229) );
  INV_X1 U9985 ( .A(n8554), .ZN(n8555) );
  AOI21_X1 U9986 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8563) );
  NAND2_X1 U9987 ( .A1(n9155), .A2(n8988), .ZN(n8559) );
  NAND2_X1 U9988 ( .A1(n9150), .A2(n9199), .ZN(n8558) );
  NAND2_X1 U9989 ( .A1(n8559), .A2(n8558), .ZN(n9342) );
  AOI22_X1 U9990 ( .A1(n9342), .A2(n8599), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8560) );
  OAI21_X1 U9991 ( .B1(n9674), .B2(n9334), .A(n8560), .ZN(n8561) );
  AOI21_X1 U9992 ( .B1(n9471), .B2(n9670), .A(n8561), .ZN(n8562) );
  OAI21_X1 U9993 ( .B1(n8563), .B2(n9665), .A(n8562), .ZN(P1_U3233) );
  AOI21_X1 U9994 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8572) );
  NAND2_X1 U9995 ( .A1(n9160), .A2(n8577), .ZN(n8568) );
  NAND2_X1 U9996 ( .A1(n9155), .A2(n9199), .ZN(n8567) );
  NAND2_X1 U9997 ( .A1(n8568), .A2(n8567), .ZN(n9301) );
  AOI22_X1 U9998 ( .A1(n9301), .A2(n8599), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8569) );
  OAI21_X1 U9999 ( .B1(n9674), .B2(n9308), .A(n8569), .ZN(n8570) );
  AOI21_X1 U10000 ( .B1(n9307), .B2(n9670), .A(n8570), .ZN(n8571) );
  OAI21_X1 U10001 ( .B1(n8572), .B2(n9665), .A(n8571), .ZN(P1_U3235) );
  NAND2_X1 U10002 ( .A1(n8574), .A2(n8573), .ZN(n8576) );
  XNOR2_X1 U10003 ( .A(n8576), .B(n8575), .ZN(n8583) );
  NAND2_X1 U10004 ( .A1(n9150), .A2(n8577), .ZN(n8579) );
  NAND2_X1 U10005 ( .A1(n9144), .A2(n9199), .ZN(n8578) );
  NAND2_X1 U10006 ( .A1(n8579), .A2(n8578), .ZN(n9370) );
  AOI22_X1 U10007 ( .A1(n9370), .A2(n8599), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n8580) );
  OAI21_X1 U10008 ( .B1(n9674), .B2(n9378), .A(n8580), .ZN(n8581) );
  AOI21_X1 U10009 ( .B1(n9377), .B2(n9670), .A(n8581), .ZN(n8582) );
  OAI21_X1 U10010 ( .B1(n8583), .B2(n9665), .A(n8582), .ZN(P1_U3238) );
  OAI21_X1 U10011 ( .B1(n8518), .B2(n8585), .A(n8584), .ZN(n8586) );
  NAND3_X1 U10012 ( .A1(n8587), .A2(n9649), .A3(n8586), .ZN(n8593) );
  AND2_X1 U10013 ( .A1(n9169), .A2(n8988), .ZN(n8588) );
  AOI21_X1 U10014 ( .B1(n9165), .B2(n9199), .A(n8588), .ZN(n9238) );
  INV_X1 U10015 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8589) );
  OAI22_X1 U10016 ( .A1(n9238), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8589), .ZN(n8590) );
  AOI21_X1 U10017 ( .B1(n9242), .B2(n8591), .A(n8590), .ZN(n8592) );
  OAI211_X1 U10018 ( .C1(n8594), .C2(n4657), .A(n8593), .B(n8592), .ZN(
        P1_U3240) );
  INV_X1 U10019 ( .A(n8595), .ZN(n8596) );
  AOI21_X1 U10020 ( .B1(n8598), .B2(n8597), .A(n8596), .ZN(n8606) );
  NAND2_X1 U10021 ( .A1(n8600), .A2(n8599), .ZN(n8602) );
  OAI211_X1 U10022 ( .C1(n9674), .C2(n8603), .A(n8602), .B(n8601), .ZN(n8604)
         );
  AOI21_X1 U10023 ( .B1(n9139), .B2(n9670), .A(n8604), .ZN(n8605) );
  OAI21_X1 U10024 ( .B1(n8606), .B2(n9665), .A(n8605), .ZN(P1_U3241) );
  NAND2_X1 U10025 ( .A1(n8607), .A2(n8730), .ZN(n8610) );
  OR2_X1 U10026 ( .A1(n8729), .A2(n8608), .ZN(n8609) );
  NAND2_X1 U10027 ( .A1(n8610), .A2(n8609), .ZN(n8740) );
  INV_X1 U10028 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8613) );
  NAND2_X1 U10029 ( .A1(n4307), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8612) );
  INV_X1 U10030 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9424) );
  OR2_X1 U10031 ( .A1(n8615), .A2(n9424), .ZN(n8611) );
  OAI211_X1 U10032 ( .C1(n4309), .C2(n8613), .A(n8612), .B(n8611), .ZN(n9196)
         );
  INV_X1 U10033 ( .A(n9196), .ZN(n8614) );
  OR2_X1 U10034 ( .A1(n8740), .A2(n8614), .ZN(n8739) );
  INV_X1 U10035 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8619) );
  INV_X1 U10036 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9420) );
  OR2_X1 U10037 ( .A1(n8615), .A2(n9420), .ZN(n8618) );
  NAND2_X1 U10038 ( .A1(n4306), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n8617) );
  OAI211_X1 U10039 ( .C1(n4308), .C2(n8619), .A(n8618), .B(n8617), .ZN(n8989)
         );
  INV_X1 U10040 ( .A(n8989), .ZN(n8734) );
  OR2_X1 U10041 ( .A1(n8739), .A2(n8734), .ZN(n8851) );
  NAND2_X1 U10042 ( .A1(n8989), .A2(n9196), .ZN(n8621) );
  NAND2_X1 U10043 ( .A1(n8740), .A2(n8621), .ZN(n8848) );
  MUX2_X1 U10044 ( .A(n8851), .B(n8848), .S(n8738), .Z(n8733) );
  INV_X1 U10045 ( .A(n9141), .ZN(n8645) );
  INV_X1 U10046 ( .A(n8744), .ZN(n8647) );
  INV_X1 U10047 ( .A(n8622), .ZN(n8624) );
  OAI21_X1 U10048 ( .B1(n9722), .B2(n8624), .A(n8623), .ZN(n8626) );
  INV_X1 U10049 ( .A(n8738), .ZN(n8704) );
  MUX2_X1 U10050 ( .A(n8626), .B(n8625), .S(n8704), .Z(n8628) );
  NAND2_X1 U10051 ( .A1(n8628), .A2(n8627), .ZN(n8631) );
  MUX2_X1 U10052 ( .A(n8755), .B(n8629), .S(n8738), .Z(n8630) );
  NAND2_X1 U10053 ( .A1(n8631), .A2(n8630), .ZN(n8636) );
  AND2_X1 U10054 ( .A1(n8638), .A2(n8632), .ZN(n8633) );
  MUX2_X1 U10055 ( .A(n8634), .B(n8633), .S(n8704), .Z(n8635) );
  NAND2_X1 U10056 ( .A1(n8636), .A2(n8635), .ZN(n8649) );
  NAND2_X1 U10057 ( .A1(n8658), .A2(n8652), .ZN(n8640) );
  INV_X1 U10058 ( .A(n8653), .ZN(n8637) );
  OR2_X1 U10059 ( .A1(n8640), .A2(n8637), .ZN(n8798) );
  AOI21_X1 U10060 ( .B1(n8649), .B2(n8638), .A(n8798), .ZN(n8642) );
  OR2_X1 U10061 ( .A1(n8640), .A2(n8639), .ZN(n8641) );
  NAND2_X1 U10062 ( .A1(n8641), .A2(n8656), .ZN(n8800) );
  OAI21_X1 U10063 ( .B1(n8642), .B2(n8800), .A(n8661), .ZN(n8643) );
  NAND3_X1 U10064 ( .A1(n8643), .A2(n4627), .A3(n8799), .ZN(n8644) );
  AND2_X1 U10065 ( .A1(n8744), .A2(n8665), .ZN(n8806) );
  NAND3_X1 U10066 ( .A1(n8644), .A2(n8806), .A3(n8803), .ZN(n8646) );
  OAI211_X1 U10067 ( .C1(n8647), .C2(n8836), .A(n8646), .B(n8838), .ZN(n8670)
         );
  NAND2_X1 U10068 ( .A1(n8649), .A2(n8648), .ZN(n8651) );
  NAND2_X1 U10069 ( .A1(n8651), .A2(n8650), .ZN(n8654) );
  NAND3_X1 U10070 ( .A1(n8654), .A2(n8653), .A3(n8652), .ZN(n8657) );
  NAND3_X1 U10071 ( .A1(n8657), .A2(n8656), .A3(n8655), .ZN(n8659) );
  NAND2_X1 U10072 ( .A1(n8659), .A2(n8658), .ZN(n8660) );
  NAND2_X1 U10073 ( .A1(n8660), .A2(n8799), .ZN(n8664) );
  INV_X1 U10074 ( .A(n8661), .ZN(n8804) );
  NOR2_X1 U10075 ( .A1(n8763), .A2(n8804), .ZN(n8663) );
  NAND2_X1 U10076 ( .A1(n8836), .A2(n8662), .ZN(n8807) );
  AOI21_X1 U10077 ( .B1(n8664), .B2(n8663), .A(n8807), .ZN(n8667) );
  INV_X1 U10078 ( .A(n8665), .ZN(n8666) );
  OAI21_X1 U10079 ( .B1(n8667), .B2(n8666), .A(n8838), .ZN(n8668) );
  NAND2_X1 U10080 ( .A1(n8668), .A2(n8744), .ZN(n8669) );
  MUX2_X1 U10081 ( .A(n8670), .B(n8669), .S(n8704), .Z(n8672) );
  INV_X1 U10082 ( .A(n9144), .ZN(n8671) );
  OR2_X1 U10083 ( .A1(n9392), .A2(n8671), .ZN(n9367) );
  NAND2_X1 U10084 ( .A1(n9392), .A2(n8671), .ZN(n9366) );
  NAND2_X1 U10085 ( .A1(n8672), .A2(n9386), .ZN(n8686) );
  INV_X1 U10086 ( .A(n9147), .ZN(n8674) );
  OR2_X1 U10087 ( .A1(n9377), .A2(n8674), .ZN(n9365) );
  NAND2_X1 U10088 ( .A1(n9365), .A2(n9367), .ZN(n8841) );
  INV_X1 U10089 ( .A(n8841), .ZN(n8673) );
  NAND2_X1 U10090 ( .A1(n8686), .A2(n8673), .ZN(n8675) );
  INV_X1 U10091 ( .A(n9150), .ZN(n8677) );
  NAND2_X1 U10092 ( .A1(n9356), .A2(n8677), .ZN(n8843) );
  NAND2_X1 U10093 ( .A1(n9377), .A2(n8674), .ZN(n9364) );
  NAND3_X1 U10094 ( .A1(n8675), .A2(n8843), .A3(n9364), .ZN(n8682) );
  INV_X1 U10095 ( .A(n9155), .ZN(n8683) );
  OR2_X1 U10096 ( .A1(n9323), .A2(n8683), .ZN(n8844) );
  INV_X1 U10097 ( .A(n9153), .ZN(n8678) );
  INV_X1 U10098 ( .A(n9356), .ZN(n9534) );
  NAND2_X1 U10099 ( .A1(n9179), .A2(n9534), .ZN(n8676) );
  NAND2_X1 U10100 ( .A1(n8676), .A2(n8738), .ZN(n8679) );
  OR2_X1 U10101 ( .A1(n9356), .A2(n8677), .ZN(n8743) );
  OR2_X1 U10102 ( .A1(n9471), .A2(n8678), .ZN(n8845) );
  NAND3_X1 U10103 ( .A1(n8679), .A2(n8743), .A3(n8845), .ZN(n8681) );
  NAND3_X1 U10104 ( .A1(n9179), .A2(n9150), .A3(n8738), .ZN(n8680) );
  NAND2_X1 U10105 ( .A1(n8681), .A2(n8680), .ZN(n8688) );
  NAND3_X1 U10106 ( .A1(n8682), .A2(n8844), .A3(n8688), .ZN(n8685) );
  NAND2_X1 U10107 ( .A1(n9323), .A2(n8683), .ZN(n8742) );
  NAND2_X1 U10108 ( .A1(n8742), .A2(n9179), .ZN(n8684) );
  NAND2_X1 U10109 ( .A1(n8685), .A2(n9180), .ZN(n8693) );
  NAND2_X1 U10110 ( .A1(n9364), .A2(n9366), .ZN(n8840) );
  INV_X1 U10111 ( .A(n8840), .ZN(n8769) );
  NAND2_X1 U10112 ( .A1(n8686), .A2(n8769), .ZN(n8687) );
  AND2_X1 U10113 ( .A1(n8743), .A2(n9365), .ZN(n8810) );
  NAND2_X1 U10114 ( .A1(n8687), .A2(n8810), .ZN(n8689) );
  NAND2_X1 U10115 ( .A1(n8689), .A2(n8688), .ZN(n8691) );
  AND2_X1 U10116 ( .A1(n8844), .A2(n8845), .ZN(n8812) );
  INV_X1 U10117 ( .A(n8742), .ZN(n8690) );
  AOI21_X1 U10118 ( .B1(n8691), .B2(n8812), .A(n8690), .ZN(n8692) );
  INV_X1 U10119 ( .A(n9157), .ZN(n8694) );
  OR2_X1 U10120 ( .A1(n9307), .A2(n8694), .ZN(n9181) );
  NAND2_X1 U10121 ( .A1(n9307), .A2(n8694), .ZN(n9182) );
  NAND2_X1 U10122 ( .A1(n9181), .A2(n9182), .ZN(n9299) );
  NAND2_X1 U10123 ( .A1(n8741), .A2(n9181), .ZN(n8782) );
  NAND2_X1 U10124 ( .A1(n9291), .A2(n8695), .ZN(n9265) );
  NAND2_X1 U10125 ( .A1(n9265), .A2(n9182), .ZN(n8816) );
  INV_X1 U10126 ( .A(n9162), .ZN(n8697) );
  NAND2_X1 U10127 ( .A1(n9275), .A2(n8697), .ZN(n8818) );
  NAND2_X1 U10128 ( .A1(n9185), .A2(n8818), .ZN(n9266) );
  INV_X1 U10129 ( .A(n9266), .ZN(n8699) );
  MUX2_X1 U10130 ( .A(n9265), .B(n8741), .S(n8738), .Z(n8698) );
  MUX2_X1 U10131 ( .A(n9185), .B(n8818), .S(n8738), .Z(n8701) );
  INV_X1 U10132 ( .A(n8884), .ZN(n8713) );
  NAND2_X1 U10133 ( .A1(n9241), .A2(n8713), .ZN(n9189) );
  NAND2_X1 U10134 ( .A1(n9257), .A2(n8702), .ZN(n9186) );
  NAND3_X1 U10135 ( .A1(n9189), .A2(n8704), .A3(n9186), .ZN(n8703) );
  AOI21_X1 U10136 ( .B1(n8709), .B2(n9187), .A(n8703), .ZN(n8708) );
  INV_X1 U10137 ( .A(n9169), .ZN(n8706) );
  NOR2_X1 U10138 ( .A1(n9241), .A2(n8713), .ZN(n9190) );
  NAND2_X1 U10139 ( .A1(n9190), .A2(n8704), .ZN(n8705) );
  NAND2_X1 U10140 ( .A1(n8779), .A2(n8705), .ZN(n8707) );
  INV_X1 U10141 ( .A(n9200), .ZN(n9170) );
  NAND2_X1 U10142 ( .A1(n9212), .A2(n9170), .ZN(n9193) );
  NAND2_X1 U10143 ( .A1(n9228), .A2(n8706), .ZN(n9191) );
  AND2_X1 U10144 ( .A1(n9193), .A2(n9191), .ZN(n8712) );
  OAI21_X1 U10145 ( .B1(n8708), .B2(n8707), .A(n8712), .ZN(n8719) );
  INV_X1 U10146 ( .A(n9186), .ZN(n8819) );
  NAND2_X1 U10147 ( .A1(n9187), .A2(n8738), .ZN(n8710) );
  NOR2_X1 U10148 ( .A1(n9190), .A2(n8710), .ZN(n8711) );
  INV_X1 U10149 ( .A(n8712), .ZN(n8824) );
  NAND2_X1 U10150 ( .A1(n8824), .A2(n8738), .ZN(n8715) );
  NAND3_X1 U10151 ( .A1(n9241), .A2(n8713), .A3(n8738), .ZN(n8714) );
  OAI21_X1 U10152 ( .B1(n8824), .B2(n8779), .A(n8777), .ZN(n8717) );
  AOI22_X1 U10153 ( .A1(n8719), .A2(n8718), .B1(n8738), .B2(n8717), .ZN(n8726)
         );
  NAND2_X1 U10154 ( .A1(n8720), .A2(n8730), .ZN(n8723) );
  OR2_X1 U10155 ( .A1(n8729), .A2(n8721), .ZN(n8722) );
  INV_X1 U10156 ( .A(n8724), .ZN(n8725) );
  NAND2_X1 U10157 ( .A1(n9428), .A2(n8725), .ZN(n8826) );
  MUX2_X1 U10158 ( .A(n8826), .B(n8778), .S(n8738), .Z(n8727) );
  NAND4_X1 U10159 ( .A1(n8728), .A2(n8727), .A3(n8848), .A4(n8851), .ZN(n8732)
         );
  AND2_X1 U10160 ( .A1(n9496), .A2(n8989), .ZN(n8871) );
  INV_X1 U10161 ( .A(n8871), .ZN(n8831) );
  NAND2_X1 U10162 ( .A1(n8735), .A2(n8734), .ZN(n8867) );
  OAI211_X1 U10163 ( .C1(n8738), .C2(n8737), .A(n8853), .B(n8980), .ZN(n8776)
         );
  NAND2_X1 U10164 ( .A1(n8867), .A2(n8739), .ZN(n8832) );
  NOR2_X1 U10165 ( .A1(n9500), .A2(n9196), .ZN(n8829) );
  NAND2_X1 U10166 ( .A1(n8777), .A2(n9193), .ZN(n9207) );
  AND2_X2 U10167 ( .A1(n8779), .A2(n9191), .ZN(n9221) );
  AND2_X1 U10168 ( .A1(n9187), .A2(n9186), .ZN(n9249) );
  INV_X1 U10169 ( .A(n9299), .ZN(n9304) );
  NOR2_X1 U10170 ( .A1(n8745), .A2(n9747), .ZN(n8751) );
  NOR2_X1 U10171 ( .A1(n8746), .A2(n6772), .ZN(n8750) );
  NOR2_X1 U10172 ( .A1(n8747), .A2(n8786), .ZN(n8748) );
  NAND4_X1 U10173 ( .A1(n8751), .A2(n8750), .A3(n8749), .A4(n8748), .ZN(n8752)
         );
  NOR2_X1 U10174 ( .A1(n8752), .A2(n9730), .ZN(n8757) );
  INV_X1 U10175 ( .A(n8753), .ZN(n8756) );
  NAND4_X1 U10176 ( .A1(n8757), .A2(n8756), .A3(n8755), .A4(n8754), .ZN(n8759)
         );
  NOR2_X1 U10177 ( .A1(n8759), .A2(n8758), .ZN(n8760) );
  NAND4_X1 U10178 ( .A1(n8762), .A2(n4635), .A3(n8761), .A4(n8760), .ZN(n8764)
         );
  NOR2_X1 U10179 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  NAND3_X1 U10180 ( .A1(n9414), .A2(n8766), .A3(n8765), .ZN(n8767) );
  NOR2_X1 U10181 ( .A1(n8841), .A2(n8767), .ZN(n8768) );
  AND4_X1 U10182 ( .A1(n9341), .A2(n8769), .A3(n9353), .A4(n8768), .ZN(n8770)
         );
  NAND4_X1 U10183 ( .A1(n9295), .A2(n9304), .A3(n9317), .A4(n8770), .ZN(n8771)
         );
  NOR2_X1 U10184 ( .A1(n9266), .A2(n8771), .ZN(n8773) );
  NOR2_X1 U10185 ( .A1(n9241), .A2(n8884), .ZN(n9167) );
  NAND2_X1 U10186 ( .A1(n9241), .A2(n8884), .ZN(n9168) );
  INV_X1 U10187 ( .A(n9168), .ZN(n8772) );
  OR2_X1 U10188 ( .A1(n9167), .A2(n8772), .ZN(n9236) );
  NAND4_X1 U10189 ( .A1(n9221), .A2(n9249), .A3(n8773), .A4(n9236), .ZN(n8774)
         );
  NAND2_X1 U10190 ( .A1(n8778), .A2(n8777), .ZN(n8828) );
  INV_X1 U10191 ( .A(n9190), .ZN(n8780) );
  NAND2_X1 U10192 ( .A1(n8780), .A2(n8779), .ZN(n8822) );
  INV_X1 U10193 ( .A(n9185), .ZN(n8781) );
  AOI21_X1 U10194 ( .B1(n9265), .B2(n8782), .A(n8781), .ZN(n8784) );
  INV_X1 U10195 ( .A(n8818), .ZN(n8783) );
  OAI21_X1 U10196 ( .B1(n8784), .B2(n8783), .A(n9187), .ZN(n8815) );
  NOR3_X1 U10197 ( .A1(n8828), .A2(n8822), .A3(n8815), .ZN(n8846) );
  INV_X1 U10198 ( .A(n8785), .ZN(n8797) );
  AND4_X1 U10199 ( .A1(n8789), .A2(n8788), .A3(n8787), .A4(n8786), .ZN(n8793)
         );
  NAND4_X1 U10200 ( .A1(n8793), .A2(n8792), .A3(n8791), .A4(n8790), .ZN(n8796)
         );
  INV_X1 U10201 ( .A(n8794), .ZN(n8795) );
  AOI21_X1 U10202 ( .B1(n8797), .B2(n8796), .A(n8795), .ZN(n8802) );
  INV_X1 U10203 ( .A(n8798), .ZN(n8801) );
  AOI211_X1 U10204 ( .C1(n8802), .C2(n8801), .A(n4633), .B(n8800), .ZN(n8805)
         );
  NOR3_X1 U10205 ( .A1(n8805), .A2(n8804), .A3(n4632), .ZN(n8808) );
  OAI21_X1 U10206 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8809) );
  AOI21_X1 U10207 ( .B1(n8809), .B2(n8838), .A(n8841), .ZN(n8811) );
  OAI21_X1 U10208 ( .B1(n8811), .B2(n8840), .A(n8810), .ZN(n8814) );
  INV_X1 U10209 ( .A(n8812), .ZN(n8813) );
  AOI21_X1 U10210 ( .B1(n8814), .B2(n8843), .A(n8813), .ZN(n8830) );
  INV_X1 U10211 ( .A(n8815), .ZN(n8821) );
  INV_X1 U10212 ( .A(n8816), .ZN(n8817) );
  NAND3_X1 U10213 ( .A1(n8818), .A2(n8817), .A3(n9180), .ZN(n8820) );
  AOI21_X1 U10214 ( .B1(n8821), .B2(n8820), .A(n8819), .ZN(n8823) );
  AOI21_X1 U10215 ( .B1(n8823), .B2(n9189), .A(n8822), .ZN(n8825) );
  NOR2_X1 U10216 ( .A1(n8825), .A2(n8824), .ZN(n8827) );
  AOI211_X1 U10217 ( .C1(n8846), .C2(n8830), .A(n8829), .B(n8847), .ZN(n8833)
         );
  NAND2_X1 U10218 ( .A1(n9400), .A2(n9414), .ZN(n8839) );
  NAND2_X1 U10219 ( .A1(n8841), .A2(n9364), .ZN(n8842) );
  NAND4_X1 U10220 ( .A1(n8846), .A2(n9340), .A3(n8845), .A4(n8844), .ZN(n8850)
         );
  INV_X1 U10221 ( .A(n8847), .ZN(n8849) );
  NAND3_X1 U10222 ( .A1(n8850), .A2(n8849), .A3(n8848), .ZN(n8852) );
  AOI21_X1 U10223 ( .B1(n8852), .B2(n8851), .A(n8871), .ZN(n8856) );
  INV_X1 U10224 ( .A(n8867), .ZN(n8855) );
  NAND2_X1 U10225 ( .A1(n8853), .A2(n8866), .ZN(n8858) );
  NOR4_X1 U10226 ( .A1(n8856), .A2(n8855), .A3(n8854), .A4(n8858), .ZN(n8861)
         );
  INV_X1 U10227 ( .A(n8857), .ZN(n8859) );
  NOR2_X1 U10228 ( .A1(n8859), .A2(n8858), .ZN(n8860) );
  INV_X1 U10229 ( .A(n8864), .ZN(n8865) );
  OAI21_X1 U10230 ( .B1(n8867), .B2(n8866), .A(n8865), .ZN(n8880) );
  INV_X1 U10231 ( .A(n8882), .ZN(n8869) );
  NAND2_X1 U10232 ( .A1(n8869), .A2(n8868), .ZN(n8874) );
  AOI211_X1 U10233 ( .C1(n8871), .C2(n8980), .A(n8870), .B(n8874), .ZN(n8879)
         );
  NOR2_X1 U10234 ( .A1(n8873), .A2(n8872), .ZN(n8876) );
  INV_X1 U10235 ( .A(P1_B_REG_SCAN_IN), .ZN(n9019) );
  INV_X1 U10236 ( .A(n8874), .ZN(n8875) );
  AOI211_X1 U10237 ( .C1(n8877), .C2(n8876), .A(n9019), .B(n8875), .ZN(n8878)
         );
  AOI21_X1 U10238 ( .B1(n8880), .B2(n8879), .A(n8878), .ZN(n8881) );
  OAI21_X1 U10239 ( .B1(n8883), .B2(n8882), .A(n8881), .ZN(P1_U3242) );
  MUX2_X1 U10240 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n8989), .S(P1_U3973), .Z(
        P1_U3585) );
  MUX2_X1 U10241 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10242 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9200), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10243 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9169), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10244 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8884), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10245 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9165), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10246 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9162), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10247 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9160), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10248 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9157), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10249 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9155), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10250 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9153), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10251 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9150), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10252 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9147), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10253 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9144), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10254 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9141), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10255 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8885), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10256 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n8886), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10257 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8887), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10258 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8888), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10259 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n8889), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10260 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n8890), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10261 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n8891), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10262 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n8892), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10263 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n8893), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10264 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n8894), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10265 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n8895), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10266 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n8896), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10267 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n8897), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10268 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n8898), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10269 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6752), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10270 ( .C1(n8901), .C2(n8900), .A(n9695), .B(n8899), .ZN(n8910)
         );
  OAI211_X1 U10271 ( .C1(n8904), .C2(n8903), .A(n8975), .B(n8902), .ZN(n8909)
         );
  AOI22_X1 U10272 ( .A1(n9679), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n8908) );
  NAND2_X1 U10273 ( .A1(n8906), .A2(n8905), .ZN(n8907) );
  NAND4_X1 U10274 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(
        P1_U3244) );
  NAND2_X1 U10275 ( .A1(n8912), .A2(n8911), .ZN(n8914) );
  NAND2_X1 U10276 ( .A1(n8914), .A2(n8913), .ZN(n8918) );
  NOR2_X1 U10277 ( .A1(n8934), .A2(n8915), .ZN(n8916) );
  AOI21_X1 U10278 ( .B1(n8915), .B2(n8934), .A(n8916), .ZN(n8917) );
  NOR2_X1 U10279 ( .A1(n8917), .A2(n8918), .ZN(n8940) );
  AOI21_X1 U10280 ( .B1(n8918), .B2(n8917), .A(n8940), .ZN(n8932) );
  NOR2_X1 U10281 ( .A1(n8920), .A2(n8919), .ZN(n8922) );
  NAND2_X1 U10282 ( .A1(n8934), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8923) );
  OAI21_X1 U10283 ( .B1(n8934), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8923), .ZN(
        n8924) );
  AOI211_X1 U10284 ( .C1(n8925), .C2(n8924), .A(n8933), .B(n8960), .ZN(n8926)
         );
  INV_X1 U10285 ( .A(n8926), .ZN(n8931) );
  NOR2_X1 U10286 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8927), .ZN(n8929) );
  NOR2_X1 U10287 ( .A1(n9689), .A2(n8941), .ZN(n8928) );
  AOI211_X1 U10288 ( .C1(n9679), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n8929), .B(
        n8928), .ZN(n8930) );
  OAI211_X1 U10289 ( .C1(n8932), .C2(n9691), .A(n8931), .B(n8930), .ZN(
        P1_U3259) );
  AOI22_X1 U10290 ( .A1(n8957), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n5985), .B2(
        n8949), .ZN(n8935) );
  AOI221_X1 U10291 ( .B1(n8936), .B2(n8956), .C1(n8935), .C2(n8956), .A(n8960), 
        .ZN(n8937) );
  INV_X1 U10292 ( .A(n8937), .ZN(n8948) );
  NOR2_X1 U10293 ( .A1(n8957), .A2(n8938), .ZN(n8939) );
  AOI21_X1 U10294 ( .B1(n8938), .B2(n8957), .A(n8939), .ZN(n8943) );
  AOI21_X1 U10295 ( .B1(n8941), .B2(n8915), .A(n8940), .ZN(n8942) );
  NOR2_X1 U10296 ( .A1(n8942), .A2(n8943), .ZN(n8950) );
  AOI21_X1 U10297 ( .B1(n8943), .B2(n8942), .A(n8950), .ZN(n8944) );
  NOR2_X1 U10298 ( .A1(n9691), .A2(n8944), .ZN(n8945) );
  AOI211_X1 U10299 ( .C1(n9679), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n8946), .B(
        n8945), .ZN(n8947) );
  OAI211_X1 U10300 ( .C1(n9689), .C2(n8949), .A(n8948), .B(n8947), .ZN(
        P1_U3260) );
  INV_X1 U10301 ( .A(n8971), .ZN(n8967) );
  INV_X1 U10302 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9483) );
  XNOR2_X1 U10303 ( .A(n8971), .B(n9483), .ZN(n8954) );
  OR2_X1 U10304 ( .A1(n8957), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8952) );
  INV_X1 U10305 ( .A(n8950), .ZN(n8951) );
  AND2_X1 U10306 ( .A1(n8952), .A2(n8951), .ZN(n8953) );
  NAND2_X1 U10307 ( .A1(n8954), .A2(n8953), .ZN(n8973) );
  OAI211_X1 U10308 ( .C1(n8954), .C2(n8953), .A(n8975), .B(n8973), .ZN(n8966)
         );
  NOR2_X1 U10309 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8955), .ZN(n8964) );
  OR2_X1 U10310 ( .A1(n8971), .A2(n9379), .ZN(n8959) );
  NAND2_X1 U10311 ( .A1(n8971), .A2(n9379), .ZN(n8958) );
  AND2_X1 U10312 ( .A1(n8959), .A2(n8958), .ZN(n8961) );
  AOI211_X1 U10313 ( .C1(n8962), .C2(n8961), .A(n8969), .B(n8960), .ZN(n8963)
         );
  AOI211_X1 U10314 ( .C1(n9679), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n8964), .B(
        n8963), .ZN(n8965) );
  OAI211_X1 U10315 ( .C1(n9689), .C2(n8967), .A(n8966), .B(n8965), .ZN(
        P1_U3261) );
  INV_X1 U10316 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8985) );
  AND2_X1 U10317 ( .A1(n8971), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n8968) );
  OR2_X1 U10318 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  XNOR2_X1 U10319 ( .A(n8970), .B(n9358), .ZN(n8976) );
  NAND2_X1 U10320 ( .A1(n8971), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8972) );
  NAND2_X1 U10321 ( .A1(n8973), .A2(n8972), .ZN(n8974) );
  XNOR2_X1 U10322 ( .A(n8974), .B(n9478), .ZN(n8977) );
  AOI22_X1 U10323 ( .A1(n8976), .A2(n9695), .B1(n8975), .B2(n8977), .ZN(n8982)
         );
  INV_X1 U10324 ( .A(n8976), .ZN(n8979) );
  OAI21_X1 U10325 ( .B1(n9691), .B2(n8977), .A(n9689), .ZN(n8978) );
  AOI21_X1 U10326 ( .B1(n8979), .B2(n9695), .A(n8978), .ZN(n8981) );
  MUX2_X1 U10327 ( .A(n8982), .B(n8981), .S(n8980), .Z(n8984) );
  NAND2_X1 U10328 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n8983) );
  OAI211_X1 U10329 ( .C1(n8985), .C2(n9699), .A(n8984), .B(n8983), .ZN(
        P1_U3262) );
  INV_X1 U10330 ( .A(n9428), .ZN(n9178) );
  INV_X1 U10331 ( .A(n9377), .ZN(n9538) );
  INV_X1 U10332 ( .A(n9471), .ZN(n9338) );
  NAND2_X1 U10333 ( .A1(n9500), .A2(n9173), .ZN(n9133) );
  XNOR2_X1 U10334 ( .A(n9496), .B(n9133), .ZN(n8986) );
  NAND2_X1 U10335 ( .A1(n8986), .A2(n9750), .ZN(n9419) );
  OR2_X1 U10336 ( .A1(n9677), .A2(n9019), .ZN(n8987) );
  AND2_X1 U10337 ( .A1(n8988), .A2(n8987), .ZN(n9197) );
  NAND2_X1 U10338 ( .A1(n8989), .A2(n9197), .ZN(n9422) );
  NOR2_X1 U10339 ( .A1(n9422), .A2(n9758), .ZN(n9135) );
  NOR2_X1 U10340 ( .A1(n9496), .A2(n9744), .ZN(n8990) );
  AOI211_X1 U10341 ( .C1(n9758), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9135), .B(
        n8990), .ZN(n8991) );
  OAI21_X1 U10342 ( .B1(n9419), .B2(n9413), .A(n8991), .ZN(n9132) );
  INV_X1 U10343 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n8993) );
  AOI22_X1 U10344 ( .A1(n8993), .A2(keyinput30), .B1(keyinput59), .B2(n6890), 
        .ZN(n8992) );
  OAI221_X1 U10345 ( .B1(n8993), .B2(keyinput30), .C1(n6890), .C2(keyinput59), 
        .A(n8992), .ZN(n8999) );
  INV_X1 U10346 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8995) );
  AOI22_X1 U10347 ( .A1(n5176), .A2(keyinput6), .B1(n8995), .B2(keyinput29), 
        .ZN(n8994) );
  OAI221_X1 U10348 ( .B1(n5176), .B2(keyinput6), .C1(n8995), .C2(keyinput29), 
        .A(n8994), .ZN(n8998) );
  AOI22_X1 U10349 ( .A1(n9740), .A2(keyinput43), .B1(keyinput37), .B2(n4791), 
        .ZN(n8996) );
  OAI221_X1 U10350 ( .B1(n9740), .B2(keyinput43), .C1(n4791), .C2(keyinput37), 
        .A(n8996), .ZN(n8997) );
  NOR3_X1 U10351 ( .A1(n8999), .A2(n8998), .A3(n8997), .ZN(n9016) );
  INV_X1 U10352 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9844) );
  AOI22_X1 U10353 ( .A1(n9103), .A2(keyinput20), .B1(keyinput36), .B2(n9844), 
        .ZN(n9000) );
  OAI221_X1 U10354 ( .B1(n9103), .B2(keyinput20), .C1(n9844), .C2(keyinput36), 
        .A(n9000), .ZN(n9004) );
  INV_X1 U10355 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9002) );
  AOI22_X1 U10356 ( .A1(n9002), .A2(keyinput14), .B1(n5985), .B2(keyinput25), 
        .ZN(n9001) );
  OAI221_X1 U10357 ( .B1(n9002), .B2(keyinput14), .C1(n5985), .C2(keyinput25), 
        .A(n9001), .ZN(n9003) );
  NOR2_X1 U10358 ( .A1(n9004), .A2(n9003), .ZN(n9015) );
  INV_X1 U10359 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9923) );
  AOI22_X1 U10360 ( .A1(n9102), .A2(keyinput46), .B1(keyinput10), .B2(n9923), 
        .ZN(n9005) );
  OAI221_X1 U10361 ( .B1(n9102), .B2(keyinput46), .C1(n9923), .C2(keyinput10), 
        .A(n9005), .ZN(n9008) );
  INV_X1 U10362 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10099) );
  INV_X1 U10363 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U10364 ( .A1(n10099), .A2(keyinput13), .B1(keyinput22), .B2(n10094), 
        .ZN(n9006) );
  OAI221_X1 U10365 ( .B1(n10099), .B2(keyinput13), .C1(n10094), .C2(keyinput22), .A(n9006), .ZN(n9007) );
  NOR2_X1 U10366 ( .A1(n9008), .A2(n9007), .ZN(n9014) );
  XNOR2_X1 U10367 ( .A(n9009), .B(keyinput21), .ZN(n9012) );
  XNOR2_X1 U10368 ( .A(n9010), .B(keyinput61), .ZN(n9011) );
  NOR2_X1 U10369 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  NAND4_X1 U10370 ( .A1(n9016), .A2(n9015), .A3(n9014), .A4(n9013), .ZN(n9078)
         );
  AOI22_X1 U10371 ( .A1(n9760), .A2(keyinput42), .B1(keyinput58), .B2(n4907), 
        .ZN(n9017) );
  OAI221_X1 U10372 ( .B1(n9760), .B2(keyinput42), .C1(n4907), .C2(keyinput58), 
        .A(n9017), .ZN(n9024) );
  AOI22_X1 U10373 ( .A1(n9020), .A2(keyinput38), .B1(n9019), .B2(keyinput24), 
        .ZN(n9018) );
  OAI221_X1 U10374 ( .B1(n9020), .B2(keyinput38), .C1(n9019), .C2(keyinput24), 
        .A(n9018), .ZN(n9023) );
  INV_X1 U10375 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n9098) );
  AOI22_X1 U10376 ( .A1(n9424), .A2(keyinput27), .B1(n9098), .B2(keyinput0), 
        .ZN(n9021) );
  OAI221_X1 U10377 ( .B1(n9424), .B2(keyinput27), .C1(n9098), .C2(keyinput0), 
        .A(n9021), .ZN(n9022) );
  NOR3_X1 U10378 ( .A1(n9024), .A2(n9023), .A3(n9022), .ZN(n9042) );
  INV_X1 U10379 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10100) );
  INV_X1 U10380 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9026) );
  AOI22_X1 U10381 ( .A1(n10100), .A2(keyinput34), .B1(n9026), .B2(keyinput33), 
        .ZN(n9025) );
  OAI221_X1 U10382 ( .B1(n10100), .B2(keyinput34), .C1(n9026), .C2(keyinput33), 
        .A(n9025), .ZN(n9033) );
  INV_X1 U10383 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9607) );
  XNOR2_X1 U10384 ( .A(n9607), .B(keyinput60), .ZN(n9032) );
  XNOR2_X1 U10385 ( .A(keyinput39), .B(P2_IR_REG_29__SCAN_IN), .ZN(n9030) );
  XNOR2_X1 U10386 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput26), .ZN(n9029) );
  XNOR2_X1 U10387 ( .A(keyinput63), .B(P1_REG0_REG_4__SCAN_IN), .ZN(n9028) );
  XNOR2_X1 U10388 ( .A(keyinput32), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n9027) );
  NAND4_X1 U10389 ( .A1(n9030), .A2(n9029), .A3(n9028), .A4(n9027), .ZN(n9031)
         );
  NOR3_X1 U10390 ( .A1(n9033), .A2(n9032), .A3(n9031), .ZN(n9041) );
  AOI22_X1 U10391 ( .A1(n9035), .A2(keyinput54), .B1(keyinput15), .B2(n7748), 
        .ZN(n9034) );
  OAI221_X1 U10392 ( .B1(n9035), .B2(keyinput54), .C1(n7748), .C2(keyinput15), 
        .A(n9034), .ZN(n9039) );
  INV_X1 U10393 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U10394 ( .A1(n10027), .A2(keyinput12), .B1(n9037), .B2(keyinput7), 
        .ZN(n9036) );
  OAI221_X1 U10395 ( .B1(n10027), .B2(keyinput12), .C1(n9037), .C2(keyinput7), 
        .A(n9036), .ZN(n9038) );
  NOR2_X1 U10396 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  NAND3_X1 U10397 ( .A1(n9042), .A2(n9041), .A3(n9040), .ZN(n9077) );
  AOI22_X1 U10398 ( .A1(n9044), .A2(keyinput16), .B1(keyinput17), .B2(n9095), 
        .ZN(n9043) );
  OAI221_X1 U10399 ( .B1(n9044), .B2(keyinput16), .C1(n9095), .C2(keyinput17), 
        .A(n9043), .ZN(n9050) );
  XNOR2_X1 U10400 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput19), .ZN(n9048) );
  XNOR2_X1 U10401 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(keyinput8), .ZN(n9047) );
  XNOR2_X1 U10402 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput45), .ZN(n9046) );
  XNOR2_X1 U10403 ( .A(SI_29_), .B(keyinput4), .ZN(n9045) );
  NAND4_X1 U10404 ( .A1(n9048), .A2(n9047), .A3(n9046), .A4(n9045), .ZN(n9049)
         );
  NOR2_X1 U10405 ( .A1(n9050), .A2(n9049), .ZN(n9075) );
  XNOR2_X1 U10406 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput11), .ZN(n9054) );
  XNOR2_X1 U10407 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput48), .ZN(n9053) );
  XNOR2_X1 U10408 ( .A(SI_17_), .B(keyinput52), .ZN(n9052) );
  XNOR2_X1 U10409 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput3), .ZN(n9051) );
  NAND4_X1 U10410 ( .A1(n9054), .A2(n9053), .A3(n9052), .A4(n9051), .ZN(n9060)
         );
  XNOR2_X1 U10411 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput31), .ZN(n9058) );
  XNOR2_X1 U10412 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput50), .ZN(n9057) );
  XNOR2_X1 U10413 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput5), .ZN(n9056) );
  XNOR2_X1 U10414 ( .A(P1_REG1_REG_19__SCAN_IN), .B(keyinput49), .ZN(n9055) );
  NAND4_X1 U10415 ( .A1(n9058), .A2(n9057), .A3(n9056), .A4(n9055), .ZN(n9059)
         );
  NOR2_X1 U10416 ( .A1(n9060), .A2(n9059), .ZN(n9074) );
  INV_X1 U10417 ( .A(keyinput62), .ZN(n9061) );
  XNOR2_X1 U10418 ( .A(n9762), .B(n9061), .ZN(n9073) );
  XNOR2_X1 U10419 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput2), .ZN(n9065) );
  XNOR2_X1 U10420 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput18), .ZN(n9064) );
  XNOR2_X1 U10421 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput23), .ZN(n9063) );
  XNOR2_X1 U10422 ( .A(SI_0_), .B(keyinput28), .ZN(n9062) );
  NAND4_X1 U10423 ( .A1(n9065), .A2(n9064), .A3(n9063), .A4(n9062), .ZN(n9071)
         );
  XNOR2_X1 U10424 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput9), .ZN(n9069) );
  XNOR2_X1 U10425 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput41), .ZN(n9068) );
  XNOR2_X1 U10426 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput51), .ZN(n9067) );
  XNOR2_X1 U10427 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput53), .ZN(n9066) );
  NAND4_X1 U10428 ( .A1(n9069), .A2(n9068), .A3(n9067), .A4(n9066), .ZN(n9070)
         );
  NOR2_X1 U10429 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  NAND4_X1 U10430 ( .A1(n9075), .A2(n9074), .A3(n9073), .A4(n9072), .ZN(n9076)
         );
  NOR3_X1 U10431 ( .A1(n9078), .A2(n9077), .A3(n9076), .ZN(n9090) );
  INV_X1 U10432 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9567) );
  AOI22_X1 U10433 ( .A1(n4918), .A2(keyinput44), .B1(keyinput55), .B2(n9567), 
        .ZN(n9079) );
  OAI221_X1 U10434 ( .B1(n4918), .B2(keyinput44), .C1(n9567), .C2(keyinput55), 
        .A(n9079), .ZN(n9088) );
  INV_X1 U10435 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9615) );
  AOI22_X1 U10436 ( .A1(n9081), .A2(keyinput57), .B1(keyinput47), .B2(n9615), 
        .ZN(n9080) );
  OAI221_X1 U10437 ( .B1(n9081), .B2(keyinput57), .C1(n9615), .C2(keyinput47), 
        .A(n9080), .ZN(n9087) );
  AOI22_X1 U10438 ( .A1(n9083), .A2(keyinput1), .B1(n6190), .B2(keyinput40), 
        .ZN(n9082) );
  OAI221_X1 U10439 ( .B1(n9083), .B2(keyinput1), .C1(n6190), .C2(keyinput40), 
        .A(n9082), .ZN(n9086) );
  AOI22_X1 U10440 ( .A1(n9759), .A2(keyinput35), .B1(n9761), .B2(keyinput56), 
        .ZN(n9084) );
  OAI221_X1 U10441 ( .B1(n9759), .B2(keyinput35), .C1(n9761), .C2(keyinput56), 
        .A(n9084), .ZN(n9085) );
  NOR4_X1 U10442 ( .A1(n9088), .A2(n9087), .A3(n9086), .A4(n9085), .ZN(n9089)
         );
  NAND2_X1 U10443 ( .A1(n9090), .A2(n9089), .ZN(n9130) );
  NAND4_X1 U10444 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .A3(P2_IR_REG_0__SCAN_IN), .A4(P1_REG1_REG_30__SCAN_IN), .ZN(n9094) );
  NAND4_X1 U10445 ( .A1(P1_REG0_REG_12__SCAN_IN), .A2(P1_REG0_REG_4__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .A4(P2_ADDR_REG_18__SCAN_IN), .ZN(n9093)
         );
  NAND4_X1 U10446 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(P2_REG0_REG_3__SCAN_IN), .A4(P2_REG2_REG_31__SCAN_IN), .ZN(n9092)
         );
  NAND4_X1 U10447 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_23__SCAN_IN), .A4(P2_REG0_REG_8__SCAN_IN), .ZN(n9091)
         );
  NOR4_X1 U10448 ( .A1(n9094), .A2(n9093), .A3(n9092), .A4(n9091), .ZN(n9128)
         );
  NAND4_X1 U10449 ( .A1(n9098), .A2(n9097), .A3(n9096), .A4(n9095), .ZN(n9101)
         );
  INV_X1 U10450 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9099) );
  NAND4_X1 U10451 ( .A1(n8993), .A2(n9099), .A3(P1_IR_REG_17__SCAN_IN), .A4(
        P1_IR_REG_26__SCAN_IN), .ZN(n9100) );
  NOR2_X1 U10452 ( .A1(n9101), .A2(n9100), .ZN(n9115) );
  NAND4_X1 U10453 ( .A1(SI_17_), .A2(n9104), .A3(n9103), .A4(n9102), .ZN(n9106) );
  NAND4_X1 U10454 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_RD_REG_SCAN_IN), .A3(
        P1_B_REG_SCAN_IN), .A4(P1_D_REG_1__SCAN_IN), .ZN(n9105) );
  NOR2_X1 U10455 ( .A1(n9106), .A2(n9105), .ZN(n9108) );
  NOR4_X1 U10456 ( .A1(P1_REG0_REG_20__SCAN_IN), .A2(P1_REG1_REG_19__SCAN_IN), 
        .A3(P1_REG2_REG_1__SCAN_IN), .A4(P2_REG2_REG_7__SCAN_IN), .ZN(n9107)
         );
  NAND4_X1 U10457 ( .A1(n9109), .A2(n9108), .A3(n10094), .A4(n9107), .ZN(n9113) );
  INV_X1 U10458 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9110) );
  NAND2_X1 U10459 ( .A1(n9111), .A2(n9110), .ZN(n9112) );
  NOR2_X1 U10460 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  NAND4_X1 U10461 ( .A1(n9115), .A2(P1_ADDR_REG_3__SCAN_IN), .A3(n9114), .A4(
        n9923), .ZN(n9117) );
  NAND4_X1 U10462 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(n9761), .ZN(n9116) );
  NOR2_X1 U10463 ( .A1(n9117), .A2(n9116), .ZN(n9125) );
  NAND4_X1 U10464 ( .A1(SI_0_), .A2(SI_31_), .A3(n9118), .A4(n4918), .ZN(n9122) );
  NAND4_X1 U10465 ( .A1(n9026), .A2(n9119), .A3(P1_IR_REG_23__SCAN_IN), .A4(
        P1_IR_REG_19__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U10466 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), 
        .ZN(n9120) );
  NOR3_X1 U10467 ( .A1(n9122), .A2(n9121), .A3(n9120), .ZN(n9123) );
  AND4_X1 U10468 ( .A1(n9125), .A2(n10098), .A3(n9124), .A4(n9123), .ZN(n9127)
         );
  NOR4_X1 U10469 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .A3(
        P2_REG0_REG_24__SCAN_IN), .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n9126) );
  NAND3_X1 U10470 ( .A1(n9128), .A2(n9127), .A3(n9126), .ZN(n9129) );
  XNOR2_X1 U10471 ( .A(n9130), .B(n9129), .ZN(n9131) );
  XNOR2_X1 U10472 ( .A(n9132), .B(n9131), .ZN(P1_U3263) );
  OAI211_X1 U10473 ( .C1(n9500), .C2(n9173), .A(n9750), .B(n9133), .ZN(n9423)
         );
  NOR2_X1 U10474 ( .A1(n9500), .A2(n9744), .ZN(n9134) );
  AOI211_X1 U10475 ( .C1(n9758), .C2(P1_REG2_REG_30__SCAN_IN), .A(n9135), .B(
        n9134), .ZN(n9136) );
  OAI21_X1 U10476 ( .B1(n9413), .B2(n9423), .A(n9136), .ZN(P1_U3264) );
  NAND2_X1 U10477 ( .A1(n4457), .A2(n9141), .ZN(n9142) );
  OR2_X1 U10478 ( .A1(n9392), .A2(n9144), .ZN(n9143) );
  NAND2_X1 U10479 ( .A1(n9385), .A2(n9143), .ZN(n9146) );
  NAND2_X1 U10480 ( .A1(n9392), .A2(n9144), .ZN(n9145) );
  OR2_X1 U10481 ( .A1(n9377), .A2(n9147), .ZN(n9148) );
  NAND2_X1 U10482 ( .A1(n9356), .A2(n9150), .ZN(n9151) );
  OR2_X1 U10483 ( .A1(n9471), .A2(n9153), .ZN(n9154) );
  NAND2_X1 U10484 ( .A1(n9323), .A2(n9155), .ZN(n9156) );
  NAND2_X1 U10485 ( .A1(n9305), .A2(n9299), .ZN(n9159) );
  NAND2_X1 U10486 ( .A1(n9307), .A2(n9157), .ZN(n9158) );
  OR2_X1 U10487 ( .A1(n9291), .A2(n9160), .ZN(n9161) );
  NOR2_X1 U10488 ( .A1(n9275), .A2(n9162), .ZN(n9164) );
  NAND2_X1 U10489 ( .A1(n9275), .A2(n9162), .ZN(n9163) );
  AND2_X1 U10490 ( .A1(n9257), .A2(n9165), .ZN(n9166) );
  NAND2_X1 U10491 ( .A1(n9212), .A2(n9200), .ZN(n9171) );
  INV_X1 U10492 ( .A(n9214), .ZN(n9174) );
  AOI211_X1 U10493 ( .C1(n9428), .C2(n9174), .A(n9403), .B(n9173), .ZN(n9427)
         );
  INV_X1 U10494 ( .A(n9175), .ZN(n9176) );
  AOI22_X1 U10495 ( .A1(n9758), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9335), .B2(
        n9176), .ZN(n9177) );
  OAI21_X1 U10496 ( .B1(n9178), .B2(n9744), .A(n9177), .ZN(n9202) );
  NAND2_X1 U10497 ( .A1(n9340), .A2(n9341), .ZN(n9339) );
  INV_X1 U10498 ( .A(n9265), .ZN(n9183) );
  NOR2_X1 U10499 ( .A1(n9266), .A2(n9183), .ZN(n9184) );
  NAND2_X1 U10500 ( .A1(n9268), .A2(n9185), .ZN(n9251) );
  INV_X1 U10501 ( .A(n9191), .ZN(n9192) );
  OAI21_X1 U10502 ( .B1(n4305), .B2(n9415), .A(n9203), .ZN(P1_U3356) );
  NAND2_X1 U10503 ( .A1(n9204), .A2(n4614), .ZN(n9205) );
  NAND2_X1 U10504 ( .A1(n9206), .A2(n9205), .ZN(n9435) );
  XNOR2_X1 U10505 ( .A(n9208), .B(n9207), .ZN(n9210) );
  AOI21_X1 U10506 ( .B1(n9210), .B2(n9738), .A(n9209), .ZN(n9433) );
  OAI21_X1 U10507 ( .B1(n9741), .B2(n9211), .A(n9433), .ZN(n9218) );
  AND2_X1 U10508 ( .A1(n9226), .A2(n9212), .ZN(n9213) );
  NOR2_X1 U10509 ( .A1(n9432), .A2(n9413), .ZN(n9217) );
  OAI22_X1 U10510 ( .A1(n9503), .A2(n9744), .B1(n9215), .B2(n9394), .ZN(n9216)
         );
  AOI211_X1 U10511 ( .C1(n9218), .C2(n9394), .A(n9217), .B(n9216), .ZN(n9219)
         );
  OAI21_X1 U10512 ( .B1(n9435), .B2(n9415), .A(n9219), .ZN(P1_U3265) );
  XNOR2_X1 U10513 ( .A(n9220), .B(n9221), .ZN(n9438) );
  INV_X1 U10514 ( .A(n9438), .ZN(n9234) );
  XNOR2_X1 U10515 ( .A(n9222), .B(n9221), .ZN(n9223) );
  NAND2_X1 U10516 ( .A1(n9223), .A2(n9738), .ZN(n9225) );
  NAND2_X1 U10517 ( .A1(n9225), .A2(n9224), .ZN(n9436) );
  INV_X1 U10518 ( .A(n9226), .ZN(n9227) );
  AOI211_X1 U10519 ( .C1(n9228), .C2(n4659), .A(n9403), .B(n9227), .ZN(n9437)
         );
  NAND2_X1 U10520 ( .A1(n9437), .A2(n9754), .ZN(n9231) );
  AOI22_X1 U10521 ( .A1(n9758), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9335), .B2(
        n9229), .ZN(n9230) );
  OAI211_X1 U10522 ( .C1(n9507), .C2(n9744), .A(n9231), .B(n9230), .ZN(n9232)
         );
  AOI21_X1 U10523 ( .B1(n9436), .B2(n9394), .A(n9232), .ZN(n9233) );
  OAI21_X1 U10524 ( .B1(n9234), .B2(n9415), .A(n9233), .ZN(P1_U3266) );
  XOR2_X1 U10525 ( .A(n9235), .B(n9236), .Z(n9442) );
  INV_X1 U10526 ( .A(n9442), .ZN(n9247) );
  XNOR2_X1 U10527 ( .A(n9237), .B(n9236), .ZN(n9239) );
  OAI21_X1 U10528 ( .B1(n9239), .B2(n9706), .A(n9238), .ZN(n9440) );
  AOI211_X1 U10529 ( .C1(n9241), .C2(n9255), .A(n9403), .B(n9240), .ZN(n9441)
         );
  NAND2_X1 U10530 ( .A1(n9441), .A2(n9754), .ZN(n9244) );
  AOI22_X1 U10531 ( .A1(n9242), .A2(n9335), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9758), .ZN(n9243) );
  OAI211_X1 U10532 ( .C1(n4657), .C2(n9744), .A(n9244), .B(n9243), .ZN(n9245)
         );
  AOI21_X1 U10533 ( .B1(n9440), .B2(n9394), .A(n9245), .ZN(n9246) );
  OAI21_X1 U10534 ( .B1(n9247), .B2(n9415), .A(n9246), .ZN(P1_U3267) );
  XNOR2_X1 U10535 ( .A(n9248), .B(n9249), .ZN(n9447) );
  INV_X1 U10536 ( .A(n9447), .ZN(n9263) );
  INV_X1 U10537 ( .A(n9249), .ZN(n9250) );
  XNOR2_X1 U10538 ( .A(n9251), .B(n9250), .ZN(n9252) );
  NAND2_X1 U10539 ( .A1(n9252), .A2(n9738), .ZN(n9254) );
  NAND2_X1 U10540 ( .A1(n9254), .A2(n9253), .ZN(n9445) );
  INV_X1 U10541 ( .A(n9255), .ZN(n9256) );
  AOI211_X1 U10542 ( .C1(n9257), .C2(n9272), .A(n9403), .B(n9256), .ZN(n9446)
         );
  NAND2_X1 U10543 ( .A1(n9446), .A2(n9754), .ZN(n9260) );
  AOI22_X1 U10544 ( .A1(n9258), .A2(n9335), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9758), .ZN(n9259) );
  OAI211_X1 U10545 ( .C1(n9514), .C2(n9744), .A(n9260), .B(n9259), .ZN(n9261)
         );
  AOI21_X1 U10546 ( .B1(n9445), .B2(n9394), .A(n9261), .ZN(n9262) );
  OAI21_X1 U10547 ( .B1(n9263), .B2(n9415), .A(n9262), .ZN(P1_U3268) );
  XNOR2_X1 U10548 ( .A(n9264), .B(n9266), .ZN(n9452) );
  INV_X1 U10549 ( .A(n9452), .ZN(n9281) );
  NAND2_X1 U10550 ( .A1(n9283), .A2(n9265), .ZN(n9267) );
  NAND2_X1 U10551 ( .A1(n9267), .A2(n9266), .ZN(n9269) );
  NAND3_X1 U10552 ( .A1(n9269), .A2(n9738), .A3(n9268), .ZN(n9271) );
  NAND2_X1 U10553 ( .A1(n9271), .A2(n9270), .ZN(n9450) );
  INV_X1 U10554 ( .A(n9289), .ZN(n9274) );
  INV_X1 U10555 ( .A(n9272), .ZN(n9273) );
  AOI211_X1 U10556 ( .C1(n9275), .C2(n9274), .A(n9403), .B(n9273), .ZN(n9451)
         );
  NAND2_X1 U10557 ( .A1(n9451), .A2(n9754), .ZN(n9278) );
  AOI22_X1 U10558 ( .A1(n9276), .A2(n9335), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9758), .ZN(n9277) );
  OAI211_X1 U10559 ( .C1(n9518), .C2(n9744), .A(n9278), .B(n9277), .ZN(n9279)
         );
  AOI21_X1 U10560 ( .B1(n9450), .B2(n9394), .A(n9279), .ZN(n9280) );
  OAI21_X1 U10561 ( .B1(n9281), .B2(n9415), .A(n9280), .ZN(P1_U3269) );
  INV_X1 U10562 ( .A(n9282), .ZN(n9288) );
  OAI21_X1 U10563 ( .B1(n9295), .B2(n9284), .A(n9283), .ZN(n9285) );
  NAND2_X1 U10564 ( .A1(n9285), .A2(n9738), .ZN(n9287) );
  NAND2_X1 U10565 ( .A1(n9287), .A2(n9286), .ZN(n9455) );
  AOI21_X1 U10566 ( .B1(n9288), .B2(n9335), .A(n9455), .ZN(n9298) );
  INV_X1 U10567 ( .A(n9306), .ZN(n9290) );
  AOI211_X1 U10568 ( .C1(n9291), .C2(n9290), .A(n9403), .B(n9289), .ZN(n9456)
         );
  OAI22_X1 U10569 ( .A1(n9522), .A2(n9744), .B1(n9292), .B2(n9394), .ZN(n9293)
         );
  AOI21_X1 U10570 ( .B1(n9456), .B2(n9754), .A(n9293), .ZN(n9297) );
  XNOR2_X1 U10571 ( .A(n9294), .B(n9295), .ZN(n9457) );
  NAND2_X1 U10572 ( .A1(n9457), .A2(n9755), .ZN(n9296) );
  OAI211_X1 U10573 ( .C1(n9298), .C2(n9758), .A(n9297), .B(n9296), .ZN(
        P1_U3270) );
  XNOR2_X1 U10574 ( .A(n9300), .B(n9299), .ZN(n9303) );
  INV_X1 U10575 ( .A(n9301), .ZN(n9302) );
  OAI21_X1 U10576 ( .B1(n9303), .B2(n9706), .A(n9302), .ZN(n9460) );
  INV_X1 U10577 ( .A(n9460), .ZN(n9313) );
  XNOR2_X1 U10578 ( .A(n9305), .B(n9304), .ZN(n9462) );
  NAND2_X1 U10579 ( .A1(n9462), .A2(n9755), .ZN(n9312) );
  AOI211_X1 U10580 ( .C1(n9307), .C2(n9321), .A(n9403), .B(n9306), .ZN(n9461)
         );
  INV_X1 U10581 ( .A(n9307), .ZN(n9526) );
  NOR2_X1 U10582 ( .A1(n9526), .A2(n9744), .ZN(n9310) );
  OAI22_X1 U10583 ( .A1(n9394), .A2(n9026), .B1(n9308), .B2(n9741), .ZN(n9309)
         );
  AOI211_X1 U10584 ( .C1(n9461), .C2(n9754), .A(n9310), .B(n9309), .ZN(n9311)
         );
  OAI211_X1 U10585 ( .C1(n9758), .C2(n9313), .A(n9312), .B(n9311), .ZN(
        P1_U3271) );
  XOR2_X1 U10586 ( .A(n9314), .B(n9317), .Z(n9467) );
  INV_X1 U10587 ( .A(n9467), .ZN(n9329) );
  OAI21_X1 U10588 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9318) );
  NAND2_X1 U10589 ( .A1(n9318), .A2(n9738), .ZN(n9320) );
  NAND2_X1 U10590 ( .A1(n9320), .A2(n9319), .ZN(n9465) );
  INV_X1 U10591 ( .A(n9321), .ZN(n9322) );
  AOI211_X1 U10592 ( .C1(n9323), .C2(n9331), .A(n9403), .B(n9322), .ZN(n9466)
         );
  NAND2_X1 U10593 ( .A1(n9466), .A2(n9754), .ZN(n9326) );
  AOI22_X1 U10594 ( .A1(n9758), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9324), .B2(
        n9335), .ZN(n9325) );
  OAI211_X1 U10595 ( .C1(n4650), .C2(n9744), .A(n9326), .B(n9325), .ZN(n9327)
         );
  AOI21_X1 U10596 ( .B1(n9465), .B2(n9394), .A(n9327), .ZN(n9328) );
  OAI21_X1 U10597 ( .B1(n9329), .B2(n9415), .A(n9328), .ZN(P1_U3272) );
  XOR2_X1 U10598 ( .A(n9330), .B(n9341), .Z(n9474) );
  INV_X1 U10599 ( .A(n9354), .ZN(n9333) );
  INV_X1 U10600 ( .A(n9331), .ZN(n9332) );
  AOI211_X1 U10601 ( .C1(n9471), .C2(n9333), .A(n9403), .B(n9332), .ZN(n9470)
         );
  INV_X1 U10602 ( .A(n9334), .ZN(n9336) );
  AOI22_X1 U10603 ( .A1(n9758), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9336), .B2(
        n9335), .ZN(n9337) );
  OAI21_X1 U10604 ( .B1(n9338), .B2(n9744), .A(n9337), .ZN(n9345) );
  OAI21_X1 U10605 ( .B1(n9341), .B2(n9340), .A(n9339), .ZN(n9343) );
  AOI21_X1 U10606 ( .B1(n9343), .B2(n9738), .A(n9342), .ZN(n9473) );
  NOR2_X1 U10607 ( .A1(n9473), .A2(n9758), .ZN(n9344) );
  AOI211_X1 U10608 ( .C1(n9470), .C2(n9754), .A(n9345), .B(n9344), .ZN(n9346)
         );
  OAI21_X1 U10609 ( .B1(n9415), .B2(n9474), .A(n9346), .ZN(P1_U3273) );
  XNOR2_X1 U10610 ( .A(n9347), .B(n9353), .ZN(n9348) );
  NAND2_X1 U10611 ( .A1(n9348), .A2(n9738), .ZN(n9351) );
  INV_X1 U10612 ( .A(n9349), .ZN(n9350) );
  NAND2_X1 U10613 ( .A1(n9351), .A2(n9350), .ZN(n9475) );
  INV_X1 U10614 ( .A(n9475), .ZN(n9363) );
  XOR2_X1 U10615 ( .A(n9352), .B(n9353), .Z(n9477) );
  NAND2_X1 U10616 ( .A1(n9477), .A2(n9755), .ZN(n9362) );
  INV_X1 U10617 ( .A(n9375), .ZN(n9355) );
  AOI211_X1 U10618 ( .C1(n9356), .C2(n9355), .A(n9403), .B(n9354), .ZN(n9476)
         );
  NOR2_X1 U10619 ( .A1(n9534), .A2(n9744), .ZN(n9360) );
  OAI22_X1 U10620 ( .A1(n9394), .A2(n9358), .B1(n9357), .B2(n9741), .ZN(n9359)
         );
  AOI211_X1 U10621 ( .C1(n9476), .C2(n9754), .A(n9360), .B(n9359), .ZN(n9361)
         );
  OAI211_X1 U10622 ( .C1(n9758), .C2(n9363), .A(n9362), .B(n9361), .ZN(
        P1_U3274) );
  NAND2_X1 U10623 ( .A1(n9365), .A2(n9364), .ZN(n9374) );
  INV_X1 U10624 ( .A(n9366), .ZN(n9368) );
  OAI21_X1 U10625 ( .B1(n9387), .B2(n9368), .A(n9367), .ZN(n9369) );
  XOR2_X1 U10626 ( .A(n9374), .B(n9369), .Z(n9372) );
  INV_X1 U10627 ( .A(n9370), .ZN(n9371) );
  OAI21_X1 U10628 ( .B1(n9372), .B2(n9706), .A(n9371), .ZN(n9480) );
  INV_X1 U10629 ( .A(n9480), .ZN(n9384) );
  XOR2_X1 U10630 ( .A(n9374), .B(n4301), .Z(n9482) );
  NAND2_X1 U10631 ( .A1(n9482), .A2(n9755), .ZN(n9383) );
  INV_X1 U10632 ( .A(n9391), .ZN(n9376) );
  AOI211_X1 U10633 ( .C1(n9377), .C2(n9376), .A(n9403), .B(n9375), .ZN(n9481)
         );
  NOR2_X1 U10634 ( .A1(n9538), .A2(n9744), .ZN(n9381) );
  OAI22_X1 U10635 ( .A1(n9394), .A2(n9379), .B1(n9378), .B2(n9741), .ZN(n9380)
         );
  AOI211_X1 U10636 ( .C1(n9481), .C2(n9754), .A(n9381), .B(n9380), .ZN(n9382)
         );
  OAI211_X1 U10637 ( .C1(n9758), .C2(n9384), .A(n9383), .B(n9382), .ZN(
        P1_U3275) );
  XNOR2_X1 U10638 ( .A(n4304), .B(n9386), .ZN(n9487) );
  INV_X1 U10639 ( .A(n9487), .ZN(n9399) );
  XOR2_X1 U10640 ( .A(n9387), .B(n9386), .Z(n9390) );
  INV_X1 U10641 ( .A(n9388), .ZN(n9389) );
  OAI21_X1 U10642 ( .B1(n9390), .B2(n9706), .A(n9389), .ZN(n9485) );
  NAND2_X1 U10643 ( .A1(n9485), .A2(n9394), .ZN(n9398) );
  AOI211_X1 U10644 ( .C1(n9392), .C2(n9405), .A(n9403), .B(n9391), .ZN(n9486)
         );
  NOR2_X1 U10645 ( .A1(n9543), .A2(n9744), .ZN(n9396) );
  OAI22_X1 U10646 ( .A1(n9394), .A2(n5985), .B1(n9393), .B2(n9741), .ZN(n9395)
         );
  AOI211_X1 U10647 ( .C1(n9486), .C2(n9754), .A(n9396), .B(n9395), .ZN(n9397)
         );
  OAI211_X1 U10648 ( .C1(n9399), .C2(n9415), .A(n9398), .B(n9397), .ZN(
        P1_U3276) );
  XOR2_X1 U10649 ( .A(n9400), .B(n9414), .Z(n9402) );
  OAI21_X1 U10650 ( .B1(n9402), .B2(n9706), .A(n9401), .ZN(n9635) );
  AOI21_X1 U10651 ( .B1(n9404), .B2(n4457), .A(n9403), .ZN(n9406) );
  NAND2_X1 U10652 ( .A1(n9406), .A2(n9405), .ZN(n9634) );
  NAND2_X1 U10653 ( .A1(n9758), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9407) );
  OAI21_X1 U10654 ( .B1(n9741), .B2(n9408), .A(n9407), .ZN(n9409) );
  AOI21_X1 U10655 ( .B1(n4457), .B2(n9410), .A(n9409), .ZN(n9412) );
  OAI21_X1 U10656 ( .B1(n9634), .B2(n9413), .A(n9412), .ZN(n9417) );
  AND2_X1 U10657 ( .A1(n4402), .A2(n9414), .ZN(n9633) );
  NOR3_X1 U10658 ( .A1(n9140), .A2(n9633), .A3(n9415), .ZN(n9416) );
  AOI211_X1 U10659 ( .C1(n9394), .C2(n9635), .A(n9417), .B(n9416), .ZN(n9418)
         );
  INV_X1 U10660 ( .A(n9418), .ZN(P1_U3277) );
  INV_X1 U10661 ( .A(n9853), .ZN(n9492) );
  NAND2_X1 U10662 ( .A1(n9879), .A2(n9492), .ZN(n9489) );
  AND2_X1 U10663 ( .A1(n9419), .A2(n9422), .ZN(n9493) );
  MUX2_X1 U10664 ( .A(n9420), .B(n9493), .S(n9879), .Z(n9421) );
  OAI21_X1 U10665 ( .B1(n9496), .B2(n9489), .A(n9421), .ZN(P1_U3553) );
  AND2_X1 U10666 ( .A1(n9423), .A2(n9422), .ZN(n9497) );
  MUX2_X1 U10667 ( .A(n9424), .B(n9497), .S(n9879), .Z(n9425) );
  OAI21_X1 U10668 ( .B1(n9500), .B2(n9489), .A(n9425), .ZN(P1_U3552) );
  AOI21_X1 U10669 ( .B1(n9492), .B2(n9428), .A(n9427), .ZN(n9429) );
  OAI21_X1 U10670 ( .B1(n9431), .B2(n9632), .A(n9430), .ZN(n9501) );
  MUX2_X1 U10671 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9501), .S(n9879), .Z(
        P1_U3551) );
  INV_X1 U10672 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9439) );
  AOI211_X1 U10673 ( .C1(n9438), .C2(n9850), .A(n9437), .B(n9436), .ZN(n9504)
         );
  INV_X1 U10674 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9443) );
  AOI211_X1 U10675 ( .C1(n9442), .C2(n9850), .A(n9441), .B(n9440), .ZN(n9508)
         );
  MUX2_X1 U10676 ( .A(n9443), .B(n9508), .S(n9879), .Z(n9444) );
  OAI21_X1 U10677 ( .B1(n4657), .B2(n9489), .A(n9444), .ZN(P1_U3548) );
  AOI211_X1 U10678 ( .C1(n9447), .C2(n9850), .A(n9446), .B(n9445), .ZN(n9512)
         );
  INV_X1 U10679 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9448) );
  MUX2_X1 U10680 ( .A(n9512), .B(n9448), .S(n9877), .Z(n9449) );
  OAI21_X1 U10681 ( .B1(n9514), .B2(n9489), .A(n9449), .ZN(P1_U3547) );
  INV_X1 U10682 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9453) );
  AOI211_X1 U10683 ( .C1(n9452), .C2(n9850), .A(n9451), .B(n9450), .ZN(n9515)
         );
  MUX2_X1 U10684 ( .A(n9453), .B(n9515), .S(n9879), .Z(n9454) );
  OAI21_X1 U10685 ( .B1(n9518), .B2(n9489), .A(n9454), .ZN(P1_U3546) );
  INV_X1 U10686 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9458) );
  AOI211_X1 U10687 ( .C1(n9457), .C2(n9850), .A(n9456), .B(n9455), .ZN(n9519)
         );
  MUX2_X1 U10688 ( .A(n9458), .B(n9519), .S(n9879), .Z(n9459) );
  OAI21_X1 U10689 ( .B1(n9522), .B2(n9489), .A(n9459), .ZN(P1_U3545) );
  AOI211_X1 U10690 ( .C1(n9462), .C2(n9850), .A(n9461), .B(n9460), .ZN(n9523)
         );
  MUX2_X1 U10691 ( .A(n9463), .B(n9523), .S(n9879), .Z(n9464) );
  OAI21_X1 U10692 ( .B1(n9526), .B2(n9489), .A(n9464), .ZN(P1_U3544) );
  AOI211_X1 U10693 ( .C1(n9467), .C2(n9850), .A(n9466), .B(n9465), .ZN(n9527)
         );
  MUX2_X1 U10694 ( .A(n9468), .B(n9527), .S(n9879), .Z(n9469) );
  OAI21_X1 U10695 ( .B1(n4650), .B2(n9489), .A(n9469), .ZN(P1_U3543) );
  AOI21_X1 U10696 ( .B1(n9492), .B2(n9471), .A(n9470), .ZN(n9472) );
  OAI211_X1 U10697 ( .C1(n9474), .C2(n9632), .A(n9473), .B(n9472), .ZN(n9530)
         );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9530), .S(n9879), .Z(
        P1_U3542) );
  AOI211_X1 U10699 ( .C1(n9477), .C2(n9850), .A(n9476), .B(n9475), .ZN(n9531)
         );
  MUX2_X1 U10700 ( .A(n9478), .B(n9531), .S(n9879), .Z(n9479) );
  OAI21_X1 U10701 ( .B1(n9534), .B2(n9489), .A(n9479), .ZN(P1_U3541) );
  AOI211_X1 U10702 ( .C1(n9482), .C2(n9850), .A(n9481), .B(n9480), .ZN(n9535)
         );
  MUX2_X1 U10703 ( .A(n9483), .B(n9535), .S(n9879), .Z(n9484) );
  OAI21_X1 U10704 ( .B1(n9538), .B2(n9489), .A(n9484), .ZN(P1_U3540) );
  AOI211_X1 U10705 ( .C1(n9487), .C2(n9850), .A(n9486), .B(n9485), .ZN(n9539)
         );
  MUX2_X1 U10706 ( .A(n8938), .B(n9539), .S(n9879), .Z(n9488) );
  OAI21_X1 U10707 ( .B1(n9543), .B2(n9489), .A(n9488), .ZN(P1_U3539) );
  AND2_X2 U10708 ( .A1(n9491), .A2(n9490), .ZN(n9862) );
  NAND2_X1 U10709 ( .A1(n9862), .A2(n9492), .ZN(n9542) );
  INV_X1 U10710 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U10711 ( .A(n9494), .B(n9493), .S(n9862), .Z(n9495) );
  OAI21_X1 U10712 ( .B1(n9496), .B2(n9542), .A(n9495), .ZN(P1_U3521) );
  INV_X1 U10713 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9498) );
  MUX2_X1 U10714 ( .A(n9498), .B(n9497), .S(n9862), .Z(n9499) );
  OAI21_X1 U10715 ( .B1(n9500), .B2(n9542), .A(n9499), .ZN(P1_U3520) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9501), .S(n9862), .Z(
        P1_U3519) );
  MUX2_X1 U10717 ( .A(n9505), .B(n9504), .S(n9862), .Z(n9506) );
  MUX2_X1 U10718 ( .A(n9509), .B(n9508), .S(n9862), .Z(n9510) );
  OAI21_X1 U10719 ( .B1(n4657), .B2(n9542), .A(n9510), .ZN(P1_U3516) );
  MUX2_X1 U10720 ( .A(n9512), .B(n9511), .S(n9860), .Z(n9513) );
  OAI21_X1 U10721 ( .B1(n9514), .B2(n9542), .A(n9513), .ZN(P1_U3515) );
  MUX2_X1 U10722 ( .A(n9516), .B(n9515), .S(n9862), .Z(n9517) );
  OAI21_X1 U10723 ( .B1(n9518), .B2(n9542), .A(n9517), .ZN(P1_U3514) );
  INV_X1 U10724 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9520) );
  MUX2_X1 U10725 ( .A(n9520), .B(n9519), .S(n9862), .Z(n9521) );
  OAI21_X1 U10726 ( .B1(n9522), .B2(n9542), .A(n9521), .ZN(P1_U3513) );
  MUX2_X1 U10727 ( .A(n9524), .B(n9523), .S(n9862), .Z(n9525) );
  OAI21_X1 U10728 ( .B1(n9526), .B2(n9542), .A(n9525), .ZN(P1_U3512) );
  INV_X1 U10729 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U10730 ( .A(n9528), .B(n9527), .S(n9862), .Z(n9529) );
  OAI21_X1 U10731 ( .B1(n4650), .B2(n9542), .A(n9529), .ZN(P1_U3511) );
  MUX2_X1 U10732 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9530), .S(n9862), .Z(
        P1_U3510) );
  INV_X1 U10733 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9532) );
  MUX2_X1 U10734 ( .A(n9532), .B(n9531), .S(n9862), .Z(n9533) );
  OAI21_X1 U10735 ( .B1(n9534), .B2(n9542), .A(n9533), .ZN(P1_U3509) );
  MUX2_X1 U10736 ( .A(n9536), .B(n9535), .S(n9862), .Z(n9537) );
  OAI21_X1 U10737 ( .B1(n9538), .B2(n9542), .A(n9537), .ZN(P1_U3507) );
  INV_X1 U10738 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9540) );
  MUX2_X1 U10739 ( .A(n9540), .B(n9539), .S(n9862), .Z(n9541) );
  OAI21_X1 U10740 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(P1_U3504) );
  MUX2_X1 U10741 ( .A(P1_D_REG_0__SCAN_IN), .B(n9544), .S(n9763), .Z(P1_U3439)
         );
  INV_X1 U10742 ( .A(n9545), .ZN(n9548) );
  NAND3_X1 U10743 ( .A1(n9546), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9547) );
  OAI22_X1 U10744 ( .A1(n9548), .A2(n9547), .B1(n6846), .B2(n9554), .ZN(n9549)
         );
  INV_X1 U10745 ( .A(n9549), .ZN(n9550) );
  OAI21_X1 U10746 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(P1_U3324) );
  OAI222_X1 U10747 ( .A1(n9555), .A2(P1_U3086), .B1(n9554), .B2(n8721), .C1(
        n9553), .C2(n9562), .ZN(P1_U3326) );
  OAI222_X1 U10748 ( .A1(P1_U3086), .A2(n9563), .B1(n9562), .B2(n9561), .C1(
        n9560), .C2(n9559), .ZN(P1_U3329) );
  MUX2_X1 U10749 ( .A(n9564), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U10750 ( .A1(n9566), .A2(n9565), .ZN(n9618) );
  NOR2_X1 U10751 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9614) );
  NOR2_X1 U10752 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9610) );
  NOR2_X1 U10753 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9606) );
  NOR2_X1 U10754 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9602) );
  NOR2_X1 U10755 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9600) );
  NOR2_X1 U10756 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9598) );
  NOR2_X1 U10757 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9595) );
  NOR2_X1 U10758 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9591) );
  NOR2_X1 U10759 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9587) );
  NOR2_X1 U10760 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n9584) );
  NOR2_X1 U10761 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n9582) );
  NOR2_X1 U10762 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n9580) );
  NOR2_X1 U10763 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n9576) );
  NOR2_X1 U10764 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n9574) );
  NAND2_X1 U10765 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9571) );
  INV_X1 U10766 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n9904) );
  AOI22_X1 U10767 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n9904), .B2(n9567), .ZN(n10133) );
  NAND2_X1 U10768 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9569) );
  NOR2_X1 U10769 ( .A1(n10098), .A2(P1_ADDR_REG_1__SCAN_IN), .ZN(n10097) );
  AOI21_X1 U10770 ( .B1(n10098), .B2(P1_ADDR_REG_1__SCAN_IN), .A(
        P2_ADDR_REG_1__SCAN_IN), .ZN(n10093) );
  NOR2_X1 U10771 ( .A1(n10097), .A2(n10093), .ZN(n10131) );
  XOR2_X1 U10772 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10130) );
  NAND2_X1 U10773 ( .A1(n10131), .A2(n10130), .ZN(n9568) );
  NAND2_X1 U10774 ( .A1(n9569), .A2(n9568), .ZN(n10132) );
  NAND2_X1 U10775 ( .A1(n10133), .A2(n10132), .ZN(n9570) );
  NAND2_X1 U10776 ( .A1(n9571), .A2(n9570), .ZN(n10135) );
  AOI22_X1 U10777 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9572), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n9923), .ZN(n10134) );
  NOR2_X1 U10778 ( .A1(n10135), .A2(n10134), .ZN(n9573) );
  NOR2_X1 U10779 ( .A1(n9574), .A2(n9573), .ZN(n10123) );
  XNOR2_X1 U10780 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10122) );
  NOR2_X1 U10781 ( .A1(n10123), .A2(n10122), .ZN(n9575) );
  NOR2_X1 U10782 ( .A1(n9576), .A2(n9575), .ZN(n10121) );
  INV_X1 U10783 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9578) );
  INV_X1 U10784 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n9577) );
  AOI22_X1 U10785 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n9578), .B1(
        P1_ADDR_REG_6__SCAN_IN), .B2(n9577), .ZN(n10120) );
  NOR2_X1 U10786 ( .A1(n10121), .A2(n10120), .ZN(n9579) );
  NOR2_X1 U10787 ( .A1(n9580), .A2(n9579), .ZN(n10127) );
  XNOR2_X1 U10788 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10126) );
  NOR2_X1 U10789 ( .A1(n10127), .A2(n10126), .ZN(n9581) );
  NOR2_X1 U10790 ( .A1(n9582), .A2(n9581), .ZN(n10129) );
  XNOR2_X1 U10791 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10128) );
  NOR2_X1 U10792 ( .A1(n10129), .A2(n10128), .ZN(n9583) );
  NOR2_X1 U10793 ( .A1(n9584), .A2(n9583), .ZN(n10125) );
  AOI22_X1 U10794 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n6356), .B1(
        P1_ADDR_REG_9__SCAN_IN), .B2(n9585), .ZN(n10124) );
  NOR2_X1 U10795 ( .A1(n10125), .A2(n10124), .ZN(n9586) );
  NOR2_X1 U10796 ( .A1(n9587), .A2(n9586), .ZN(n10119) );
  INV_X1 U10797 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9589) );
  AOI22_X1 U10798 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(n9589), .B1(
        P1_ADDR_REG_10__SCAN_IN), .B2(n9588), .ZN(n10118) );
  NOR2_X1 U10799 ( .A1(n10119), .A2(n10118), .ZN(n9590) );
  NOR2_X1 U10800 ( .A1(n9591), .A2(n9590), .ZN(n10117) );
  INV_X1 U10801 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9593) );
  AOI22_X1 U10802 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n9593), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n9592), .ZN(n10116) );
  NOR2_X1 U10803 ( .A1(n10117), .A2(n10116), .ZN(n9594) );
  NOR2_X1 U10804 ( .A1(n9595), .A2(n9594), .ZN(n10115) );
  INV_X1 U10805 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9698) );
  AOI22_X1 U10806 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9698), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n9596), .ZN(n10114) );
  NOR2_X1 U10807 ( .A1(n10115), .A2(n10114), .ZN(n9597) );
  NOR2_X1 U10808 ( .A1(n9598), .A2(n9597), .ZN(n10113) );
  XNOR2_X1 U10809 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10112) );
  NOR2_X1 U10810 ( .A1(n10113), .A2(n10112), .ZN(n9599) );
  NOR2_X1 U10811 ( .A1(n9600), .A2(n9599), .ZN(n10111) );
  XNOR2_X1 U10812 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10110) );
  NOR2_X1 U10813 ( .A1(n10111), .A2(n10110), .ZN(n9601) );
  NOR2_X1 U10814 ( .A1(n9602), .A2(n9601), .ZN(n10109) );
  INV_X1 U10815 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9604) );
  AOI22_X1 U10816 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9604), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9603), .ZN(n10108) );
  NOR2_X1 U10817 ( .A1(n10109), .A2(n10108), .ZN(n9605) );
  NOR2_X1 U10818 ( .A1(n9606), .A2(n9605), .ZN(n10107) );
  INV_X1 U10819 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9608) );
  AOI22_X1 U10820 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9608), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n9607), .ZN(n10106) );
  NOR2_X1 U10821 ( .A1(n10107), .A2(n10106), .ZN(n9609) );
  NOR2_X1 U10822 ( .A1(n9610), .A2(n9609), .ZN(n10105) );
  INV_X1 U10823 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9612) );
  AOI22_X1 U10824 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9612), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9611), .ZN(n10104) );
  NOR2_X1 U10825 ( .A1(n10105), .A2(n10104), .ZN(n9613) );
  NOR2_X1 U10826 ( .A1(n9614), .A2(n9613), .ZN(n10102) );
  NOR2_X1 U10827 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10102), .ZN(n9616) );
  NAND2_X1 U10828 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10102), .ZN(n10101) );
  OAI21_X1 U10829 ( .B1(n9616), .B2(n9615), .A(n10101), .ZN(n9617) );
  XOR2_X1 U10830 ( .A(n9618), .B(n9617), .Z(ADD_1068_U4) );
  INV_X1 U10831 ( .A(n9619), .ZN(n9620) );
  OAI22_X1 U10832 ( .A1(n9621), .A2(n10061), .B1(n9620), .B2(n10054), .ZN(
        n9622) );
  NOR2_X1 U10833 ( .A1(n9623), .A2(n9622), .ZN(n9628) );
  AOI22_X1 U10834 ( .A1(n10092), .A2(n9628), .B1(n5263), .B2(n10090), .ZN(
        P2_U3473) );
  NOR2_X1 U10835 ( .A1(n9624), .A2(n10061), .ZN(n9626) );
  AOI211_X1 U10836 ( .C1(n10073), .C2(n9627), .A(n9626), .B(n9625), .ZN(n9630)
         );
  AOI22_X1 U10837 ( .A1(n10092), .A2(n9630), .B1(n5250), .B2(n10090), .ZN(
        P2_U3472) );
  INV_X1 U10838 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9629) );
  AOI22_X1 U10839 ( .A1(n10076), .A2(n9629), .B1(n9628), .B2(n10074), .ZN(
        P2_U3432) );
  INV_X1 U10840 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9631) );
  AOI22_X1 U10841 ( .A1(n10076), .A2(n9631), .B1(n9630), .B2(n10074), .ZN(
        P2_U3429) );
  NOR2_X1 U10842 ( .A1(n9633), .A2(n9632), .ZN(n9638) );
  OAI21_X1 U10843 ( .B1(n4652), .B2(n9853), .A(n9634), .ZN(n9636) );
  AOI211_X1 U10844 ( .C1(n9638), .C2(n4297), .A(n9636), .B(n9635), .ZN(n9645)
         );
  AOI22_X1 U10845 ( .A1(n9879), .A2(n9645), .B1(n8915), .B2(n9877), .ZN(
        P1_U3538) );
  OAI211_X1 U10846 ( .C1(n9641), .C2(n9853), .A(n9640), .B(n9639), .ZN(n9642)
         );
  AOI21_X1 U10847 ( .B1(n9643), .B2(n9850), .A(n9642), .ZN(n9647) );
  AOI22_X1 U10848 ( .A1(n9879), .A2(n9647), .B1(n5947), .B2(n9877), .ZN(
        P1_U3537) );
  INV_X1 U10849 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9644) );
  AOI22_X1 U10850 ( .A1(n9862), .A2(n9645), .B1(n9644), .B2(n9860), .ZN(
        P1_U3501) );
  INV_X1 U10851 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9646) );
  AOI22_X1 U10852 ( .A1(n9862), .A2(n9647), .B1(n9646), .B2(n9860), .ZN(
        P1_U3498) );
  XNOR2_X1 U10853 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI22_X1 U10854 ( .A1(n9648), .A2(n9660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5779), .ZN(n9655) );
  OAI211_X1 U10855 ( .C1(n9652), .C2(n9651), .A(n9650), .B(n9649), .ZN(n9653)
         );
  INV_X1 U10856 ( .A(n9653), .ZN(n9654) );
  AOI211_X1 U10857 ( .C1(n9656), .C2(n9670), .A(n9655), .B(n9654), .ZN(n9657)
         );
  OAI21_X1 U10858 ( .B1(n9674), .B2(n9658), .A(n9657), .ZN(P1_U3213) );
  OAI21_X1 U10859 ( .B1(n9787), .B2(n9660), .A(n9659), .ZN(n9669) );
  INV_X1 U10860 ( .A(n9661), .ZN(n9667) );
  AOI21_X1 U10861 ( .B1(n9664), .B2(n9663), .A(n9662), .ZN(n9666) );
  NOR3_X1 U10862 ( .A1(n9667), .A2(n9666), .A3(n9665), .ZN(n9668) );
  AOI211_X1 U10863 ( .C1(n9671), .C2(n9670), .A(n9669), .B(n9668), .ZN(n9672)
         );
  OAI21_X1 U10864 ( .B1(n9674), .B2(n9673), .A(n9672), .ZN(P1_U3230) );
  AOI21_X1 U10865 ( .B1(n9677), .B2(n9676), .A(n9675), .ZN(n9678) );
  XNOR2_X1 U10866 ( .A(n9678), .B(P1_IR_REG_0__SCAN_IN), .ZN(n9682) );
  AOI22_X1 U10867 ( .A1(n9679), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9680) );
  OAI21_X1 U10868 ( .B1(n9682), .B2(n9681), .A(n9680), .ZN(P1_U3243) );
  OAI21_X1 U10869 ( .B1(n9685), .B2(n9684), .A(n9683), .ZN(n9694) );
  AOI21_X1 U10870 ( .B1(n9688), .B2(n9687), .A(n9686), .ZN(n9692) );
  OAI22_X1 U10871 ( .A1(n9692), .A2(n9691), .B1(n9690), .B2(n9689), .ZN(n9693)
         );
  AOI21_X1 U10872 ( .B1(n9695), .B2(n9694), .A(n9693), .ZN(n9697) );
  OAI211_X1 U10873 ( .C1(n9699), .C2(n9698), .A(n9697), .B(n9696), .ZN(
        P1_U3255) );
  XNOR2_X1 U10874 ( .A(n9700), .B(n9703), .ZN(n9817) );
  NAND2_X1 U10875 ( .A1(n9702), .A2(n9701), .ZN(n9704) );
  XNOR2_X1 U10876 ( .A(n9704), .B(n9703), .ZN(n9707) );
  OAI21_X1 U10877 ( .B1(n9707), .B2(n9706), .A(n9705), .ZN(n9708) );
  AOI21_X1 U10878 ( .B1(n9709), .B2(n9817), .A(n9708), .ZN(n9814) );
  NOR2_X1 U10879 ( .A1(n9741), .A2(n9710), .ZN(n9711) );
  AOI21_X1 U10880 ( .B1(n9758), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9711), .ZN(
        n9712) );
  OAI21_X1 U10881 ( .B1(n9744), .B2(n9813), .A(n9712), .ZN(n9713) );
  INV_X1 U10882 ( .A(n9713), .ZN(n9721) );
  INV_X1 U10883 ( .A(n9714), .ZN(n9717) );
  INV_X1 U10884 ( .A(n9715), .ZN(n9716) );
  OAI211_X1 U10885 ( .C1(n9813), .C2(n9717), .A(n9716), .B(n9750), .ZN(n9812)
         );
  INV_X1 U10886 ( .A(n9812), .ZN(n9718) );
  AOI22_X1 U10887 ( .A1(n9817), .A2(n9719), .B1(n9754), .B2(n9718), .ZN(n9720)
         );
  OAI211_X1 U10888 ( .C1(n9758), .C2(n9814), .A(n9721), .B(n9720), .ZN(
        P1_U3285) );
  XNOR2_X1 U10889 ( .A(n9722), .B(n9730), .ZN(n9724) );
  AOI21_X1 U10890 ( .B1(n9724), .B2(n9738), .A(n9723), .ZN(n9800) );
  NOR2_X1 U10891 ( .A1(n9741), .A2(n9725), .ZN(n9726) );
  AOI21_X1 U10892 ( .B1(n9758), .B2(P1_REG2_REG_6__SCAN_IN), .A(n9726), .ZN(
        n9727) );
  OAI21_X1 U10893 ( .B1(n9744), .B2(n9799), .A(n9727), .ZN(n9728) );
  INV_X1 U10894 ( .A(n9728), .ZN(n9735) );
  XNOR2_X1 U10895 ( .A(n9729), .B(n9730), .ZN(n9803) );
  OAI211_X1 U10896 ( .C1(n9732), .C2(n9799), .A(n9731), .B(n9750), .ZN(n9798)
         );
  INV_X1 U10897 ( .A(n9798), .ZN(n9733) );
  AOI22_X1 U10898 ( .A1(n9803), .A2(n9755), .B1(n9754), .B2(n9733), .ZN(n9734)
         );
  OAI211_X1 U10899 ( .C1(n9758), .C2(n9800), .A(n9735), .B(n9734), .ZN(
        P1_U3287) );
  XOR2_X1 U10900 ( .A(n9747), .B(n9736), .Z(n9739) );
  AOI21_X1 U10901 ( .B1(n9739), .B2(n9738), .A(n9737), .ZN(n9776) );
  NOR2_X1 U10902 ( .A1(n9741), .A2(n9740), .ZN(n9742) );
  AOI21_X1 U10903 ( .B1(n9758), .B2(P1_REG2_REG_2__SCAN_IN), .A(n9742), .ZN(
        n9743) );
  OAI21_X1 U10904 ( .B1(n9744), .B2(n9775), .A(n9743), .ZN(n9745) );
  INV_X1 U10905 ( .A(n9745), .ZN(n9757) );
  XNOR2_X1 U10906 ( .A(n9747), .B(n9746), .ZN(n9779) );
  INV_X1 U10907 ( .A(n9748), .ZN(n9752) );
  INV_X1 U10908 ( .A(n9749), .ZN(n9751) );
  OAI211_X1 U10909 ( .C1(n9775), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9774)
         );
  INV_X1 U10910 ( .A(n9774), .ZN(n9753) );
  AOI22_X1 U10911 ( .A1(n9779), .A2(n9755), .B1(n9754), .B2(n9753), .ZN(n9756)
         );
  OAI211_X1 U10912 ( .C1(n9758), .C2(n9776), .A(n9757), .B(n9756), .ZN(
        P1_U3291) );
  AND2_X1 U10913 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9764), .ZN(P1_U3294) );
  AND2_X1 U10914 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9764), .ZN(P1_U3295) );
  AND2_X1 U10915 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9764), .ZN(P1_U3296) );
  AND2_X1 U10916 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9764), .ZN(P1_U3297) );
  AND2_X1 U10917 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9764), .ZN(P1_U3298) );
  AND2_X1 U10918 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9764), .ZN(P1_U3299) );
  AND2_X1 U10919 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9764), .ZN(P1_U3300) );
  AND2_X1 U10920 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9764), .ZN(P1_U3301) );
  NOR2_X1 U10921 ( .A1(n9763), .A2(n9759), .ZN(P1_U3302) );
  AND2_X1 U10922 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9764), .ZN(P1_U3303) );
  AND2_X1 U10923 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9764), .ZN(P1_U3304) );
  NOR2_X1 U10924 ( .A1(n9763), .A2(n9760), .ZN(P1_U3305) );
  AND2_X1 U10925 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9764), .ZN(P1_U3306) );
  AND2_X1 U10926 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9764), .ZN(P1_U3307) );
  AND2_X1 U10927 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9764), .ZN(P1_U3308) );
  NOR2_X1 U10928 ( .A1(n9763), .A2(n9761), .ZN(P1_U3309) );
  AND2_X1 U10929 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9764), .ZN(P1_U3310) );
  AND2_X1 U10930 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9764), .ZN(P1_U3311) );
  NOR2_X1 U10931 ( .A1(n9763), .A2(n9762), .ZN(P1_U3312) );
  AND2_X1 U10932 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9764), .ZN(P1_U3313) );
  AND2_X1 U10933 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9764), .ZN(P1_U3314) );
  AND2_X1 U10934 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9764), .ZN(P1_U3315) );
  AND2_X1 U10935 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9764), .ZN(P1_U3316) );
  AND2_X1 U10936 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9764), .ZN(P1_U3317) );
  AND2_X1 U10937 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9764), .ZN(P1_U3318) );
  AND2_X1 U10938 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9764), .ZN(P1_U3319) );
  AND2_X1 U10939 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9764), .ZN(P1_U3320) );
  AND2_X1 U10940 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9764), .ZN(P1_U3321) );
  AND2_X1 U10941 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9764), .ZN(P1_U3322) );
  AND2_X1 U10942 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9764), .ZN(P1_U3323) );
  INV_X1 U10943 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9765) );
  AOI22_X1 U10944 ( .A1(n9862), .A2(n9766), .B1(n9765), .B2(n9860), .ZN(
        P1_U3453) );
  INV_X1 U10945 ( .A(n9767), .ZN(n9856) );
  OAI21_X1 U10946 ( .B1(n9769), .B2(n9853), .A(n9768), .ZN(n9771) );
  AOI211_X1 U10947 ( .C1(n9856), .C2(n9772), .A(n9771), .B(n9770), .ZN(n9863)
         );
  INV_X1 U10948 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9773) );
  AOI22_X1 U10949 ( .A1(n9862), .A2(n9863), .B1(n9773), .B2(n9860), .ZN(
        P1_U3456) );
  OAI21_X1 U10950 ( .B1(n9775), .B2(n9853), .A(n9774), .ZN(n9778) );
  INV_X1 U10951 ( .A(n9776), .ZN(n9777) );
  AOI211_X1 U10952 ( .C1(n9850), .C2(n9779), .A(n9778), .B(n9777), .ZN(n9864)
         );
  INV_X1 U10953 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9780) );
  AOI22_X1 U10954 ( .A1(n9862), .A2(n9864), .B1(n9780), .B2(n9860), .ZN(
        P1_U3459) );
  OAI211_X1 U10955 ( .C1(n9783), .C2(n9853), .A(n9782), .B(n9781), .ZN(n9784)
         );
  AOI21_X1 U10956 ( .B1(n9850), .B2(n9785), .A(n9784), .ZN(n9865) );
  INV_X1 U10957 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10958 ( .A1(n9862), .A2(n9865), .B1(n9786), .B2(n9860), .ZN(
        P1_U3462) );
  OAI211_X1 U10959 ( .C1(n9789), .C2(n9853), .A(n9788), .B(n9787), .ZN(n9791)
         );
  AOI211_X1 U10960 ( .C1(n9850), .C2(n9792), .A(n9791), .B(n9790), .ZN(n9866)
         );
  AOI22_X1 U10961 ( .A1(n9862), .A2(n9866), .B1(n5711), .B2(n9860), .ZN(
        P1_U3465) );
  OAI21_X1 U10962 ( .B1(n9794), .B2(n9853), .A(n9793), .ZN(n9796) );
  AOI211_X1 U10963 ( .C1(n9850), .C2(n9797), .A(n9796), .B(n9795), .ZN(n9867)
         );
  AOI22_X1 U10964 ( .A1(n9862), .A2(n9867), .B1(n5737), .B2(n9860), .ZN(
        P1_U3468) );
  OAI21_X1 U10965 ( .B1(n9799), .B2(n9853), .A(n9798), .ZN(n9802) );
  INV_X1 U10966 ( .A(n9800), .ZN(n9801) );
  AOI211_X1 U10967 ( .C1(n9850), .C2(n9803), .A(n9802), .B(n9801), .ZN(n9869)
         );
  AOI22_X1 U10968 ( .A1(n9862), .A2(n9869), .B1(n5754), .B2(n9860), .ZN(
        P1_U3471) );
  INV_X1 U10969 ( .A(n9804), .ZN(n9805) );
  NAND2_X1 U10970 ( .A1(n9805), .A2(n9856), .ZN(n9807) );
  OAI211_X1 U10971 ( .C1(n9808), .C2(n9853), .A(n9807), .B(n9806), .ZN(n9809)
         );
  NOR2_X1 U10972 ( .A1(n9810), .A2(n9809), .ZN(n9870) );
  INV_X1 U10973 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U10974 ( .A1(n9862), .A2(n9870), .B1(n9811), .B2(n9860), .ZN(
        P1_U3474) );
  OAI21_X1 U10975 ( .B1(n9813), .B2(n9853), .A(n9812), .ZN(n9816) );
  INV_X1 U10976 ( .A(n9814), .ZN(n9815) );
  AOI211_X1 U10977 ( .C1(n9856), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9871)
         );
  INV_X1 U10978 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9818) );
  AOI22_X1 U10979 ( .A1(n9862), .A2(n9871), .B1(n9818), .B2(n9860), .ZN(
        P1_U3477) );
  AND2_X1 U10980 ( .A1(n9819), .A2(n9850), .ZN(n9823) );
  OAI21_X1 U10981 ( .B1(n9821), .B2(n9853), .A(n9820), .ZN(n9822) );
  NOR3_X1 U10982 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n9872) );
  INV_X1 U10983 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9825) );
  AOI22_X1 U10984 ( .A1(n9862), .A2(n9872), .B1(n9825), .B2(n9860), .ZN(
        P1_U3480) );
  OAI211_X1 U10985 ( .C1(n9828), .C2(n9853), .A(n9827), .B(n9826), .ZN(n9829)
         );
  AOI21_X1 U10986 ( .B1(n9850), .B2(n9830), .A(n9829), .ZN(n9873) );
  INV_X1 U10987 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U10988 ( .A1(n9862), .A2(n9873), .B1(n9831), .B2(n9860), .ZN(
        P1_U3483) );
  OAI21_X1 U10989 ( .B1(n9833), .B2(n9853), .A(n9832), .ZN(n9834) );
  AOI21_X1 U10990 ( .B1(n9835), .B2(n9856), .A(n9834), .ZN(n9836) );
  INV_X1 U10991 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U10992 ( .A1(n9862), .A2(n9874), .B1(n9838), .B2(n9860), .ZN(
        P1_U3486) );
  OAI211_X1 U10993 ( .C1(n9841), .C2(n9853), .A(n9840), .B(n9839), .ZN(n9842)
         );
  AOI21_X1 U10994 ( .B1(n9850), .B2(n9843), .A(n9842), .ZN(n9875) );
  AOI22_X1 U10995 ( .A1(n9862), .A2(n9875), .B1(n9844), .B2(n9860), .ZN(
        P1_U3489) );
  OAI211_X1 U10996 ( .C1(n9847), .C2(n9853), .A(n9846), .B(n9845), .ZN(n9848)
         );
  AOI21_X1 U10997 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9876) );
  INV_X1 U10998 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9851) );
  AOI22_X1 U10999 ( .A1(n9862), .A2(n9876), .B1(n9851), .B2(n9860), .ZN(
        P1_U3492) );
  OAI21_X1 U11000 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  AOI21_X1 U11001 ( .B1(n9857), .B2(n9856), .A(n9855), .ZN(n9858) );
  AND2_X1 U11002 ( .A1(n9859), .A2(n9858), .ZN(n9878) );
  INV_X1 U11003 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9861) );
  AOI22_X1 U11004 ( .A1(n9862), .A2(n9878), .B1(n9861), .B2(n9860), .ZN(
        P1_U3495) );
  AOI22_X1 U11005 ( .A1(n9879), .A2(n9863), .B1(n6306), .B2(n9877), .ZN(
        P1_U3523) );
  AOI22_X1 U11006 ( .A1(n9879), .A2(n9864), .B1(n6307), .B2(n9877), .ZN(
        P1_U3524) );
  AOI22_X1 U11007 ( .A1(n9879), .A2(n9865), .B1(n6321), .B2(n9877), .ZN(
        P1_U3525) );
  AOI22_X1 U11008 ( .A1(n9879), .A2(n9866), .B1(n6323), .B2(n9877), .ZN(
        P1_U3526) );
  AOI22_X1 U11009 ( .A1(n9879), .A2(n9867), .B1(n6318), .B2(n9877), .ZN(
        P1_U3527) );
  AOI22_X1 U11010 ( .A1(n9879), .A2(n9869), .B1(n9868), .B2(n9877), .ZN(
        P1_U3528) );
  AOI22_X1 U11011 ( .A1(n9879), .A2(n9870), .B1(n6343), .B2(n9877), .ZN(
        P1_U3529) );
  AOI22_X1 U11012 ( .A1(n9879), .A2(n9871), .B1(n6342), .B2(n9877), .ZN(
        P1_U3530) );
  AOI22_X1 U11013 ( .A1(n9879), .A2(n9872), .B1(n5803), .B2(n9877), .ZN(
        P1_U3531) );
  AOI22_X1 U11014 ( .A1(n9879), .A2(n9873), .B1(n6414), .B2(n9877), .ZN(
        P1_U3532) );
  AOI22_X1 U11015 ( .A1(n9879), .A2(n9874), .B1(n6612), .B2(n9877), .ZN(
        P1_U3533) );
  AOI22_X1 U11016 ( .A1(n9879), .A2(n9875), .B1(n5883), .B2(n9877), .ZN(
        P1_U3534) );
  AOI22_X1 U11017 ( .A1(n9879), .A2(n9876), .B1(n5907), .B2(n9877), .ZN(
        P1_U3535) );
  AOI22_X1 U11018 ( .A1(n9879), .A2(n9878), .B1(n6952), .B2(n9877), .ZN(
        P1_U3536) );
  AOI22_X1 U11019 ( .A1(n9959), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n9887) );
  NOR2_X1 U11020 ( .A1(n9882), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9880) );
  AOI211_X1 U11021 ( .C1(n9882), .C2(n9881), .A(P2_IR_REG_0__SCAN_IN), .B(
        n9880), .ZN(n9883) );
  OAI22_X1 U11022 ( .A1(n9885), .A2(n9970), .B1(n9884), .B2(n9883), .ZN(n9886)
         );
  OAI211_X1 U11023 ( .C1(n9980), .C2(n4791), .A(n9887), .B(n9886), .ZN(
        P2_U3182) );
  INV_X1 U11024 ( .A(n9888), .ZN(n9897) );
  AOI21_X1 U11025 ( .B1(n5097), .B2(n9890), .A(n9889), .ZN(n9894) );
  AOI21_X1 U11026 ( .B1(n6551), .B2(n9892), .A(n9891), .ZN(n9893) );
  OAI22_X1 U11027 ( .A1(n9974), .A2(n9894), .B1(n9893), .B2(n9965), .ZN(n9895)
         );
  AOI211_X1 U11028 ( .C1(n9897), .C2(n9914), .A(n9896), .B(n9895), .ZN(n9903)
         );
  OAI21_X1 U11029 ( .B1(n9900), .B2(n9899), .A(n9898), .ZN(n9901) );
  NAND2_X1 U11030 ( .A1(n9901), .A2(n9970), .ZN(n9902) );
  OAI211_X1 U11031 ( .C1(n9904), .C2(n9924), .A(n9903), .B(n9902), .ZN(
        P2_U3185) );
  AOI21_X1 U11032 ( .B1(n9907), .B2(n9906), .A(n9905), .ZN(n9911) );
  AOI21_X1 U11033 ( .B1(n9909), .B2(n9908), .A(n4410), .ZN(n9910) );
  OAI22_X1 U11034 ( .A1(n9974), .A2(n9911), .B1(n9910), .B2(n9965), .ZN(n9912)
         );
  AOI211_X1 U11035 ( .C1(n9915), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9922)
         );
  AOI211_X1 U11036 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9916), .ZN(n9920)
         );
  INV_X1 U11037 ( .A(n9920), .ZN(n9921) );
  OAI211_X1 U11038 ( .C1(n9924), .C2(n9923), .A(n9922), .B(n9921), .ZN(
        P2_U3186) );
  AOI21_X1 U11039 ( .B1(n9926), .B2(n5124), .A(n9925), .ZN(n9927) );
  OAI22_X1 U11040 ( .A1(n9980), .A2(n9928), .B1(n9965), .B2(n9927), .ZN(n9929)
         );
  AOI21_X1 U11041 ( .B1(n9959), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9929), .ZN(
        n9939) );
  INV_X1 U11042 ( .A(n9930), .ZN(n9938) );
  XOR2_X1 U11043 ( .A(n9932), .B(n9931), .Z(n9933) );
  NAND2_X1 U11044 ( .A1(n9933), .A2(n9970), .ZN(n9937) );
  OAI21_X1 U11045 ( .B1(n4408), .B2(P2_REG1_REG_5__SCAN_IN), .A(n9934), .ZN(
        n9935) );
  NAND2_X1 U11046 ( .A1(n9951), .A2(n9935), .ZN(n9936) );
  NAND4_X1 U11047 ( .A1(n9939), .A2(n9938), .A3(n9937), .A4(n9936), .ZN(
        P2_U3187) );
  AOI21_X1 U11048 ( .B1(n9941), .B2(n6890), .A(n9940), .ZN(n9943) );
  OAI22_X1 U11049 ( .A1(n9943), .A2(n9965), .B1(n9980), .B2(n9942), .ZN(n9944)
         );
  AOI21_X1 U11050 ( .B1(n9959), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n9944), .ZN(
        n9957) );
  OAI21_X1 U11051 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(n9948) );
  NAND2_X1 U11052 ( .A1(n9948), .A2(n9970), .ZN(n9955) );
  INV_X1 U11053 ( .A(n9949), .ZN(n9950) );
  NOR2_X1 U11054 ( .A1(n9950), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9952) );
  OAI21_X1 U11055 ( .B1(n9953), .B2(n9952), .A(n9951), .ZN(n9954) );
  NAND4_X1 U11056 ( .A1(n9957), .A2(n9956), .A3(n9955), .A4(n9954), .ZN(
        P2_U3189) );
  AOI22_X1 U11057 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n9959), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n9978) );
  AOI21_X1 U11058 ( .B1(n4346), .B2(n9961), .A(n9960), .ZN(n9975) );
  AOI21_X1 U11059 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9966) );
  OR2_X1 U11060 ( .A1(n9966), .A2(n9965), .ZN(n9973) );
  OAI21_X1 U11061 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(n9971) );
  NAND2_X1 U11062 ( .A1(n9971), .A2(n9970), .ZN(n9972) );
  OAI211_X1 U11063 ( .C1(n9975), .C2(n9974), .A(n9973), .B(n9972), .ZN(n9976)
         );
  INV_X1 U11064 ( .A(n9976), .ZN(n9977) );
  OAI211_X1 U11065 ( .C1(n9980), .C2(n9979), .A(n9978), .B(n9977), .ZN(
        P2_U3196) );
  XOR2_X1 U11066 ( .A(n9990), .B(n9981), .Z(n9986) );
  AOI222_X1 U11067 ( .A1(n9987), .A2(n9986), .B1(n9985), .B2(n9984), .C1(n9983), .C2(n9982), .ZN(n10042) );
  NAND2_X1 U11068 ( .A1(n9989), .A2(n9988), .ZN(n9991) );
  XNOR2_X1 U11069 ( .A(n9991), .B(n9990), .ZN(n10040) );
  INV_X1 U11070 ( .A(n9992), .ZN(n9995) );
  AOI222_X1 U11071 ( .A1(n10040), .A2(n9996), .B1(n9995), .B2(n9994), .C1(
        n10039), .C2(n9993), .ZN(n9997) );
  OAI221_X1 U11072 ( .B1(n8334), .B2(n10042), .C1(n10016), .C2(n9998), .A(
        n9997), .ZN(P2_U3227) );
  OAI21_X1 U11073 ( .B1(n9999), .B2(n10005), .A(n10000), .ZN(n10021) );
  OAI22_X1 U11074 ( .A1(n10018), .A2(n10003), .B1(n10002), .B2(n10001), .ZN(
        n10014) );
  XNOR2_X1 U11075 ( .A(n10004), .B(n10005), .ZN(n10012) );
  OAI22_X1 U11076 ( .A1(n10008), .A2(n10007), .B1(n10006), .B2(n8307), .ZN(
        n10009) );
  AOI21_X1 U11077 ( .B1(n10021), .B2(n10010), .A(n10009), .ZN(n10011) );
  OAI21_X1 U11078 ( .B1(n10013), .B2(n10012), .A(n10011), .ZN(n10019) );
  AOI211_X1 U11079 ( .C1(n10015), .C2(n10021), .A(n10014), .B(n10019), .ZN(
        n10017) );
  AOI22_X1 U11080 ( .A1(n8334), .A2(n5077), .B1(n10017), .B2(n10016), .ZN(
        P2_U3231) );
  INV_X1 U11081 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U11082 ( .A1(n10018), .A2(n10054), .ZN(n10020) );
  AOI211_X1 U11083 ( .C1(n10046), .C2(n10021), .A(n10020), .B(n10019), .ZN(
        n10077) );
  AOI22_X1 U11084 ( .A1(n10076), .A2(n10022), .B1(n10077), .B2(n10074), .ZN(
        P2_U3396) );
  OAI21_X1 U11085 ( .B1(n10024), .B2(n10054), .A(n10023), .ZN(n10025) );
  AOI21_X1 U11086 ( .B1(n10026), .B2(n10068), .A(n10025), .ZN(n10078) );
  AOI22_X1 U11087 ( .A1(n10076), .A2(n10027), .B1(n10078), .B2(n10074), .ZN(
        P2_U3399) );
  INV_X1 U11088 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10033) );
  INV_X1 U11089 ( .A(n10028), .ZN(n10032) );
  OAI21_X1 U11090 ( .B1(n10030), .B2(n10054), .A(n10029), .ZN(n10031) );
  AOI21_X1 U11091 ( .B1(n10032), .B2(n10068), .A(n10031), .ZN(n10079) );
  AOI22_X1 U11092 ( .A1(n10076), .A2(n10033), .B1(n10079), .B2(n10074), .ZN(
        P2_U3402) );
  INV_X1 U11093 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10038) );
  NOR2_X1 U11094 ( .A1(n10034), .A2(n10054), .ZN(n10036) );
  AOI211_X1 U11095 ( .C1(n10037), .C2(n10068), .A(n10036), .B(n10035), .ZN(
        n10081) );
  AOI22_X1 U11096 ( .A1(n10076), .A2(n10038), .B1(n10081), .B2(n10074), .ZN(
        P2_U3405) );
  AOI22_X1 U11097 ( .A1(n10040), .A2(n10068), .B1(n10073), .B2(n10039), .ZN(
        n10041) );
  AND2_X1 U11098 ( .A1(n10042), .A2(n10041), .ZN(n10083) );
  AOI22_X1 U11099 ( .A1(n10076), .A2(n5144), .B1(n10083), .B2(n10074), .ZN(
        P2_U3408) );
  INV_X1 U11100 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U11101 ( .A1(n10043), .A2(n10054), .ZN(n10045) );
  AOI211_X1 U11102 ( .C1(n10047), .C2(n10046), .A(n10045), .B(n10044), .ZN(
        n10084) );
  AOI22_X1 U11103 ( .A1(n10076), .A2(n10048), .B1(n10084), .B2(n10074), .ZN(
        P2_U3411) );
  INV_X1 U11104 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10053) );
  OAI22_X1 U11105 ( .A1(n10050), .A2(n10056), .B1(n10049), .B2(n10054), .ZN(
        n10051) );
  NOR2_X1 U11106 ( .A1(n10052), .A2(n10051), .ZN(n10086) );
  AOI22_X1 U11107 ( .A1(n10076), .A2(n10053), .B1(n10086), .B2(n10074), .ZN(
        P2_U3417) );
  INV_X1 U11108 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10060) );
  OAI22_X1 U11109 ( .A1(n10057), .A2(n10056), .B1(n10055), .B2(n10054), .ZN(
        n10058) );
  NOR2_X1 U11110 ( .A1(n10059), .A2(n10058), .ZN(n10087) );
  AOI22_X1 U11111 ( .A1(n10076), .A2(n10060), .B1(n10087), .B2(n10074), .ZN(
        P2_U3420) );
  INV_X1 U11112 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U11113 ( .A1(n10062), .A2(n10061), .ZN(n10064) );
  AOI211_X1 U11114 ( .C1(n10073), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10089) );
  AOI22_X1 U11115 ( .A1(n10076), .A2(n10066), .B1(n10089), .B2(n10074), .ZN(
        P2_U3423) );
  INV_X1 U11116 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10075) );
  AND3_X1 U11117 ( .A1(n10069), .A2(n10068), .A3(n10067), .ZN(n10071) );
  AOI211_X1 U11118 ( .C1(n10073), .C2(n10072), .A(n10071), .B(n10070), .ZN(
        n10091) );
  AOI22_X1 U11119 ( .A1(n10076), .A2(n10075), .B1(n10091), .B2(n10074), .ZN(
        P2_U3426) );
  AOI22_X1 U11120 ( .A1(n10092), .A2(n10077), .B1(n6571), .B2(n10090), .ZN(
        P2_U3461) );
  AOI22_X1 U11121 ( .A1(n10092), .A2(n10078), .B1(n5097), .B2(n10090), .ZN(
        P2_U3462) );
  AOI22_X1 U11122 ( .A1(n10092), .A2(n10079), .B1(n6579), .B2(n10090), .ZN(
        P2_U3463) );
  AOI22_X1 U11123 ( .A1(n10092), .A2(n10081), .B1(n10080), .B2(n10090), .ZN(
        P2_U3464) );
  AOI22_X1 U11124 ( .A1(n10092), .A2(n10083), .B1(n10082), .B2(n10090), .ZN(
        P2_U3465) );
  AOI22_X1 U11125 ( .A1(n10092), .A2(n10084), .B1(n5157), .B2(n10090), .ZN(
        P2_U3466) );
  AOI22_X1 U11126 ( .A1(n10092), .A2(n10086), .B1(n10085), .B2(n10090), .ZN(
        P2_U3468) );
  AOI22_X1 U11127 ( .A1(n10092), .A2(n10087), .B1(n5208), .B2(n10090), .ZN(
        P2_U3469) );
  AOI22_X1 U11128 ( .A1(n10092), .A2(n10089), .B1(n10088), .B2(n10090), .ZN(
        P2_U3470) );
  AOI22_X1 U11129 ( .A1(n10092), .A2(n10091), .B1(n7254), .B2(n10090), .ZN(
        P2_U3471) );
  INV_X1 U11130 ( .A(n10093), .ZN(n10096) );
  AOI21_X1 U11131 ( .B1(P1_ADDR_REG_1__SCAN_IN), .B2(n10098), .A(n10097), .ZN(
        n10095) );
  OAI22_X1 U11132 ( .A1(n10097), .A2(n10096), .B1(n10095), .B2(n10094), .ZN(
        ADD_1068_U5) );
  AOI21_X1 U11133 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(ADD_1068_U46) );
  OAI21_X1 U11134 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n10102), .A(n10101), 
        .ZN(n10103) );
  XNOR2_X1 U11135 ( .A(n10103), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  XNOR2_X1 U11136 ( .A(n10105), .B(n10104), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11137 ( .A(n10107), .B(n10106), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11138 ( .A(n10109), .B(n10108), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11139 ( .A(n10111), .B(n10110), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11140 ( .A(n10113), .B(n10112), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11141 ( .A(n10115), .B(n10114), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11142 ( .A(n10117), .B(n10116), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11143 ( .A(n10119), .B(n10118), .ZN(ADD_1068_U63) );
  XNOR2_X1 U11144 ( .A(n10121), .B(n10120), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11145 ( .A(n10123), .B(n10122), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11146 ( .A(n10125), .B(n10124), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11147 ( .A(n10127), .B(n10126), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11148 ( .A(n10129), .B(n10128), .ZN(ADD_1068_U48) );
  XOR2_X1 U11149 ( .A(n10131), .B(n10130), .Z(ADD_1068_U54) );
  XOR2_X1 U11150 ( .A(n10133), .B(n10132), .Z(ADD_1068_U53) );
  XNOR2_X1 U11151 ( .A(n10135), .B(n10134), .ZN(ADD_1068_U52) );
  NAND2_X1 U4825 ( .A1(n5352), .A2(n5351), .ZN(n5366) );
  CLKBUF_X1 U4805 ( .A(n5798), .Z(n4299) );
  CLKBUF_X1 U4855 ( .A(n5088), .Z(n5305) );
  INV_X1 U4973 ( .A(n8737), .ZN(n8786) );
  CLKBUF_X2 U5068 ( .A(n8620), .Z(n4308) );
  CLKBUF_X1 U7180 ( .A(n9431), .Z(n4305) );
endmodule

