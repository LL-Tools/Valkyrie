

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362;

  INV_X1 U4790 ( .A(n8874), .ZN(n10102) );
  CLKBUF_X2 U4791 ( .A(n7096), .Z(n7204) );
  CLKBUF_X2 U4792 ( .A(n7096), .Z(n8406) );
  INV_X1 U4793 ( .A(n6976), .ZN(n6127) );
  OR2_X1 U4794 ( .A1(n9371), .A2(n8235), .ZN(n8154) );
  AND3_X1 U4795 ( .A1(n5083), .A2(n5082), .A3(n5081), .ZN(n7862) );
  NAND4_X1 U4796 ( .A1(n5070), .A2(n5069), .A3(n5068), .A4(n5067), .ZN(n5084)
         );
  INV_X1 U4797 ( .A(n5065), .ZN(n5579) );
  CLKBUF_X2 U4798 ( .A(n5578), .Z(n4290) );
  AND2_X1 U4799 ( .A1(n4565), .A2(n4324), .ZN(n4564) );
  NAND2_X1 U4800 ( .A1(n6542), .A2(n6541), .ZN(n6732) );
  AND2_X1 U4801 ( .A1(n8212), .A2(n8019), .ZN(n6384) );
  INV_X1 U4802 ( .A(n4999), .ZN(n5002) );
  INV_X1 U4803 ( .A(n8403), .ZN(n7260) );
  AND2_X1 U4804 ( .A1(n4289), .A2(n4292), .ZN(n5576) );
  NAND2_X1 U4805 ( .A1(n6568), .A2(n6700), .ZN(n7825) );
  MUX2_X1 U4806 ( .A(n8746), .B(n8745), .S(n8744), .Z(n8747) );
  NAND2_X1 U4807 ( .A1(n4907), .A2(n4905), .ZN(n4909) );
  AND3_X1 U4808 ( .A1(n5126), .A2(n5125), .A3(n5124), .ZN(n10057) );
  AOI22_X1 U4809 ( .A1(n8578), .A2(n8579), .B1(n6502), .B2(n6470), .ZN(n6476)
         );
  OAI21_X1 U4810 ( .B1(n8437), .B2(n4937), .A(n4935), .ZN(n8506) );
  AND2_X1 U4811 ( .A1(n6163), .A2(n6162), .ZN(n8788) );
  NOR2_X1 U4812 ( .A1(n7758), .A2(n7759), .ZN(n7809) );
  AND2_X1 U4813 ( .A1(n5554), .A2(n5553), .ZN(n8404) );
  AND2_X1 U4814 ( .A1(n6374), .A2(n6373), .ZN(n9572) );
  INV_X1 U4815 ( .A(n5640), .ZN(n7334) );
  INV_X1 U4817 ( .A(n5000), .ZN(n9987) );
  INV_X1 U4818 ( .A(n6385), .ZN(n6341) );
  OAI21_X1 U4819 ( .B1(n9268), .B2(n9267), .A(n9302), .ZN(n9273) );
  INV_X1 U4820 ( .A(n8404), .ZN(n5555) );
  NAND4_X2 U4821 ( .A1(n5110), .A2(n5109), .A3(n5108), .A4(n5107), .ZN(n9372)
         );
  AND2_X1 U4823 ( .A1(n4795), .A2(n4794), .ZN(n4284) );
  NAND2_X1 U4824 ( .A1(n9987), .A2(n5002), .ZN(n5578) );
  INV_X2 U4825 ( .A(n5929), .ZN(n9084) );
  NAND2_X1 U4826 ( .A1(n10002), .A2(n5674), .ZN(n5053) );
  NAND2_X2 U4827 ( .A1(n5929), .A2(n5930), .ZN(n5957) );
  MUX2_X2 U4828 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5751), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5752) );
  NAND2_X2 U4829 ( .A1(n5755), .A2(n4749), .ZN(n4396) );
  CLKBUF_X1 U4830 ( .A(n7344), .Z(n4285) );
  BUF_X4 U4831 ( .A(n7344), .Z(n4286) );
  NAND2_X1 U4832 ( .A1(n5009), .A2(n5008), .ZN(n7344) );
  NAND2_X2 U4833 ( .A1(n5810), .A2(n5809), .ZN(n7484) );
  INV_X1 U4834 ( .A(n5748), .ZN(n5755) );
  OAI222_X1 U4835 ( .A1(n7492), .A2(P2_U3151), .B1(n9093), .B2(n7357), .C1(
        n7356), .C2(n9097), .ZN(P2_U3293) );
  NOR2_X2 U4836 ( .A1(n8739), .A2(n8738), .ZN(n8743) );
  INV_X1 U4837 ( .A(n6539), .ZN(n5672) );
  AOI22_X2 U4838 ( .A1(n7048), .A2(n6228), .B1(n7053), .B2(n8759), .ZN(n7021)
         );
  AOI21_X2 U4839 ( .B1(n8756), .B2(n6948), .A(n6955), .ZN(n7048) );
  NAND2_X2 U4840 ( .A1(n8703), .A2(n4630), .ZN(n5830) );
  NAND2_X2 U4841 ( .A1(n5922), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5731) );
  NAND2_X2 U4842 ( .A1(n5732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5734) );
  XNOR2_X2 U4843 ( .A(n5759), .B(n7473), .ZN(n7467) );
  OAI22_X2 U4844 ( .A1(n7467), .A2(n7644), .B1(n5759), .B2(n7473), .ZN(n8617)
         );
  AOI21_X2 U4845 ( .B1(n7487), .B2(n7488), .A(n4352), .ZN(n5759) );
  XNOR2_X2 U4846 ( .A(n5812), .B(n7473), .ZN(n7468) );
  OAI21_X1 U4847 ( .B1(n5824), .B2(n4627), .A(n4316), .ZN(n4626) );
  XNOR2_X2 U4848 ( .A(n4732), .B(n4731), .ZN(n8635) );
  XNOR2_X2 U4849 ( .A(n5802), .B(n5801), .ZN(n8019) );
  AOI22_X2 U4850 ( .A1(n7499), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n7503), .B2(
        n5764), .ZN(n7616) );
  XNOR2_X2 U4851 ( .A(n5764), .B(n5987), .ZN(n7499) );
  XNOR2_X2 U4852 ( .A(n4996), .B(n4995), .ZN(n5000) );
  NAND2_X2 U4853 ( .A1(n9982), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4996) );
  INV_X4 U4854 ( .A(n6308), .ZN(n5895) );
  NAND2_X1 U4855 ( .A1(n8311), .A2(n8310), .ZN(n8309) );
  AOI21_X1 U4856 ( .B1(n4555), .B2(n4552), .A(n4342), .ZN(n4551) );
  NOR3_X1 U4857 ( .A1(n9727), .A2(n4765), .A3(n9662), .ZN(n4763) );
  AND2_X1 U4858 ( .A1(n5536), .A2(n5535), .ZN(n7272) );
  AOI21_X1 U4859 ( .B1(n7691), .B2(n4314), .A(n4626), .ZN(n5825) );
  NAND2_X1 U4860 ( .A1(n5312), .A2(n5311), .ZN(n9870) );
  NAND2_X1 U4861 ( .A1(n4747), .A2(n4746), .ZN(n7765) );
  OR2_X1 U4862 ( .A1(n7608), .A2(n7609), .ZN(n7512) );
  OR2_X1 U4863 ( .A1(n9370), .A2(n8249), .ZN(n6765) );
  INV_X1 U4864 ( .A(n6761), .ZN(n7933) );
  INV_X1 U4865 ( .A(n7624), .ZN(n7627) );
  INV_X1 U4866 ( .A(n7825), .ZN(n6759) );
  INV_X1 U4867 ( .A(n6454), .ZN(n6471) );
  NAND2_X1 U4868 ( .A1(n5683), .A2(n7862), .ZN(n7846) );
  OR2_X1 U4869 ( .A1(n7615), .A2(n4739), .ZN(n4735) );
  CLKBUF_X2 U4870 ( .A(P1_U3973), .Z(n9390) );
  AND4_X1 U4871 ( .A1(n5006), .A2(n5005), .A3(n5004), .A4(n5003), .ZN(n7071)
         );
  NAND2_X1 U4872 ( .A1(n8620), .A2(n5815), .ZN(n5816) );
  NAND4_X2 U4873 ( .A1(n5090), .A2(n5089), .A3(n5088), .A4(n5087), .ZN(n9373)
         );
  INV_X2 U4874 ( .A(n8615), .ZN(n6247) );
  INV_X2 U4875 ( .A(n6980), .ZN(n6988) );
  NAND2_X1 U4876 ( .A1(n7629), .A2(n7645), .ZN(n6850) );
  NAND2_X2 U4877 ( .A1(n6385), .A2(n7036), .ZN(n6980) );
  BUF_X2 U4878 ( .A(n5950), .Z(n6966) );
  NAND2_X1 U4879 ( .A1(n7062), .A2(n8188), .ZN(n9801) );
  INV_X1 U4880 ( .A(n7836), .ZN(n7715) );
  INV_X2 U4881 ( .A(n5053), .ZN(n7441) );
  INV_X2 U4882 ( .A(n7345), .ZN(n7473) );
  XNOR2_X1 U4883 ( .A(n5839), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7487) );
  CLKBUF_X3 U4884 ( .A(n4286), .Z(n7342) );
  INV_X1 U4885 ( .A(n4286), .ZN(n5118) );
  OR2_X1 U4886 ( .A1(n5756), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5761) );
  NAND2_X2 U4887 ( .A1(n5009), .A2(n5008), .ZN(n4292) );
  NAND3_X1 U4888 ( .A1(n5748), .A2(n5693), .A3(n5692), .ZN(n5760) );
  AOI21_X1 U4889 ( .B1(n9580), .B2(n10344), .A(n9579), .ZN(n9581) );
  AND2_X1 U4890 ( .A1(n9590), .A2(n4434), .ZN(n9906) );
  AND2_X1 U4891 ( .A1(n6377), .A2(n9778), .ZN(n4423) );
  INV_X1 U4892 ( .A(n4438), .ZN(n4386) );
  OR2_X1 U4893 ( .A1(n8436), .A2(n9963), .ZN(n4433) );
  OR2_X1 U4894 ( .A1(n8436), .A2(n9872), .ZN(n6370) );
  AND3_X1 U4895 ( .A1(n4616), .A2(n4639), .A3(n7037), .ZN(n4459) );
  NAND2_X1 U4896 ( .A1(n7266), .A2(n7265), .ZN(n9320) );
  AOI21_X1 U4897 ( .B1(n9583), .B2(n10061), .A(n5918), .ZN(n4434) );
  AOI21_X1 U4898 ( .B1(n4728), .B2(n10096), .A(n4725), .ZN(n8987) );
  AND2_X1 U4899 ( .A1(n4886), .A2(n6295), .ZN(n7041) );
  NOR2_X1 U4900 ( .A1(n6821), .A2(n6794), .ZN(n6795) );
  AND2_X1 U4901 ( .A1(n8395), .A2(n9807), .ZN(n8391) );
  AND2_X1 U4902 ( .A1(n4648), .A2(n4394), .ZN(n6975) );
  NAND2_X1 U4903 ( .A1(n4803), .A2(n4801), .ZN(n9112) );
  XNOR2_X1 U4904 ( .A(n6527), .B(n6685), .ZN(n6528) );
  OR2_X1 U4905 ( .A1(n7239), .A2(n4804), .ZN(n4803) );
  NOR2_X1 U4906 ( .A1(n6937), .A2(n4346), .ZN(n4394) );
  NAND2_X1 U4907 ( .A1(n8716), .A2(n5831), .ZN(n8728) );
  NAND2_X1 U4908 ( .A1(n4708), .A2(n6273), .ZN(n8833) );
  AOI21_X1 U4909 ( .B1(n4551), .B2(n4553), .A(n4548), .ZN(n4547) );
  AOI21_X1 U4910 ( .B1(n4810), .B2(n4813), .A(n4809), .ZN(n4808) );
  AOI21_X1 U4911 ( .B1(n4814), .B2(n4812), .A(n4811), .ZN(n4810) );
  AND2_X1 U4912 ( .A1(n9637), .A2(n6645), .ZN(n9652) );
  NAND2_X1 U4913 ( .A1(n4463), .A2(n4461), .ZN(n5560) );
  NAND2_X1 U4914 ( .A1(n4502), .A2(n4914), .ZN(n7748) );
  NAND2_X1 U4915 ( .A1(n6147), .A2(n6146), .ZN(n9025) );
  NAND2_X1 U4916 ( .A1(n5412), .A2(n5411), .ZN(n7218) );
  AND2_X1 U4917 ( .A1(n7105), .A2(n4300), .ZN(n4796) );
  NAND2_X1 U4918 ( .A1(n5330), .A2(n5329), .ZN(n9861) );
  NAND2_X1 U4919 ( .A1(n6137), .A2(n6136), .ZN(n6277) );
  NAND2_X1 U4920 ( .A1(n5823), .A2(n7699), .ZN(n5824) );
  NAND2_X1 U4921 ( .A1(n5399), .A2(n5398), .ZN(n9843) );
  AND2_X1 U4922 ( .A1(n7918), .A2(n7916), .ZN(n7105) );
  NAND2_X1 U4923 ( .A1(n6070), .A2(n6069), .ZN(n9065) );
  NAND2_X1 U4924 ( .A1(n10099), .A2(n10098), .ZN(n10097) );
  NAND2_X1 U4925 ( .A1(n5388), .A2(n5387), .ZN(n9847) );
  NAND2_X1 U4926 ( .A1(n5258), .A2(n5257), .ZN(n8354) );
  NAND2_X1 U4927 ( .A1(n6059), .A2(n6058), .ZN(n8972) );
  NAND2_X1 U4928 ( .A1(n6050), .A2(n6049), .ZN(n8563) );
  NAND2_X1 U4929 ( .A1(n9259), .A2(n7143), .ZN(n6592) );
  NAND2_X1 U4930 ( .A1(n5858), .A2(n7514), .ZN(n7677) );
  OAI21_X1 U4931 ( .B1(n5395), .B2(n5394), .A(n5393), .ZN(n5430) );
  NAND2_X1 U4932 ( .A1(n5290), .A2(n5289), .ZN(n9967) );
  CLKBUF_X1 U4933 ( .A(n9259), .Z(n4435) );
  NAND2_X1 U4934 ( .A1(n5241), .A2(n5240), .ZN(n9885) );
  NAND2_X1 U4935 ( .A1(n6765), .A2(n6576), .ZN(n8241) );
  NAND2_X1 U4936 ( .A1(n6037), .A2(n6036), .ZN(n8976) );
  NAND2_X1 U4937 ( .A1(n5219), .A2(n5218), .ZN(n9133) );
  NAND2_X1 U4938 ( .A1(n5200), .A2(n5199), .ZN(n9259) );
  NAND2_X1 U4939 ( .A1(n7672), .A2(n7673), .ZN(n7671) );
  XNOR2_X1 U4940 ( .A(n4403), .B(n4977), .ZN(n7393) );
  AND2_X1 U4941 ( .A1(n5168), .A2(n5167), .ZN(n8249) );
  AND2_X1 U4942 ( .A1(n5147), .A2(n5146), .ZN(n8235) );
  OR2_X1 U4943 ( .A1(n6138), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U4944 ( .A1(n5816), .A2(n7503), .ZN(n5817) );
  XNOR2_X1 U4945 ( .A(n5816), .B(n5987), .ZN(n7498) );
  NAND2_X1 U4946 ( .A1(n6245), .A2(n7454), .ZN(n6837) );
  INV_X1 U4947 ( .A(n10124), .ZN(n7654) );
  INV_X2 U4948 ( .A(n7381), .ZN(n7400) );
  AND3_X1 U4949 ( .A1(n5102), .A2(n5101), .A3(n5100), .ZN(n7854) );
  OR2_X1 U4950 ( .A1(n7465), .A2(n7466), .ZN(n8626) );
  AND4_X1 U4951 ( .A1(n5185), .A2(n5184), .A3(n5183), .A4(n5182), .ZN(n7134)
         );
  AND2_X1 U4952 ( .A1(n7066), .A2(n7935), .ZN(n4439) );
  NAND4_X1 U4953 ( .A1(n5136), .A2(n5135), .A3(n5134), .A4(n5133), .ZN(n9371)
         );
  INV_X1 U4954 ( .A(n7273), .ZN(n7096) );
  NAND4_X1 U4955 ( .A1(n5999), .A2(n5998), .A3(n5997), .A4(n5996), .ZN(n10079)
         );
  NAND2_X1 U4956 ( .A1(n5814), .A2(n5813), .ZN(n8621) );
  INV_X1 U4957 ( .A(n5686), .ZN(n7065) );
  OAI211_X1 U4958 ( .C1(n6229), .C2(n7355), .A(n4605), .B(n4299), .ZN(n7454)
         );
  AND2_X2 U4959 ( .A1(n5624), .A2(n5623), .ZN(n7070) );
  AOI21_X1 U4960 ( .B1(n4866), .B2(n4868), .A(n4864), .ZN(n4863) );
  XNOR2_X1 U4961 ( .A(n5600), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U4962 ( .A1(n4444), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5259) );
  NAND2_X1 U4963 ( .A1(n5629), .A2(n5633), .ZN(n8188) );
  XNOR2_X1 U4964 ( .A(n5386), .B(n5592), .ZN(n6539) );
  INV_X1 U4965 ( .A(n6969), .ZN(n5926) );
  NAND2_X2 U4966 ( .A1(n6316), .A2(n4292), .ZN(n6976) );
  AND2_X1 U4967 ( .A1(n5713), .A2(n5732), .ZN(n7365) );
  XNOR2_X1 U4968 ( .A(n5628), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7062) );
  INV_X1 U4969 ( .A(n5222), .ZN(n4444) );
  NAND2_X1 U4970 ( .A1(n5385), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5386) );
  NOR2_X1 U4971 ( .A1(n5191), .A2(n4870), .ZN(n4869) );
  NAND2_X1 U4972 ( .A1(n5178), .A2(n5190), .ZN(n5191) );
  NAND2_X1 U4973 ( .A1(n4445), .A2(n4336), .ZN(n5222) );
  INV_X2 U4974 ( .A(n9082), .ZN(n9093) );
  NAND2_X1 U4975 ( .A1(n5363), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5384) );
  INV_X1 U4976 ( .A(n5202), .ZN(n4445) );
  NAND2_X1 U4977 ( .A1(n9080), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U4978 ( .A1(n5011), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5013) );
  NAND2_X1 U4979 ( .A1(n4389), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5925) );
  NAND2_X2 U4980 ( .A1(n7342), .A2(P1_U3086), .ZN(n9994) );
  NAND2_X1 U4981 ( .A1(n5808), .A2(n5807), .ZN(n7579) );
  INV_X1 U4982 ( .A(n7492), .ZN(n5839) );
  NAND2_X1 U4983 ( .A1(n5758), .A2(n5761), .ZN(n7345) );
  NAND3_X2 U4984 ( .A1(n4396), .A2(n5756), .A3(n4750), .ZN(n7492) );
  INV_X1 U4985 ( .A(n5760), .ZN(n4677) );
  AND2_X1 U4986 ( .A1(n4980), .A2(n5733), .ZN(n4910) );
  NAND2_X2 U4987 ( .A1(n5752), .A2(n5755), .ZN(n7587) );
  NAND3_X1 U4988 ( .A1(n5906), .A2(n4458), .A3(n4457), .ZN(n5009) );
  AND4_X1 U4989 ( .A1(n5695), .A2(n5696), .A3(n5697), .A4(n5723), .ZN(n4674)
         );
  INV_X1 U4990 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5590) );
  INV_X1 U4991 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5710) );
  INV_X1 U4992 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5708) );
  NOR2_X1 U4993 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5700) );
  NOR2_X1 U4994 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5699) );
  INV_X1 U4995 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U4996 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4759) );
  NOR2_X1 U4997 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n4760) );
  NOR2_X1 U4998 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4761) );
  NOR2_X1 U4999 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4762) );
  INV_X4 U5000 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U5001 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5694) );
  INV_X4 U5002 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5003 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5906) );
  INV_X1 U5004 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5120) );
  NOR2_X1 U5005 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5693) );
  INV_X1 U5006 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4458) );
  INV_X1 U5007 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4457) );
  CLKBUF_X1 U5008 ( .A(n7610), .Z(n4287) );
  AOI21_X1 U5009 ( .B1(n4294), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n4453), .ZN(
        n4452) );
  NAND2_X2 U5010 ( .A1(n7610), .A2(n5818), .ZN(n5819) );
  OAI21_X2 U5011 ( .B1(n7498), .B2(n4620), .A(n4619), .ZN(n7610) );
  NAND2_X1 U5012 ( .A1(n4439), .A2(n7067), .ZN(n4288) );
  OAI21_X2 U5013 ( .B1(n9179), .B2(n9178), .A(n9177), .ZN(n9180) );
  NAND2_X2 U5014 ( .A1(n7483), .A2(n5811), .ZN(n5812) );
  NAND2_X1 U5015 ( .A1(n10002), .A2(n5674), .ZN(n4289) );
  BUF_X2 U5016 ( .A(n5578), .Z(n4291) );
  OAI211_X1 U5017 ( .C1(n6316), .C2(n7492), .A(n5955), .B(n5954), .ZN(n10118)
         );
  INV_X1 U5018 ( .A(n5838), .ZN(n6308) );
  NOR2_X4 U5019 ( .A1(n5099), .A2(n4987), .ZN(n5138) );
  XNOR2_X2 U5020 ( .A(n5928), .B(n9077), .ZN(n5927) );
  AOI21_X2 U5021 ( .B1(n5817), .B2(n5982), .A(n4622), .ZN(n4619) );
  NOR2_X2 U5022 ( .A1(n5413), .A2(n10221), .ZN(n4446) );
  OR2_X2 U5023 ( .A1(n5400), .A2(n9270), .ZN(n5413) );
  NAND4_X2 U5024 ( .A1(n4597), .A2(n4778), .A3(n4779), .A4(n4941), .ZN(n5099)
         );
  INV_X4 U5025 ( .A(n6229), .ZN(n5988) );
  NAND2_X1 U5026 ( .A1(n4940), .A2(n4452), .ZN(n5640) );
  AND2_X1 U5027 ( .A1(n4289), .A2(n5118), .ZN(n4294) );
  OR2_X1 U5028 ( .A1(n9861), .A2(n9335), .ZN(n6614) );
  AND2_X1 U5029 ( .A1(n5699), .A2(n5694), .ZN(n4675) );
  INV_X1 U5030 ( .A(n5190), .ZN(n4868) );
  NOR2_X1 U5031 ( .A1(n6975), .A2(n6962), .ZN(n6991) );
  NOR2_X1 U5032 ( .A1(n6961), .A2(n4365), .ZN(n6962) );
  XNOR2_X1 U5033 ( .A(n5928), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U5034 ( .A1(n9084), .A2(n5930), .ZN(n5950) );
  OR2_X1 U5035 ( .A1(n8460), .A2(n8551), .ZN(n7004) );
  AOI21_X1 U5036 ( .B1(n4718), .B2(n4717), .A(n4303), .ZN(n4716) );
  INV_X1 U5037 ( .A(n6287), .ZN(n4717) );
  NAND2_X1 U5038 ( .A1(n8776), .A2(n4533), .ZN(n6942) );
  INV_X1 U5039 ( .A(n8995), .ZN(n4533) );
  INV_X1 U5040 ( .A(n9290), .ZN(n4805) );
  NAND2_X1 U5041 ( .A1(n8324), .A2(n8325), .ZN(n4819) );
  NOR2_X1 U5042 ( .A1(n4557), .A2(n9652), .ZN(n4555) );
  AND2_X1 U5043 ( .A1(n4546), .A2(n4363), .ZN(n4544) );
  INV_X1 U5044 ( .A(n4825), .ZN(n4824) );
  INV_X1 U5045 ( .A(n8776), .ZN(n6502) );
  NOR2_X1 U5046 ( .A1(n8603), .A2(n4492), .ZN(n4490) );
  INV_X1 U5047 ( .A(n5957), .ZN(n6231) );
  NAND2_X1 U5048 ( .A1(n6948), .A2(n6292), .ZN(n8758) );
  NAND2_X1 U5049 ( .A1(n4671), .A2(n5712), .ZN(n4389) );
  INV_X1 U5050 ( .A(n6660), .ZN(n4835) );
  NOR2_X1 U5051 ( .A1(n6784), .A2(n4837), .ZN(n4836) );
  INV_X1 U5052 ( .A(n5520), .ZN(n4837) );
  NAND2_X1 U5053 ( .A1(n4558), .A2(n6755), .ZN(n4557) );
  NAND2_X1 U5054 ( .A1(n4972), .A2(n4559), .ZN(n4558) );
  INV_X1 U5055 ( .A(n6757), .ZN(n4559) );
  NAND2_X1 U5056 ( .A1(n6591), .A2(n6597), .ZN(n4416) );
  AND2_X1 U5057 ( .A1(n6596), .A2(n6710), .ZN(n4454) );
  NAND2_X1 U5058 ( .A1(n6661), .A2(n6663), .ZN(n4456) );
  AOI211_X1 U5059 ( .C1(n6936), .C2(n6949), .A(n6935), .B(n8758), .ZN(n6937)
         );
  NOR4_X1 U5060 ( .A1(n6244), .A2(n7524), .A3(n7624), .A4(n6385), .ZN(n7002)
         );
  OR2_X1 U5061 ( .A1(n7184), .A2(n4788), .ZN(n4786) );
  NAND2_X1 U5062 ( .A1(n6587), .A2(n6577), .ZN(n6583) );
  INV_X1 U5063 ( .A(n5337), .ZN(n5338) );
  OAI21_X1 U5064 ( .B1(n4869), .B2(n4868), .A(n4977), .ZN(n4867) );
  INV_X1 U5065 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6111) );
  AND2_X1 U5066 ( .A1(n8075), .A2(n4697), .ZN(n4696) );
  NAND2_X1 U5067 ( .A1(n4310), .A2(n6264), .ZN(n4697) );
  NAND2_X1 U5068 ( .A1(n7630), .A2(n8615), .ZN(n6842) );
  NAND2_X1 U5069 ( .A1(n10118), .A2(n6247), .ZN(n6843) );
  NAND2_X1 U5070 ( .A1(n5936), .A2(n5935), .ZN(n6839) );
  OAI22_X1 U5071 ( .A1(n6326), .A2(P2_D_REG_0__SCAN_IN), .B1(n7361), .B2(n7365), .ZN(n6387) );
  NOR2_X1 U5072 ( .A1(n4328), .A2(n4873), .ZN(n4872) );
  INV_X1 U5073 ( .A(n6284), .ZN(n4873) );
  AND2_X1 U5074 ( .A1(n4709), .A2(n8823), .ZN(n4706) );
  OR2_X1 U5075 ( .A1(n9019), .A2(n8496), .ZN(n8790) );
  AOI21_X1 U5076 ( .B1(n7219), .B2(n7199), .A(n9184), .ZN(n7228) );
  NOR2_X1 U5077 ( .A1(n4818), .A2(n7163), .ZN(n4814) );
  AOI21_X1 U5078 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9527), .A(n10008), .ZN(
        n9529) );
  OR2_X1 U5079 ( .A1(n6668), .A2(n7272), .ZN(n6807) );
  NAND2_X1 U5080 ( .A1(n7321), .A2(n4947), .ZN(n6699) );
  NAND2_X1 U5081 ( .A1(n8432), .A2(n9349), .ZN(n6748) );
  OR2_X1 U5082 ( .A1(n8432), .A2(n9349), .ZN(n6809) );
  INV_X1 U5083 ( .A(n4775), .ZN(n4773) );
  NAND2_X1 U5084 ( .A1(n4944), .A2(n4942), .ZN(n9612) );
  INV_X1 U5085 ( .A(n4943), .ZN(n4942) );
  OAI21_X1 U5086 ( .B1(n5665), .B2(n4945), .A(n9607), .ZN(n4943) );
  OR2_X1 U5087 ( .A1(n9922), .A2(n9292), .ZN(n6642) );
  AND2_X1 U5088 ( .A1(n9776), .A2(n6614), .ZN(n4952) );
  NAND2_X1 U5089 ( .A1(n6569), .A2(n6703), .ZN(n6761) );
  NAND2_X1 U5090 ( .A1(n6539), .A2(n8188), .ZN(n5686) );
  AND2_X1 U5091 ( .A1(n5563), .A2(n5528), .ZN(n5538) );
  AND2_X1 U5092 ( .A1(n5524), .A2(n5510), .ZN(n5522) );
  AND2_X1 U5093 ( .A1(n5506), .A2(n5488), .ZN(n5504) );
  INV_X1 U5094 ( .A(SI_19_), .ZN(n5379) );
  AOI21_X1 U5095 ( .B1(n4496), .B2(n4495), .A(n4353), .ZN(n4494) );
  AOI21_X1 U5096 ( .B1(n4876), .B2(n4878), .A(n4875), .ZN(n4874) );
  INV_X1 U5097 ( .A(n5362), .ZN(n4875) );
  INV_X1 U5098 ( .A(n4881), .ZN(n4876) );
  AOI21_X1 U5099 ( .B1(n4856), .B2(n4859), .A(n4351), .ZN(n4853) );
  XNOR2_X1 U5100 ( .A(n6396), .B(n7454), .ZN(n6388) );
  NOR2_X1 U5101 ( .A1(n4927), .A2(n4333), .ZN(n4926) );
  NOR2_X1 U5102 ( .A1(n6466), .A2(n4930), .ZN(n4927) );
  OR2_X1 U5103 ( .A1(n6982), .A2(n6981), .ZN(n6983) );
  NAND2_X1 U5104 ( .A1(n4647), .A2(n7028), .ZN(n4646) );
  INV_X1 U5105 ( .A(n8212), .ZN(n7031) );
  INV_X1 U5106 ( .A(n7768), .ZN(n4746) );
  NAND2_X1 U5107 ( .A1(n8655), .A2(n8654), .ZN(n8653) );
  NOR2_X1 U5108 ( .A1(n8883), .A2(n4906), .ZN(n4905) );
  INV_X1 U5109 ( .A(n6903), .ZN(n4906) );
  AND4_X1 U5110 ( .A1(n6033), .A2(n6032), .A3(n6031), .A4(n6030), .ZN(n8551)
         );
  NAND2_X1 U5111 ( .A1(n10097), .A2(n4614), .ZN(n4912) );
  NOR2_X1 U5112 ( .A1(n6858), .A2(n4615), .ZN(n4614) );
  INV_X1 U5113 ( .A(n6859), .ZN(n4615) );
  NAND2_X1 U5114 ( .A1(n6492), .A2(n7430), .ZN(n6495) );
  OR2_X1 U5115 ( .A1(n6980), .A2(n6480), .ZN(n8896) );
  AND2_X1 U5116 ( .A1(n4892), .A2(n6953), .ZN(n4893) );
  NAND2_X1 U5117 ( .A1(n6942), .A2(n6941), .ZN(n4892) );
  NOR2_X1 U5118 ( .A1(n6293), .A2(n4884), .ZN(n4883) );
  INV_X1 U5119 ( .A(n6291), .ZN(n4884) );
  NAND2_X1 U5120 ( .A1(n6942), .A2(n6953), .ZN(n8766) );
  OR2_X1 U5121 ( .A1(n8590), .A2(n8510), .ZN(n6903) );
  INV_X1 U5122 ( .A(n8898), .ZN(n10093) );
  NAND2_X1 U5123 ( .A1(n5712), .A2(n4910), .ZN(n5922) );
  NOR2_X1 U5124 ( .A1(n5724), .A2(n4518), .ZN(n4517) );
  NAND2_X1 U5125 ( .A1(n4522), .A2(n5718), .ZN(n4518) );
  XNOR2_X1 U5126 ( .A(n5620), .B(n5619), .ZN(n7442) );
  NAND2_X1 U5127 ( .A1(n5626), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5620) );
  OR2_X1 U5128 ( .A1(n7238), .A2(n4805), .ZN(n4802) );
  AND2_X1 U5129 ( .A1(n7238), .A2(n4805), .ZN(n4804) );
  OAI21_X1 U5130 ( .B1(n7110), .B2(n7334), .A(n7074), .ZN(n7075) );
  INV_X1 U5131 ( .A(n9324), .ZN(n9336) );
  AND2_X1 U5132 ( .A1(n7443), .A2(n5674), .ZN(n9324) );
  XNOR2_X1 U5133 ( .A(n9552), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9563) );
  AOI21_X1 U5134 ( .B1(n4572), .B2(n4571), .A(n4570), .ZN(n4569) );
  INV_X1 U5135 ( .A(n9551), .ZN(n4570) );
  NOR2_X1 U5136 ( .A1(n4775), .A2(n4777), .ZN(n4774) );
  NAND2_X1 U5137 ( .A1(n9605), .A2(n5501), .ZN(n5503) );
  INV_X1 U5138 ( .A(n5298), .ZN(n4828) );
  NAND2_X1 U5139 ( .A1(n6809), .A2(n6748), .ZN(n6786) );
  NAND2_X1 U5140 ( .A1(n6642), .A2(n6727), .ZN(n9642) );
  INV_X1 U5141 ( .A(n4555), .ZN(n4553) );
  INV_X1 U5142 ( .A(n4560), .ZN(n4552) );
  NAND2_X1 U5143 ( .A1(n4544), .A2(n4825), .ZN(n4543) );
  AOI21_X1 U5144 ( .B1(n7427), .B2(n5605), .A(n7429), .ZN(n7327) );
  NAND2_X1 U5145 ( .A1(n5673), .A2(n6824), .ZN(n9778) );
  NAND2_X1 U5146 ( .A1(n6515), .A2(n6514), .ZN(n6522) );
  AND2_X1 U5147 ( .A1(n5467), .A2(n5452), .ZN(n5465) );
  NAND2_X1 U5148 ( .A1(n6398), .A2(n6397), .ZN(n7649) );
  NAND2_X1 U5149 ( .A1(n4523), .A2(n4931), .ZN(n6459) );
  AND2_X1 U5150 ( .A1(n6216), .A2(n6215), .ZN(n8584) );
  NAND2_X1 U5151 ( .A1(n6227), .A2(n6226), .ZN(n8759) );
  OR2_X1 U5152 ( .A1(n10006), .A2(n7554), .ZN(n10034) );
  AND2_X1 U5153 ( .A1(n8155), .A2(n6703), .ZN(n4388) );
  OR2_X1 U5154 ( .A1(n6870), .A2(n6869), .ZN(n6873) );
  NAND2_X1 U5155 ( .A1(n6599), .A2(n6826), .ZN(n4414) );
  NOR2_X1 U5156 ( .A1(n4400), .A2(n7971), .ZN(n4399) );
  NAND2_X1 U5157 ( .A1(n4402), .A2(n4401), .ZN(n4400) );
  NOR2_X1 U5158 ( .A1(n7786), .A2(n7796), .ZN(n4402) );
  INV_X1 U5159 ( .A(n7993), .ZN(n4398) );
  AND2_X1 U5160 ( .A1(n6675), .A2(n6672), .ZN(n4413) );
  AOI21_X1 U5161 ( .B1(n6551), .B2(n4441), .A(n4440), .ZN(n6674) );
  NOR2_X1 U5162 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  NAND2_X1 U5163 ( .A1(n6549), .A2(n6550), .ZN(n4440) );
  NAND2_X1 U5164 ( .A1(n6807), .A2(n6826), .ZN(n4442) );
  INV_X1 U5165 ( .A(n7778), .ZN(n4627) );
  NOR2_X1 U5166 ( .A1(n4719), .A2(n4714), .ZN(n4713) );
  INV_X1 U5167 ( .A(n6286), .ZN(n4714) );
  INV_X1 U5168 ( .A(n6802), .ZN(n4961) );
  AND2_X1 U5169 ( .A1(n4992), .A2(n10207), .ZN(n4822) );
  INV_X1 U5170 ( .A(n5321), .ZN(n5324) );
  INV_X1 U5171 ( .A(SI_15_), .ZN(n5323) );
  AOI21_X1 U5172 ( .B1(n4858), .B2(n4857), .A(n5285), .ZN(n4856) );
  INV_X1 U5173 ( .A(n4861), .ZN(n4857) );
  INV_X1 U5174 ( .A(n5145), .ZN(n4851) );
  AND2_X1 U5175 ( .A1(n8534), .A2(n6450), .ZN(n4934) );
  OR2_X1 U5176 ( .A1(n6220), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6230) );
  NOR2_X1 U5177 ( .A1(n6168), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6178) );
  INV_X1 U5178 ( .A(n6113), .ZN(n6112) );
  INV_X1 U5179 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4540) );
  AND2_X1 U5180 ( .A1(n6071), .A2(n4537), .ZN(n4536) );
  INV_X1 U5181 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4537) );
  INV_X1 U5182 ( .A(n6073), .ZN(n6072) );
  NAND2_X1 U5183 ( .A1(n4679), .A2(n4681), .ZN(n10081) );
  AOI21_X1 U5184 ( .B1(n7786), .B2(n4682), .A(n4347), .ZN(n4681) );
  NOR2_X1 U5185 ( .A1(n6326), .A2(n6340), .ZN(n6352) );
  OR2_X1 U5186 ( .A1(n6980), .A2(n6384), .ZN(n6491) );
  AOI21_X1 U5187 ( .B1(n4603), .B2(n6932), .A(n4601), .ZN(n4600) );
  OR2_X1 U5188 ( .A1(n9001), .A2(n6469), .ZN(n6938) );
  NAND2_X1 U5189 ( .A1(n4904), .A2(n6924), .ZN(n4901) );
  NOR2_X1 U5190 ( .A1(n6929), .A2(n4903), .ZN(n4902) );
  INV_X1 U5191 ( .A(n6924), .ZN(n4903) );
  NAND2_X1 U5192 ( .A1(n9025), .A2(n6456), .ZN(n6925) );
  INV_X1 U5193 ( .A(n9025), .ZN(n4848) );
  OR2_X1 U5194 ( .A1(n8861), .A2(n6274), .ZN(n4708) );
  OR2_X1 U5195 ( .A1(n9059), .A2(n8897), .ZN(n6901) );
  INV_X1 U5196 ( .A(n4890), .ZN(n4889) );
  OAI21_X1 U5197 ( .B1(n8193), .B2(n4891), .A(n6079), .ZN(n4890) );
  INV_X1 U5198 ( .A(n6068), .ZN(n4891) );
  OR2_X1 U5199 ( .A1(n7305), .A2(n6352), .ZN(n6497) );
  NAND2_X1 U5200 ( .A1(n6325), .A2(n7365), .ZN(n6326) );
  INV_X1 U5201 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5701) );
  AND2_X1 U5202 ( .A1(n5718), .A2(n5801), .ZN(n4521) );
  INV_X1 U5203 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4522) );
  INV_X1 U5204 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5718) );
  INV_X1 U5205 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5722) );
  INV_X1 U5206 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5746) );
  NOR2_X1 U5207 ( .A1(n5766), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U5208 ( .A1(n4677), .A2(n5694), .ZN(n5766) );
  AND2_X1 U5209 ( .A1(n4975), .A2(n4785), .ZN(n4784) );
  NAND2_X1 U5210 ( .A1(n4787), .A2(n4786), .ZN(n4785) );
  NAND2_X1 U5211 ( .A1(n7215), .A2(n7214), .ZN(n7216) );
  AND2_X1 U5212 ( .A1(n4792), .A2(n9206), .ZN(n4791) );
  OR2_X1 U5213 ( .A1(n4793), .A2(n9237), .ZN(n4792) );
  INV_X1 U5214 ( .A(n7253), .ZN(n4793) );
  OR2_X1 U5215 ( .A1(n5179), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5213) );
  INV_X1 U5216 ( .A(n7287), .ZN(n7443) );
  NAND2_X1 U5217 ( .A1(n6765), .A2(n6766), .ZN(n5647) );
  NAND2_X1 U5218 ( .A1(n4404), .A2(n4325), .ZN(n6768) );
  INV_X1 U5219 ( .A(n6583), .ZN(n4404) );
  NAND2_X1 U5220 ( .A1(n6592), .A2(n8158), .ZN(n6764) );
  OR2_X1 U5221 ( .A1(n9259), .A2(n7143), .ZN(n6587) );
  AOI21_X1 U5222 ( .B1(n7933), .B2(n4956), .A(n4955), .ZN(n4954) );
  INV_X1 U5223 ( .A(n6568), .ZN(n4956) );
  NAND2_X1 U5224 ( .A1(n7818), .A2(n7817), .ZN(n5643) );
  INV_X1 U5225 ( .A(n9621), .ZN(n4946) );
  OR2_X1 U5226 ( .A1(n9847), .A2(n9313), .ZN(n6630) );
  OR2_X1 U5227 ( .A1(n8354), .A2(n8304), .ZN(n6597) );
  NAND2_X1 U5228 ( .A1(n5560), .A2(n5563), .ZN(n6511) );
  AND2_X1 U5229 ( .A1(n5561), .A2(n5565), .ZN(n6510) );
  NAND2_X1 U5230 ( .A1(n4986), .A2(n5120), .ZN(n4987) );
  INV_X1 U5231 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4986) );
  INV_X1 U5232 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4597) );
  INV_X1 U5233 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4779) );
  INV_X1 U5234 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n4941) );
  AOI21_X1 U5235 ( .B1(n5522), .B2(n4466), .A(n4465), .ZN(n4464) );
  INV_X1 U5236 ( .A(n5524), .ZN(n4465) );
  INV_X1 U5237 ( .A(n5506), .ZN(n4466) );
  INV_X1 U5238 ( .A(n5522), .ZN(n4467) );
  AOI21_X1 U5239 ( .B1(n4475), .B2(n4477), .A(n4472), .ZN(n4471) );
  INV_X1 U5240 ( .A(n5467), .ZN(n4472) );
  AND2_X1 U5241 ( .A1(n5483), .A2(n5471), .ZN(n5481) );
  NAND2_X1 U5242 ( .A1(n5450), .A2(n5449), .ZN(n5467) );
  INV_X1 U5243 ( .A(SI_23_), .ZN(n5449) );
  INV_X1 U5244 ( .A(n5446), .ZN(n4482) );
  INV_X1 U5245 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5592) );
  NAND4_X1 U5246 ( .A1(n4988), .A2(n5138), .A3(n5346), .A4(n4822), .ZN(n5595)
         );
  INV_X1 U5247 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5346) );
  OR2_X1 U5248 ( .A1(n5252), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n5253) );
  INV_X1 U5249 ( .A(SI_11_), .ZN(n5234) );
  NAND2_X1 U5250 ( .A1(n5176), .A2(n5175), .ZN(n5190) );
  INV_X1 U5251 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n4985) );
  INV_X1 U5252 ( .A(n6462), .ZN(n8523) );
  NOR2_X1 U5253 ( .A1(n6466), .A2(n4929), .ZN(n4928) );
  INV_X1 U5254 ( .A(n8543), .ZN(n4929) );
  OR2_X1 U5255 ( .A1(n6980), .A2(n6242), .ZN(n6496) );
  AND2_X1 U5256 ( .A1(n8593), .A2(n6435), .ZN(n4938) );
  AND4_X1 U5257 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n8102)
         );
  AOI21_X1 U5258 ( .B1(n7587), .B2(n5754), .A(n5753), .ZN(n7581) );
  NAND2_X1 U5259 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n4624), .ZN(n4623) );
  OR2_X1 U5260 ( .A1(n5773), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U5261 ( .A1(n7765), .A2(n5780), .ZN(n5783) );
  XNOR2_X1 U5262 ( .A(n5796), .B(n4628), .ZN(n8670) );
  NAND2_X1 U5263 ( .A1(n8670), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U5264 ( .A1(n8653), .A2(n5827), .ZN(n5828) );
  NAND2_X1 U5265 ( .A1(n8717), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U5266 ( .A1(n6178), .A2(n4532), .ZN(n6199) );
  NAND2_X1 U5267 ( .A1(n6112), .A2(n4306), .ZN(n6130) );
  AOI21_X1 U5268 ( .B1(n4689), .B2(n4687), .A(n4315), .ZN(n4686) );
  INV_X1 U5269 ( .A(n6269), .ZN(n4687) );
  INV_X1 U5270 ( .A(n4696), .ZN(n4695) );
  AOI21_X1 U5271 ( .B1(n4696), .B2(n4694), .A(n4340), .ZN(n4693) );
  INV_X1 U5272 ( .A(n6264), .ZN(n4694) );
  AND4_X1 U5273 ( .A1(n6056), .A2(n6055), .A3(n6054), .A4(n6053), .ZN(n8455)
         );
  OR2_X1 U5274 ( .A1(n6019), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U5275 ( .A1(n7626), .A2(n7624), .ZN(n6249) );
  NAND2_X1 U5276 ( .A1(n5940), .A2(n5939), .ZN(n4655) );
  OR2_X1 U5277 ( .A1(n6980), .A2(n6483), .ZN(n8898) );
  OR2_X1 U5278 ( .A1(n4318), .A2(n8758), .ZN(n4729) );
  NAND2_X1 U5279 ( .A1(n8759), .A2(n10091), .ZN(n4727) );
  NAND2_X1 U5280 ( .A1(n4602), .A2(n4600), .ZN(n8782) );
  NAND2_X1 U5281 ( .A1(n4701), .A2(n4699), .ZN(n6285) );
  AOI21_X1 U5282 ( .B1(n4702), .B2(n4705), .A(n4700), .ZN(n4699) );
  INV_X1 U5283 ( .A(n8811), .ZN(n4700) );
  NOR2_X1 U5284 ( .A1(n8794), .A2(n6997), .ZN(n8802) );
  INV_X1 U5285 ( .A(n4706), .ZN(n4705) );
  AND2_X1 U5286 ( .A1(n4703), .A2(n4711), .ZN(n4702) );
  NAND2_X1 U5287 ( .A1(n4706), .A2(n4704), .ZN(n4703) );
  AND2_X1 U5288 ( .A1(n6282), .A2(n6281), .ZN(n4711) );
  INV_X1 U5289 ( .A(n6273), .ZN(n4704) );
  AND2_X1 U5290 ( .A1(n6275), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U5291 ( .A1(n6274), .A2(n6273), .ZN(n4710) );
  NAND2_X1 U5292 ( .A1(n8861), .A2(n6273), .ZN(n4707) );
  NAND2_X1 U5293 ( .A1(n6277), .A2(n6451), .ZN(n6924) );
  NAND2_X1 U5294 ( .A1(n6927), .A2(n6924), .ZN(n8835) );
  AOI21_X1 U5295 ( .B1(n4611), .B2(n4613), .A(n6918), .ZN(n4609) );
  NAND2_X1 U5296 ( .A1(n4909), .A2(n4611), .ZN(n4610) );
  INV_X1 U5297 ( .A(n4612), .ZN(n4611) );
  NAND2_X1 U5298 ( .A1(n6917), .A2(n6916), .ZN(n8844) );
  OR2_X1 U5299 ( .A1(n8948), .A2(n8568), .ZN(n8859) );
  NAND2_X1 U5300 ( .A1(n6093), .A2(n6092), .ZN(n8590) );
  NAND2_X1 U5301 ( .A1(n8189), .A2(n8193), .ZN(n8191) );
  OAI21_X1 U5302 ( .B1(n6044), .B2(n7005), .A(n7003), .ZN(n6045) );
  NAND2_X1 U5303 ( .A1(n5712), .A2(n4939), .ZN(n5714) );
  NOR2_X1 U5304 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4939) );
  XNOR2_X1 U5305 ( .A(n5728), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7036) );
  NAND2_X1 U5306 ( .A1(n6240), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5726) );
  INV_X1 U5307 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5794) );
  AND2_X1 U5308 ( .A1(n9114), .A2(n4802), .ZN(n4801) );
  AND2_X1 U5309 ( .A1(n9218), .A2(n9217), .ZN(n9148) );
  INV_X1 U5310 ( .A(n5491), .ZN(n5493) );
  OAI22_X1 U5311 ( .A1(n9974), .A2(n7273), .B1(n7143), .B2(n8403), .ZN(n9248)
         );
  NAND2_X1 U5312 ( .A1(n4446), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5457) );
  INV_X1 U5313 ( .A(n9355), .ZN(n9118) );
  NAND2_X1 U5314 ( .A1(n8340), .A2(n7065), .ZN(n7066) );
  INV_X1 U5315 ( .A(n7162), .ZN(n4811) );
  INV_X1 U5316 ( .A(n4820), .ZN(n4812) );
  INV_X1 U5317 ( .A(n4814), .ZN(n4813) );
  INV_X1 U5318 ( .A(n9152), .ZN(n4390) );
  INV_X1 U5319 ( .A(n8200), .ZN(n4798) );
  NAND2_X1 U5320 ( .A1(n9147), .A2(n9146), .ZN(n9215) );
  NAND2_X1 U5321 ( .A1(n7064), .A2(n7062), .ZN(n7287) );
  AND2_X1 U5322 ( .A1(n5463), .A2(n5462), .ZN(n9292) );
  OR2_X1 U5323 ( .A1(n6530), .A2(n5066), .ZN(n5067) );
  INV_X1 U5324 ( .A(n7548), .ZN(n4593) );
  INV_X1 U5325 ( .A(n7547), .ZN(n4589) );
  OAI21_X1 U5326 ( .B1(n9415), .B2(n4593), .A(n9425), .ZN(n4592) );
  NOR2_X1 U5327 ( .A1(n5216), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5238) );
  CLKBUF_X1 U5328 ( .A(n5138), .Z(n5139) );
  OR2_X1 U5329 ( .A1(n4587), .A2(n10029), .ZN(n4586) );
  NAND2_X1 U5330 ( .A1(n4586), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U5331 ( .A1(n9548), .A2(n9547), .ZN(n4575) );
  NAND2_X1 U5332 ( .A1(n9598), .A2(n9908), .ZN(n6379) );
  NOR2_X1 U5333 ( .A1(n4840), .A2(n5521), .ZN(n4839) );
  INV_X1 U5334 ( .A(n5502), .ZN(n4840) );
  NOR2_X1 U5335 ( .A1(n4561), .A2(n6757), .ZN(n4560) );
  INV_X1 U5336 ( .A(n5406), .ZN(n4561) );
  NOR2_X1 U5337 ( .A1(n4951), .A2(n4949), .ZN(n4948) );
  INV_X1 U5338 ( .A(n9738), .ZN(n4949) );
  INV_X1 U5339 ( .A(n5299), .ZN(n4831) );
  NAND2_X1 U5340 ( .A1(n8302), .A2(n6713), .ZN(n8359) );
  AOI21_X1 U5341 ( .B1(n7892), .B2(n7896), .A(n5150), .ZN(n5151) );
  OR2_X1 U5342 ( .A1(n9369), .A2(n9172), .ZN(n5187) );
  NAND2_X1 U5343 ( .A1(n9797), .A2(n8188), .ZN(n9784) );
  NAND2_X1 U5344 ( .A1(n6568), .A2(n7820), .ZN(n7926) );
  NAND2_X1 U5345 ( .A1(n5643), .A2(n6759), .ZN(n7820) );
  INV_X1 U5346 ( .A(n9778), .ZN(n9757) );
  OR2_X1 U5347 ( .A1(n6534), .A2(n5016), .ZN(n5017) );
  INV_X1 U5348 ( .A(n7445), .ZN(n7296) );
  NAND2_X1 U5349 ( .A1(n7322), .A2(n6760), .ZN(n7321) );
  AND2_X1 U5350 ( .A1(n8340), .A2(n8301), .ZN(n9797) );
  NAND2_X1 U5351 ( .A1(n6517), .A2(n6516), .ZN(n9567) );
  INV_X1 U5352 ( .A(n4551), .ZN(n4549) );
  OR2_X1 U5353 ( .A1(n6757), .A2(n6756), .ZN(n9674) );
  NOR2_X1 U5354 ( .A1(n5405), .A2(n5404), .ZN(n4972) );
  AND2_X1 U5355 ( .A1(n6630), .A2(n6690), .ZN(n9705) );
  AOI21_X1 U5356 ( .B1(n4824), .B2(n4826), .A(n4335), .ZN(n4546) );
  AND2_X1 U5357 ( .A1(n9721), .A2(n6627), .ZN(n9738) );
  AND2_X1 U5358 ( .A1(n6611), .A2(n9752), .ZN(n9776) );
  AND2_X1 U5359 ( .A1(n7825), .A2(n6761), .ZN(n5127) );
  OR2_X1 U5360 ( .A1(n7710), .A2(n7070), .ZN(n7445) );
  AND2_X1 U5361 ( .A1(n5604), .A2(n5621), .ZN(n7427) );
  XNOR2_X1 U5362 ( .A(n6522), .B(n6521), .ZN(n8424) );
  NAND2_X1 U5363 ( .A1(n5573), .A2(SI_29_), .ZN(n6515) );
  XNOR2_X1 U5364 ( .A(n6511), .B(n6510), .ZN(n8396) );
  NAND2_X1 U5365 ( .A1(n5507), .A2(n5506), .ZN(n5523) );
  NOR2_X1 U5366 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n4990) );
  AOI21_X1 U5367 ( .B1(n4480), .B2(n5429), .A(n4479), .ZN(n4478) );
  INV_X1 U5368 ( .A(n5445), .ZN(n4479) );
  OAI21_X1 U5369 ( .B1(n5430), .B2(n5429), .A(n5428), .ZN(n5447) );
  XNOR2_X1 U5370 ( .A(n5410), .B(n5409), .ZN(n6145) );
  NAND2_X1 U5371 ( .A1(n4498), .A2(n4874), .ZN(n5378) );
  NAND2_X1 U5372 ( .A1(n5305), .A2(n4499), .ZN(n4498) );
  NAND2_X1 U5373 ( .A1(n4880), .A2(n5339), .ZN(n5361) );
  NAND2_X1 U5374 ( .A1(n5326), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U5375 ( .A1(n4489), .A2(n4863), .ZN(n5233) );
  NAND2_X1 U5376 ( .A1(n4852), .A2(n5145), .ZN(n5163) );
  NAND2_X1 U5377 ( .A1(n5143), .A2(n5142), .ZN(n4852) );
  NAND2_X1 U5378 ( .A1(n9983), .A2(n4985), .ZN(n4596) );
  NAND2_X1 U5379 ( .A1(n5038), .A2(n4985), .ZN(n5039) );
  NOR2_X1 U5380 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5038) );
  AND4_X1 U5381 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n7533)
         );
  INV_X1 U5382 ( .A(n8871), .ZN(n8469) );
  NAND2_X1 U5383 ( .A1(n4286), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4606) );
  AND2_X1 U5384 ( .A1(n6185), .A2(n6184), .ZN(n8526) );
  NAND2_X1 U5385 ( .A1(n8506), .A2(n6441), .ZN(n8516) );
  NAND2_X1 U5386 ( .A1(n7649), .A2(n6404), .ZN(n7650) );
  NAND2_X1 U5387 ( .A1(n7432), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U5388 ( .A1(n4916), .A2(n4917), .ZN(n8574) );
  AND2_X1 U5389 ( .A1(n8569), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U5390 ( .A1(n8516), .A2(n8570), .ZN(n4916) );
  NAND2_X1 U5391 ( .A1(n8517), .A2(n8570), .ZN(n4918) );
  NAND2_X1 U5392 ( .A1(n4921), .A2(n4920), .ZN(n8578) );
  AOI21_X1 U5393 ( .B1(n4301), .B2(n4925), .A(n4327), .ZN(n4920) );
  NAND2_X1 U5394 ( .A1(n6479), .A2(n8874), .ZN(n8586) );
  INV_X1 U5395 ( .A(n8586), .ZN(n8602) );
  AND2_X1 U5396 ( .A1(n8019), .A2(n6994), .ZN(n4638) );
  NAND2_X1 U5397 ( .A1(n4313), .A2(n8019), .ZN(n4645) );
  NAND2_X1 U5398 ( .A1(n4617), .A2(n4968), .ZN(n4460) );
  XNOR2_X1 U5399 ( .A(n7029), .B(n7028), .ZN(n4617) );
  NAND2_X1 U5400 ( .A1(n4534), .A2(n6204), .ZN(n8776) );
  NAND2_X1 U5401 ( .A1(n8771), .A2(n6231), .ZN(n4534) );
  INV_X1 U5402 ( .A(n8526), .ZN(n8803) );
  INV_X1 U5403 ( .A(n8788), .ZN(n8812) );
  NAND2_X1 U5404 ( .A1(n6173), .A2(n6172), .ZN(n8825) );
  NAND2_X1 U5405 ( .A1(n6144), .A2(n6143), .ZN(n8850) );
  INV_X1 U5406 ( .A(n8551), .ZN(n8609) );
  XNOR2_X1 U5407 ( .A(n5828), .B(n4628), .ZN(n8683) );
  NAND2_X1 U5408 ( .A1(n8683), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U5409 ( .A1(n8705), .A2(n8704), .ZN(n8703) );
  AND2_X1 U5410 ( .A1(n7459), .A2(n5895), .ZN(n8723) );
  INV_X1 U5411 ( .A(n8747), .ZN(n4756) );
  INV_X1 U5412 ( .A(n4755), .ZN(n4754) );
  AOI21_X1 U5413 ( .B1(n8736), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8735), .ZN(
        n4755) );
  NAND2_X1 U5414 ( .A1(n4909), .A2(n4297), .ZN(n8950) );
  AND2_X1 U5415 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  NAND2_X1 U5416 ( .A1(n6236), .A2(n8967), .ZN(n6364) );
  NAND2_X1 U5417 ( .A1(n6207), .A2(n6206), .ZN(n8989) );
  NAND2_X1 U5418 ( .A1(n4715), .A2(n4718), .ZN(n6290) );
  NAND2_X1 U5419 ( .A1(n6157), .A2(n6156), .ZN(n9013) );
  NAND2_X1 U5420 ( .A1(n6239), .A2(n6240), .ZN(n8212) );
  OR2_X1 U5421 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  INV_X1 U5422 ( .A(n9345), .ZN(n9302) );
  NAND2_X1 U5423 ( .A1(n6793), .A2(n6792), .ZN(n6794) );
  OR2_X1 U5424 ( .A1(n5372), .A2(n5371), .ZN(n9359) );
  NAND2_X1 U5425 ( .A1(n9437), .A2(n4331), .ZN(n9451) );
  AOI21_X1 U5426 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n9540), .A(n9538), .ZN(
        n9548) );
  OAI21_X1 U5427 ( .B1(n9561), .B2(n10034), .A(n10043), .ZN(n4409) );
  OAI22_X1 U5428 ( .A1(n9563), .A2(n10034), .B1(n9562), .B2(n10022), .ZN(n4578) );
  NOR2_X1 U5429 ( .A1(n8434), .A2(n8433), .ZN(n4421) );
  AOI21_X1 U5430 ( .B1(n5916), .B2(n9778), .A(n7295), .ZN(n9590) );
  NAND2_X1 U5431 ( .A1(n9596), .A2(n9595), .ZN(n9812) );
  NAND2_X1 U5432 ( .A1(n5503), .A2(n5502), .ZN(n9591) );
  CLKBUF_X1 U5433 ( .A(n9712), .Z(n10337) );
  XNOR2_X1 U5434 ( .A(n5587), .B(n6786), .ZN(n8436) );
  AOI21_X1 U5435 ( .B1(n9572), .B2(n10061), .A(n9573), .ZN(n4438) );
  NOR2_X1 U5436 ( .A1(n9812), .A2(n4383), .ZN(n9909) );
  NAND2_X1 U5437 ( .A1(n4385), .A2(n4384), .ZN(n4383) );
  NAND2_X1 U5438 ( .A1(n9814), .A2(n10064), .ZN(n4384) );
  INV_X1 U5439 ( .A(n9813), .ZN(n4385) );
  NAND2_X1 U5440 ( .A1(n5454), .A2(n5453), .ZN(n9922) );
  INV_X1 U5441 ( .A(n7062), .ZN(n8301) );
  CLKBUF_X1 U5442 ( .A(n6539), .Z(n9564) );
  NOR2_X1 U5443 ( .A1(n8131), .A2(n8130), .ZN(n10189) );
  NOR2_X1 U5444 ( .A1(n8137), .A2(n8136), .ZN(n10183) );
  NAND2_X1 U5445 ( .A1(n4667), .A2(n4665), .ZN(n6840) );
  OAI21_X1 U5446 ( .B1(n6838), .B2(n8342), .A(n6839), .ZN(n4667) );
  NAND2_X1 U5447 ( .A1(n4666), .A2(n6988), .ZN(n4665) );
  INV_X1 U5448 ( .A(n6839), .ZN(n4666) );
  OR2_X1 U5449 ( .A1(n6573), .A2(n6679), .ZN(n4417) );
  MUX2_X1 U5450 ( .A(n6881), .B(n6880), .S(n6980), .Z(n6882) );
  INV_X1 U5451 ( .A(n6999), .ZN(n4663) );
  NOR2_X1 U5452 ( .A1(n4661), .A2(n4660), .ZN(n4659) );
  INV_X1 U5453 ( .A(n6902), .ZN(n4660) );
  AND2_X1 U5454 ( .A1(n8906), .A2(n4662), .ZN(n4661) );
  INV_X1 U5455 ( .A(n4636), .ZN(n4635) );
  OAI21_X1 U5456 ( .B1(n6921), .B2(n4296), .A(n6928), .ZN(n4636) );
  AOI21_X1 U5457 ( .B1(n6947), .B2(n6948), .A(n4528), .ZN(n4527) );
  NOR2_X1 U5458 ( .A1(n6948), .A2(n6980), .ZN(n4528) );
  NAND2_X1 U5459 ( .A1(n6946), .A2(n6292), .ZN(n4529) );
  OAI21_X1 U5460 ( .B1(n8766), .B2(n6945), .A(n6944), .ZN(n6946) );
  OR2_X1 U5461 ( .A1(n6941), .A2(n6980), .ZN(n6945) );
  NOR2_X1 U5462 ( .A1(n4601), .A2(n8794), .ZN(n4651) );
  NOR2_X1 U5463 ( .A1(n6954), .A2(n6955), .ZN(n4649) );
  NAND2_X1 U5464 ( .A1(n7020), .A2(n6957), .ZN(n6960) );
  NOR2_X1 U5465 ( .A1(n8054), .A2(n4397), .ZN(n7008) );
  NOR2_X1 U5466 ( .A1(n4680), .A2(n6003), .ZN(n4678) );
  INV_X1 U5467 ( .A(n6254), .ZN(n4680) );
  INV_X1 U5468 ( .A(n6255), .ZN(n4682) );
  AND2_X1 U5469 ( .A1(n6186), .A2(n6995), .ZN(n4603) );
  INV_X1 U5470 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5719) );
  INV_X1 U5471 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5721) );
  NOR2_X2 U5472 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5723) );
  NOR2_X1 U5473 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5692) );
  AND2_X1 U5474 ( .A1(n7184), .A2(n4788), .ZN(n4787) );
  NAND2_X1 U5475 ( .A1(n6673), .A2(n4412), .ZN(n4411) );
  NOR2_X1 U5476 ( .A1(n6732), .A2(n6543), .ZN(n6740) );
  AND2_X1 U5477 ( .A1(n6635), .A2(n9672), .ZN(n6733) );
  INV_X1 U5478 ( .A(n6569), .ZN(n4955) );
  AOI21_X1 U5479 ( .B1(n4481), .B2(n4478), .A(n4476), .ZN(n4475) );
  INV_X1 U5480 ( .A(n5465), .ZN(n4476) );
  INV_X1 U5481 ( .A(n4478), .ZN(n4477) );
  NAND2_X1 U5482 ( .A1(n5469), .A2(n5468), .ZN(n5483) );
  INV_X1 U5483 ( .A(n5420), .ZN(n5426) );
  INV_X1 U5484 ( .A(n4499), .ZN(n4495) );
  NOR2_X1 U5485 ( .A1(n5360), .A2(n4879), .ZN(n4878) );
  INV_X1 U5486 ( .A(n5339), .ZN(n4879) );
  INV_X1 U5487 ( .A(SI_17_), .ZN(n5342) );
  AND2_X1 U5488 ( .A1(n4338), .A2(n5304), .ZN(n4501) );
  AND2_X1 U5489 ( .A1(n4866), .A2(n5232), .ZN(n4483) );
  AND2_X1 U5490 ( .A1(n6463), .A2(n8527), .ZN(n6465) );
  INV_X1 U5491 ( .A(n6963), .ZN(n4492) );
  NAND2_X1 U5492 ( .A1(n8616), .A2(n4334), .ZN(n5764) );
  NOR2_X1 U5493 ( .A1(n4738), .A2(n7510), .ZN(n4734) );
  AOI21_X1 U5494 ( .B1(n7963), .B2(n7962), .A(n4428), .ZN(n5826) );
  NOR2_X1 U5495 ( .A1(n7961), .A2(n8973), .ZN(n4428) );
  NAND2_X1 U5496 ( .A1(n8687), .A2(n4752), .ZN(n5798) );
  NAND2_X1 U5497 ( .A1(n4631), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4752) );
  NOR2_X1 U5498 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n4532) );
  AND2_X1 U5499 ( .A1(n8883), .A2(n4690), .ZN(n4689) );
  AND2_X1 U5500 ( .A1(n6003), .A2(n6862), .ZN(n4911) );
  INV_X1 U5501 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5979) );
  INV_X1 U5502 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U5503 ( .A1(n5926), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4654) );
  NAND2_X1 U5504 ( .A1(n6958), .A2(n8605), .ZN(n7020) );
  NAND2_X1 U5505 ( .A1(n6196), .A2(n6952), .ZN(n4895) );
  OR2_X1 U5506 ( .A1(n8989), .A2(n8584), .ZN(n6948) );
  NAND2_X1 U5507 ( .A1(n6287), .A2(n6288), .ZN(n4720) );
  INV_X1 U5508 ( .A(n8821), .ZN(n6280) );
  OAI21_X1 U5509 ( .B1(n4297), .B2(n4613), .A(n6835), .ZN(n4612) );
  INV_X1 U5510 ( .A(n8844), .ZN(n8846) );
  CLKBUF_X1 U5511 ( .A(n7974), .Z(n7975) );
  NOR2_X1 U5512 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4676) );
  INV_X1 U5513 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5739) );
  NOR2_X1 U5514 ( .A1(n5777), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U5515 ( .A1(n5769), .A2(n5718), .ZN(n5773) );
  AND2_X1 U5516 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5104) );
  NOR2_X1 U5517 ( .A1(n7149), .A2(n4821), .ZN(n4820) );
  INV_X1 U5518 ( .A(n8325), .ZN(n4821) );
  NOR2_X1 U5519 ( .A1(n5367), .A2(n5366), .ZN(n4448) );
  AND2_X1 U5520 ( .A1(n7224), .A2(n7223), .ZN(n9152) );
  NOR2_X1 U5521 ( .A1(n5291), .A2(n9105), .ZN(n4447) );
  OR2_X1 U5522 ( .A1(n5065), .A2(n10001), .ZN(n5005) );
  OR2_X1 U5523 ( .A1(n6534), .A2(n5001), .ZN(n5004) );
  INV_X1 U5524 ( .A(n9550), .ZN(n4574) );
  INV_X1 U5525 ( .A(n9547), .ZN(n4571) );
  NAND2_X1 U5526 ( .A1(n4776), .A2(n9602), .ZN(n4775) );
  NOR2_X1 U5527 ( .A1(n8419), .A2(n6668), .ZN(n4776) );
  AND2_X1 U5528 ( .A1(n5670), .A2(n4960), .ZN(n4959) );
  NAND2_X1 U5529 ( .A1(n6784), .A2(n4961), .ZN(n4960) );
  NOR2_X1 U5530 ( .A1(n9843), .A2(n9847), .ZN(n4766) );
  NAND2_X1 U5531 ( .A1(n4766), .A2(n9933), .ZN(n4765) );
  NAND2_X1 U5532 ( .A1(n4448), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5400) );
  NOR2_X1 U5533 ( .A1(n9787), .A2(n9861), .ZN(n9741) );
  NOR3_X1 U5534 ( .A1(n8066), .A2(n4768), .A3(n9967), .ZN(n8365) );
  NAND2_X1 U5535 ( .A1(n4769), .A2(n9287), .ZN(n4768) );
  INV_X1 U5536 ( .A(n4770), .ZN(n4769) );
  NAND2_X1 U5537 ( .A1(n9204), .A2(n4771), .ZN(n4770) );
  AND2_X1 U5538 ( .A1(n8235), .A2(n10057), .ZN(n4772) );
  OR2_X1 U5539 ( .A1(n5578), .A2(n7333), .ZN(n5020) );
  AOI21_X1 U5540 ( .B1(n4959), .B2(n5537), .A(n4443), .ZN(n4957) );
  INV_X1 U5541 ( .A(n9642), .ZN(n4548) );
  NOR2_X1 U5542 ( .A1(n9727), .A2(n9847), .ZN(n9709) );
  AOI21_X1 U5543 ( .B1(n4464), .B2(n4467), .A(n4462), .ZN(n4461) );
  INV_X1 U5544 ( .A(n5538), .ZN(n4462) );
  INV_X1 U5545 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5546 ( .A1(n5617), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5625) );
  INV_X1 U5547 ( .A(SI_20_), .ZN(n5422) );
  NOR2_X1 U5548 ( .A1(n4877), .A2(n4500), .ZN(n4499) );
  INV_X1 U5549 ( .A(n4501), .ZN(n4500) );
  INV_X1 U5550 ( .A(n4878), .ZN(n4877) );
  NOR2_X1 U5551 ( .A1(n5340), .A2(n4882), .ZN(n4881) );
  INV_X1 U5552 ( .A(n5325), .ZN(n4882) );
  NOR2_X1 U5553 ( .A1(n5270), .A2(n4862), .ZN(n4861) );
  INV_X1 U5554 ( .A(n5249), .ZN(n4862) );
  INV_X1 U5555 ( .A(n4859), .ZN(n4858) );
  OAI21_X1 U5556 ( .B1(n5270), .B2(n4860), .A(n5269), .ZN(n4859) );
  NAND2_X1 U5557 ( .A1(n5250), .A2(n5249), .ZN(n4860) );
  INV_X1 U5558 ( .A(n5209), .ZN(n4864) );
  NAND2_X1 U5559 ( .A1(n5174), .A2(n4866), .ZN(n4489) );
  INV_X1 U5560 ( .A(n5173), .ZN(n4870) );
  AOI21_X1 U5561 ( .B1(n5162), .B2(n4851), .A(n4350), .ZN(n4850) );
  INV_X1 U5562 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5007) );
  NOR2_X1 U5563 ( .A1(n8463), .A2(n4525), .ZN(n4524) );
  INV_X1 U5564 ( .A(n6446), .ZN(n4525) );
  AOI21_X1 U5565 ( .B1(n6385), .B2(n8212), .A(n6384), .ZN(n4526) );
  AND2_X1 U5566 ( .A1(n6417), .A2(n4513), .ZN(n4512) );
  AND2_X1 U5567 ( .A1(n8554), .A2(n6416), .ZN(n6417) );
  NAND2_X1 U5568 ( .A1(n4978), .A2(n4516), .ZN(n4513) );
  INV_X1 U5569 ( .A(n4978), .ZN(n4514) );
  NAND2_X1 U5570 ( .A1(n8465), .A2(n4934), .ZN(n8533) );
  AND2_X1 U5571 ( .A1(n4932), .A2(n8492), .ZN(n4931) );
  OR2_X1 U5572 ( .A1(n4934), .A2(n4933), .ZN(n4932) );
  NAND2_X1 U5573 ( .A1(n4919), .A2(n6442), .ZN(n8572) );
  INV_X1 U5574 ( .A(n8516), .ZN(n4919) );
  NAND2_X1 U5575 ( .A1(n4926), .A2(n4924), .ZN(n4923) );
  INV_X1 U5576 ( .A(n4928), .ZN(n4924) );
  INV_X1 U5577 ( .A(n4926), .ZN(n4925) );
  AND2_X1 U5578 ( .A1(n6499), .A2(n6498), .ZN(n7431) );
  INV_X1 U5579 ( .A(n7025), .ZN(n7026) );
  AND2_X1 U5580 ( .A1(n6973), .A2(n6972), .ZN(n8603) );
  OAI21_X1 U5581 ( .B1(n7492), .B2(n5806), .A(n4618), .ZN(n7485) );
  NAND2_X1 U5582 ( .A1(n7492), .A2(n5806), .ZN(n4618) );
  NAND2_X1 U5583 ( .A1(n7484), .A2(n7485), .ZN(n7483) );
  NAND2_X1 U5584 ( .A1(n8617), .A2(n8618), .ZN(n8616) );
  NAND2_X1 U5585 ( .A1(n8621), .A2(n8622), .ZN(n8620) );
  NAND2_X1 U5586 ( .A1(n5862), .A2(n7674), .ZN(n7696) );
  NAND2_X1 U5587 ( .A1(n7699), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4748) );
  NAND2_X1 U5588 ( .A1(n5776), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5589 ( .A1(n4355), .A2(n6035), .ZN(n4745) );
  NAND2_X1 U5590 ( .A1(n5870), .A2(n7770), .ZN(n7907) );
  XNOR2_X1 U5591 ( .A(n5825), .B(n6048), .ZN(n7903) );
  OAI22_X1 U5592 ( .A1(n7903), .A2(n8088), .B1(n6048), .B2(n5825), .ZN(n7963)
         );
  XNOR2_X1 U5593 ( .A(n5826), .B(n7543), .ZN(n8636) );
  NAND2_X1 U5594 ( .A1(n5879), .A2(n8637), .ZN(n8659) );
  OAI22_X1 U5595 ( .A1(n8636), .A2(n8966), .B1(n7543), .B2(n5826), .ZN(n8655)
         );
  NAND2_X1 U5596 ( .A1(n8669), .A2(n5797), .ZN(n8689) );
  NAND2_X1 U5597 ( .A1(n8689), .A2(n8688), .ZN(n8687) );
  NAND2_X1 U5598 ( .A1(n5887), .A2(n8671), .ZN(n8693) );
  XNOR2_X1 U5599 ( .A(n5798), .B(n4629), .ZN(n8709) );
  XNOR2_X1 U5600 ( .A(n5830), .B(n4629), .ZN(n8717) );
  NAND2_X1 U5601 ( .A1(n4631), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4630) );
  INV_X1 U5602 ( .A(n6230), .ZN(n8380) );
  NAND2_X1 U5603 ( .A1(n6208), .A2(n10199), .ZN(n6220) );
  NAND2_X1 U5604 ( .A1(n6178), .A2(n4530), .ZN(n6209) );
  AND2_X1 U5605 ( .A1(n4532), .A2(n4531), .ZN(n4530) );
  INV_X1 U5606 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4531) );
  NAND2_X1 U5607 ( .A1(n6178), .A2(n6177), .ZN(n6189) );
  OR2_X1 U5608 ( .A1(n6166), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U5609 ( .A1(n6149), .A2(n6148), .ZN(n6166) );
  INV_X1 U5610 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6148) );
  INV_X1 U5611 ( .A(n6150), .ZN(n6149) );
  AND2_X1 U5612 ( .A1(n4306), .A2(n4539), .ZN(n4538) );
  INV_X1 U5613 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4539) );
  NAND2_X1 U5614 ( .A1(n6112), .A2(n6111), .ZN(n6120) );
  INV_X1 U5615 ( .A(n4689), .ZN(n4688) );
  INV_X1 U5616 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4535) );
  OR2_X1 U5617 ( .A1(n6104), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U5618 ( .A1(n6072), .A2(n4536), .ZN(n6094) );
  NAND2_X1 U5619 ( .A1(n6072), .A2(n6071), .ZN(n6083) );
  AOI21_X1 U5620 ( .B1(n4354), .B2(n4693), .A(n4302), .ZN(n4691) );
  NAND2_X1 U5621 ( .A1(n6061), .A2(n6060), .ZN(n6073) );
  INV_X1 U5622 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6060) );
  INV_X1 U5623 ( .A(n6062), .ZN(n6061) );
  OR2_X1 U5624 ( .A1(n6051), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6062) );
  OR2_X1 U5625 ( .A1(n8976), .A2(n8055), .ZN(n8050) );
  NAND2_X1 U5626 ( .A1(n6027), .A2(n10300), .ZN(n6028) );
  INV_X1 U5627 ( .A(n6039), .ZN(n6027) );
  OR2_X1 U5628 ( .A1(n6028), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6051) );
  INV_X1 U5629 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U5630 ( .A1(n6007), .A2(n6006), .ZN(n6019) );
  INV_X1 U5631 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6006) );
  INV_X1 U5632 ( .A(n6017), .ZN(n6007) );
  NAND4_X1 U5633 ( .A1(n5968), .A2(n5969), .A3(n5979), .A4(n4541), .ZN(n6017)
         );
  INV_X1 U5634 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n4541) );
  NAND2_X1 U5635 ( .A1(n5969), .A2(n5968), .ZN(n5980) );
  AND2_X1 U5636 ( .A1(n8212), .A2(n7028), .ZN(n6354) );
  OR2_X1 U5637 ( .A1(n6966), .A2(n7644), .ZN(n5963) );
  NAND2_X1 U5638 ( .A1(n6244), .A2(n7734), .ZN(n4672) );
  NAND2_X1 U5639 ( .A1(n4673), .A2(n7530), .ZN(n7734) );
  NAND2_X1 U5640 ( .A1(n7735), .A2(n5945), .ZN(n7732) );
  NAND2_X1 U5641 ( .A1(n6987), .A2(n7020), .ZN(n7016) );
  AND2_X1 U5642 ( .A1(n6353), .A2(n6491), .ZN(n7306) );
  NAND2_X1 U5643 ( .A1(n6964), .A2(n6963), .ZN(n4493) );
  AND2_X1 U5644 ( .A1(n6996), .A2(n6995), .ZN(n8795) );
  NAND2_X1 U5645 ( .A1(n4899), .A2(n4897), .ZN(n8809) );
  INV_X1 U5646 ( .A(n4898), .ZN(n4897) );
  OAI21_X1 U5647 ( .B1(n4901), .B2(n6929), .A(n6928), .ZN(n4898) );
  AND2_X1 U5648 ( .A1(n6901), .A2(n6900), .ZN(n8906) );
  AOI21_X1 U5649 ( .B1(n4889), .B2(n4891), .A(n4345), .ZN(n4888) );
  AND2_X1 U5650 ( .A1(n8059), .A2(n6321), .ZN(n10146) );
  INV_X1 U5651 ( .A(n10135), .ZN(n10151) );
  AND2_X1 U5652 ( .A1(n6343), .A2(n6342), .ZN(n6489) );
  NOR2_X1 U5653 ( .A1(n6497), .A2(n6495), .ZN(n6485) );
  NAND2_X1 U5654 ( .A1(n6341), .A2(n8342), .ZN(n10135) );
  NAND2_X1 U5655 ( .A1(n5712), .A2(n4980), .ZN(n5732) );
  NAND2_X1 U5656 ( .A1(n5714), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U5657 ( .A1(n5703), .A2(n5710), .ZN(n5704) );
  NAND2_X1 U5658 ( .A1(n5714), .A2(n5717), .ZN(n6500) );
  NAND2_X1 U5659 ( .A1(n5712), .A2(n5701), .ZN(n5715) );
  NAND2_X1 U5660 ( .A1(n5725), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  NOR2_X1 U5661 ( .A1(n5724), .A2(n4520), .ZN(n4519) );
  NAND2_X1 U5662 ( .A1(n4522), .A2(n4521), .ZN(n4520) );
  INV_X1 U5663 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5801) );
  INV_X1 U5664 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5789) );
  OR2_X1 U5665 ( .A1(n5787), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5741) );
  AND2_X1 U5666 ( .A1(n5781), .A2(n5739), .ZN(n5784) );
  NAND2_X1 U5667 ( .A1(n4815), .A2(n4817), .ZN(n9126) );
  INV_X1 U5668 ( .A(n4818), .ZN(n4817) );
  NAND2_X1 U5669 ( .A1(n8328), .A2(n4820), .ZN(n4815) );
  AND2_X1 U5670 ( .A1(n9185), .A2(n7230), .ZN(n7231) );
  INV_X1 U5671 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10221) );
  INV_X1 U5672 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U5673 ( .A1(n7917), .A2(n7109), .ZN(n4797) );
  OR2_X1 U5674 ( .A1(n5331), .A2(n9222), .ZN(n5353) );
  NAND2_X1 U5675 ( .A1(n9236), .A2(n9237), .ZN(n9235) );
  OR2_X1 U5676 ( .A1(n8328), .A2(n8324), .ZN(n4816) );
  NAND2_X1 U5677 ( .A1(n7393), .A2(n5397), .ZN(n5200) );
  INV_X1 U5678 ( .A(n4446), .ZN(n5438) );
  INV_X1 U5679 ( .A(n9322), .ZN(n9337) );
  NAND2_X1 U5680 ( .A1(n5351), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5367) );
  INV_X1 U5681 ( .A(n5353), .ZN(n5351) );
  INV_X1 U5682 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5366) );
  INV_X1 U5683 ( .A(n4448), .ZN(n5389) );
  AND2_X1 U5684 ( .A1(n7443), .A2(n9386), .ZN(n9322) );
  AOI21_X1 U5685 ( .B1(n4791), .B2(n4793), .A(n4344), .ZN(n4790) );
  INV_X1 U5686 ( .A(n4447), .ZN(n5314) );
  NAND2_X1 U5687 ( .A1(n4447), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5331) );
  AND3_X1 U5688 ( .A1(n6791), .A2(n6688), .A3(n4983), .ZN(n6815) );
  AND2_X1 U5689 ( .A1(n6687), .A2(n6686), .ZN(n6827) );
  OR2_X1 U5690 ( .A1(n9574), .A2(n4291), .ZN(n5554) );
  AND2_X1 U5691 ( .A1(n5480), .A2(n5479), .ZN(n9119) );
  AND4_X1 U5692 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8287)
         );
  AND4_X1 U5693 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n8304)
         );
  AND4_X1 U5694 ( .A1(n5246), .A2(n5245), .A3(n5244), .A4(n5243), .ZN(n8288)
         );
  AND4_X1 U5695 ( .A1(n5227), .A2(n5226), .A3(n5225), .A4(n5224), .ZN(n7153)
         );
  AND4_X1 U5696 ( .A1(n5207), .A2(n5206), .A3(n5205), .A4(n5204), .ZN(n7143)
         );
  NAND4_X1 U5697 ( .A1(n5025), .A2(n5024), .A3(n5023), .A4(n5022), .ZN(n5642)
         );
  OR2_X1 U5698 ( .A1(n6534), .A2(n8171), .ZN(n5024) );
  OR2_X1 U5699 ( .A1(n4290), .A2(n9393), .ZN(n5023) );
  OR2_X1 U5700 ( .A1(n5213), .A2(n5212), .ZN(n5216) );
  NAND2_X1 U5701 ( .A1(n9498), .A2(n4339), .ZN(n7599) );
  INV_X1 U5702 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7602) );
  OR2_X1 U5703 ( .A1(n7590), .A2(n7591), .ZN(n4583) );
  NOR2_X1 U5704 ( .A1(n9524), .A2(n4581), .ZN(n10009) );
  AND2_X1 U5705 ( .A1(n9525), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4581) );
  AND2_X1 U5706 ( .A1(n4585), .A2(n4584), .ZN(n9533) );
  NAND2_X1 U5707 ( .A1(n6747), .A2(n6742), .ZN(n6665) );
  NOR2_X1 U5708 ( .A1(n9727), .A2(n4764), .ZN(n9678) );
  INV_X1 U5709 ( .A(n4766), .ZN(n4764) );
  CLKBUF_X1 U5710 ( .A(n9741), .Z(n9767) );
  NAND2_X1 U5711 ( .A1(n8365), .A2(n5684), .ZN(n9787) );
  INV_X1 U5712 ( .A(n9870), .ZN(n5684) );
  NAND2_X1 U5713 ( .A1(n9775), .A2(n9776), .ZN(n9774) );
  INV_X1 U5714 ( .A(n8365), .ZN(n9785) );
  INV_X1 U5715 ( .A(n8310), .ZN(n5654) );
  NOR2_X1 U5716 ( .A1(n8066), .A2(n9885), .ZN(n8291) );
  INV_X1 U5717 ( .A(n5649), .ZN(n8005) );
  NAND2_X1 U5718 ( .A1(n8239), .A2(n8241), .ZN(n8255) );
  INV_X1 U5719 ( .A(n8235), .ZN(n8219) );
  NAND2_X1 U5720 ( .A1(n7939), .A2(n4772), .ZN(n8248) );
  CLKBUF_X1 U5721 ( .A(n7886), .Z(n8157) );
  NAND2_X1 U5722 ( .A1(n7939), .A2(n10057), .ZN(n7938) );
  AND2_X2 U5723 ( .A1(n6699), .A2(n6697), .ZN(n7840) );
  NAND2_X1 U5724 ( .A1(n5639), .A2(n9802), .ZN(n8264) );
  AND2_X1 U5725 ( .A1(n9797), .A2(n7282), .ZN(n7332) );
  INV_X1 U5726 ( .A(n5685), .ZN(n6380) );
  NAND2_X1 U5727 ( .A1(n5512), .A2(n5511), .ZN(n9814) );
  NAND2_X1 U5728 ( .A1(n4946), .A2(n5665), .ZN(n9609) );
  AND2_X1 U5729 ( .A1(n4950), .A2(n6617), .ZN(n9737) );
  NAND2_X1 U5730 ( .A1(n5275), .A2(n5274), .ZN(n9880) );
  AND2_X1 U5731 ( .A1(n8159), .A2(n4847), .ZN(n4844) );
  NAND2_X1 U5732 ( .A1(n8000), .A2(n8001), .ZN(n8003) );
  AND2_X1 U5733 ( .A1(n7279), .A2(n7284), .ZN(n5920) );
  INV_X1 U5734 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4997) );
  INV_X1 U5735 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4962) );
  OAI21_X1 U5736 ( .B1(n5507), .B2(n4467), .A(n4464), .ZN(n5539) );
  XNOR2_X1 U5737 ( .A(n5603), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5621) );
  OR2_X1 U5738 ( .A1(n7442), .A2(P1_U3086), .ZN(n7444) );
  NAND2_X1 U5739 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  XNOR2_X1 U5740 ( .A(n5395), .B(n5394), .ZN(n8018) );
  AND2_X1 U5741 ( .A1(n5272), .A2(n5256), .ZN(n7592) );
  OAI21_X1 U5742 ( .B1(n5251), .B2(n5250), .A(n5249), .ZN(n5271) );
  XNOR2_X1 U5743 ( .A(n5171), .B(n5169), .ZN(n7373) );
  NAND3_X1 U5744 ( .A1(n7366), .A2(n7361), .A3(n7365), .ZN(n6492) );
  NAND2_X1 U5745 ( .A1(n7746), .A2(n6409), .ZN(n7871) );
  NAND2_X1 U5746 ( .A1(n8574), .A2(n4524), .ZN(n8465) );
  NAND2_X1 U5747 ( .A1(n8574), .A2(n6446), .ZN(n8464) );
  NAND2_X1 U5748 ( .A1(n6219), .A2(n6218), .ZN(n8480) );
  AND2_X1 U5749 ( .A1(n7869), .A2(n6412), .ZN(n8106) );
  INV_X1 U5750 ( .A(n7450), .ZN(n6391) );
  NAND2_X1 U5751 ( .A1(n8533), .A2(n6453), .ZN(n8493) );
  NAND2_X1 U5752 ( .A1(n8542), .A2(n4928), .ZN(n4922) );
  INV_X1 U5753 ( .A(n4936), .ZN(n4935) );
  OAI21_X1 U5754 ( .B1(n4938), .B2(n4937), .A(n8507), .ZN(n4936) );
  INV_X1 U5755 ( .A(n6438), .ZN(n4937) );
  NAND2_X1 U5756 ( .A1(n8592), .A2(n6438), .ZN(n8508) );
  NAND2_X1 U5757 ( .A1(n7650), .A2(n7719), .ZN(n4913) );
  INV_X1 U5758 ( .A(n8528), .ZN(n4504) );
  NAND2_X1 U5759 ( .A1(n4507), .A2(n4506), .ZN(n4505) );
  OR2_X1 U5760 ( .A1(n8528), .A2(n4509), .ZN(n4506) );
  NAND2_X1 U5761 ( .A1(n8528), .A2(n4343), .ZN(n4507) );
  NAND2_X1 U5762 ( .A1(n8528), .A2(n4510), .ZN(n4508) );
  AND4_X1 U5763 ( .A1(n6013), .A2(n6012), .A3(n6011), .A4(n6010), .ZN(n8033)
         );
  INV_X1 U5764 ( .A(n8597), .ZN(n8580) );
  NAND2_X1 U5765 ( .A1(n4915), .A2(n6406), .ZN(n4914) );
  NAND2_X1 U5766 ( .A1(n7650), .A2(n4329), .ZN(n4502) );
  INV_X1 U5767 ( .A(n7720), .ZN(n4915) );
  INV_X1 U5768 ( .A(n8606), .ZN(n8897) );
  NAND2_X1 U5769 ( .A1(n8437), .A2(n4938), .ZN(n8592) );
  AND2_X1 U5770 ( .A1(n8437), .A2(n6435), .ZN(n8594) );
  NAND2_X1 U5771 ( .A1(n7431), .A2(n8345), .ZN(n8599) );
  INV_X1 U5772 ( .A(n8584), .ZN(n8768) );
  NAND2_X1 U5773 ( .A1(n6195), .A2(n6194), .ZN(n8767) );
  NAND2_X1 U5774 ( .A1(n6126), .A2(n6125), .ZN(n8871) );
  NOR2_X1 U5775 ( .A1(n5949), .A2(n5948), .ZN(n5952) );
  INV_X1 U5776 ( .A(n7612), .ZN(n4622) );
  NAND2_X1 U5777 ( .A1(n5817), .A2(n4621), .ZN(n7611) );
  NAND2_X1 U5778 ( .A1(n7498), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4621) );
  XNOR2_X1 U5779 ( .A(n5819), .B(n6014), .ZN(n7509) );
  NAND2_X1 U5780 ( .A1(n7685), .A2(n7686), .ZN(n7684) );
  XNOR2_X1 U5781 ( .A(n5776), .B(n6035), .ZN(n7692) );
  NAND2_X1 U5782 ( .A1(n5824), .A2(n4625), .ZN(n7779) );
  NAND2_X1 U5783 ( .A1(n7691), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4625) );
  INV_X1 U5784 ( .A(n4747), .ZN(n7767) );
  AND2_X1 U5785 ( .A1(n5783), .A2(n7910), .ZN(n4405) );
  NAND2_X1 U5786 ( .A1(n8682), .A2(n5829), .ZN(n8705) );
  NOR2_X1 U5787 ( .A1(n8744), .A2(n8865), .ZN(n4432) );
  OAI21_X1 U5788 ( .B1(n5910), .B2(n8694), .A(n5909), .ZN(n5911) );
  NOR2_X1 U5789 ( .A1(n8744), .A2(n8945), .ZN(n4406) );
  NAND2_X1 U5790 ( .A1(n4965), .A2(n6320), .ZN(n8379) );
  OR2_X1 U5791 ( .A1(n7312), .A2(n8917), .ZN(n7316) );
  NAND2_X1 U5792 ( .A1(n4909), .A2(n6905), .ZN(n8879) );
  NAND2_X1 U5793 ( .A1(n6110), .A2(n6109), .ZN(n8948) );
  OAI21_X1 U5794 ( .B1(n8053), .B2(n4695), .A(n4693), .ZN(n8192) );
  NAND2_X1 U5795 ( .A1(n4912), .A2(n6862), .ZN(n7784) );
  NAND2_X1 U5796 ( .A1(n4683), .A2(n6255), .ZN(n7785) );
  NAND2_X1 U5797 ( .A1(n7795), .A2(n6254), .ZN(n4683) );
  NAND2_X1 U5798 ( .A1(n6002), .A2(n6001), .ZN(n7790) );
  NAND2_X1 U5799 ( .A1(n10097), .A2(n6859), .ZN(n7793) );
  OR2_X1 U5800 ( .A1(n10135), .A2(n6354), .ZN(n8778) );
  OR2_X1 U5801 ( .A1(n6478), .A2(n6495), .ZN(n8874) );
  OR2_X1 U5802 ( .A1(n7313), .A2(n8778), .ZN(n8901) );
  INV_X1 U5803 ( .A(n8917), .ZN(n10104) );
  NOR2_X1 U5804 ( .A1(n10166), .A2(n8921), .ZN(n4724) );
  INV_X1 U5805 ( .A(n4493), .ZN(n8983) );
  AOI21_X1 U5806 ( .B1(n8424), .B2(n5988), .A(n6977), .ZN(n8986) );
  INV_X1 U5807 ( .A(n8480), .ZN(n7053) );
  NAND2_X1 U5808 ( .A1(n4727), .A2(n4726), .ZN(n4725) );
  NAND2_X1 U5809 ( .A1(n4886), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5810 ( .A1(n8776), .A2(n10093), .ZN(n4726) );
  NAND2_X1 U5811 ( .A1(n6198), .A2(n6197), .ZN(n8995) );
  NAND2_X1 U5812 ( .A1(n4894), .A2(n6952), .ZN(n8764) );
  OR2_X1 U5813 ( .A1(n8782), .A2(n6196), .ZN(n4894) );
  NAND2_X1 U5814 ( .A1(n6188), .A2(n6187), .ZN(n9001) );
  NAND2_X1 U5815 ( .A1(n6176), .A2(n6175), .ZN(n9007) );
  NAND2_X1 U5816 ( .A1(n6285), .A2(n6284), .ZN(n8801) );
  NAND2_X1 U5817 ( .A1(n6165), .A2(n6164), .ZN(n9019) );
  NAND2_X1 U5818 ( .A1(n4698), .A2(n4702), .ZN(n8810) );
  OR2_X1 U5819 ( .A1(n8861), .A2(n4705), .ZN(n4698) );
  NAND2_X1 U5820 ( .A1(n6145), .A2(n5988), .ZN(n6147) );
  NAND2_X1 U5821 ( .A1(n4707), .A2(n4709), .ZN(n8822) );
  NAND2_X1 U5822 ( .A1(n4900), .A2(n6924), .ZN(n8820) );
  OR2_X1 U5823 ( .A1(n8832), .A2(n4904), .ZN(n4900) );
  NAND2_X1 U5824 ( .A1(n8950), .A2(n7011), .ZN(n8843) );
  NAND2_X1 U5825 ( .A1(n6119), .A2(n6118), .ZN(n9041) );
  NAND2_X1 U5826 ( .A1(n6103), .A2(n6102), .ZN(n9048) );
  NAND2_X1 U5827 ( .A1(n4907), .A2(n6903), .ZN(n8882) );
  INV_X1 U5828 ( .A(n8590), .ZN(n9056) );
  NAND2_X1 U5829 ( .A1(n6082), .A2(n6081), .ZN(n9059) );
  NAND2_X1 U5830 ( .A1(n8191), .A2(n6068), .ZN(n8320) );
  OR2_X1 U5831 ( .A1(n10154), .A2(n10146), .ZN(n9074) );
  OAI21_X1 U5832 ( .B1(n8053), .B2(n4310), .A(n6264), .ZN(n8077) );
  NAND2_X1 U5833 ( .A1(n6026), .A2(n6025), .ZN(n8460) );
  INV_X2 U5834 ( .A(n10154), .ZN(n10152) );
  NAND2_X1 U5835 ( .A1(n4669), .A2(n5712), .ZN(n9080) );
  AND2_X1 U5836 ( .A1(n4910), .A2(n4670), .ZN(n4669) );
  AND2_X1 U5837 ( .A1(n5730), .A2(n5924), .ZN(n4670) );
  INV_X1 U5838 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9095) );
  INV_X1 U5839 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9098) );
  XNOR2_X1 U5840 ( .A(n5702), .B(n5708), .ZN(n6323) );
  NAND2_X1 U5841 ( .A1(n5704), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5702) );
  INV_X1 U5842 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8375) );
  NAND2_X1 U5843 ( .A1(n5705), .A2(n5704), .ZN(n6322) );
  OR2_X1 U5844 ( .A1(n5703), .A2(n5710), .ZN(n5705) );
  INV_X1 U5845 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8344) );
  INV_X1 U5846 ( .A(n7036), .ZN(n8342) );
  INV_X1 U5847 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10233) );
  INV_X1 U5848 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8210) );
  INV_X1 U5849 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10259) );
  INV_X1 U5850 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7946) );
  INV_X1 U5851 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10253) );
  INV_X1 U5852 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7745) );
  INV_X1 U5853 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7426) );
  INV_X1 U5854 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7419) );
  INV_X1 U5855 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10261) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10289) );
  INV_X1 U5857 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7380) );
  INV_X1 U5858 ( .A(n5987), .ZN(n7503) );
  NAND2_X1 U5859 ( .A1(n5761), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U5860 ( .A1(n7442), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7710) );
  INV_X1 U5861 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8329) );
  AND2_X1 U5862 ( .A1(n7274), .A2(n9302), .ZN(n4782) );
  INV_X1 U5863 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9105) );
  AND2_X1 U5864 ( .A1(n4803), .A2(n4802), .ZN(n9113) );
  NAND2_X1 U5865 ( .A1(n9235), .A2(n7253), .ZN(n9205) );
  NAND2_X1 U5866 ( .A1(n5490), .A2(n5489), .ZN(n9211) );
  NAND2_X1 U5867 ( .A1(n4393), .A2(n7221), .ZN(n4392) );
  NAND2_X1 U5868 ( .A1(n9214), .A2(n9151), .ZN(n4393) );
  NAND2_X1 U5869 ( .A1(n9136), .A2(n7105), .ZN(n7917) );
  XNOR2_X1 U5870 ( .A(n7239), .B(n7238), .ZN(n9289) );
  OR2_X1 U5871 ( .A1(n8328), .A2(n4813), .ZN(n4807) );
  NAND2_X1 U5872 ( .A1(n4799), .A2(n4300), .ZN(n4795) );
  OR2_X1 U5873 ( .A1(n7298), .A2(n7297), .ZN(n9326) );
  INV_X1 U5874 ( .A(n9331), .ZN(n9343) );
  OR2_X1 U5875 ( .A1(n7298), .A2(n7281), .ZN(n9345) );
  INV_X1 U5876 ( .A(n7272), .ZN(n9350) );
  INV_X1 U5877 ( .A(n9292), .ZN(n9354) );
  OR2_X1 U5878 ( .A1(n9663), .A2(n4290), .ZN(n5444) );
  INV_X1 U5879 ( .A(n7134), .ZN(n9369) );
  OR2_X1 U5880 ( .A1(n5583), .A2(n5064), .ZN(n5069) );
  MUX2_X1 U5881 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5021), .S(n9396), .Z(n9399)
         );
  NAND2_X1 U5882 ( .A1(n9414), .A2(n9415), .ZN(n9413) );
  NAND2_X1 U5883 ( .A1(n9400), .A2(n7547), .ZN(n9414) );
  NOR2_X1 U5884 ( .A1(n4593), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U5885 ( .A1(n9413), .A2(n7548), .ZN(n9424) );
  NAND2_X1 U5886 ( .A1(n9438), .A2(n9439), .ZN(n9437) );
  NAND2_X1 U5887 ( .A1(n9450), .A2(n4332), .ZN(n9464) );
  NAND2_X1 U5888 ( .A1(n9464), .A2(n9465), .ZN(n9463) );
  NOR2_X1 U5889 ( .A1(n7550), .A2(n7551), .ZN(n7588) );
  AOI21_X1 U5890 ( .B1(n9893), .B2(n7594), .A(n7593), .ZN(n9487) );
  NAND2_X1 U5891 ( .A1(n9500), .A2(n9499), .ZN(n9498) );
  INV_X1 U5892 ( .A(n4583), .ZN(n7658) );
  AND2_X1 U5893 ( .A1(n7446), .A2(n7553), .ZN(n10004) );
  AOI21_X1 U5894 ( .B1(n7665), .B2(n10196), .A(n7664), .ZN(n7667) );
  AND2_X1 U5895 ( .A1(n4583), .A2(n4582), .ZN(n7661) );
  NAND2_X1 U5896 ( .A1(n7665), .A2(n8294), .ZN(n4582) );
  AND2_X1 U5897 ( .A1(n7661), .A2(n7660), .ZN(n9524) );
  NOR2_X1 U5898 ( .A1(n9530), .A2(n4585), .ZN(n10025) );
  NAND2_X1 U5899 ( .A1(n4575), .A2(n9550), .ZN(n10036) );
  NAND2_X1 U5900 ( .A1(n4575), .A2(n4572), .ZN(n10045) );
  INV_X1 U5901 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9566) );
  NOR2_X1 U5902 ( .A1(n9568), .A2(n9784), .ZN(n9809) );
  INV_X1 U5903 ( .A(n9814), .ZN(n9602) );
  AND2_X1 U5904 ( .A1(n5546), .A2(n5514), .ZN(n9599) );
  NAND2_X1 U5905 ( .A1(n6803), .A2(n6737), .ZN(n9656) );
  NAND2_X1 U5906 ( .A1(n4556), .A2(n4554), .ZN(n9653) );
  INV_X1 U5907 ( .A(n4557), .ZN(n4554) );
  NAND2_X1 U5908 ( .A1(n9703), .A2(n4560), .ZN(n4556) );
  CLKBUF_X1 U5909 ( .A(n9704), .Z(n9706) );
  NAND2_X1 U5910 ( .A1(n5365), .A2(n5364), .ZN(n9852) );
  OR2_X1 U5911 ( .A1(n8363), .A2(n4829), .ZN(n4823) );
  NAND2_X1 U5912 ( .A1(n8153), .A2(n8159), .ZN(n8152) );
  NAND2_X1 U5913 ( .A1(n4846), .A2(n5189), .ZN(n8153) );
  NAND2_X1 U5914 ( .A1(n7926), .A2(n7933), .ZN(n7925) );
  INV_X1 U5915 ( .A(n7854), .ZN(n8044) );
  INV_X1 U5916 ( .A(n9715), .ZN(n10331) );
  NAND2_X1 U5917 ( .A1(n7321), .A2(n5641), .ZN(n7833) );
  NAND2_X1 U5918 ( .A1(n7937), .A2(n9564), .ZN(n10341) );
  NAND2_X1 U5919 ( .A1(n7296), .A2(n7285), .ZN(n9780) );
  NAND2_X1 U5920 ( .A1(n7937), .A2(n7332), .ZN(n9715) );
  INV_X1 U5921 ( .A(n9211), .ZN(n9913) );
  NAND2_X1 U5922 ( .A1(n5473), .A2(n5472), .ZN(n9920) );
  OAI21_X1 U5923 ( .B1(n9703), .B2(n4553), .A(n4551), .ZN(n9643) );
  INV_X1 U5924 ( .A(n7218), .ZN(n9933) );
  AOI21_X1 U5925 ( .B1(n9703), .B2(n5406), .A(n4972), .ZN(n9670) );
  NAND2_X1 U5926 ( .A1(n5350), .A2(n5349), .ZN(n9951) );
  NAND2_X1 U5927 ( .A1(n4545), .A2(n4546), .ZN(n9736) );
  OR2_X1 U5928 ( .A1(n8363), .A2(n4825), .ZN(n4545) );
  NAND2_X1 U5929 ( .A1(n4832), .A2(n5299), .ZN(n9772) );
  NAND2_X1 U5930 ( .A1(n8363), .A2(n5298), .ZN(n4832) );
  INV_X1 U5931 ( .A(n4435), .ZN(n9974) );
  NAND2_X1 U5932 ( .A1(n7824), .A2(n5127), .ZN(n7894) );
  NAND2_X1 U5933 ( .A1(n5576), .A2(n4608), .ZN(n4940) );
  AND2_X1 U5934 ( .A1(n8374), .A2(n9997), .ZN(n7429) );
  INV_X1 U5935 ( .A(n10051), .ZN(n10052) );
  XNOR2_X1 U5936 ( .A(n6526), .B(n6525), .ZN(n9981) );
  OAI22_X1 U5937 ( .A1(n6522), .A2(n6521), .B1(SI_30_), .B2(n6520), .ZN(n6526)
         );
  NOR2_X1 U5938 ( .A1(n4993), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n4833) );
  INV_X1 U5939 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10191) );
  XNOR2_X1 U5940 ( .A(n5591), .B(n5590), .ZN(n8378) );
  INV_X1 U5941 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8373) );
  XNOR2_X1 U5942 ( .A(n5466), .B(n5465), .ZN(n6155) );
  INV_X1 U5943 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8341) );
  INV_X1 U5944 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8300) );
  INV_X1 U5945 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8187) );
  INV_X1 U5946 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10314) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7868) );
  INV_X1 U5948 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7742) );
  INV_X1 U5949 ( .A(n7592), .ZN(n7665) );
  INV_X1 U5950 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7421) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7397) );
  INV_X1 U5952 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7394) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U5954 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4598) );
  NOR2_X1 U5955 ( .A1(n8133), .A2(n8132), .ZN(n10187) );
  NOR2_X1 U5956 ( .A1(n8139), .A2(n8138), .ZN(n10181) );
  OAI21_X1 U5957 ( .B1(n6505), .B2(n8602), .A(n6504), .ZN(n6506) );
  INV_X1 U5958 ( .A(n4644), .ZN(n4643) );
  OAI21_X1 U5959 ( .B1(n8730), .B2(n4298), .A(n8701), .ZN(n4757) );
  AND3_X1 U5960 ( .A1(n4321), .A2(n4965), .A3(n6320), .ZN(n6365) );
  OAI21_X1 U5961 ( .B1(n8987), .B2(n10164), .A(n4721), .ZN(P2_U3486) );
  INV_X1 U5962 ( .A(n4722), .ZN(n4721) );
  OAI21_X1 U5963 ( .B1(n8992), .B2(n8975), .A(n4723), .ZN(n4722) );
  NOR2_X1 U5964 ( .A1(n4375), .A2(n4724), .ZN(n4723) );
  INV_X1 U5965 ( .A(n6831), .ZN(n6832) );
  AOI21_X1 U5966 ( .B1(n4578), .B2(n9564), .A(n4577), .ZN(n4576) );
  OAI21_X1 U5967 ( .B1(n10050), .B2(n9566), .A(n9565), .ZN(n4577) );
  INV_X1 U5968 ( .A(n4420), .ZN(n4419) );
  NAND2_X1 U5969 ( .A1(n8435), .A2(n10344), .ZN(n4418) );
  OAI21_X1 U5970 ( .B1(n8436), .B2(n9793), .A(n4421), .ZN(n4420) );
  OAI22_X1 U5971 ( .A1(n9578), .A2(n9902), .B1(n10073), .B2(n7057), .ZN(n7058)
         );
  NOR2_X1 U5972 ( .A1(n4376), .A2(n4450), .ZN(n4449) );
  NOR2_X1 U5973 ( .A1(n10073), .A2(n5921), .ZN(n4450) );
  NAND2_X1 U5974 ( .A1(n4431), .A2(n9858), .ZN(n4429) );
  NOR2_X1 U5975 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  NOR2_X1 U5976 ( .A1(n10070), .A2(n9907), .ZN(n4567) );
  NOR2_X1 U5977 ( .A1(n9908), .A2(n9978), .ZN(n4568) );
  NAND2_X1 U5978 ( .A1(n4431), .A2(n9952), .ZN(n4430) );
  AND4_X1 U5979 ( .A1(n4834), .A2(n4562), .A3(n4565), .A4(n4988), .ZN(n4295)
         );
  INV_X2 U5980 ( .A(n6966), .ZN(n6211) );
  INV_X2 U5981 ( .A(n5091), .ZN(n5397) );
  AND2_X1 U5982 ( .A1(n6926), .A2(n6980), .ZN(n4296) );
  AOI21_X1 U5983 ( .B1(n9981), .B2(n5397), .A(n4966), .ZN(n6685) );
  OAI21_X1 U5984 ( .B1(n5305), .B2(n4497), .A(n4494), .ZN(n5395) );
  INV_X1 U5985 ( .A(n9912), .ZN(n4431) );
  AND2_X1 U5986 ( .A1(n4908), .A2(n6905), .ZN(n4297) );
  AND2_X1 U5987 ( .A1(n8732), .A2(n4358), .ZN(n4298) );
  OR2_X1 U5988 ( .A1(n6316), .A2(n7587), .ZN(n4299) );
  INV_X1 U5989 ( .A(n4313), .ZN(n4647) );
  OR2_X1 U5990 ( .A1(n7113), .A2(n4798), .ZN(n4300) );
  AND2_X1 U5991 ( .A1(n6467), .A2(n4923), .ZN(n4301) );
  AOI21_X1 U5992 ( .B1(n4830), .B2(n4828), .A(n4341), .ZN(n4827) );
  INV_X1 U5993 ( .A(n4827), .ZN(n4826) );
  INV_X1 U5994 ( .A(n4993), .ZN(n4565) );
  NOR2_X1 U5995 ( .A1(n8972), .A2(n8607), .ZN(n4302) );
  NAND2_X1 U5996 ( .A1(n4357), .A2(n6289), .ZN(n4303) );
  AND2_X1 U5997 ( .A1(n7278), .A2(n9302), .ZN(n4304) );
  NAND2_X1 U5998 ( .A1(n6515), .A2(n5575), .ZN(n8386) );
  INV_X1 U5999 ( .A(n8386), .ZN(n5577) );
  AND2_X1 U6000 ( .A1(n6903), .A2(n6910), .ZN(n8892) );
  INV_X1 U6001 ( .A(n8892), .ZN(n4657) );
  AND2_X1 U6002 ( .A1(n6410), .A2(n6409), .ZN(n4305) );
  AOI21_X1 U6003 ( .B1(n5577), .B2(n5988), .A(n4382), .ZN(n6958) );
  AND2_X1 U6004 ( .A1(n6111), .A2(n4540), .ZN(n4306) );
  AND2_X1 U6005 ( .A1(n4797), .A2(n7113), .ZN(n4307) );
  AND2_X1 U6006 ( .A1(n4505), .A2(n8591), .ZN(n4308) );
  INV_X1 U6007 ( .A(n7743), .ZN(n4631) );
  INV_X1 U6008 ( .A(n5958), .ZN(n6097) );
  INV_X1 U6009 ( .A(n6014), .ZN(n4742) );
  BUF_X1 U6010 ( .A(n5065), .Z(n6530) );
  NAND2_X2 U6011 ( .A1(n5000), .A2(n5002), .ZN(n5065) );
  INV_X2 U6012 ( .A(n6534), .ZN(n5153) );
  NAND2_X1 U6013 ( .A1(n4474), .A2(n4478), .ZN(n5466) );
  NAND2_X1 U6014 ( .A1(n4816), .A2(n8325), .ZN(n9164) );
  INV_X1 U6015 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4624) );
  NAND2_X1 U6016 ( .A1(n8972), .A2(n8607), .ZN(n4309) );
  INV_X1 U6017 ( .A(n6679), .ZN(n6826) );
  AND2_X2 U6018 ( .A1(n4288), .A2(n7270), .ZN(n7110) );
  INV_X2 U6019 ( .A(n7110), .ZN(n8398) );
  NOR2_X1 U6020 ( .A1(n8460), .A2(n8609), .ZN(n4310) );
  INV_X1 U6021 ( .A(n4594), .ZN(n9396) );
  OR2_X1 U6022 ( .A1(n5040), .A2(n4595), .ZN(n4594) );
  INV_X1 U6023 ( .A(n7070), .ZN(n7067) );
  NAND2_X1 U6024 ( .A1(n4610), .A2(n4609), .ZN(n8832) );
  INV_X1 U6025 ( .A(n8249), .ZN(n10063) );
  NAND2_X1 U6026 ( .A1(n4827), .A2(n4823), .ZN(n9762) );
  AND2_X1 U6027 ( .A1(n4922), .A2(n4926), .ZN(n4311) );
  OR2_X1 U6028 ( .A1(n8523), .A2(n8812), .ZN(n4312) );
  OAI21_X1 U6029 ( .B1(n8786), .B2(n6288), .A(n6287), .ZN(n8774) );
  AND2_X1 U6030 ( .A1(n6964), .A2(n4490), .ZN(n4313) );
  NAND2_X1 U6031 ( .A1(n4473), .A2(n4471), .ZN(n5482) );
  NAND2_X1 U6032 ( .A1(n6129), .A2(n6128), .ZN(n6447) );
  AND2_X1 U6033 ( .A1(n7778), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4314) );
  AND2_X1 U6034 ( .A1(n9048), .A2(n8870), .ZN(n4315) );
  INV_X1 U6035 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9077) );
  OR2_X1 U6036 ( .A1(n7777), .A2(n8214), .ZN(n4316) );
  NAND2_X1 U6037 ( .A1(n7614), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4317) );
  INV_X1 U6038 ( .A(n6668), .ZN(n9908) );
  NAND2_X1 U6039 ( .A1(n5530), .A2(n5529), .ZN(n6668) );
  AND2_X1 U6040 ( .A1(n4885), .A2(n6291), .ZN(n4318) );
  AND3_X1 U6041 ( .A1(n5593), .A2(n4989), .A3(n4990), .ZN(n4319) );
  INV_X1 U6042 ( .A(n7011), .ZN(n4613) );
  AND3_X1 U6043 ( .A1(n4676), .A2(n5700), .A3(n5698), .ZN(n4320) );
  OR2_X1 U6044 ( .A1(n8385), .A2(n6321), .ZN(n4321) );
  OR2_X1 U6045 ( .A1(n6905), .A2(n6988), .ZN(n4322) );
  AND2_X1 U6046 ( .A1(n6759), .A2(n7933), .ZN(n4323) );
  AND2_X1 U6047 ( .A1(n4994), .A2(n4962), .ZN(n4324) );
  AND2_X1 U6048 ( .A1(n6576), .A2(n8155), .ZN(n4325) );
  OR2_X1 U6049 ( .A1(n9727), .A2(n4765), .ZN(n4326) );
  AND2_X1 U6050 ( .A1(n6468), .A2(n6469), .ZN(n4327) );
  NAND2_X1 U6051 ( .A1(n5544), .A2(n5543), .ZN(n8419) );
  NOR2_X1 U6052 ( .A1(n9013), .A2(n8812), .ZN(n4328) );
  INV_X1 U6053 ( .A(n7355), .ZN(n4608) );
  AND2_X1 U6054 ( .A1(n6406), .A2(n7719), .ZN(n4329) );
  OR2_X1 U6055 ( .A1(n5118), .A2(n5117), .ZN(n4330) );
  OR2_X1 U6056 ( .A1(n7563), .A2(n7564), .ZN(n4331) );
  OR2_X1 U6057 ( .A1(n7565), .A2(n7566), .ZN(n4332) );
  OR2_X1 U6058 ( .A1(n6465), .A2(n6464), .ZN(n4333) );
  OR2_X1 U6059 ( .A1(n8630), .A2(n10106), .ZN(n4334) );
  INV_X1 U6060 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4751) );
  INV_X1 U6061 ( .A(n6453), .ZN(n4933) );
  AND2_X1 U6062 ( .A1(n9861), .A2(n9361), .ZN(n4335) );
  AND2_X1 U6063 ( .A1(n6807), .A2(n6743), .ZN(n6784) );
  INV_X1 U6064 ( .A(n6784), .ZN(n5537) );
  AND2_X1 U6065 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_9__SCAN_IN), 
        .ZN(n4336) );
  AND2_X1 U6066 ( .A1(n5958), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4337) );
  OR2_X1 U6067 ( .A1(n5324), .A2(n5323), .ZN(n4338) );
  OR2_X1 U6068 ( .A1(n8419), .A2(n8404), .ZN(n6747) );
  INV_X1 U6069 ( .A(n6747), .ZN(n4443) );
  OR2_X1 U6070 ( .A1(n7597), .A2(n7598), .ZN(n4339) );
  INV_X1 U6071 ( .A(n6931), .ZN(n4637) );
  AND2_X1 U6072 ( .A1(n8563), .A2(n8608), .ZN(n4340) );
  AND2_X1 U6073 ( .A1(n9870), .A2(n9362), .ZN(n4341) );
  INV_X1 U6074 ( .A(n9843), .ZN(n9700) );
  INV_X1 U6075 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5923) );
  INV_X1 U6076 ( .A(n4738), .ZN(n4737) );
  NOR2_X1 U6077 ( .A1(n4317), .A2(n6014), .ZN(n4738) );
  OR2_X1 U6078 ( .A1(n9007), .A2(n8526), .ZN(n6996) );
  INV_X1 U6079 ( .A(n6996), .ZN(n4601) );
  AND2_X1 U6080 ( .A1(n9931), .A2(n9118), .ZN(n4342) );
  AND2_X1 U6081 ( .A1(n6685), .A2(n9347), .ZN(n6754) );
  OR2_X1 U6082 ( .A1(n4509), .A2(n4312), .ZN(n4343) );
  INV_X1 U6083 ( .A(n4719), .ZN(n4718) );
  NAND2_X1 U6084 ( .A1(n8775), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U6085 ( .A1(n7259), .A2(n7258), .ZN(n4344) );
  NOR2_X1 U6086 ( .A1(n9065), .A2(n8442), .ZN(n4345) );
  INV_X1 U6087 ( .A(n4516), .ZN(n4515) );
  NAND2_X1 U6088 ( .A1(n6412), .A2(n8107), .ZN(n4516) );
  AND2_X1 U6089 ( .A1(n4529), .A2(n4527), .ZN(n4346) );
  AND2_X1 U6090 ( .A1(n7790), .A2(n10079), .ZN(n4347) );
  OR2_X1 U6091 ( .A1(n9149), .A2(n4392), .ZN(n4391) );
  INV_X1 U6092 ( .A(n9931), .ZN(n9662) );
  AND2_X1 U6093 ( .A1(n5436), .A2(n5435), .ZN(n9931) );
  OR2_X1 U6094 ( .A1(n5773), .A2(n5724), .ZN(n4348) );
  INV_X1 U6095 ( .A(n8878), .ZN(n4908) );
  AND3_X1 U6096 ( .A1(n7002), .A2(n10098), .A3(n7641), .ZN(n4349) );
  NAND2_X1 U6097 ( .A1(n4848), .A2(n8837), .ZN(n6928) );
  AND2_X1 U6098 ( .A1(n5164), .A2(SI_6_), .ZN(n4350) );
  AND2_X1 U6099 ( .A1(n5287), .A2(SI_13_), .ZN(n4351) );
  AND2_X1 U6100 ( .A1(n7492), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4352) );
  INV_X1 U6101 ( .A(n6461), .ZN(n4930) );
  AND2_X1 U6102 ( .A1(n5377), .A2(SI_18_), .ZN(n4353) );
  AND2_X1 U6103 ( .A1(n4695), .A2(n4309), .ZN(n4354) );
  INV_X1 U6104 ( .A(n4497), .ZN(n4496) );
  NAND2_X1 U6105 ( .A1(n4874), .A2(n5375), .ZN(n4497) );
  INV_X1 U6106 ( .A(n4481), .ZN(n4480) );
  NAND2_X1 U6107 ( .A1(n5428), .A2(n4482), .ZN(n4481) );
  OAI21_X1 U6108 ( .B1(n8200), .B2(n4800), .A(n7109), .ZN(n4799) );
  OAI21_X1 U6109 ( .B1(n4635), .B2(n6931), .A(n6930), .ZN(n4632) );
  INV_X1 U6110 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U6111 ( .A1(n6035), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4355) );
  AND2_X1 U6112 ( .A1(n4693), .A2(n4309), .ZN(n4356) );
  OR2_X1 U6113 ( .A1(n8995), .A2(n8776), .ZN(n4357) );
  AND2_X1 U6114 ( .A1(n8733), .A2(n8731), .ZN(n4358) );
  INV_X1 U6115 ( .A(n8159), .ZN(n4845) );
  AND2_X1 U6116 ( .A1(n6737), .A2(n9652), .ZN(n4359) );
  AND2_X1 U6117 ( .A1(n4524), .A2(n6453), .ZN(n4360) );
  AND2_X1 U6118 ( .A1(n4988), .A2(n4565), .ZN(n4361) );
  AND2_X1 U6119 ( .A1(n6934), .A2(n4637), .ZN(n4362) );
  AND2_X1 U6120 ( .A1(n6577), .A2(n8158), .ZN(n8258) );
  INV_X1 U6121 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U6122 ( .A1(n9951), .A2(n9360), .ZN(n4363) );
  AND2_X1 U6123 ( .A1(n4624), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4364) );
  INV_X1 U6124 ( .A(n8823), .ZN(n8819) );
  NAND2_X1 U6125 ( .A1(n6928), .A2(n6925), .ZN(n8823) );
  AND2_X1 U6126 ( .A1(n6960), .A2(n6959), .ZN(n4365) );
  INV_X1 U6127 ( .A(n4830), .ZN(n4829) );
  NOR2_X1 U6128 ( .A1(n4831), .A2(n5320), .ZN(n4830) );
  AND2_X1 U6129 ( .A1(n8465), .A2(n6450), .ZN(n4366) );
  OR2_X1 U6130 ( .A1(n4664), .A2(n4663), .ZN(n4367) );
  AND2_X1 U6131 ( .A1(n4772), .A2(n8249), .ZN(n4368) );
  AND2_X1 U6132 ( .A1(n4895), .A2(n6942), .ZN(n4369) );
  NAND2_X1 U6133 ( .A1(n8906), .A2(n4367), .ZN(n4370) );
  AND2_X1 U6134 ( .A1(n4632), .A2(n6934), .ZN(n4371) );
  INV_X1 U6135 ( .A(n9606), .ZN(n4945) );
  OR2_X1 U6136 ( .A1(n9920), .A2(n9119), .ZN(n9606) );
  OAI21_X1 U6137 ( .B1(n9908), .B2(n9331), .A(n7302), .ZN(n7303) );
  NAND2_X1 U6138 ( .A1(n6964), .A2(n4491), .ZN(n4372) );
  INV_X1 U6139 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5012) );
  INV_X1 U6140 ( .A(n8678), .ZN(n4628) );
  NAND2_X1 U6141 ( .A1(n6474), .A2(n6473), .ZN(n8591) );
  INV_X1 U6142 ( .A(n10075), .ZN(n4401) );
  INV_X1 U6143 ( .A(n9963), .ZN(n9952) );
  NAND2_X1 U6144 ( .A1(n7869), .A2(n4515), .ZN(n8028) );
  AND2_X1 U6145 ( .A1(n4810), .A2(n4807), .ZN(n4373) );
  AOI21_X1 U6146 ( .B1(n5577), .B2(n5576), .A(n4976), .ZN(n8432) );
  INV_X1 U6147 ( .A(n8432), .ZN(n4777) );
  NAND2_X1 U6148 ( .A1(n7848), .A2(n5085), .ZN(n7824) );
  AND2_X1 U6149 ( .A1(n5672), .A2(n8188), .ZN(n7063) );
  OR2_X1 U6150 ( .A1(n7961), .A2(n5786), .ZN(n4374) );
  AND2_X1 U6151 ( .A1(n8989), .A2(n8967), .ZN(n4375) );
  NOR2_X1 U6152 ( .A1(n8066), .A2(n4770), .ZN(n8292) );
  AND2_X1 U6153 ( .A1(n5775), .A2(n5777), .ZN(n6035) );
  INV_X1 U6154 ( .A(n6035), .ZN(n7699) );
  NOR2_X1 U6155 ( .A1(n9908), .A2(n9902), .ZN(n4376) );
  AND2_X1 U6156 ( .A1(n7109), .A2(n4800), .ZN(n4377) );
  AND2_X1 U6157 ( .A1(n4913), .A2(n7720), .ZN(n4378) );
  INV_X1 U6158 ( .A(n4767), .ZN(n8364) );
  NOR2_X1 U6159 ( .A1(n8066), .A2(n4768), .ZN(n4767) );
  INV_X1 U6160 ( .A(n4510), .ZN(n4509) );
  NAND2_X1 U6161 ( .A1(n8523), .A2(n8812), .ZN(n4510) );
  AND2_X1 U6162 ( .A1(n7917), .A2(n4377), .ZN(n4379) );
  AND2_X1 U6163 ( .A1(n6368), .A2(n6367), .ZN(n4380) );
  AND2_X1 U6164 ( .A1(n4536), .A2(n4535), .ZN(n4381) );
  INV_X1 U6165 ( .A(n6617), .ZN(n4951) );
  INV_X1 U6166 ( .A(n7543), .ZN(n4731) );
  INV_X1 U6167 ( .A(n8720), .ZN(n4629) );
  INV_X1 U6168 ( .A(n9885), .ZN(n4771) );
  AND2_X2 U6169 ( .A1(n5638), .A2(n5920), .ZN(n10070) );
  AND3_X2 U6170 ( .A1(n5920), .A2(n7327), .A3(n7328), .ZN(n10073) );
  NOR2_X1 U6171 ( .A1(n6976), .A2(n9085), .ZN(n4382) );
  AND2_X1 U6172 ( .A1(n7459), .A2(n6308), .ZN(n8701) );
  INV_X1 U6173 ( .A(n10043), .ZN(n10030) );
  INV_X1 U6174 ( .A(n9194), .ZN(n4809) );
  INV_X1 U6175 ( .A(n4573), .ZN(n4572) );
  OR2_X1 U6176 ( .A1(n10035), .A2(n4574), .ZN(n4573) );
  NOR2_X1 U6177 ( .A1(n4655), .A2(n4653), .ZN(n7737) );
  INV_X1 U6178 ( .A(n7737), .ZN(n4673) );
  INV_X1 U6179 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4995) );
  INV_X1 U6180 ( .A(n8019), .ZN(n7028) );
  INV_X1 U6181 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4778) );
  INV_X1 U6182 ( .A(n7071), .ZN(n6693) );
  NAND2_X1 U6183 ( .A1(n5660), .A2(n6690), .ZN(n9671) );
  AOI21_X1 U6184 ( .B1(n8728), .B2(n8729), .A(n4406), .ZN(n5832) );
  OAI21_X1 U6185 ( .B1(n9906), .B2(n7060), .A(n4449), .ZN(P1_U3549) );
  OAI21_X1 U6186 ( .B1(n9906), .B2(n6383), .A(n4566), .ZN(P1_U3517) );
  NAND2_X1 U6187 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  NAND2_X1 U6188 ( .A1(n4422), .A2(n8412), .ZN(n9580) );
  NAND2_X1 U6189 ( .A1(n8649), .A2(n5792), .ZN(n5796) );
  NOR2_X2 U6190 ( .A1(n7950), .A2(n7951), .ZN(n7949) );
  NAND2_X1 U6191 ( .A1(n4758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5014) );
  NAND2_X1 U6192 ( .A1(n4599), .A2(n4893), .ZN(n8756) );
  NAND2_X1 U6193 ( .A1(n8890), .A2(n6910), .ZN(n4907) );
  AND3_X2 U6194 ( .A1(n4674), .A2(n4675), .A3(n4320), .ZN(n4426) );
  NOR2_X2 U6195 ( .A1(n9580), .A2(n4386), .ZN(n7061) );
  NAND2_X1 U6196 ( .A1(n4387), .A2(n8154), .ZN(n6573) );
  NAND2_X1 U6197 ( .A1(n6572), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U6198 ( .A1(n4411), .A2(n6676), .ZN(n6680) );
  NAND2_X1 U6199 ( .A1(n4469), .A2(n6385), .ZN(n4468) );
  NAND2_X1 U6200 ( .A1(n4865), .A2(n5190), .ZN(n4403) );
  AOI21_X2 U6201 ( .B1(n8076), .B2(n8078), .A(n6057), .ZN(n8189) );
  OAI211_X1 U6202 ( .C1(n6574), .C2(n6826), .A(n4417), .B(n6575), .ZN(n6582)
         );
  NAND2_X1 U6203 ( .A1(n4416), .A2(n6679), .ZN(n4415) );
  NAND2_X1 U6204 ( .A1(n4415), .A2(n4414), .ZN(n6604) );
  AOI21_X1 U6205 ( .B1(n6638), .B2(n6637), .A(n6636), .ZN(n6641) );
  AOI21_X1 U6206 ( .B1(n6689), .B2(n6688), .A(n8340), .ZN(n6796) );
  AOI21_X1 U6207 ( .B1(n6651), .B2(n9652), .A(n6650), .ZN(n6658) );
  NAND2_X1 U6208 ( .A1(n5915), .A2(n6784), .ZN(n6375) );
  INV_X1 U6209 ( .A(n4592), .ZN(n4591) );
  NAND2_X1 U6210 ( .A1(n4580), .A2(n5672), .ZN(n4579) );
  AND2_X2 U6211 ( .A1(n4391), .A2(n4390), .ZN(n9179) );
  NAND2_X1 U6212 ( .A1(n4841), .A2(n4843), .ZN(n8001) );
  NAND3_X2 U6213 ( .A1(n4543), .A2(n4542), .A3(n5359), .ZN(n9719) );
  NAND2_X2 U6214 ( .A1(n8309), .A2(n5284), .ZN(n8363) );
  AND2_X1 U6215 ( .A1(n5188), .A2(n5187), .ZN(n5189) );
  NAND3_X1 U6216 ( .A1(n4395), .A2(n4380), .A3(n6370), .ZN(P1_U3551) );
  NAND2_X2 U6217 ( .A1(n8004), .A2(n6594), .ZN(n8062) );
  NAND2_X2 U6218 ( .A1(n4950), .A2(n4948), .ZN(n9720) );
  AOI21_X2 U6219 ( .B1(n5682), .B2(n9778), .A(n5681), .ZN(n8427) );
  NAND2_X1 U6220 ( .A1(n6369), .A2(n10073), .ZN(n4395) );
  AOI21_X1 U6221 ( .B1(n4659), .B2(n4370), .A(n4657), .ZN(n4656) );
  OR2_X1 U6222 ( .A1(n6993), .A2(n4640), .ZN(n4616) );
  NAND2_X1 U6223 ( .A1(n4863), .A2(n5229), .ZN(n4486) );
  INV_X1 U6224 ( .A(n4867), .ZN(n4866) );
  NOR2_X1 U6225 ( .A1(n6897), .A2(n6898), .ZN(n4662) );
  NAND2_X1 U6226 ( .A1(n5251), .A2(n4861), .ZN(n4855) );
  NAND2_X1 U6227 ( .A1(n4855), .A2(n4858), .ZN(n5286) );
  AOI21_X1 U6228 ( .B1(n4633), .B2(n4427), .A(n4371), .ZN(n6949) );
  MUX2_X1 U6229 ( .A(n6868), .B(n6867), .S(n6980), .Z(n6872) );
  NAND2_X1 U6230 ( .A1(n7001), .A2(n6385), .ZN(n6838) );
  NAND2_X1 U6231 ( .A1(n5938), .A2(n4654), .ZN(n4653) );
  NAND2_X4 U6232 ( .A1(n5927), .A2(n5929), .ZN(n6969) );
  NAND2_X1 U6233 ( .A1(n4424), .A2(n6907), .ZN(n6915) );
  NAND2_X1 U6234 ( .A1(n4652), .A2(n4651), .ZN(n4650) );
  NOR2_X1 U6235 ( .A1(n6922), .A2(n4296), .ZN(n4634) );
  OAI21_X1 U6236 ( .B1(n6985), .B2(n6984), .A(n6983), .ZN(n6993) );
  NAND2_X2 U6237 ( .A1(n7684), .A2(n5822), .ZN(n5823) );
  XNOR2_X2 U6238 ( .A(n5750), .B(n5749), .ZN(n7348) );
  NAND3_X1 U6239 ( .A1(n4349), .A2(n4399), .A3(n4398), .ZN(n4397) );
  NAND2_X1 U6240 ( .A1(n6378), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U6241 ( .A1(n4451), .A2(n4374), .ZN(n4732) );
  AOI21_X2 U6242 ( .B1(n7902), .B2(P2_REG2_REG_11__SCAN_IN), .A(n4405), .ZN(
        n7950) );
  XNOR2_X2 U6243 ( .A(n5783), .B(n6048), .ZN(n7902) );
  NAND2_X1 U6244 ( .A1(n5821), .A2(n5820), .ZN(n7685) );
  NAND2_X1 U6245 ( .A1(n4408), .A2(n4407), .ZN(n4580) );
  NAND2_X1 U6246 ( .A1(n9562), .A2(n10037), .ZN(n4407) );
  INV_X1 U6247 ( .A(n4409), .ZN(n4408) );
  NAND2_X1 U6248 ( .A1(n4579), .A2(n4576), .ZN(P1_U3262) );
  NAND2_X1 U6249 ( .A1(n9520), .A2(n9519), .ZN(n9539) );
  NOR2_X1 U6250 ( .A1(n10021), .A2(n9518), .ZN(n9520) );
  OAI21_X1 U6251 ( .B1(n5038), .B2(n4598), .A(n4596), .ZN(n4595) );
  NAND3_X1 U6252 ( .A1(n4410), .A2(n4324), .A3(n5012), .ZN(n4563) );
  INV_X1 U6253 ( .A(n4987), .ZN(n4410) );
  OAI21_X1 U6254 ( .B1(n4826), .B2(n4830), .A(n9753), .ZN(n4825) );
  NAND2_X1 U6255 ( .A1(n5503), .A2(n4839), .ZN(n4838) );
  AND2_X1 U6256 ( .A1(n6674), .A2(n4413), .ZN(n4412) );
  NAND2_X1 U6257 ( .A1(n4854), .A2(n4853), .ZN(n5302) );
  NAND2_X1 U6258 ( .A1(n4419), .A2(n4418), .ZN(P1_U3356) );
  OAI21_X4 U6259 ( .B1(n9719), .B2(n5373), .A(n5374), .ZN(n9703) );
  NAND2_X1 U6260 ( .A1(n5116), .A2(n5115), .ZN(n5143) );
  NAND2_X1 U6261 ( .A1(n9671), .A2(n6733), .ZN(n6801) );
  NAND2_X2 U6262 ( .A1(n8062), .A2(n8071), .ZN(n8284) );
  NAND2_X1 U6263 ( .A1(n4736), .A2(n4317), .ZN(n4743) );
  NAND2_X1 U6264 ( .A1(n6801), .A2(n4359), .ZN(n9636) );
  NAND2_X1 U6265 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(n8709), .ZN(n8732) );
  NOR2_X1 U6266 ( .A1(n8730), .A2(n4432), .ZN(n5803) );
  NAND3_X1 U6267 ( .A1(n4668), .A2(n4322), .A3(n4908), .ZN(n4424) );
  NAND2_X1 U6268 ( .A1(n4425), .A2(n5837), .ZN(n7481) );
  NAND2_X1 U6269 ( .A1(n7577), .A2(n7578), .ZN(n4425) );
  NAND2_X2 U6270 ( .A1(n5876), .A2(n7954), .ZN(n8640) );
  NAND2_X2 U6271 ( .A1(n5884), .A2(n8656), .ZN(n8674) );
  AND2_X4 U6272 ( .A1(n4426), .A2(n4677), .ZN(n5712) );
  NAND2_X1 U6273 ( .A1(n6951), .A2(n8793), .ZN(n4652) );
  AOI21_X1 U6274 ( .B1(n4650), .B2(n4649), .A(n4365), .ZN(n4648) );
  AND2_X1 U6275 ( .A1(n4634), .A2(n4362), .ZN(n4427) );
  INV_X1 U6276 ( .A(n6308), .ZN(n7032) );
  NAND2_X1 U6277 ( .A1(n9816), .A2(n4429), .ZN(P1_U3548) );
  NAND2_X1 U6278 ( .A1(n9911), .A2(n4430), .ZN(P1_U3516) );
  XNOR2_X2 U6279 ( .A(n7073), .B(n7334), .ZN(n6760) );
  AOI21_X2 U6280 ( .B1(n8732), .B2(n8733), .A(n8731), .ZN(n8730) );
  OAI21_X1 U6281 ( .B1(n4313), .B2(n4470), .A(n4468), .ZN(n7027) );
  OAI211_X1 U6282 ( .C1(n4643), .C2(n4642), .A(n4460), .B(n4459), .ZN(P2_U3296) );
  NAND2_X2 U6283 ( .A1(n5664), .A2(n6727), .ZN(n9621) );
  XNOR2_X2 U6284 ( .A(n5192), .B(n5191), .ZN(n7378) );
  NAND3_X1 U6285 ( .A1(n5691), .A2(n5690), .A3(n4433), .ZN(P1_U3519) );
  NAND2_X1 U6286 ( .A1(n5668), .A2(n6802), .ZN(n5915) );
  NAND2_X1 U6287 ( .A1(n4953), .A2(n4954), .ZN(n7886) );
  NAND2_X1 U6288 ( .A1(n4958), .A2(n4957), .ZN(n5671) );
  INV_X1 U6289 ( .A(n7615), .ZN(n4736) );
  INV_X1 U6290 ( .A(n7949), .ZN(n4451) );
  NAND2_X1 U6291 ( .A1(n5174), .A2(n4869), .ZN(n4865) );
  INV_X2 U6292 ( .A(n5936), .ZN(n6245) );
  NAND2_X2 U6293 ( .A1(n5934), .A2(n4436), .ZN(n5936) );
  NOR2_X2 U6294 ( .A1(n4337), .A2(n4437), .ZN(n4436) );
  NAND2_X1 U6295 ( .A1(n5933), .A2(n5932), .ZN(n4437) );
  NAND2_X1 U6296 ( .A1(n8786), .A2(n6287), .ZN(n4715) );
  NAND2_X1 U6297 ( .A1(n4685), .A2(n4684), .ZN(n6272) );
  NAND2_X1 U6298 ( .A1(n4692), .A2(n4691), .ZN(n8314) );
  NAND2_X4 U6299 ( .A1(n4439), .A2(n7067), .ZN(n8403) );
  INV_X2 U6300 ( .A(n9351), .ZN(n6540) );
  NOR2_X2 U6301 ( .A1(n5474), .A2(n9241), .ZN(n5491) );
  OAI21_X1 U6302 ( .B1(n7149), .B2(n4819), .A(n7148), .ZN(n4818) );
  OAI21_X2 U6303 ( .B1(n7183), .B2(n4787), .A(n4786), .ZN(n9144) );
  NAND2_X1 U6304 ( .A1(n8651), .A2(n8650), .ZN(n8649) );
  NAND2_X1 U6305 ( .A1(n4741), .A2(n4740), .ZN(n7672) );
  NAND2_X1 U6306 ( .A1(n5805), .A2(n8701), .ZN(n5914) );
  NAND2_X2 U6307 ( .A1(n5866), .A2(n7693), .ZN(n7773) );
  NOR2_X1 U6308 ( .A1(n4756), .A2(n4754), .ZN(n4753) );
  NOR2_X1 U6309 ( .A1(n5053), .A2(n7557), .ZN(n4453) );
  NAND2_X1 U6310 ( .A1(n6589), .A2(n4454), .ZN(n6590) );
  NAND3_X1 U6311 ( .A1(n6662), .A2(n6664), .A3(n4455), .ZN(n6673) );
  NOR2_X1 U6312 ( .A1(n4456), .A2(n6665), .ZN(n4455) );
  NAND2_X2 U6313 ( .A1(n5171), .A2(n5170), .ZN(n5174) );
  NAND2_X2 U6314 ( .A1(n5181), .A2(n5180), .ZN(n9172) );
  NAND2_X1 U6315 ( .A1(n5507), .A2(n4464), .ZN(n4463) );
  NAND3_X1 U6316 ( .A1(n4372), .A2(n7022), .A3(n4604), .ZN(n4469) );
  NAND4_X1 U6317 ( .A1(n7018), .A2(n7017), .A3(n7047), .A4(n7024), .ZN(n4470)
         );
  NAND2_X1 U6318 ( .A1(n5430), .A2(n4475), .ZN(n4473) );
  NAND2_X1 U6319 ( .A1(n5430), .A2(n4480), .ZN(n4474) );
  NAND2_X1 U6320 ( .A1(n5174), .A2(n4483), .ZN(n4484) );
  INV_X1 U6321 ( .A(n4486), .ZN(n4488) );
  NAND3_X1 U6322 ( .A1(n4485), .A2(n4856), .A3(n4484), .ZN(n4854) );
  NAND2_X1 U6323 ( .A1(n4486), .A2(n5232), .ZN(n4485) );
  NAND2_X1 U6324 ( .A1(n4487), .A2(n5232), .ZN(n5251) );
  NAND2_X1 U6325 ( .A1(n4488), .A2(n4489), .ZN(n4487) );
  AOI21_X1 U6326 ( .B1(n8986), .B2(n8603), .A(n4492), .ZN(n4491) );
  NAND2_X1 U6327 ( .A1(n4493), .A2(n8603), .ZN(n7023) );
  NAND2_X1 U6328 ( .A1(n5305), .A2(n4501), .ZN(n5326) );
  NAND2_X1 U6329 ( .A1(n5305), .A2(n5304), .ZN(n5322) );
  XNOR2_X1 U6330 ( .A(n8524), .B(n8523), .ZN(n8525) );
  OAI211_X1 U6331 ( .C1(n8524), .C2(n4508), .A(n4308), .B(n4503), .ZN(n4511)
         );
  NAND3_X1 U6332 ( .A1(n8524), .A2(n4504), .A3(n4312), .ZN(n4503) );
  NAND2_X1 U6333 ( .A1(n4511), .A2(n8532), .ZN(P2_U3169) );
  OAI21_X1 U6334 ( .B1(n7869), .B2(n4514), .A(n4512), .ZN(n6424) );
  AND2_X1 U6335 ( .A1(n5769), .A2(n4517), .ZN(n5799) );
  NAND2_X1 U6336 ( .A1(n5769), .A2(n4519), .ZN(n5725) );
  NAND2_X1 U6337 ( .A1(n8574), .A2(n4360), .ZN(n4523) );
  NAND2_X2 U6338 ( .A1(n6432), .A2(n6431), .ZN(n8437) );
  OAI21_X2 U6339 ( .B1(n6387), .B2(n6386), .A(n4526), .ZN(n6396) );
  XNOR2_X2 U6340 ( .A(n5726), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U6341 ( .A1(n6072), .A2(n4381), .ZN(n6104) );
  NAND2_X1 U6342 ( .A1(n6112), .A2(n4538), .ZN(n6138) );
  NAND3_X1 U6343 ( .A1(n5979), .A2(n5969), .A3(n5968), .ZN(n5993) );
  NAND2_X1 U6344 ( .A1(n4544), .A2(n8363), .ZN(n4542) );
  INV_X1 U6345 ( .A(n9703), .ZN(n4550) );
  OAI21_X2 U6346 ( .B1(n4550), .B2(n4549), .A(n4547), .ZN(n9641) );
  AND2_X1 U6347 ( .A1(n5186), .A2(n8241), .ZN(n4847) );
  NOR2_X1 U6348 ( .A1(n4563), .A2(n5099), .ZN(n4562) );
  NAND3_X1 U6349 ( .A1(n5307), .A2(n4564), .A3(n4834), .ZN(n5011) );
  AND2_X2 U6350 ( .A1(n5138), .A2(n4988), .ZN(n5307) );
  INV_X1 U6351 ( .A(n4834), .ZN(n5588) );
  OAI21_X1 U6352 ( .B1(n9548), .B2(n4573), .A(n4569), .ZN(n9552) );
  INV_X1 U6353 ( .A(n9530), .ZN(n4584) );
  NAND2_X1 U6354 ( .A1(n4584), .A2(n4586), .ZN(n10026) );
  INV_X1 U6355 ( .A(n9529), .ZN(n4587) );
  NAND2_X1 U6356 ( .A1(n9400), .A2(n4588), .ZN(n4590) );
  NAND2_X1 U6357 ( .A1(n4590), .A2(n4591), .ZN(n9423) );
  MUX2_X1 U6358 ( .A(n8171), .B(P1_REG2_REG_2__SCAN_IN), .S(n4594), .Z(n9402)
         );
  NAND3_X1 U6359 ( .A1(n4369), .A2(n4600), .A3(n4602), .ZN(n4599) );
  NAND2_X1 U6360 ( .A1(n8809), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U6361 ( .A1(n7021), .A2(n7020), .ZN(n4604) );
  OR2_X1 U6362 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  INV_X2 U6363 ( .A(n6316), .ZN(n4607) );
  NAND2_X1 U6364 ( .A1(n6316), .A2(n5118), .ZN(n6229) );
  INV_X1 U6365 ( .A(n7735), .ZN(n6244) );
  AND2_X2 U6366 ( .A1(n6839), .A2(n6837), .ZN(n7735) );
  INV_X1 U6367 ( .A(n5817), .ZN(n4620) );
  NAND2_X1 U6368 ( .A1(n5748), .A2(n4751), .ZN(n5756) );
  NAND2_X1 U6369 ( .A1(n5748), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U6370 ( .A1(n5748), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5754) );
  NOR2_X1 U6371 ( .A1(n5748), .A2(n4623), .ZN(n5753) );
  NAND2_X1 U6372 ( .A1(n5755), .A2(n4364), .ZN(n5807) );
  XNOR2_X2 U6373 ( .A(n5823), .B(n6035), .ZN(n7691) );
  INV_X1 U6374 ( .A(n6923), .ZN(n4633) );
  NAND3_X1 U6375 ( .A1(n6993), .A2(n6992), .A3(n4638), .ZN(n4639) );
  NAND2_X1 U6376 ( .A1(n4641), .A2(n6994), .ZN(n4640) );
  INV_X1 U6377 ( .A(n4646), .ZN(n4641) );
  INV_X1 U6378 ( .A(n6994), .ZN(n4642) );
  OAI21_X1 U6379 ( .B1(n6992), .B2(n4646), .A(n4645), .ZN(n4644) );
  NAND2_X1 U6380 ( .A1(n4658), .A2(n4656), .ZN(n6911) );
  NAND2_X1 U6381 ( .A1(n6899), .A2(n4659), .ZN(n4658) );
  INV_X1 U6382 ( .A(n6897), .ZN(n4664) );
  NAND3_X1 U6383 ( .A1(n6904), .A2(n6988), .A3(n6905), .ZN(n4668) );
  AND2_X1 U6384 ( .A1(n4910), .A2(n5730), .ZN(n4671) );
  NAND2_X2 U6385 ( .A1(n6842), .A2(n6843), .ZN(n7624) );
  NAND2_X1 U6386 ( .A1(n4672), .A2(n6246), .ZN(n7626) );
  NAND2_X1 U6387 ( .A1(n7795), .A2(n4678), .ZN(n4679) );
  OAI21_X1 U6388 ( .B1(n8891), .B2(n4688), .A(n4686), .ZN(n8869) );
  AOI21_X1 U6389 ( .B1(n4686), .B2(n4688), .A(n4908), .ZN(n4684) );
  NAND2_X1 U6390 ( .A1(n8891), .A2(n4686), .ZN(n4685) );
  OAI21_X1 U6391 ( .B1(n8891), .B2(n6270), .A(n6269), .ZN(n8884) );
  NAND2_X1 U6392 ( .A1(n6270), .A2(n6269), .ZN(n4690) );
  NAND2_X1 U6393 ( .A1(n8053), .A2(n4356), .ZN(n4692) );
  NAND2_X1 U6394 ( .A1(n8861), .A2(n4702), .ZN(n4701) );
  NAND2_X1 U6395 ( .A1(n4871), .A2(n4713), .ZN(n4712) );
  NAND2_X1 U6396 ( .A1(n4871), .A2(n6286), .ZN(n8786) );
  NAND2_X1 U6397 ( .A1(n4712), .A2(n4716), .ZN(n4885) );
  OR2_X1 U6398 ( .A1(n6976), .A2(n7356), .ZN(n5955) );
  AND2_X1 U6399 ( .A1(n5926), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5949) );
  OAI22_X1 U6400 ( .A1(n7642), .A2(n6250), .B1(n7629), .B2(n10121), .ZN(n10090) );
  NAND2_X2 U6401 ( .A1(n5952), .A2(n5951), .ZN(n8615) );
  OAI21_X1 U6402 ( .B1(n10081), .B2(n6257), .A(n6256), .ZN(n7974) );
  INV_X1 U6403 ( .A(n4886), .ZN(n8757) );
  NAND2_X1 U6404 ( .A1(n4896), .A2(n6349), .ZN(n6351) );
  OAI21_X2 U6405 ( .B1(n8635), .B2(n8323), .A(n4730), .ZN(n8651) );
  NAND2_X1 U6406 ( .A1(n4732), .A2(n4731), .ZN(n4730) );
  NAND3_X1 U6407 ( .A1(n4735), .A2(n4734), .A3(n4733), .ZN(n4741) );
  NAND2_X1 U6408 ( .A1(n7615), .A2(n4742), .ZN(n4733) );
  NAND3_X1 U6409 ( .A1(n4735), .A2(n4737), .A3(n4733), .ZN(n7511) );
  NAND2_X1 U6410 ( .A1(n4317), .A2(n6014), .ZN(n4739) );
  NAND2_X1 U6411 ( .A1(n4743), .A2(n4742), .ZN(n4740) );
  OAI21_X2 U6412 ( .B1(n5776), .B2(n4748), .A(n4744), .ZN(n4747) );
  NOR2_X1 U6413 ( .A1(n5923), .A2(n4751), .ZN(n4749) );
  NAND2_X1 U6414 ( .A1(n5923), .A2(n4751), .ZN(n4750) );
  OAI211_X1 U6415 ( .C1(n8749), .C2(n8748), .A(n4757), .B(n4753), .ZN(P2_U3200) );
  NAND4_X1 U6416 ( .A1(n4834), .A2(n4833), .A3(n5138), .A4(n4988), .ZN(n4758)
         );
  AND4_X2 U6417 ( .A1(n4762), .A2(n4761), .A3(n4760), .A4(n4759), .ZN(n4988)
         );
  INV_X1 U6418 ( .A(n4763), .ZN(n9660) );
  AND2_X2 U6419 ( .A1(n4368), .A2(n7939), .ZN(n8267) );
  AND2_X1 U6420 ( .A1(n9597), .A2(n4773), .ZN(n5685) );
  AND2_X1 U6421 ( .A1(n9597), .A2(n9602), .ZN(n9598) );
  NAND2_X1 U6422 ( .A1(n9597), .A2(n4774), .ZN(n6509) );
  NAND2_X1 U6423 ( .A1(n4781), .A2(n4780), .ZN(P1_U3214) );
  AOI21_X1 U6424 ( .B1(n9320), .B2(n4304), .A(n7303), .ZN(n4780) );
  NAND2_X1 U6425 ( .A1(n7275), .A2(n4782), .ZN(n4781) );
  NAND2_X1 U6426 ( .A1(n9320), .A2(n7278), .ZN(n8422) );
  NAND2_X1 U6427 ( .A1(n4783), .A2(n4784), .ZN(n7232) );
  NAND2_X1 U6428 ( .A1(n7183), .A2(n4786), .ZN(n4783) );
  NAND2_X1 U6429 ( .A1(n7183), .A2(n7184), .ZN(n9101) );
  OR2_X1 U6430 ( .A1(n7183), .A2(n7184), .ZN(n9102) );
  INV_X1 U6431 ( .A(n9104), .ZN(n4788) );
  NAND2_X1 U6432 ( .A1(n4789), .A2(n4790), .ZN(n9318) );
  NAND2_X1 U6433 ( .A1(n9236), .A2(n4791), .ZN(n4789) );
  NAND2_X1 U6434 ( .A1(n4796), .A2(n9136), .ZN(n4794) );
  INV_X1 U6435 ( .A(n7113), .ZN(n4800) );
  NAND2_X1 U6436 ( .A1(n4806), .A2(n4808), .ZN(n7171) );
  NAND2_X1 U6437 ( .A1(n8328), .A2(n4810), .ZN(n4806) );
  AND3_X1 U6438 ( .A1(n5138), .A2(n4988), .A3(n4822), .ZN(n5347) );
  NAND3_X1 U6439 ( .A1(n5139), .A2(n4988), .A3(n10207), .ZN(n5309) );
  AND2_X2 U6440 ( .A1(n4319), .A2(n4991), .ZN(n4834) );
  NAND3_X1 U6441 ( .A1(n4834), .A2(n4361), .A3(n5139), .ZN(n5602) );
  NAND2_X1 U6442 ( .A1(n4838), .A2(n5520), .ZN(n5917) );
  AOI21_X2 U6443 ( .B1(n4838), .B2(n4836), .A(n4835), .ZN(n6371) );
  INV_X1 U6444 ( .A(n4842), .ZN(n4841) );
  OAI21_X1 U6445 ( .B1(n5189), .B2(n4845), .A(n5208), .ZN(n4842) );
  NAND2_X1 U6446 ( .A1(n4844), .A2(n8239), .ZN(n4843) );
  NAND2_X1 U6447 ( .A1(n8239), .A2(n4847), .ZN(n4846) );
  NAND3_X1 U6448 ( .A1(n7824), .A2(n5127), .A3(n7896), .ZN(n5152) );
  NAND3_X1 U6449 ( .A1(n10002), .A2(n5674), .A3(n9409), .ZN(n5081) );
  XNOR2_X2 U6450 ( .A(n5014), .B(n4994), .ZN(n10002) );
  NAND2_X1 U6451 ( .A1(n4849), .A2(n4850), .ZN(n5171) );
  NAND3_X1 U6452 ( .A1(n5143), .A2(n5142), .A3(n5162), .ZN(n4849) );
  NAND2_X1 U6453 ( .A1(n5174), .A2(n5173), .ZN(n5192) );
  NAND2_X1 U6454 ( .A1(n6285), .A2(n4872), .ZN(n4871) );
  NAND2_X1 U6455 ( .A1(n5326), .A2(n5325), .ZN(n5341) );
  NAND2_X1 U6456 ( .A1(n4885), .A2(n4883), .ZN(n4886) );
  NAND2_X1 U6457 ( .A1(n6290), .A2(n6289), .ZN(n8765) );
  NAND2_X1 U6458 ( .A1(n4887), .A2(n4888), .ZN(n8905) );
  NAND2_X1 U6459 ( .A1(n8189), .A2(n4889), .ZN(n4887) );
  NAND4_X1 U6460 ( .A1(n4965), .A2(n4321), .A3(n6320), .A4(n10152), .ZN(n4896)
         );
  NAND2_X1 U6461 ( .A1(n8832), .A2(n4902), .ZN(n4899) );
  INV_X1 U6462 ( .A(n6927), .ZN(n4904) );
  NAND2_X1 U6463 ( .A1(n4912), .A2(n4911), .ZN(n7990) );
  NAND2_X1 U6464 ( .A1(n8542), .A2(n4301), .ZN(n4921) );
  AOI21_X1 U6465 ( .B1(n8542), .B2(n8543), .A(n6461), .ZN(n8524) );
  NAND2_X1 U6466 ( .A1(n7746), .A2(n4305), .ZN(n7869) );
  INV_X1 U6467 ( .A(n5576), .ZN(n5091) );
  AND2_X4 U6468 ( .A1(n5053), .A2(n5118), .ZN(n5137) );
  NAND2_X1 U6469 ( .A1(n9621), .A2(n9606), .ZN(n4944) );
  AND2_X1 U6470 ( .A1(n4981), .A2(n5641), .ZN(n4947) );
  NAND2_X1 U6471 ( .A1(n9773), .A2(n4952), .ZN(n4950) );
  NAND2_X1 U6472 ( .A1(n5643), .A2(n4323), .ZN(n4953) );
  NAND2_X1 U6473 ( .A1(n5668), .A2(n4959), .ZN(n4958) );
  OAI21_X1 U6474 ( .B1(n5668), .B2(n5537), .A(n4959), .ZN(n6377) );
  NAND2_X1 U6475 ( .A1(n6238), .A2(n6237), .ZN(n6240) );
  OAI21_X1 U6476 ( .B1(n6796), .B2(n8301), .A(n6795), .ZN(n6834) );
  INV_X1 U6477 ( .A(n6815), .ZN(n6793) );
  XNOR2_X1 U6478 ( .A(n5523), .B(n5522), .ZN(n9094) );
  NAND2_X1 U6479 ( .A1(n7232), .A2(n7231), .ZN(n9186) );
  OR2_X1 U6480 ( .A1(n5625), .A2(n5618), .ZN(n5627) );
  NAND2_X1 U6481 ( .A1(n5625), .A2(n5618), .ZN(n5626) );
  OR2_X1 U6482 ( .A1(n5578), .A2(n7718), .ZN(n5003) );
  MUX2_X1 U6483 ( .A(n6680), .B(n6679), .S(n9567), .Z(n6682) );
  MUX2_X1 U6484 ( .A(n6826), .B(n6680), .S(n9567), .Z(n6678) );
  INV_X1 U6485 ( .A(n7016), .ZN(n6294) );
  INV_X1 U6486 ( .A(n7019), .ZN(n7022) );
  INV_X1 U6487 ( .A(n5058), .ZN(n5059) );
  NAND2_X1 U6488 ( .A1(n7318), .A2(n7073), .ZN(n5058) );
  NAND2_X1 U6489 ( .A1(n7079), .A2(n7078), .ZN(n7080) );
  NAND2_X1 U6490 ( .A1(n6528), .A2(n9764), .ZN(n8395) );
  NAND2_X1 U6491 ( .A1(n6958), .A2(n6988), .ZN(n6959) );
  OR2_X1 U6492 ( .A1(n4289), .A2(n4594), .ZN(n5041) );
  NAND2_X1 U6493 ( .A1(n9372), .A2(n10057), .ZN(n6703) );
  NAND2_X1 U6494 ( .A1(n8823), .A2(n6280), .ZN(n6282) );
  NAND2_X1 U6495 ( .A1(n6508), .A2(n6507), .ZN(P2_U3154) );
  INV_X1 U6496 ( .A(n6322), .ZN(n7361) );
  NAND2_X1 U6497 ( .A1(n6373), .A2(n5556), .ZN(n5587) );
  AND2_X1 U6498 ( .A1(n7990), .A2(n7989), .ZN(n10074) );
  NAND2_X1 U6499 ( .A1(n6145), .A2(n5397), .ZN(n5412) );
  NAND2_X2 U6501 ( .A1(n6272), .A2(n6271), .ZN(n8861) );
  CLKBUF_X1 U6502 ( .A(n9773), .Z(n9775) );
  OR2_X1 U6503 ( .A1(n6277), .A2(n6451), .ZN(n6927) );
  AND2_X1 U6504 ( .A1(n6316), .A2(n6309), .ZN(n6480) );
  XNOR2_X1 U6505 ( .A(n7021), .B(n7016), .ZN(n8385) );
  OAI21_X1 U6506 ( .B1(n5430), .B2(n5422), .A(n5423), .ZN(n5408) );
  XNOR2_X1 U6507 ( .A(n5430), .B(n5396), .ZN(n8186) );
  OR2_X1 U6508 ( .A1(n4295), .A2(n9983), .ZN(n4998) );
  AND2_X1 U6509 ( .A1(n7342), .A2(P2_U3151), .ZN(n9091) );
  OAI211_X1 U6510 ( .C1(n4292), .C2(P1_DATAO_REG_2__SCAN_IN), .A(n5073), .B(
        SI_2_), .ZN(n5079) );
  OAI21_X1 U6511 ( .B1(n5072), .B2(n4292), .A(n5071), .ZN(n5095) );
  NAND2_X1 U6512 ( .A1(n4285), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5071) );
  XNOR2_X1 U6513 ( .A(n5671), .B(n6786), .ZN(n5682) );
  AND2_X1 U6514 ( .A1(n7315), .A2(n7314), .ZN(n4963) );
  AND2_X1 U6515 ( .A1(n7316), .A2(n4963), .ZN(n4964) );
  OR2_X1 U6516 ( .A1(n8385), .A2(n8059), .ZN(n4965) );
  AND2_X1 U6517 ( .A1(n7313), .A2(n8874), .ZN(n10107) );
  NAND2_X1 U6518 ( .A1(n10166), .A2(n10151), .ZN(n8961) );
  AND3_X2 U6519 ( .A1(n7306), .A2(n6362), .A3(n7304), .ZN(n10166) );
  INV_X1 U6520 ( .A(n7679), .ZN(n5771) );
  AND2_X1 U6521 ( .A1(n6354), .A2(n8342), .ZN(n10141) );
  INV_X1 U6522 ( .A(n10073), .ZN(n7060) );
  INV_X1 U6523 ( .A(n9902), .ZN(n6366) );
  NAND2_X1 U6524 ( .A1(n7331), .A2(n9780), .ZN(n7937) );
  AND2_X1 U6525 ( .A1(n5137), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n4966) );
  AND2_X1 U6526 ( .A1(n5913), .A2(n5912), .ZN(n4967) );
  AND2_X1 U6527 ( .A1(n7031), .A2(n7030), .ZN(n4968) );
  NOR2_X1 U6528 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4969) );
  OR2_X1 U6529 ( .A1(n9578), .A2(n9978), .ZN(n4970) );
  AND2_X1 U6530 ( .A1(n6364), .A2(n6363), .ZN(n4971) );
  AND3_X1 U6531 ( .A1(n5720), .A2(n5719), .A3(n5746), .ZN(n4973) );
  AND4_X1 U6532 ( .A1(n5723), .A2(n5722), .A3(n5739), .A4(n5721), .ZN(n4974)
         );
  AND3_X1 U6533 ( .A1(n7228), .A2(n7213), .A3(n7221), .ZN(n4975) );
  AND2_X1 U6534 ( .A1(n5137), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6535 ( .A1(n6301), .A2(n6300), .ZN(n10096) );
  AND2_X1 U6536 ( .A1(n5209), .A2(n5195), .ZN(n4977) );
  AND2_X1 U6537 ( .A1(n8452), .A2(n8109), .ZN(n4978) );
  INV_X1 U6538 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5072) );
  INV_X1 U6539 ( .A(n9584), .ZN(n5918) );
  INV_X1 U6540 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5924) );
  AND2_X1 U6541 ( .A1(n6827), .A2(n6826), .ZN(n4979) );
  NAND2_X1 U6542 ( .A1(n7064), .A2(n6539), .ZN(n7068) );
  AND4_X1 U6543 ( .A1(n5711), .A2(n5710), .A3(n5709), .A4(n5708), .ZN(n4980)
         );
  OR2_X1 U6544 ( .A1(n5642), .A2(n8172), .ZN(n4981) );
  AND3_X1 U6545 ( .A1(n7004), .A2(n7968), .A3(n8050), .ZN(n4982) );
  AND4_X1 U6546 ( .A1(n6790), .A2(n6789), .A3(n6788), .A4(n6787), .ZN(n4983)
         );
  AND2_X1 U6547 ( .A1(n4970), .A2(n6382), .ZN(n4984) );
  INV_X1 U6548 ( .A(n10070), .ZN(n6383) );
  NAND2_X1 U6549 ( .A1(n6943), .A2(n6988), .ZN(n6944) );
  NOR4_X1 U6551 ( .A1(n7016), .A2(n8758), .A3(n8766), .A4(n7015), .ZN(n7018)
         );
  NOR2_X1 U6552 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5695) );
  OR2_X1 U6553 ( .A1(n9007), .A2(n8803), .ZN(n6287) );
  INV_X1 U6554 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5709) );
  NOR2_X1 U6555 ( .A1(n6786), .A2(n6785), .ZN(n6790) );
  INV_X1 U6556 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n4992) );
  INV_X1 U6557 ( .A(n7786), .ZN(n6003) );
  INV_X1 U6558 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n4994) );
  INV_X1 U6559 ( .A(n7872), .ZN(n6410) );
  OAI21_X1 U6560 ( .B1(n8983), .B2(n7024), .A(n7023), .ZN(n7025) );
  INV_X1 U6561 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n5786) );
  NOR2_X1 U6562 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  INV_X1 U6563 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U6564 ( .A1(n4973), .A2(n4974), .ZN(n5724) );
  BUF_X4 U6565 ( .A(n8398), .Z(n7246) );
  OR2_X1 U6566 ( .A1(n7235), .A2(n7234), .ZN(n7236) );
  INV_X1 U6567 ( .A(SI_9_), .ZN(n10301) );
  INV_X1 U6568 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10256) );
  INV_X1 U6569 ( .A(n7845), .ZN(n5683) );
  INV_X1 U6570 ( .A(SI_27_), .ZN(n5525) );
  INV_X1 U6571 ( .A(SI_24_), .ZN(n5468) );
  INV_X1 U6572 ( .A(SI_22_), .ZN(n5431) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5119) );
  INV_X1 U6574 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5733) );
  INV_X1 U6575 ( .A(n8767), .ZN(n6469) );
  OR2_X1 U6576 ( .A1(n7777), .A2(n5779), .ZN(n5780) );
  AND2_X1 U6577 ( .A1(n7028), .A2(n7036), .ZN(n6342) );
  INV_X1 U6578 ( .A(n8850), .ZN(n6451) );
  INV_X1 U6579 ( .A(n6480), .ZN(n6483) );
  AND2_X1 U6580 ( .A1(n5622), .A2(n5621), .ZN(n5623) );
  XNOR2_X1 U6581 ( .A(n7216), .B(n7270), .ZN(n7235) );
  NAND2_X1 U6582 ( .A1(n5455), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5474) );
  NAND2_X1 U6583 ( .A1(n5491), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U6584 ( .A1(n5276), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5291) );
  NOR2_X2 U6585 ( .A1(n9644), .A2(n9920), .ZN(n9628) );
  NAND2_X1 U6586 ( .A1(n5526), .A2(n5525), .ZN(n5563) );
  INV_X1 U6587 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5596) );
  INV_X1 U6588 ( .A(n8825), .ZN(n8496) );
  INV_X1 U6589 ( .A(n10129), .ZN(n7725) );
  INV_X1 U6590 ( .A(n8595), .ZN(n8583) );
  OR2_X1 U6591 ( .A1(P2_U3150), .A2(n5905), .ZN(n7953) );
  OR2_X1 U6592 ( .A1(n6359), .A2(n6358), .ZN(n6360) );
  OR2_X1 U6593 ( .A1(n10135), .A2(n7310), .ZN(n6478) );
  INV_X1 U6594 ( .A(n6950), .ZN(n8794) );
  INV_X1 U6595 ( .A(n6045), .ZN(n6046) );
  INV_X1 U6596 ( .A(n10096), .ZN(n8894) );
  NAND2_X1 U6597 ( .A1(n6243), .A2(n6496), .ZN(n8059) );
  INV_X1 U6598 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6237) );
  INV_X1 U6599 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9270) );
  OR2_X1 U6600 ( .A1(n6828), .A2(n4979), .ZN(n6829) );
  INV_X1 U6601 ( .A(n4291), .ZN(n5531) );
  INV_X1 U6602 ( .A(n5674), .ZN(n9386) );
  INV_X1 U6603 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9304) );
  OR2_X1 U6604 ( .A1(n10006), .A2(n9386), .ZN(n10043) );
  INV_X1 U6605 ( .A(n9363), .ZN(n9338) );
  INV_X1 U6606 ( .A(n7284), .ZN(n7285) );
  INV_X1 U6607 ( .A(n8419), .ZN(n9578) );
  INV_X1 U6608 ( .A(n9978), .ZN(n5687) );
  INV_X1 U6609 ( .A(n5650), .ZN(n8071) );
  NAND2_X1 U6610 ( .A1(n9797), .A2(n7063), .ZN(n7284) );
  AND2_X1 U6611 ( .A1(n6500), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7430) );
  INV_X1 U6612 ( .A(n7953), .ZN(n8736) );
  AND2_X1 U6613 ( .A1(n7973), .A2(n8051), .ZN(n7982) );
  AND2_X1 U6614 ( .A1(n10078), .A2(n10077), .ZN(n10142) );
  INV_X1 U6615 ( .A(n8896), .ZN(n10091) );
  INV_X1 U6616 ( .A(n8901), .ZN(n10101) );
  INV_X1 U6617 ( .A(n8961), .ZN(n8967) );
  NAND2_X1 U6618 ( .A1(n6361), .A2(n6360), .ZN(n7304) );
  INV_X1 U6619 ( .A(n9055), .ZN(n9066) );
  INV_X1 U6620 ( .A(n10146), .ZN(n10139) );
  OR2_X1 U6621 ( .A1(n6477), .A2(n6346), .ZN(n6347) );
  INV_X1 U6622 ( .A(n6323), .ZN(n7366) );
  INV_X1 U6623 ( .A(n9326), .ZN(n9339) );
  NAND2_X1 U6624 ( .A1(n7294), .A2(n7293), .ZN(n9328) );
  NAND2_X1 U6625 ( .A1(n6821), .A2(n6819), .ZN(n6822) );
  OR2_X1 U6626 ( .A1(n9614), .A2(n4290), .ZN(n5500) );
  AND4_X1 U6627 ( .A1(n5336), .A2(n5335), .A3(n5334), .A4(n5333), .ZN(n9335)
         );
  OR2_X1 U6628 ( .A1(n10006), .A2(n7572), .ZN(n10022) );
  INV_X1 U6629 ( .A(n10034), .ZN(n9501) );
  INV_X1 U6630 ( .A(n10022), .ZN(n10037) );
  INV_X1 U6631 ( .A(n9784), .ZN(n9764) );
  AND2_X1 U6632 ( .A1(n6541), .A2(n6543), .ZN(n9607) );
  INV_X1 U6633 ( .A(n9793), .ZN(n10333) );
  INV_X1 U6634 ( .A(n10341), .ZN(n9788) );
  INV_X1 U6635 ( .A(n5919), .ZN(n7328) );
  INV_X1 U6636 ( .A(n9872), .ZN(n9858) );
  NAND2_X1 U6637 ( .A1(n8264), .A2(n10067), .ZN(n10061) );
  MUX2_X1 U6638 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5632), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5633) );
  INV_X1 U6639 ( .A(n7430), .ZN(n7364) );
  INV_X1 U6640 ( .A(n8599), .ZN(n8560) );
  INV_X1 U6641 ( .A(n8591), .ZN(n8588) );
  INV_X1 U6642 ( .A(P2_U3893), .ZN(n8614) );
  INV_X1 U6643 ( .A(n8701), .ZN(n8734) );
  INV_X1 U6644 ( .A(n8723), .ZN(n8748) );
  INV_X1 U6645 ( .A(n7982), .ZN(n8979) );
  AND3_X1 U6646 ( .A1(n10085), .A2(n10084), .A3(n10083), .ZN(n10144) );
  OR2_X1 U6647 ( .A1(n10107), .A2(n7311), .ZN(n8917) );
  NAND2_X1 U6648 ( .A1(n10166), .A2(n10139), .ZN(n8975) );
  INV_X1 U6649 ( .A(n10166), .ZN(n10164) );
  OR2_X1 U6650 ( .A1(n10154), .A2(n10135), .ZN(n9055) );
  AND2_X1 U6651 ( .A1(n10144), .A2(n10143), .ZN(n10163) );
  AND2_X1 U6652 ( .A1(n6348), .A2(n6347), .ZN(n10154) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U6654 ( .A1(n5793), .A2(n5791), .ZN(n8663) );
  INV_X1 U6655 ( .A(n9328), .ZN(n9341) );
  AND2_X1 U6656 ( .A1(n7286), .A2(n9780), .ZN(n9331) );
  INV_X1 U6657 ( .A(n9119), .ZN(n9353) );
  INV_X1 U6658 ( .A(n7153), .ZN(n9367) );
  INV_X1 U6659 ( .A(n7143), .ZN(n9368) );
  INV_X1 U6660 ( .A(n7073), .ZN(n9375) );
  INV_X1 U6661 ( .A(n10004), .ZN(n10050) );
  INV_X1 U6662 ( .A(n7937), .ZN(n9712) );
  NAND2_X1 U6663 ( .A1(n7937), .A2(n7936), .ZN(n9793) );
  INV_X1 U6664 ( .A(n7058), .ZN(n7059) );
  NAND2_X1 U6665 ( .A1(n10073), .A2(n10061), .ZN(n9872) );
  AND2_X1 U6666 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NAND2_X1 U6667 ( .A1(n10070), .A2(n10061), .ZN(n9963) );
  NOR2_X1 U6668 ( .A1(n7427), .A2(n7445), .ZN(n10051) );
  INV_X1 U6669 ( .A(n7064), .ZN(n8340) );
  INV_X1 U6670 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8389) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7423) );
  NOR2_X1 U6672 ( .A1(n8129), .A2(n8128), .ZN(n10352) );
  NOR2_X1 U6673 ( .A1(n8135), .A2(n8134), .ZN(n10185) );
  NOR2_X2 U6674 ( .A1(n6492), .A2(n7364), .ZN(P2_U3893) );
  NAND2_X1 U6675 ( .A1(n5914), .A2(n4967), .ZN(P2_U3201) );
  NOR2_X1 U6676 ( .A1(n7067), .A2(n7710), .ZN(P1_U3973) );
  NOR3_X1 U6677 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n4991) );
  NOR2_X2 U6678 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5593) );
  NOR2_X1 U6679 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4989) );
  NAND3_X1 U6680 ( .A1(n4992), .A2(n10207), .A3(n5590), .ZN(n4993) );
  NAND2_X1 U6681 ( .A1(n4295), .A2(n4997), .ZN(n9982) );
  XNOR2_X2 U6682 ( .A(n4998), .B(n4997), .ZN(n4999) );
  AND2_X2 U6683 ( .A1(n5000), .A2(n4999), .ZN(n5063) );
  NAND2_X1 U6684 ( .A1(n5063), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5006) );
  INV_X1 U6685 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10001) );
  NAND2_X4 U6686 ( .A1(n9987), .A2(n4999), .ZN(n6534) );
  INV_X1 U6687 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5001) );
  INV_X1 U6688 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7718) );
  NAND3_X1 U6689 ( .A1(n5007), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U6690 ( .A1(n4292), .A2(SI_0_), .ZN(n5010) );
  XNOR2_X1 U6691 ( .A(n5010), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9999) );
  XNOR2_X2 U6692 ( .A(n5013), .B(n5012), .ZN(n5674) );
  MUX2_X1 U6693 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9999), .S(n5053), .Z(n7836) );
  NAND2_X1 U6694 ( .A1(n6693), .A2(n7836), .ZN(n7318) );
  INV_X1 U6695 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7333) );
  NAND2_X1 U6696 ( .A1(n5063), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5019) );
  INV_X1 U6697 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5015) );
  OR2_X1 U6698 ( .A1(n5065), .A2(n5015), .ZN(n5018) );
  INV_X1 U6699 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5016) );
  AND4_X4 U6700 ( .A1(n5020), .A2(n5019), .A3(n5018), .A4(n5017), .ZN(n7073)
         );
  NAND2_X1 U6701 ( .A1(n5063), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5025) );
  INV_X1 U6702 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9393) );
  INV_X1 U6703 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5021) );
  OR2_X1 U6704 ( .A1(n6530), .A2(n5021), .ZN(n5022) );
  NAND2_X1 U6705 ( .A1(n5058), .A2(n9374), .ZN(n5044) );
  NAND2_X1 U6706 ( .A1(n5137), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6707 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5048) );
  INV_X1 U6708 ( .A(SI_1_), .ZN(n5049) );
  NAND2_X1 U6709 ( .A1(n5048), .A2(n5049), .ZN(n5026) );
  NAND2_X1 U6710 ( .A1(n5026), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5029) );
  INV_X1 U6711 ( .A(n5048), .ZN(n5027) );
  NAND2_X1 U6712 ( .A1(n5027), .A2(SI_1_), .ZN(n5028) );
  NAND2_X1 U6713 ( .A1(n5029), .A2(n5028), .ZN(n5030) );
  NAND2_X1 U6714 ( .A1(n4292), .A2(n5030), .ZN(n5035) );
  INV_X1 U6715 ( .A(n4286), .ZN(n5047) );
  NOR2_X1 U6716 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6717 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6718 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5031) );
  OAI21_X1 U6719 ( .B1(n5032), .B2(n5045), .A(n5031), .ZN(n5033) );
  NAND2_X1 U6720 ( .A1(n5047), .A2(n5033), .ZN(n5034) );
  NAND2_X1 U6721 ( .A1(n5035), .A2(n5034), .ZN(n5076) );
  XNOR2_X1 U6722 ( .A(n5076), .B(SI_2_), .ZN(n5037) );
  MUX2_X1 U6723 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4292), .Z(n5036) );
  XNOR2_X1 U6724 ( .A(n5037), .B(n5036), .ZN(n5953) );
  NAND2_X1 U6725 ( .A1(n5576), .A2(n5953), .ZN(n5042) );
  INV_X1 U6726 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9983) );
  INV_X1 U6727 ( .A(n5039), .ZN(n5040) );
  AND3_X2 U6728 ( .A1(n5043), .A2(n5042), .A3(n5041), .ZN(n8172) );
  NAND2_X1 U6729 ( .A1(n5044), .A2(n8172), .ZN(n5062) );
  INV_X1 U6730 ( .A(n8172), .ZN(n7813) );
  INV_X1 U6731 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6732 ( .A1(n5118), .A2(n5046), .ZN(n5943) );
  OAI21_X1 U6733 ( .B1(n5048), .B2(n5118), .A(n5943), .ZN(n5050) );
  XNOR2_X1 U6734 ( .A(n5050), .B(n5049), .ZN(n5052) );
  MUX2_X1 U6735 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(P1_DATAO_REG_1__SCAN_IN), 
        .S(n5118), .Z(n5051) );
  XNOR2_X1 U6736 ( .A(n5052), .B(n5051), .ZN(n7355) );
  NAND2_X1 U6737 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5054) );
  MUX2_X1 U6738 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5054), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5056) );
  INV_X1 U6739 ( .A(n5038), .ZN(n5055) );
  NAND2_X1 U6740 ( .A1(n5056), .A2(n5055), .ZN(n7557) );
  INV_X1 U6741 ( .A(n7557), .ZN(n9381) );
  AOI21_X1 U6742 ( .B1(n5642), .B2(n7813), .A(n4293), .ZN(n5057) );
  OAI21_X1 U6743 ( .B1(n7318), .B2(n7073), .A(n5057), .ZN(n5061) );
  NAND2_X1 U6744 ( .A1(n5059), .A2(n7084), .ZN(n5060) );
  NAND3_X1 U6745 ( .A1(n5062), .A2(n5061), .A3(n5060), .ZN(n7850) );
  OR2_X1 U6746 ( .A1(n4291), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5070) );
  INV_X2 U6747 ( .A(n5063), .ZN(n5583) );
  INV_X1 U6748 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U6749 ( .A1(n5153), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5068) );
  INV_X1 U6750 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5066) );
  XNOR2_X1 U6751 ( .A(n5095), .B(SI_3_), .ZN(n5092) );
  INV_X1 U6752 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7350) );
  NAND2_X1 U6753 ( .A1(n4292), .A2(n7350), .ZN(n5073) );
  INV_X1 U6754 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U6755 ( .A1(n4286), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5075) );
  INV_X1 U6756 ( .A(SI_2_), .ZN(n5074) );
  OAI211_X1 U6757 ( .C1(n4286), .C2(n7356), .A(n5075), .B(n5074), .ZN(n5077)
         );
  NAND2_X1 U6758 ( .A1(n5077), .A2(n5076), .ZN(n5078) );
  NAND2_X1 U6759 ( .A1(n5079), .A2(n5078), .ZN(n5093) );
  XNOR2_X1 U6760 ( .A(n5092), .B(n5093), .ZN(n5964) );
  NAND2_X1 U6761 ( .A1(n5576), .A2(n5964), .ZN(n5083) );
  NAND2_X1 U6762 ( .A1(n5137), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6763 ( .A1(n5039), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6764 ( .A(n5080), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9409) );
  OR2_X2 U6765 ( .A1(n5084), .A2(n7862), .ZN(n7817) );
  NAND2_X1 U6766 ( .A1(n5084), .A2(n7862), .ZN(n6696) );
  NAND2_X1 U6767 ( .A1(n7817), .A2(n6696), .ZN(n7849) );
  NAND2_X1 U6768 ( .A1(n7850), .A2(n7849), .ZN(n7848) );
  INV_X1 U6769 ( .A(n5084), .ZN(n7812) );
  NAND2_X1 U6770 ( .A1(n7812), .A2(n7862), .ZN(n5085) );
  NAND2_X1 U6771 ( .A1(n5579), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5090) );
  INV_X1 U6772 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5086) );
  OR2_X1 U6773 ( .A1(n5583), .A2(n5086), .ZN(n5089) );
  INV_X1 U6774 ( .A(n5104), .ZN(n5105) );
  OAI21_X1 U6775 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n5105), .ZN(n8041) );
  OR2_X1 U6776 ( .A1(n4291), .A2(n8041), .ZN(n5088) );
  NAND2_X1 U6777 ( .A1(n5153), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5087) );
  INV_X1 U6778 ( .A(n5092), .ZN(n5094) );
  NAND2_X1 U6779 ( .A1(n5094), .A2(n5093), .ZN(n5097) );
  NAND2_X1 U6780 ( .A1(n5095), .A2(SI_3_), .ZN(n5096) );
  NAND2_X1 U6781 ( .A1(n5097), .A2(n5096), .ZN(n5112) );
  INV_X1 U6782 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7349) );
  INV_X1 U6783 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7352) );
  MUX2_X1 U6784 ( .A(n7349), .B(n7352), .S(n4292), .Z(n5113) );
  XNOR2_X1 U6785 ( .A(n5113), .B(SI_4_), .ZN(n5111) );
  INV_X1 U6786 ( .A(n5111), .ZN(n5098) );
  XNOR2_X1 U6787 ( .A(n5112), .B(n5098), .ZN(n7347) );
  NAND2_X1 U6788 ( .A1(n5576), .A2(n7347), .ZN(n5102) );
  NAND2_X1 U6789 ( .A1(n5137), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5101) );
  NAND2_X1 U6790 ( .A1(n5099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5121) );
  XNOR2_X1 U6791 ( .A(n5121), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U6792 ( .A1(n7441), .A2(n9422), .ZN(n5100) );
  OR2_X2 U6793 ( .A1(n9373), .A2(n7854), .ZN(n6568) );
  NAND2_X1 U6794 ( .A1(n9373), .A2(n7854), .ZN(n6700) );
  NAND2_X1 U6795 ( .A1(n5579), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5110) );
  INV_X1 U6796 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5103) );
  OR2_X1 U6797 ( .A1(n5583), .A2(n5103), .ZN(n5109) );
  NAND2_X1 U6798 ( .A1(n5104), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5130) );
  INV_X1 U6799 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U6800 ( .A1(n5105), .A2(n8203), .ZN(n5106) );
  NAND2_X1 U6801 ( .A1(n5130), .A2(n5106), .ZN(n8209) );
  OR2_X1 U6802 ( .A1(n4291), .A2(n8209), .ZN(n5108) );
  INV_X1 U6803 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7549) );
  OR2_X1 U6804 ( .A1(n6534), .A2(n7549), .ZN(n5107) );
  NAND2_X1 U6805 ( .A1(n5112), .A2(n5111), .ZN(n5116) );
  INV_X1 U6806 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6807 ( .A1(n5114), .A2(SI_4_), .ZN(n5115) );
  INV_X1 U6808 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5117) );
  OAI21_X1 U6809 ( .B1(n4286), .B2(n5119), .A(n4330), .ZN(n5144) );
  XNOR2_X1 U6810 ( .A(n5144), .B(SI_5_), .ZN(n5141) );
  XNOR2_X1 U6811 ( .A(n5143), .B(n5141), .ZN(n7358) );
  NAND2_X1 U6812 ( .A1(n5576), .A2(n7358), .ZN(n5126) );
  NAND2_X1 U6813 ( .A1(n5137), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6814 ( .A1(n5121), .A2(n5120), .ZN(n5122) );
  NAND2_X1 U6815 ( .A1(n5122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5123) );
  XNOR2_X1 U6816 ( .A(n5123), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U6817 ( .A1(n7441), .A2(n9436), .ZN(n5124) );
  OR2_X2 U6818 ( .A1(n9372), .A2(n10057), .ZN(n6569) );
  NAND2_X1 U6819 ( .A1(n5579), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5136) );
  NAND2_X1 U6820 ( .A1(n5153), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5135) );
  INV_X1 U6821 ( .A(n5130), .ZN(n5128) );
  NAND2_X1 U6822 ( .A1(n5128), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5154) );
  INV_X1 U6823 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6824 ( .A1(n5130), .A2(n5129), .ZN(n5131) );
  NAND2_X1 U6825 ( .A1(n5154), .A2(n5131), .ZN(n8229) );
  OR2_X1 U6826 ( .A1(n4290), .A2(n8229), .ZN(n5134) );
  INV_X1 U6827 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5132) );
  OR2_X1 U6828 ( .A1(n5583), .A2(n5132), .ZN(n5133) );
  OR2_X1 U6829 ( .A1(n5139), .A2(n9983), .ZN(n5140) );
  XNOR2_X1 U6830 ( .A(n5140), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9449) );
  AOI22_X1 U6831 ( .A1(n5137), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n7441), .B2(
        n9449), .ZN(n5147) );
  INV_X1 U6832 ( .A(n5141), .ZN(n5142) );
  NAND2_X1 U6833 ( .A1(n5144), .A2(SI_5_), .ZN(n5145) );
  MUX2_X1 U6834 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4286), .Z(n5164) );
  XNOR2_X1 U6835 ( .A(n5164), .B(SI_6_), .ZN(n5161) );
  XNOR2_X1 U6836 ( .A(n5163), .B(n5161), .ZN(n7369) );
  NAND2_X1 U6837 ( .A1(n7369), .A2(n5397), .ZN(n5146) );
  NAND2_X1 U6838 ( .A1(n9371), .A2(n8235), .ZN(n8155) );
  NAND2_X1 U6839 ( .A1(n8154), .A2(n8155), .ZN(n7896) );
  NOR2_X1 U6840 ( .A1(n9373), .A2(n8044), .ZN(n7931) );
  NAND2_X1 U6841 ( .A1(n6761), .A2(n7931), .ZN(n5149) );
  INV_X1 U6842 ( .A(n9372), .ZN(n7111) );
  NAND2_X1 U6843 ( .A1(n7111), .A2(n10057), .ZN(n5148) );
  NAND2_X1 U6844 ( .A1(n5149), .A2(n5148), .ZN(n7892) );
  NOR2_X1 U6845 ( .A1(n9371), .A2(n8219), .ZN(n5150) );
  NAND2_X1 U6846 ( .A1(n5152), .A2(n5151), .ZN(n8239) );
  NAND2_X1 U6847 ( .A1(n5153), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U6848 ( .A1(n5579), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5159) );
  OR2_X2 U6849 ( .A1(n5154), .A2(n8329), .ZN(n5202) );
  NAND2_X1 U6850 ( .A1(n5154), .A2(n8329), .ZN(n5155) );
  NAND2_X1 U6851 ( .A1(n5202), .A2(n5155), .ZN(n8331) );
  OR2_X1 U6852 ( .A1(n4291), .A2(n8331), .ZN(n5158) );
  INV_X1 U6853 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5156) );
  OR2_X1 U6854 ( .A1(n5583), .A2(n5156), .ZN(n5157) );
  NAND4_X1 U6855 ( .A1(n5160), .A2(n5159), .A3(n5158), .A4(n5157), .ZN(n9370)
         );
  INV_X1 U6856 ( .A(n5161), .ZN(n5162) );
  MUX2_X1 U6857 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4286), .Z(n5172) );
  XNOR2_X1 U6858 ( .A(n5172), .B(SI_7_), .ZN(n5169) );
  NAND2_X1 U6859 ( .A1(n7373), .A2(n5397), .ZN(n5168) );
  INV_X1 U6860 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6861 ( .A1(n5139), .A2(n5165), .ZN(n5179) );
  NAND2_X1 U6862 ( .A1(n5179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6863 ( .A(n5166), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9462) );
  AOI22_X1 U6864 ( .A1(n5137), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n7441), .B2(
        n9462), .ZN(n5167) );
  NAND2_X1 U6865 ( .A1(n8249), .A2(n9370), .ZN(n6576) );
  INV_X1 U6866 ( .A(n5169), .ZN(n5170) );
  NAND2_X1 U6867 ( .A1(n5172), .A2(SI_7_), .ZN(n5173) );
  MUX2_X1 U6868 ( .A(n7380), .B(n10190), .S(n4292), .Z(n5176) );
  INV_X1 U6869 ( .A(SI_8_), .ZN(n5175) );
  INV_X1 U6870 ( .A(n5176), .ZN(n5177) );
  NAND2_X1 U6871 ( .A1(n5177), .A2(SI_8_), .ZN(n5178) );
  NAND2_X1 U6872 ( .A1(n7378), .A2(n5397), .ZN(n5181) );
  NAND2_X1 U6873 ( .A1(n5213), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5196) );
  XNOR2_X1 U6874 ( .A(n5196), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9475) );
  AOI22_X1 U6875 ( .A1(n5137), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n7441), .B2(
        n9475), .ZN(n5180) );
  NAND2_X1 U6876 ( .A1(n5579), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5185) );
  INV_X1 U6877 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9976) );
  OR2_X1 U6878 ( .A1(n5583), .A2(n9976), .ZN(n5184) );
  INV_X1 U6879 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9169) );
  XNOR2_X1 U6880 ( .A(n5202), .B(n9169), .ZN(n9175) );
  OR2_X1 U6881 ( .A1(n4290), .A2(n9175), .ZN(n5183) );
  INV_X1 U6882 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8265) );
  OR2_X1 U6883 ( .A1(n6534), .A2(n8265), .ZN(n5182) );
  OR2_X1 U6884 ( .A1(n9172), .A2(n7134), .ZN(n6577) );
  NAND2_X1 U6885 ( .A1(n9172), .A2(n7134), .ZN(n8158) );
  INV_X1 U6886 ( .A(n8258), .ZN(n5186) );
  NOR2_X1 U6887 ( .A1(n9370), .A2(n10063), .ZN(n8253) );
  NAND2_X1 U6888 ( .A1(n5186), .A2(n8253), .ZN(n5188) );
  MUX2_X1 U6889 ( .A(n10289), .B(n7394), .S(n4292), .Z(n5193) );
  NAND2_X1 U6890 ( .A1(n5193), .A2(n10301), .ZN(n5209) );
  INV_X1 U6891 ( .A(n5193), .ZN(n5194) );
  NAND2_X1 U6892 ( .A1(n5194), .A2(SI_9_), .ZN(n5195) );
  INV_X1 U6893 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6894 ( .A1(n5196), .A2(n5211), .ZN(n5197) );
  NAND2_X1 U6895 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6896 ( .A(n5198), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7556) );
  AOI22_X1 U6897 ( .A1(n5137), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n7441), .B2(
        n7556), .ZN(n5199) );
  NAND2_X1 U6898 ( .A1(n5063), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5207) );
  INV_X1 U6899 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n8164) );
  OR2_X1 U6900 ( .A1(n6534), .A2(n8164), .ZN(n5206) );
  INV_X1 U6901 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9893) );
  OR2_X1 U6902 ( .A1(n6530), .A2(n9893), .ZN(n5205) );
  INV_X1 U6903 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5201) );
  OAI21_X1 U6904 ( .B1(n5202), .B2(n9169), .A(n5201), .ZN(n5203) );
  NAND2_X1 U6905 ( .A1(n5203), .A2(n5222), .ZN(n9262) );
  OR2_X1 U6906 ( .A1(n4290), .A2(n9262), .ZN(n5204) );
  NAND2_X1 U6907 ( .A1(n6587), .A2(n6592), .ZN(n8159) );
  OR2_X1 U6908 ( .A1(n4435), .A2(n9368), .ZN(n5208) );
  MUX2_X1 U6909 ( .A(n10261), .B(n7397), .S(n4292), .Z(n5230) );
  XNOR2_X1 U6910 ( .A(n5230), .B(SI_10_), .ZN(n5229) );
  XNOR2_X1 U6911 ( .A(n5233), .B(n5229), .ZN(n7396) );
  NAND2_X1 U6912 ( .A1(n7396), .A2(n5397), .ZN(n5219) );
  INV_X1 U6913 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6914 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6915 ( .A1(n5216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5214) );
  MUX2_X1 U6916 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5214), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5215) );
  INV_X1 U6917 ( .A(n5215), .ZN(n5217) );
  NOR2_X1 U6918 ( .A1(n5217), .A2(n5238), .ZN(n9494) );
  AOI22_X1 U6919 ( .A1(n5137), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7441), .B2(
        n9494), .ZN(n5218) );
  NAND2_X1 U6920 ( .A1(n5579), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5227) );
  INV_X1 U6921 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6922 ( .A1(n5583), .A2(n5220), .ZN(n5226) );
  INV_X1 U6923 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U6924 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  NAND2_X1 U6925 ( .A1(n5259), .A2(n5223), .ZN(n9130) );
  OR2_X1 U6926 ( .A1(n4290), .A2(n9130), .ZN(n5225) );
  INV_X1 U6927 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7589) );
  OR2_X1 U6928 ( .A1(n6534), .A2(n7589), .ZN(n5224) );
  OR2_X1 U6929 ( .A1(n9133), .A2(n7153), .ZN(n6710) );
  NAND2_X1 U6930 ( .A1(n9133), .A2(n7153), .ZN(n6594) );
  NAND2_X1 U6931 ( .A1(n6710), .A2(n6594), .ZN(n8000) );
  OR2_X1 U6932 ( .A1(n9133), .A2(n9367), .ZN(n5228) );
  NAND2_X1 U6933 ( .A1(n8003), .A2(n5228), .ZN(n8070) );
  INV_X1 U6934 ( .A(n5230), .ZN(n5231) );
  NAND2_X1 U6935 ( .A1(n5231), .A2(SI_10_), .ZN(n5232) );
  MUX2_X1 U6936 ( .A(n7419), .B(n7421), .S(n4286), .Z(n5235) );
  NAND2_X1 U6937 ( .A1(n5235), .A2(n5234), .ZN(n5249) );
  INV_X1 U6938 ( .A(n5235), .ZN(n5236) );
  NAND2_X1 U6939 ( .A1(n5236), .A2(SI_11_), .ZN(n5237) );
  NAND2_X1 U6940 ( .A1(n5249), .A2(n5237), .ZN(n5250) );
  XNOR2_X1 U6941 ( .A(n5251), .B(n5250), .ZN(n7418) );
  NAND2_X1 U6942 ( .A1(n7418), .A2(n5397), .ZN(n5241) );
  INV_X1 U6943 ( .A(n5238), .ZN(n5252) );
  NAND2_X1 U6944 ( .A1(n5252), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5239) );
  XNOR2_X1 U6945 ( .A(n5239), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9508) );
  AOI22_X1 U6946 ( .A1(n5137), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n7441), .B2(
        n9508), .ZN(n5240) );
  NAND2_X1 U6947 ( .A1(n5153), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5246) );
  INV_X1 U6948 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7598) );
  OR2_X1 U6949 ( .A1(n5065), .A2(n7598), .ZN(n5245) );
  XNOR2_X1 U6950 ( .A(n5259), .B(n9304), .ZN(n9305) );
  OR2_X1 U6951 ( .A1(n4291), .A2(n9305), .ZN(n5244) );
  INV_X1 U6952 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5242) );
  OR2_X1 U6953 ( .A1(n5583), .A2(n5242), .ZN(n5243) );
  OR2_X1 U6954 ( .A1(n9885), .A2(n8288), .ZN(n6596) );
  NAND2_X1 U6955 ( .A1(n9885), .A2(n8288), .ZN(n8283) );
  NAND2_X1 U6956 ( .A1(n6596), .A2(n8283), .ZN(n5650) );
  NAND2_X1 U6957 ( .A1(n8070), .A2(n5650), .ZN(n5248) );
  INV_X1 U6958 ( .A(n8288), .ZN(n9366) );
  OR2_X1 U6959 ( .A1(n9885), .A2(n9366), .ZN(n5247) );
  NAND2_X1 U6960 ( .A1(n5248), .A2(n5247), .ZN(n8282) );
  MUX2_X1 U6961 ( .A(n7426), .B(n7423), .S(n4286), .Z(n5267) );
  XNOR2_X1 U6962 ( .A(n5267), .B(SI_12_), .ZN(n5266) );
  XNOR2_X1 U6963 ( .A(n5271), .B(n5266), .ZN(n7422) );
  NAND2_X1 U6964 ( .A1(n7422), .A2(n5397), .ZN(n5258) );
  NAND2_X1 U6965 ( .A1(n5253), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5255) );
  INV_X1 U6966 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U6967 ( .A1(n5255), .A2(n5254), .ZN(n5272) );
  OR2_X1 U6968 ( .A1(n5255), .A2(n5254), .ZN(n5256) );
  AOI22_X1 U6969 ( .A1(n5137), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n7441), .B2(
        n7592), .ZN(n5257) );
  NAND2_X1 U6970 ( .A1(n5063), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5264) );
  INV_X1 U6971 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8294) );
  OR2_X1 U6972 ( .A1(n6534), .A2(n8294), .ZN(n5263) );
  INV_X1 U6973 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10196) );
  OR2_X1 U6974 ( .A1(n5065), .A2(n10196), .ZN(n5262) );
  OAI21_X1 U6975 ( .B1(n5259), .B2(n9304), .A(n7602), .ZN(n5260) );
  OR3_X2 U6976 ( .A1(n5259), .A2(n9304), .A3(n7602), .ZN(n5277) );
  NAND2_X1 U6977 ( .A1(n5260), .A2(n5277), .ZN(n9198) );
  OR2_X1 U6978 ( .A1(n4290), .A2(n9198), .ZN(n5261) );
  NAND2_X1 U6979 ( .A1(n8354), .A2(n8304), .ZN(n6712) );
  NAND2_X1 U6980 ( .A1(n6597), .A2(n6712), .ZN(n8285) );
  NAND2_X1 U6981 ( .A1(n8282), .A2(n8285), .ZN(n8281) );
  INV_X1 U6982 ( .A(n8304), .ZN(n9365) );
  OR2_X1 U6983 ( .A1(n8354), .A2(n9365), .ZN(n5265) );
  NAND2_X1 U6984 ( .A1(n8281), .A2(n5265), .ZN(n8311) );
  INV_X1 U6985 ( .A(n5266), .ZN(n5270) );
  INV_X1 U6986 ( .A(n5267), .ZN(n5268) );
  NAND2_X1 U6987 ( .A1(n5268), .A2(SI_12_), .ZN(n5269) );
  MUX2_X1 U6988 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n4292), .Z(n5287) );
  XNOR2_X1 U6989 ( .A(n5287), .B(SI_13_), .ZN(n5285) );
  XNOR2_X1 U6990 ( .A(n5286), .B(n5285), .ZN(n7541) );
  NAND2_X1 U6991 ( .A1(n7541), .A2(n5397), .ZN(n5275) );
  NAND2_X1 U6992 ( .A1(n5272), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5273) );
  XNOR2_X1 U6993 ( .A(n5273), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9525) );
  AOI22_X1 U6994 ( .A1(n9525), .A2(n7441), .B1(n5137), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6995 ( .A1(n5153), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5283) );
  INV_X1 U6996 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9514) );
  OR2_X1 U6997 ( .A1(n6530), .A2(n9514), .ZN(n5282) );
  INV_X1 U6998 ( .A(n5277), .ZN(n5276) );
  INV_X1 U6999 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U7000 ( .A1(n5277), .A2(n10313), .ZN(n5278) );
  NAND2_X1 U7001 ( .A1(n5291), .A2(n5278), .ZN(n9281) );
  OR2_X1 U7002 ( .A1(n4291), .A2(n9281), .ZN(n5281) );
  INV_X1 U7003 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5279) );
  OR2_X1 U7004 ( .A1(n5583), .A2(n5279), .ZN(n5280) );
  OR2_X1 U7005 ( .A1(n9880), .A2(n8287), .ZN(n6716) );
  NAND2_X1 U7006 ( .A1(n9880), .A2(n8287), .ZN(n6713) );
  NAND2_X1 U7007 ( .A1(n6716), .A2(n6713), .ZN(n8310) );
  INV_X1 U7008 ( .A(n8287), .ZN(n9364) );
  OR2_X1 U7009 ( .A1(n9880), .A2(n9364), .ZN(n5284) );
  MUX2_X1 U7010 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7342), .Z(n5303) );
  XNOR2_X1 U7011 ( .A(n5303), .B(SI_14_), .ZN(n5300) );
  XNOR2_X1 U7012 ( .A(n5302), .B(n5300), .ZN(n7636) );
  NAND2_X1 U7013 ( .A1(n7636), .A2(n5397), .ZN(n5290) );
  OR2_X1 U7014 ( .A1(n5307), .A2(n9983), .ZN(n5288) );
  XNOR2_X1 U7015 ( .A(n5288), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U7016 ( .A1(n5137), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n7441), .B2(
        n9527), .ZN(n5289) );
  NAND2_X1 U7017 ( .A1(n5153), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5297) );
  INV_X1 U7018 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9515) );
  OR2_X1 U7019 ( .A1(n5065), .A2(n9515), .ZN(n5296) );
  NAND2_X1 U7020 ( .A1(n5291), .A2(n9105), .ZN(n5292) );
  NAND2_X1 U7021 ( .A1(n5314), .A2(n5292), .ZN(n9107) );
  OR2_X1 U7022 ( .A1(n4291), .A2(n9107), .ZN(n5295) );
  INV_X1 U7023 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5293) );
  OR2_X1 U7024 ( .A1(n5583), .A2(n5293), .ZN(n5294) );
  NAND4_X1 U7025 ( .A1(n5297), .A2(n5296), .A3(n5295), .A4(n5294), .ZN(n9363)
         );
  NAND2_X1 U7026 ( .A1(n9967), .A2(n9363), .ZN(n5298) );
  OR2_X1 U7027 ( .A1(n9967), .A2(n9363), .ZN(n5299) );
  INV_X1 U7028 ( .A(n5300), .ZN(n5301) );
  NAND2_X1 U7029 ( .A1(n5302), .A2(n5301), .ZN(n5305) );
  NAND2_X1 U7030 ( .A1(n5303), .A2(SI_14_), .ZN(n5304) );
  MUX2_X1 U7031 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n4286), .Z(n5321) );
  XNOR2_X1 U7032 ( .A(n5321), .B(SI_15_), .ZN(n5306) );
  XNOR2_X1 U7033 ( .A(n5322), .B(n5306), .ZN(n7705) );
  NAND2_X1 U7034 ( .A1(n7705), .A2(n5397), .ZN(n5312) );
  NAND2_X1 U7035 ( .A1(n5309), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5308) );
  MUX2_X1 U7036 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5308), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5310) );
  INV_X1 U7037 ( .A(n5347), .ZN(n5589) );
  AND2_X1 U7038 ( .A1(n5310), .A2(n5589), .ZN(n10029) );
  AOI22_X1 U7039 ( .A1(n5137), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n7441), .B2(
        n10029), .ZN(n5311) );
  NAND2_X1 U7040 ( .A1(n5579), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5319) );
  INV_X1 U7041 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9782) );
  OR2_X1 U7042 ( .A1(n6534), .A2(n9782), .ZN(n5318) );
  INV_X1 U7043 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U7044 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U7045 ( .A1(n5331), .A2(n5315), .ZN(n9781) );
  OR2_X1 U7046 ( .A1(n4290), .A2(n9781), .ZN(n5317) );
  INV_X1 U7047 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9961) );
  OR2_X1 U7048 ( .A1(n5583), .A2(n9961), .ZN(n5316) );
  NAND4_X1 U7049 ( .A1(n5319), .A2(n5318), .A3(n5317), .A4(n5316), .ZN(n9362)
         );
  NOR2_X1 U7050 ( .A1(n9870), .A2(n9362), .ZN(n5320) );
  NAND2_X1 U7051 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  MUX2_X1 U7052 ( .A(n7745), .B(n7742), .S(n7342), .Z(n5337) );
  XNOR2_X1 U7053 ( .A(n5337), .B(SI_16_), .ZN(n5327) );
  XNOR2_X1 U7054 ( .A(n5341), .B(n5327), .ZN(n7741) );
  NAND2_X1 U7055 ( .A1(n7741), .A2(n5397), .ZN(n5330) );
  NAND2_X1 U7056 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5328) );
  XNOR2_X1 U7057 ( .A(n5328), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U7058 ( .A1(n5137), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n7441), .B2(
        n9540), .ZN(n5329) );
  NAND2_X1 U7059 ( .A1(n5063), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5336) );
  INV_X1 U7060 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9865) );
  OR2_X1 U7061 ( .A1(n6530), .A2(n9865), .ZN(n5335) );
  NAND2_X1 U7062 ( .A1(n5331), .A2(n9222), .ZN(n5332) );
  NAND2_X1 U7063 ( .A1(n5353), .A2(n5332), .ZN(n9759) );
  OR2_X1 U7064 ( .A1(n4290), .A2(n9759), .ZN(n5334) );
  INV_X1 U7065 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9760) );
  OR2_X1 U7066 ( .A1(n6534), .A2(n9760), .ZN(n5333) );
  NAND2_X1 U7067 ( .A1(n9861), .A2(n9335), .ZN(n6691) );
  NAND2_X1 U7068 ( .A1(n6614), .A2(n6691), .ZN(n9753) );
  INV_X1 U7069 ( .A(n9335), .ZN(n9361) );
  NOR2_X1 U7070 ( .A1(n5338), .A2(SI_16_), .ZN(n5340) );
  NAND2_X1 U7071 ( .A1(n5338), .A2(SI_16_), .ZN(n5339) );
  MUX2_X1 U7072 ( .A(n10253), .B(n7868), .S(n4286), .Z(n5343) );
  NAND2_X1 U7073 ( .A1(n5343), .A2(n5342), .ZN(n5362) );
  INV_X1 U7074 ( .A(n5343), .ZN(n5344) );
  NAND2_X1 U7075 ( .A1(n5344), .A2(SI_17_), .ZN(n5345) );
  NAND2_X1 U7076 ( .A1(n5362), .A2(n5345), .ZN(n5360) );
  XNOR2_X1 U7077 ( .A(n5361), .B(n5360), .ZN(n7866) );
  NAND2_X1 U7078 ( .A1(n7866), .A2(n5397), .ZN(n5350) );
  NAND2_X1 U7079 ( .A1(n5595), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5348) );
  XNOR2_X1 U7080 ( .A(n5348), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9553) );
  AOI22_X1 U7081 ( .A1(n5137), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n7441), .B2(
        n9553), .ZN(n5349) );
  NAND2_X1 U7082 ( .A1(n5063), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5358) );
  INV_X1 U7083 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9857) );
  OR2_X1 U7084 ( .A1(n5065), .A2(n9857), .ZN(n5357) );
  INV_X1 U7085 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5352) );
  NAND2_X1 U7086 ( .A1(n5353), .A2(n5352), .ZN(n5354) );
  NAND2_X1 U7087 ( .A1(n5367), .A2(n5354), .ZN(n9744) );
  OR2_X1 U7088 ( .A1(n4291), .A2(n9744), .ZN(n5356) );
  INV_X1 U7089 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9745) );
  OR2_X1 U7090 ( .A1(n6534), .A2(n9745), .ZN(n5355) );
  NAND4_X1 U7091 ( .A1(n5358), .A2(n5357), .A3(n5356), .A4(n5355), .ZN(n9360)
         );
  OR2_X1 U7092 ( .A1(n9951), .A2(n9360), .ZN(n5359) );
  MUX2_X1 U7093 ( .A(n7946), .B(n10314), .S(n7342), .Z(n5376) );
  XNOR2_X1 U7094 ( .A(n5376), .B(SI_18_), .ZN(n5375) );
  XNOR2_X1 U7095 ( .A(n5378), .B(n5375), .ZN(n7924) );
  NAND2_X1 U7096 ( .A1(n7924), .A2(n5397), .ZN(n5365) );
  NAND2_X1 U7097 ( .A1(n5347), .A2(n4969), .ZN(n5363) );
  XNOR2_X1 U7098 ( .A(n5384), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U7099 ( .A1(n5137), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9557), .B2(
        n7441), .ZN(n5364) );
  NAND2_X1 U7100 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NAND2_X1 U7101 ( .A1(n5389), .A2(n5368), .ZN(n9729) );
  NAND2_X1 U7102 ( .A1(n5063), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5369) );
  OAI21_X1 U7103 ( .B1(n9729), .B2(n4290), .A(n5369), .ZN(n5372) );
  INV_X1 U7104 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U7105 ( .A1(n5579), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5370) );
  OAI21_X1 U7106 ( .B1(n6534), .B2(n9730), .A(n5370), .ZN(n5371) );
  NOR2_X1 U7107 ( .A1(n9852), .A2(n9359), .ZN(n5373) );
  NAND2_X1 U7108 ( .A1(n9852), .A2(n9359), .ZN(n5374) );
  INV_X1 U7109 ( .A(n5376), .ZN(n5377) );
  MUX2_X1 U7110 ( .A(n10259), .B(n8389), .S(n7342), .Z(n5380) );
  NAND2_X1 U7111 ( .A1(n5380), .A2(n5379), .ZN(n5393) );
  INV_X1 U7112 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U7113 ( .A1(n5381), .A2(SI_19_), .ZN(n5382) );
  NAND2_X1 U7114 ( .A1(n5393), .A2(n5382), .ZN(n5394) );
  NAND2_X1 U7115 ( .A1(n8018), .A2(n5397), .ZN(n5388) );
  INV_X1 U7116 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5383) );
  NAND2_X1 U7117 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  AOI22_X1 U7118 ( .A1(n5672), .A2(n7441), .B1(n5137), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n5387) );
  INV_X1 U7119 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9942) );
  INV_X1 U7120 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9159) );
  NAND2_X1 U7121 ( .A1(n5389), .A2(n9159), .ZN(n5390) );
  NAND2_X1 U7122 ( .A1(n5400), .A2(n5390), .ZN(n9710) );
  OR2_X1 U7123 ( .A1(n9710), .A2(n4291), .ZN(n5392) );
  AOI22_X1 U7124 ( .A1(n5153), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n5579), .B2(
        P1_REG1_REG_19__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U7125 ( .C1(n5583), .C2(n9942), .A(n5392), .B(n5391), .ZN(n9358)
         );
  OR2_X1 U7126 ( .A1(n9847), .A2(n9358), .ZN(n9687) );
  MUX2_X1 U7127 ( .A(n8210), .B(n8187), .S(n7342), .Z(n5423) );
  XNOR2_X1 U7128 ( .A(n5423), .B(SI_20_), .ZN(n5396) );
  NAND2_X1 U7129 ( .A1(n8186), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U7130 ( .A1(n5137), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5398) );
  INV_X1 U7131 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U7132 ( .A1(n5400), .A2(n9270), .ZN(n5401) );
  NAND2_X1 U7133 ( .A1(n5413), .A2(n5401), .ZN(n9269) );
  OR2_X1 U7134 ( .A1(n9269), .A2(n4290), .ZN(n5403) );
  AOI22_X1 U7135 ( .A1(n5153), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n5579), .B2(
        P1_REG1_REG_20__SCAN_IN), .ZN(n5402) );
  OAI211_X1 U7136 ( .C1(n5583), .C2(n9938), .A(n5403), .B(n5402), .ZN(n9357)
         );
  OR2_X1 U7137 ( .A1(n9843), .A2(n9357), .ZN(n6778) );
  AND2_X1 U7138 ( .A1(n9687), .A2(n6778), .ZN(n5406) );
  INV_X1 U7139 ( .A(n6778), .ZN(n5405) );
  NAND2_X1 U7140 ( .A1(n9843), .A2(n9357), .ZN(n6779) );
  NAND2_X1 U7141 ( .A1(n9847), .A2(n9358), .ZN(n9688) );
  AND2_X1 U7142 ( .A1(n6779), .A2(n9688), .ZN(n5404) );
  NAND2_X1 U7143 ( .A1(n5430), .A2(n5422), .ZN(n5407) );
  NAND2_X1 U7144 ( .A1(n5408), .A2(n5407), .ZN(n5410) );
  MUX2_X1 U7145 ( .A(n10233), .B(n8300), .S(n7342), .Z(n5420) );
  XNOR2_X1 U7146 ( .A(n5420), .B(SI_21_), .ZN(n5409) );
  NAND2_X1 U7147 ( .A1(n5137), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U7148 ( .A1(n5413), .A2(n10221), .ZN(n5414) );
  AND2_X1 U7149 ( .A1(n5438), .A2(n5414), .ZN(n9681) );
  NAND2_X1 U7150 ( .A1(n9681), .A2(n5531), .ZN(n5419) );
  INV_X1 U7151 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U7152 ( .A1(n5153), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7153 ( .A1(n5063), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5415) );
  OAI211_X1 U7154 ( .C1(n5065), .C2(n10274), .A(n5416), .B(n5415), .ZN(n5417)
         );
  INV_X1 U7155 ( .A(n5417), .ZN(n5418) );
  NAND2_X1 U7156 ( .A1(n5419), .A2(n5418), .ZN(n9356) );
  NOR2_X1 U7157 ( .A1(n7218), .A2(n9356), .ZN(n6757) );
  NAND2_X1 U7158 ( .A1(n7218), .A2(n9356), .ZN(n6755) );
  INV_X1 U7159 ( .A(n5423), .ZN(n5425) );
  OAI22_X1 U7160 ( .A1(SI_20_), .A2(n5425), .B1(n5426), .B2(SI_21_), .ZN(n5429) );
  INV_X1 U7161 ( .A(SI_21_), .ZN(n5421) );
  OAI21_X1 U7162 ( .B1(n5423), .B2(n5422), .A(n5421), .ZN(n5427) );
  AND2_X1 U7163 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5424) );
  AOI22_X1 U7164 ( .A1(n5427), .A2(n5426), .B1(n5425), .B2(n5424), .ZN(n5428)
         );
  MUX2_X1 U7165 ( .A(n8344), .B(n8341), .S(n7342), .Z(n5432) );
  NAND2_X1 U7166 ( .A1(n5432), .A2(n5431), .ZN(n5445) );
  INV_X1 U7167 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U7168 ( .A1(n5433), .A2(SI_22_), .ZN(n5434) );
  NAND2_X1 U7169 ( .A1(n5445), .A2(n5434), .ZN(n5446) );
  XNOR2_X1 U7170 ( .A(n5447), .B(n5446), .ZN(n8339) );
  NAND2_X1 U7171 ( .A1(n8339), .A2(n5397), .ZN(n5436) );
  NAND2_X1 U7172 ( .A1(n5137), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5435) );
  INV_X1 U7173 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U7174 ( .A1(n5438), .A2(n5437), .ZN(n5439) );
  NAND2_X1 U7175 ( .A1(n5457), .A2(n5439), .ZN(n9663) );
  INV_X1 U7176 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n9664) );
  NAND2_X1 U7177 ( .A1(n5063), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U7178 ( .A1(n5579), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5440) );
  OAI211_X1 U7179 ( .C1(n6534), .C2(n9664), .A(n5441), .B(n5440), .ZN(n5442)
         );
  INV_X1 U7180 ( .A(n5442), .ZN(n5443) );
  NAND2_X1 U7181 ( .A1(n5444), .A2(n5443), .ZN(n9355) );
  NAND2_X1 U7182 ( .A1(n9931), .A2(n9355), .ZN(n9637) );
  NAND2_X1 U7183 ( .A1(n9662), .A2(n9118), .ZN(n6645) );
  INV_X1 U7184 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5448) );
  MUX2_X1 U7185 ( .A(n8347), .B(n5448), .S(n7342), .Z(n5450) );
  INV_X1 U7186 ( .A(n5450), .ZN(n5451) );
  NAND2_X1 U7187 ( .A1(n5451), .A2(SI_23_), .ZN(n5452) );
  NAND2_X1 U7188 ( .A1(n6155), .A2(n5397), .ZN(n5454) );
  NAND2_X1 U7189 ( .A1(n5137), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5453) );
  INV_X1 U7190 ( .A(n5457), .ZN(n5455) );
  INV_X1 U7191 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U7192 ( .A1(n5457), .A2(n5456), .ZN(n5458) );
  NAND2_X1 U7193 ( .A1(n5474), .A2(n5458), .ZN(n9646) );
  OR2_X1 U7194 ( .A1(n9646), .A2(n4291), .ZN(n5463) );
  INV_X1 U7195 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9925) );
  NAND2_X1 U7196 ( .A1(n5153), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U7197 ( .A1(n5579), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5459) );
  OAI211_X1 U7198 ( .C1(n9925), .C2(n5583), .A(n5460), .B(n5459), .ZN(n5461)
         );
  INV_X1 U7199 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U7200 ( .A1(n9922), .A2(n9292), .ZN(n6727) );
  OR2_X1 U7201 ( .A1(n9922), .A2(n9354), .ZN(n5464) );
  NAND2_X1 U7202 ( .A1(n9641), .A2(n5464), .ZN(n9626) );
  MUX2_X1 U7203 ( .A(n8375), .B(n8373), .S(n7342), .Z(n5469) );
  INV_X1 U7204 ( .A(n5469), .ZN(n5470) );
  NAND2_X1 U7205 ( .A1(n5470), .A2(SI_24_), .ZN(n5471) );
  XNOR2_X1 U7206 ( .A(n5482), .B(n5481), .ZN(n8372) );
  NAND2_X1 U7207 ( .A1(n8372), .A2(n5397), .ZN(n5473) );
  NAND2_X1 U7208 ( .A1(n5137), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5472) );
  INV_X1 U7209 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9241) );
  NAND2_X1 U7210 ( .A1(n5474), .A2(n9241), .ZN(n5475) );
  AND2_X1 U7211 ( .A1(n5493), .A2(n5475), .ZN(n9631) );
  NAND2_X1 U7212 ( .A1(n9631), .A2(n5531), .ZN(n5480) );
  INV_X1 U7213 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U7214 ( .A1(n5153), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U7215 ( .A1(n5063), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5476) );
  OAI211_X1 U7216 ( .C1(n5065), .C2(n10311), .A(n5477), .B(n5476), .ZN(n5478)
         );
  INV_X1 U7217 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7218 ( .A1(n9920), .A2(n9119), .ZN(n6738) );
  NAND2_X1 U7219 ( .A1(n9606), .A2(n6738), .ZN(n9625) );
  NAND2_X1 U7220 ( .A1(n9626), .A2(n9625), .ZN(n9624) );
  OR2_X1 U7221 ( .A1(n9920), .A2(n9353), .ZN(n6644) );
  NAND2_X1 U7222 ( .A1(n9624), .A2(n6644), .ZN(n9605) );
  NAND2_X1 U7223 ( .A1(n5482), .A2(n5481), .ZN(n5484) );
  NAND2_X1 U7224 ( .A1(n5484), .A2(n5483), .ZN(n5505) );
  MUX2_X1 U7225 ( .A(n9098), .B(n10191), .S(n7342), .Z(n5486) );
  INV_X1 U7226 ( .A(SI_25_), .ZN(n5485) );
  NAND2_X1 U7227 ( .A1(n5486), .A2(n5485), .ZN(n5506) );
  INV_X1 U7228 ( .A(n5486), .ZN(n5487) );
  NAND2_X1 U7229 ( .A1(n5487), .A2(SI_25_), .ZN(n5488) );
  XNOR2_X1 U7230 ( .A(n5505), .B(n5504), .ZN(n8377) );
  NAND2_X1 U7231 ( .A1(n8377), .A2(n5397), .ZN(n5490) );
  NAND2_X1 U7232 ( .A1(n5137), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5489) );
  INV_X1 U7233 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5492) );
  NAND2_X1 U7234 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  NAND2_X1 U7235 ( .A1(n5513), .A2(n5494), .ZN(n9614) );
  INV_X1 U7236 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7237 ( .A1(n5153), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7238 ( .A1(n5579), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U7239 ( .C1(n5497), .C2(n5583), .A(n5496), .B(n5495), .ZN(n5498)
         );
  INV_X1 U7240 ( .A(n5498), .ZN(n5499) );
  NAND2_X2 U7241 ( .A1(n5500), .A2(n5499), .ZN(n9352) );
  NAND2_X1 U7242 ( .A1(n9211), .A2(n9352), .ZN(n5501) );
  OR2_X1 U7243 ( .A1(n9211), .A2(n9352), .ZN(n5502) );
  NAND2_X1 U7244 ( .A1(n5505), .A2(n5504), .ZN(n5507) );
  INV_X1 U7245 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9996) );
  MUX2_X1 U7246 ( .A(n9095), .B(n9996), .S(n7342), .Z(n5508) );
  INV_X1 U7247 ( .A(SI_26_), .ZN(n10276) );
  NAND2_X1 U7248 ( .A1(n5508), .A2(n10276), .ZN(n5524) );
  INV_X1 U7249 ( .A(n5508), .ZN(n5509) );
  NAND2_X1 U7250 ( .A1(n5509), .A2(SI_26_), .ZN(n5510) );
  NAND2_X1 U7251 ( .A1(n9094), .A2(n5397), .ZN(n5512) );
  NAND2_X1 U7252 ( .A1(n5137), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5511) );
  INV_X1 U7253 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9325) );
  OR2_X2 U7254 ( .A1(n5513), .A2(n9325), .ZN(n5546) );
  NAND2_X1 U7255 ( .A1(n5513), .A2(n9325), .ZN(n5514) );
  NAND2_X1 U7256 ( .A1(n9599), .A2(n5531), .ZN(n5519) );
  NAND2_X1 U7257 ( .A1(n5063), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7258 ( .A1(n5579), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5515) );
  OAI211_X1 U7259 ( .C1(n6534), .C2(n10297), .A(n5516), .B(n5515), .ZN(n5517)
         );
  INV_X1 U7260 ( .A(n5517), .ZN(n5518) );
  NAND2_X2 U7261 ( .A1(n5519), .A2(n5518), .ZN(n9351) );
  NOR2_X1 U7262 ( .A1(n9814), .A2(n9351), .ZN(n5521) );
  NAND2_X1 U7263 ( .A1(n9814), .A2(n9351), .ZN(n5520) );
  INV_X1 U7264 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n6205) );
  INV_X1 U7265 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9991) );
  MUX2_X1 U7266 ( .A(n6205), .B(n9991), .S(n7342), .Z(n5526) );
  INV_X1 U7267 ( .A(n5526), .ZN(n5527) );
  NAND2_X1 U7268 ( .A1(n5527), .A2(SI_27_), .ZN(n5528) );
  XNOR2_X1 U7269 ( .A(n5539), .B(n5538), .ZN(n9089) );
  NAND2_X1 U7270 ( .A1(n9089), .A2(n5576), .ZN(n5530) );
  NAND2_X1 U7271 ( .A1(n5137), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5529) );
  XNOR2_X1 U7272 ( .A(n5546), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U7273 ( .A1(n9585), .A2(n5531), .ZN(n5536) );
  INV_X1 U7274 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U7275 ( .A1(n5153), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7276 ( .A1(n5579), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5532) );
  OAI211_X1 U7277 ( .C1(n9907), .C2(n5583), .A(n5533), .B(n5532), .ZN(n5534)
         );
  INV_X1 U7278 ( .A(n5534), .ZN(n5535) );
  NAND2_X1 U7279 ( .A1(n6668), .A2(n7272), .ZN(n6743) );
  OR2_X1 U7280 ( .A1(n6668), .A2(n9350), .ZN(n6660) );
  INV_X1 U7281 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n6217) );
  INV_X1 U7282 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8397) );
  MUX2_X1 U7283 ( .A(n6217), .B(n8397), .S(n7342), .Z(n5541) );
  INV_X1 U7284 ( .A(SI_28_), .ZN(n5540) );
  NAND2_X1 U7285 ( .A1(n5541), .A2(n5540), .ZN(n5561) );
  INV_X1 U7286 ( .A(n5541), .ZN(n5542) );
  NAND2_X1 U7287 ( .A1(n5542), .A2(SI_28_), .ZN(n5565) );
  NAND2_X1 U7288 ( .A1(n8396), .A2(n5397), .ZN(n5544) );
  NAND2_X1 U7289 ( .A1(n5137), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5543) );
  INV_X1 U7290 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n7299) );
  INV_X1 U7291 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5545) );
  OAI21_X1 U7292 ( .B1(n5546), .B2(n7299), .A(n5545), .ZN(n5549) );
  INV_X1 U7293 ( .A(n5546), .ZN(n5548) );
  AND2_X1 U7294 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5547) );
  NAND2_X1 U7295 ( .A1(n5548), .A2(n5547), .ZN(n8429) );
  NAND2_X1 U7296 ( .A1(n5549), .A2(n8429), .ZN(n9574) );
  INV_X1 U7297 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10298) );
  NAND2_X1 U7298 ( .A1(n5579), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7299 ( .A1(n5153), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5550) );
  OAI211_X1 U7300 ( .C1(n5583), .C2(n10298), .A(n5551), .B(n5550), .ZN(n5552)
         );
  INV_X1 U7301 ( .A(n5552), .ZN(n5553) );
  NAND2_X1 U7302 ( .A1(n8419), .A2(n8404), .ZN(n6742) );
  NAND2_X1 U7303 ( .A1(n6371), .A2(n6665), .ZN(n6373) );
  NAND2_X1 U7304 ( .A1(n8419), .A2(n5555), .ZN(n5556) );
  INV_X1 U7305 ( .A(n5560), .ZN(n5559) );
  MUX2_X1 U7306 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7342), .Z(n5562) );
  INV_X1 U7307 ( .A(n5562), .ZN(n5557) );
  NAND2_X1 U7308 ( .A1(n5565), .A2(n5557), .ZN(n5564) );
  INV_X1 U7309 ( .A(n5564), .ZN(n5558) );
  NAND2_X1 U7310 ( .A1(n5559), .A2(n5558), .ZN(n5571) );
  NAND2_X1 U7311 ( .A1(n5561), .A2(n5562), .ZN(n5566) );
  INV_X1 U7312 ( .A(n5566), .ZN(n6512) );
  NAND3_X1 U7313 ( .A1(n5560), .A2(n6512), .A3(n5563), .ZN(n5570) );
  OAI22_X1 U7314 ( .A1(n5564), .A2(n5563), .B1(n5562), .B2(n5561), .ZN(n5568)
         );
  NOR2_X1 U7315 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  NOR2_X1 U7316 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  NAND3_X1 U7317 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n5574) );
  INV_X1 U7318 ( .A(n5574), .ZN(n5573) );
  INV_X1 U7319 ( .A(SI_29_), .ZN(n5572) );
  NAND2_X1 U7320 ( .A1(n5574), .A2(n5572), .ZN(n5575) );
  OR2_X1 U7321 ( .A1(n8429), .A2(n4290), .ZN(n5586) );
  INV_X1 U7322 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7323 ( .A1(n5579), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5581) );
  NAND2_X1 U7324 ( .A1(n5153), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5580) );
  OAI211_X1 U7325 ( .C1(n5583), .C2(n5582), .A(n5581), .B(n5580), .ZN(n5584)
         );
  INV_X1 U7326 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7327 ( .A1(n5586), .A2(n5585), .ZN(n9349) );
  OAI21_X1 U7328 ( .B1(n5589), .B2(n5588), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5591) );
  NAND2_X1 U7329 ( .A1(n8378), .A2(P1_B_REG_SCAN_IN), .ZN(n5601) );
  NOR2_X2 U7330 ( .A1(n5595), .A2(n5594), .ZN(n5630) );
  NAND2_X1 U7331 ( .A1(n5630), .A2(n5596), .ZN(n5629) );
  INV_X1 U7332 ( .A(n5629), .ZN(n5598) );
  INV_X1 U7333 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7334 ( .A1(n5598), .A2(n5597), .ZN(n5617) );
  NAND2_X1 U7335 ( .A1(n5618), .A2(n5619), .ZN(n5599) );
  OAI21_X2 U7336 ( .B1(n5617), .B2(n5599), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5600) );
  MUX2_X1 U7337 ( .A(n5601), .B(P1_B_REG_SCAN_IN), .S(n5624), .Z(n5604) );
  NAND2_X1 U7338 ( .A1(n5602), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5603) );
  INV_X1 U7339 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5605) );
  INV_X1 U7340 ( .A(n5624), .ZN(n8374) );
  INV_X1 U7341 ( .A(n5621), .ZN(n9997) );
  NOR4_X1 U7342 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5609) );
  NOR4_X1 U7343 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5608) );
  NOR4_X1 U7344 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5607) );
  NOR4_X1 U7345 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5606) );
  AND4_X1 U7346 ( .A1(n5609), .A2(n5608), .A3(n5607), .A4(n5606), .ZN(n5615)
         );
  NOR2_X1 U7347 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .ZN(
        n5613) );
  NOR4_X1 U7348 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5612) );
  NOR4_X1 U7349 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5611) );
  NOR4_X1 U7350 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5610) );
  AND4_X1 U7351 ( .A1(n5613), .A2(n5612), .A3(n5611), .A4(n5610), .ZN(n5614)
         );
  NAND2_X1 U7352 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  NAND2_X1 U7353 ( .A1(n7427), .A2(n5616), .ZN(n7280) );
  INV_X1 U7354 ( .A(n8378), .ZN(n5622) );
  AND2_X2 U7355 ( .A1(n5627), .A2(n5626), .ZN(n7064) );
  NAND2_X1 U7356 ( .A1(n5629), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5628) );
  INV_X1 U7357 ( .A(n5630), .ZN(n5631) );
  NAND2_X1 U7358 ( .A1(n5631), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5632) );
  NOR2_X1 U7359 ( .A1(n7287), .A2(n7065), .ZN(n5634) );
  NOR2_X1 U7360 ( .A1(n7445), .A2(n5634), .ZN(n5635) );
  NAND2_X1 U7361 ( .A1(n7280), .A2(n5635), .ZN(n5919) );
  NOR2_X1 U7362 ( .A1(n7327), .A2(n5919), .ZN(n5638) );
  INV_X1 U7363 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7364 ( .A1(n7427), .A2(n5636), .ZN(n5637) );
  NAND2_X1 U7365 ( .A1(n8378), .A2(n9997), .ZN(n9980) );
  NAND2_X1 U7366 ( .A1(n5637), .A2(n9980), .ZN(n7279) );
  MUX2_X1 U7367 ( .A(n9801), .B(n7065), .S(n7068), .Z(n5639) );
  INV_X1 U7368 ( .A(n9797), .ZN(n9802) );
  NAND2_X1 U7369 ( .A1(n7063), .A2(n8340), .ZN(n10067) );
  NOR2_X1 U7370 ( .A1(n6693), .A2(n7715), .ZN(n7322) );
  NAND2_X1 U7371 ( .A1(n7073), .A2(n4293), .ZN(n5641) );
  NAND2_X1 U7372 ( .A1(n9374), .A2(n8172), .ZN(n6697) );
  INV_X1 U7373 ( .A(n7849), .ZN(n6758) );
  NAND2_X1 U7374 ( .A1(n7840), .A2(n6758), .ZN(n7818) );
  NAND2_X1 U7375 ( .A1(n6765), .A2(n8154), .ZN(n5644) );
  OR2_X1 U7376 ( .A1(n6764), .A2(n5644), .ZN(n5645) );
  INV_X1 U7377 ( .A(n6765), .ZN(n8259) );
  NAND2_X1 U7378 ( .A1(n6583), .A2(n6592), .ZN(n5646) );
  NAND2_X1 U7379 ( .A1(n5647), .A2(n5646), .ZN(n6707) );
  NAND2_X1 U7380 ( .A1(n6707), .A2(n6768), .ZN(n5648) );
  OAI21_X1 U7381 ( .B1(n7886), .B2(n5645), .A(n5648), .ZN(n5649) );
  INV_X1 U7382 ( .A(n8000), .ZN(n8006) );
  NAND2_X1 U7383 ( .A1(n8005), .A2(n8006), .ZN(n8004) );
  INV_X1 U7384 ( .A(n8283), .ZN(n5651) );
  NOR2_X1 U7385 ( .A1(n8285), .A2(n5651), .ZN(n5653) );
  INV_X1 U7386 ( .A(n6597), .ZN(n5652) );
  AOI21_X2 U7387 ( .B1(n8284), .B2(n5653), .A(n5652), .ZN(n8303) );
  NAND2_X1 U7388 ( .A1(n8303), .A2(n5654), .ZN(n8302) );
  OR2_X1 U7389 ( .A1(n9967), .A2(n9338), .ZN(n6773) );
  NAND2_X1 U7390 ( .A1(n8359), .A2(n6773), .ZN(n5655) );
  NAND2_X1 U7391 ( .A1(n9967), .A2(n9338), .ZN(n6772) );
  NAND2_X1 U7392 ( .A1(n5655), .A2(n6772), .ZN(n9773) );
  INV_X1 U7393 ( .A(n9362), .ZN(n9221) );
  OR2_X1 U7394 ( .A1(n9870), .A2(n9221), .ZN(n6611) );
  NAND2_X1 U7395 ( .A1(n9870), .A2(n9221), .ZN(n9752) );
  NAND2_X1 U7396 ( .A1(n6691), .A2(n9752), .ZN(n6692) );
  NAND2_X1 U7397 ( .A1(n6692), .A2(n6614), .ZN(n6617) );
  INV_X1 U7398 ( .A(n9360), .ZN(n9312) );
  OR2_X1 U7399 ( .A1(n9951), .A2(n9312), .ZN(n9721) );
  NAND2_X1 U7400 ( .A1(n9951), .A2(n9312), .ZN(n6627) );
  INV_X1 U7401 ( .A(n9359), .ZN(n5656) );
  OR2_X1 U7402 ( .A1(n9852), .A2(n5656), .ZN(n6629) );
  NAND2_X1 U7403 ( .A1(n9852), .A2(n5656), .ZN(n6628) );
  NAND2_X1 U7404 ( .A1(n6629), .A2(n6628), .ZN(n9723) );
  INV_X1 U7405 ( .A(n9721), .ZN(n5657) );
  NOR2_X1 U7406 ( .A1(n9723), .A2(n5657), .ZN(n5658) );
  NAND2_X1 U7407 ( .A1(n9720), .A2(n5658), .ZN(n5659) );
  NAND2_X1 U7408 ( .A1(n5659), .A2(n6628), .ZN(n9704) );
  INV_X1 U7409 ( .A(n9358), .ZN(n9313) );
  NAND2_X1 U7410 ( .A1(n9847), .A2(n9313), .ZN(n6690) );
  NAND2_X1 U7411 ( .A1(n9704), .A2(n9705), .ZN(n5660) );
  INV_X1 U7412 ( .A(n9356), .ZN(n9291) );
  OR2_X1 U7413 ( .A1(n7218), .A2(n9291), .ZN(n6635) );
  INV_X1 U7414 ( .A(n9357), .ZN(n5661) );
  OR2_X1 U7415 ( .A1(n9843), .A2(n5661), .ZN(n9672) );
  NAND2_X1 U7416 ( .A1(n7218), .A2(n9291), .ZN(n6639) );
  NAND2_X1 U7417 ( .A1(n9843), .A2(n5661), .ZN(n6559) );
  NAND2_X1 U7418 ( .A1(n6639), .A2(n6559), .ZN(n6625) );
  NAND2_X1 U7419 ( .A1(n6625), .A2(n6635), .ZN(n6737) );
  INV_X1 U7420 ( .A(n9652), .ZN(n9657) );
  INV_X1 U7421 ( .A(n9637), .ZN(n5662) );
  NOR2_X1 U7422 ( .A1(n9642), .A2(n5662), .ZN(n5663) );
  NAND2_X1 U7423 ( .A1(n9636), .A2(n5663), .ZN(n5664) );
  INV_X1 U7424 ( .A(n9625), .ZN(n5665) );
  INV_X1 U7425 ( .A(n9352), .ZN(n7254) );
  OR2_X1 U7426 ( .A1(n9211), .A2(n7254), .ZN(n6541) );
  NAND2_X1 U7427 ( .A1(n9211), .A2(n7254), .ZN(n6543) );
  NAND2_X1 U7428 ( .A1(n9612), .A2(n6541), .ZN(n9592) );
  INV_X1 U7429 ( .A(n9592), .ZN(n5667) );
  XNOR2_X1 U7430 ( .A(n9814), .B(n6540), .ZN(n9593) );
  INV_X1 U7431 ( .A(n9593), .ZN(n5666) );
  NAND2_X1 U7432 ( .A1(n9814), .A2(n6540), .ZN(n6802) );
  INV_X1 U7433 ( .A(n6743), .ZN(n5669) );
  NOR2_X1 U7434 ( .A1(n6665), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U7435 ( .A1(n7064), .A2(n5672), .ZN(n5673) );
  INV_X1 U7436 ( .A(n8188), .ZN(n7282) );
  NAND2_X1 U7437 ( .A1(n7062), .A2(n7282), .ZN(n6824) );
  NAND2_X1 U7438 ( .A1(n5063), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5678) );
  INV_X1 U7439 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9810) );
  OR2_X1 U7440 ( .A1(n5065), .A2(n9810), .ZN(n5677) );
  INV_X1 U7441 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5675) );
  OR2_X1 U7442 ( .A1(n6534), .A2(n5675), .ZN(n5676) );
  AND3_X1 U7443 ( .A1(n5678), .A2(n5677), .A3(n5676), .ZN(n6750) );
  INV_X1 U7444 ( .A(P1_B_REG_SCAN_IN), .ZN(n5679) );
  OR2_X1 U7445 ( .A1(n10002), .A2(n5679), .ZN(n5680) );
  NAND2_X1 U7446 ( .A1(n9324), .A2(n5680), .ZN(n6529) );
  OAI22_X1 U7447 ( .A1(n8404), .A2(n9337), .B1(n6750), .B2(n6529), .ZN(n5681)
         );
  NAND3_X1 U7448 ( .A1(n7334), .A2(n8172), .A3(n7715), .ZN(n7845) );
  NOR2_X4 U7449 ( .A1(n7846), .A2(n8044), .ZN(n7939) );
  INV_X1 U7450 ( .A(n9172), .ZN(n9979) );
  AND2_X2 U7451 ( .A1(n8267), .A2(n9979), .ZN(n8162) );
  NAND2_X1 U7452 ( .A1(n8162), .A2(n9974), .ZN(n8009) );
  OR2_X2 U7453 ( .A1(n8009), .A2(n9133), .ZN(n8066) );
  INV_X1 U7454 ( .A(n8354), .ZN(n9204) );
  INV_X1 U7455 ( .A(n9880), .ZN(n9287) );
  INV_X1 U7456 ( .A(n9951), .ZN(n9743) );
  NAND2_X1 U7457 ( .A1(n9741), .A2(n9743), .ZN(n9742) );
  OR2_X2 U7458 ( .A1(n9742), .A2(n9852), .ZN(n9727) );
  OR2_X2 U7459 ( .A1(n9660), .A2(n9922), .ZN(n9644) );
  AND2_X2 U7460 ( .A1(n9628), .A2(n9913), .ZN(n9597) );
  OAI211_X1 U7461 ( .C1(n5685), .C2(n8432), .A(n9764), .B(n6509), .ZN(n8428)
         );
  NAND2_X1 U7462 ( .A1(n8427), .A2(n8428), .ZN(n6369) );
  NAND2_X1 U7463 ( .A1(n6369), .A2(n10070), .ZN(n5691) );
  AND2_X1 U7464 ( .A1(n9797), .A2(n5686), .ZN(n10064) );
  NAND2_X1 U7465 ( .A1(n10070), .A2(n10064), .ZN(n9978) );
  NAND2_X1 U7466 ( .A1(n4777), .A2(n5687), .ZN(n5689) );
  OR2_X1 U7467 ( .A1(n10070), .A2(n5582), .ZN(n5688) );
  NOR2_X4 U7468 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5748) );
  NOR2_X1 U7469 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5697) );
  NOR2_X1 U7470 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5696) );
  INV_X1 U7471 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5698) );
  NAND2_X1 U7472 ( .A1(n5710), .A2(n5708), .ZN(n5706) );
  OAI21_X1 U7473 ( .B1(n5714), .B2(n5706), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5707) );
  MUX2_X1 U7474 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5707), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5713) );
  NOR2_X1 U7475 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5711) );
  NAND2_X1 U7476 ( .A1(n5715), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5716) );
  MUX2_X1 U7477 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5716), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n5717) );
  NAND2_X1 U7478 ( .A1(n5789), .A2(n5794), .ZN(n5742) );
  INV_X1 U7479 ( .A(n5742), .ZN(n5720) );
  INV_X1 U7480 ( .A(n5712), .ZN(n5727) );
  NAND2_X1 U7481 ( .A1(n5727), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7482 ( .A1(n6980), .A2(n6492), .ZN(n5729) );
  NAND2_X1 U7483 ( .A1(n5729), .A2(n6500), .ZN(n5902) );
  XNOR2_X2 U7484 ( .A(n5731), .B(n5730), .ZN(n5804) );
  XNOR2_X2 U7485 ( .A(n5734), .B(n5733), .ZN(n5838) );
  NAND2_X4 U7486 ( .A1(n5804), .A2(n5838), .ZN(n6316) );
  NAND2_X1 U7487 ( .A1(n5902), .A2(n6316), .ZN(n5735) );
  NAND2_X1 U7488 ( .A1(n5735), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X1 U7489 ( .A1(n4348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U7490 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5736), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5737) );
  INV_X1 U7491 ( .A(n5737), .ZN(n5738) );
  NOR2_X1 U7492 ( .A1(n5738), .A2(n5799), .ZN(n8744) );
  INV_X1 U7493 ( .A(n8744), .ZN(n7948) );
  INV_X1 U7494 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7495 ( .A1(n5784), .A2(n5740), .ZN(n5787) );
  NAND2_X1 U7496 ( .A1(n5741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7497 ( .A1(n5742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5743) );
  NAND2_X1 U7498 ( .A1(n5790), .A2(n5743), .ZN(n5747) );
  OAI21_X1 U7499 ( .B1(n5747), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5745) );
  INV_X1 U7500 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5744) );
  XNOR2_X1 U7501 ( .A(n5745), .B(n5744), .ZN(n8720) );
  XNOR2_X1 U7502 ( .A(n5747), .B(n5746), .ZN(n7743) );
  INV_X1 U7503 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10277) );
  MUX2_X1 U7504 ( .A(n10277), .B(P2_REG2_REG_16__SCAN_IN), .S(n7743), .Z(n8688) );
  INV_X1 U7505 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5749) );
  INV_X1 U7506 ( .A(n7348), .ZN(n8630) );
  INV_X1 U7507 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10106) );
  NAND2_X1 U7508 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5751) );
  INV_X1 U7509 ( .A(n7587), .ZN(n5834) );
  INV_X1 U7510 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5937) );
  INV_X1 U7511 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5931) );
  OAI22_X1 U7512 ( .A1(n7581), .A2(n5931), .B1(n5937), .B2(n5755), .ZN(n7488)
         );
  NAND2_X1 U7513 ( .A1(n5756), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5757) );
  MUX2_X1 U7514 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5757), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5758) );
  INV_X1 U7515 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7644) );
  MUX2_X1 U7516 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n10106), .S(n7348), .Z(n8618)
         );
  OAI21_X1 U7517 ( .B1(n5761), .B2(P2_IR_REG_4__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  MUX2_X1 U7518 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5762), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5763) );
  AND2_X1 U7519 ( .A1(n5760), .A2(n5763), .ZN(n5987) );
  INV_X1 U7520 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U7521 ( .A1(n5760), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  MUX2_X1 U7522 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5765), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5767) );
  AND2_X1 U7523 ( .A1(n5767), .A2(n5766), .ZN(n6000) );
  MUX2_X1 U7524 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10286), .S(n6000), .Z(n7617)
         );
  NOR2_X2 U7525 ( .A1(n7616), .A2(n7617), .ZN(n7615) );
  INV_X1 U7526 ( .A(n6000), .ZN(n7614) );
  NAND2_X1 U7527 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5768) );
  XNOR2_X1 U7528 ( .A(n5768), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6014) );
  INV_X1 U7529 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7510) );
  INV_X1 U7530 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7996) );
  OR2_X1 U7531 ( .A1(n5769), .A2(n5923), .ZN(n5770) );
  XNOR2_X1 U7532 ( .A(n5770), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7679) );
  MUX2_X1 U7533 ( .A(n7996), .B(P2_REG2_REG_8__SCAN_IN), .S(n7679), .Z(n7673)
         );
  NAND2_X1 U7534 ( .A1(n5771), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5772) );
  NAND2_X2 U7535 ( .A1(n7671), .A2(n5772), .ZN(n5776) );
  NAND2_X1 U7536 ( .A1(n5773), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5774) );
  MUX2_X1 U7537 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5774), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n5775) );
  INV_X1 U7538 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5779) );
  NAND2_X1 U7539 ( .A1(n5777), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5778) );
  XNOR2_X1 U7540 ( .A(n5778), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7777) );
  MUX2_X1 U7541 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n5779), .S(n7777), .Z(n7768)
         );
  OR2_X1 U7542 ( .A1(n5781), .A2(n5923), .ZN(n5782) );
  XNOR2_X1 U7543 ( .A(n5782), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6048) );
  INV_X1 U7544 ( .A(n6048), .ZN(n7910) );
  OR2_X1 U7545 ( .A1(n5784), .A2(n5923), .ZN(n5785) );
  XNOR2_X1 U7546 ( .A(n5785), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7961) );
  MUX2_X1 U7547 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n5786), .S(n7961), .Z(n7951)
         );
  INV_X1 U7548 ( .A(n7961), .ZN(n7424) );
  NAND2_X1 U7549 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5788) );
  XNOR2_X1 U7550 ( .A(n5788), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7543) );
  INV_X1 U7551 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8323) );
  NAND2_X1 U7552 ( .A1(n5790), .A2(n5789), .ZN(n5793) );
  OR2_X1 U7553 ( .A1(n5790), .A2(n5789), .ZN(n5791) );
  INV_X1 U7554 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6085) );
  XNOR2_X1 U7555 ( .A(n8663), .B(n6085), .ZN(n8650) );
  NAND2_X1 U7556 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8663), .ZN(n5792) );
  NAND2_X1 U7557 ( .A1(n5793), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5795) );
  XNOR2_X1 U7558 ( .A(n5795), .B(n5794), .ZN(n8678) );
  NAND2_X1 U7559 ( .A1(n8678), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U7560 ( .A1(n8720), .A2(n5798), .ZN(n8733) );
  INV_X1 U7561 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8865) );
  XNOR2_X1 U7562 ( .A(n8744), .B(n8865), .ZN(n8731) );
  INV_X1 U7563 ( .A(n5799), .ZN(n5800) );
  NAND2_X1 U7564 ( .A1(n5800), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5802) );
  XNOR2_X1 U7565 ( .A(n8019), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n5898) );
  XNOR2_X1 U7566 ( .A(n5803), .B(n5898), .ZN(n5805) );
  NOR2_X1 U7567 ( .A1(n5804), .A2(P2_U3151), .ZN(n9086) );
  AND2_X1 U7568 ( .A1(n5902), .A2(n9086), .ZN(n7459) );
  INV_X1 U7569 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8954) );
  XNOR2_X1 U7570 ( .A(n7743), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U7571 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8663), .ZN(n5827) );
  INV_X1 U7572 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8962) );
  XNOR2_X1 U7573 ( .A(n8663), .B(n8962), .ZN(n8654) );
  INV_X1 U7574 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5806) );
  NAND2_X1 U7575 ( .A1(n7587), .A2(n5809), .ZN(n5808) );
  NAND2_X1 U7576 ( .A1(n7579), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7577 ( .A1(n7492), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5811) );
  NAND2_X1 U7578 ( .A1(n7468), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7579 ( .A1(n5812), .A2(n7345), .ZN(n5813) );
  INV_X1 U7580 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n5971) );
  MUX2_X1 U7581 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n5971), .S(n7348), .Z(n8622)
         );
  NAND2_X1 U7582 ( .A1(n7348), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5815) );
  INV_X1 U7583 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5995) );
  MUX2_X1 U7584 ( .A(n5995), .B(P2_REG1_REG_6__SCAN_IN), .S(n6000), .Z(n7612)
         );
  NAND2_X1 U7585 ( .A1(n7614), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5818) );
  NAND2_X1 U7586 ( .A1(n7509), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U7587 ( .A1(n5819), .A2(n4742), .ZN(n5820) );
  INV_X1 U7588 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6009) );
  MUX2_X1 U7589 ( .A(n6009), .B(P2_REG1_REG_8__SCAN_IN), .S(n7679), .Z(n7686)
         );
  NAND2_X1 U7590 ( .A1(n5771), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5822) );
  XNOR2_X1 U7591 ( .A(n7777), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7778) );
  INV_X1 U7592 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8214) );
  INV_X1 U7593 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8088) );
  XNOR2_X1 U7594 ( .A(n7961), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n7962) );
  INV_X1 U7595 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8966) );
  NAND2_X1 U7596 ( .A1(n8678), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U7597 ( .A1(n8720), .A2(n5830), .ZN(n5831) );
  XNOR2_X1 U7598 ( .A(n8744), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8729) );
  XNOR2_X1 U7599 ( .A(n8019), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5899) );
  XNOR2_X1 U7600 ( .A(n5832), .B(n5899), .ZN(n5833) );
  NAND2_X1 U7601 ( .A1(n5833), .A2(n8723), .ZN(n5913) );
  MUX2_X1 U7602 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5838), .Z(n5836) );
  XNOR2_X1 U7603 ( .A(n5836), .B(n5834), .ZN(n7578) );
  INV_X1 U7604 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5835) );
  MUX2_X1 U7605 ( .A(n5937), .B(n5835), .S(n5838), .Z(n7457) );
  NAND2_X1 U7606 ( .A1(n7457), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U7607 ( .A1(n5836), .A2(n7587), .ZN(n5837) );
  MUX2_X1 U7608 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n7032), .Z(n5840) );
  XNOR2_X1 U7609 ( .A(n5839), .B(n5840), .ZN(n7482) );
  NAND2_X1 U7610 ( .A1(n7481), .A2(n7482), .ZN(n5842) );
  NAND2_X1 U7611 ( .A1(n5840), .A2(n7492), .ZN(n5841) );
  NAND2_X1 U7612 ( .A1(n5842), .A2(n5841), .ZN(n7465) );
  MUX2_X1 U7613 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5895), .Z(n5843) );
  XNOR2_X1 U7614 ( .A(n5843), .B(n7345), .ZN(n7466) );
  MUX2_X1 U7615 ( .A(n10106), .B(n5971), .S(n5895), .Z(n5846) );
  XNOR2_X1 U7616 ( .A(n5846), .B(n7348), .ZN(n8628) );
  INV_X1 U7617 ( .A(n5843), .ZN(n5844) );
  NAND2_X1 U7618 ( .A1(n5844), .A2(n7473), .ZN(n8625) );
  AND2_X1 U7619 ( .A1(n8628), .A2(n8625), .ZN(n5845) );
  NAND2_X1 U7620 ( .A1(n8626), .A2(n5845), .ZN(n8627) );
  INV_X1 U7621 ( .A(n5846), .ZN(n5847) );
  NAND2_X1 U7622 ( .A1(n5847), .A2(n7348), .ZN(n5848) );
  NAND2_X1 U7623 ( .A1(n8627), .A2(n5848), .ZN(n7497) );
  MUX2_X1 U7624 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n5895), .Z(n5849) );
  XNOR2_X1 U7625 ( .A(n5849), .B(n5987), .ZN(n7496) );
  NAND2_X1 U7626 ( .A1(n7497), .A2(n7496), .ZN(n5851) );
  NAND2_X1 U7627 ( .A1(n5849), .A2(n7503), .ZN(n5850) );
  NAND2_X1 U7628 ( .A1(n5851), .A2(n5850), .ZN(n7608) );
  MUX2_X1 U7629 ( .A(n10286), .B(n5995), .S(n5895), .Z(n5852) );
  NAND2_X1 U7630 ( .A1(n5852), .A2(n6000), .ZN(n7513) );
  INV_X1 U7631 ( .A(n5852), .ZN(n5853) );
  NAND2_X1 U7632 ( .A1(n5853), .A2(n7614), .ZN(n5854) );
  NAND2_X1 U7633 ( .A1(n7513), .A2(n5854), .ZN(n7609) );
  NAND2_X1 U7634 ( .A1(n7512), .A2(n7513), .ZN(n5858) );
  INV_X1 U7635 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7508) );
  MUX2_X1 U7636 ( .A(n7510), .B(n7508), .S(n5895), .Z(n5855) );
  NAND2_X1 U7637 ( .A1(n5855), .A2(n6014), .ZN(n7676) );
  INV_X1 U7638 ( .A(n5855), .ZN(n5856) );
  NAND2_X1 U7639 ( .A1(n5856), .A2(n4742), .ZN(n5857) );
  AND2_X1 U7640 ( .A1(n7676), .A2(n5857), .ZN(n7514) );
  NAND2_X1 U7641 ( .A1(n7677), .A2(n7676), .ZN(n5862) );
  MUX2_X1 U7642 ( .A(n7996), .B(n6009), .S(n5895), .Z(n5859) );
  NAND2_X1 U7643 ( .A1(n5859), .A2(n7679), .ZN(n7695) );
  INV_X1 U7644 ( .A(n5859), .ZN(n5860) );
  NAND2_X1 U7645 ( .A1(n5860), .A2(n5771), .ZN(n5861) );
  AND2_X1 U7646 ( .A1(n7695), .A2(n5861), .ZN(n7674) );
  NAND2_X1 U7647 ( .A1(n7696), .A2(n7695), .ZN(n5866) );
  INV_X1 U7648 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7985) );
  INV_X1 U7649 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7690) );
  MUX2_X1 U7650 ( .A(n7985), .B(n7690), .S(n5895), .Z(n5863) );
  NAND2_X1 U7651 ( .A1(n5863), .A2(n6035), .ZN(n7772) );
  INV_X1 U7652 ( .A(n5863), .ZN(n5864) );
  NAND2_X1 U7653 ( .A1(n5864), .A2(n7699), .ZN(n5865) );
  AND2_X1 U7654 ( .A1(n7772), .A2(n5865), .ZN(n7693) );
  NAND2_X1 U7655 ( .A1(n7773), .A2(n7772), .ZN(n5870) );
  MUX2_X1 U7656 ( .A(n5779), .B(n8214), .S(n5895), .Z(n5867) );
  NAND2_X1 U7657 ( .A1(n5867), .A2(n7777), .ZN(n7906) );
  INV_X1 U7658 ( .A(n5867), .ZN(n5868) );
  INV_X1 U7659 ( .A(n7777), .ZN(n7398) );
  NAND2_X1 U7660 ( .A1(n5868), .A2(n7398), .ZN(n5869) );
  AND2_X1 U7661 ( .A1(n7906), .A2(n5869), .ZN(n7770) );
  NAND2_X1 U7662 ( .A1(n7907), .A2(n7906), .ZN(n5873) );
  INV_X1 U7663 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8083) );
  MUX2_X1 U7664 ( .A(n8083), .B(n8088), .S(n5895), .Z(n5871) );
  OR2_X1 U7665 ( .A1(n6048), .A2(n5871), .ZN(n5872) );
  NAND2_X1 U7666 ( .A1(n5871), .A2(n6048), .ZN(n7956) );
  AND2_X1 U7667 ( .A1(n5872), .A2(n7956), .ZN(n7904) );
  NAND2_X1 U7668 ( .A1(n5873), .A2(n7904), .ZN(n7957) );
  NAND2_X1 U7669 ( .A1(n7957), .A2(n7956), .ZN(n5876) );
  INV_X1 U7670 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8973) );
  MUX2_X1 U7671 ( .A(n5786), .B(n8973), .S(n5895), .Z(n5874) );
  OR2_X1 U7672 ( .A1(n7961), .A2(n5874), .ZN(n5875) );
  NAND2_X1 U7673 ( .A1(n7961), .A2(n5874), .ZN(n8639) );
  AND2_X1 U7674 ( .A1(n5875), .A2(n8639), .ZN(n7954) );
  NAND2_X1 U7675 ( .A1(n8640), .A2(n8639), .ZN(n5879) );
  MUX2_X1 U7676 ( .A(n8323), .B(n8966), .S(n5895), .Z(n5877) );
  NAND2_X1 U7677 ( .A1(n7543), .A2(n5877), .ZN(n8658) );
  OR2_X1 U7678 ( .A1(n7543), .A2(n5877), .ZN(n5878) );
  AND2_X1 U7679 ( .A1(n8658), .A2(n5878), .ZN(n8637) );
  NAND2_X1 U7680 ( .A1(n8659), .A2(n8658), .ZN(n5884) );
  INV_X1 U7681 ( .A(n8663), .ZN(n5880) );
  MUX2_X1 U7682 ( .A(n6085), .B(n8962), .S(n5895), .Z(n5881) );
  NAND2_X1 U7683 ( .A1(n5880), .A2(n5881), .ZN(n8673) );
  INV_X1 U7684 ( .A(n5881), .ZN(n5882) );
  NAND2_X1 U7685 ( .A1(n8663), .A2(n5882), .ZN(n5883) );
  AND2_X1 U7686 ( .A1(n8673), .A2(n5883), .ZN(n8656) );
  NAND2_X1 U7687 ( .A1(n8674), .A2(n8673), .ZN(n5887) );
  MUX2_X1 U7688 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5895), .Z(n5885) );
  OR2_X1 U7689 ( .A1(n8678), .A2(n5885), .ZN(n8692) );
  NAND2_X1 U7690 ( .A1(n8678), .A2(n5885), .ZN(n5886) );
  AND2_X1 U7691 ( .A1(n8692), .A2(n5886), .ZN(n8671) );
  NAND2_X1 U7692 ( .A1(n8693), .A2(n8692), .ZN(n5890) );
  MUX2_X1 U7693 ( .A(n10277), .B(n8954), .S(n5895), .Z(n5888) );
  NAND2_X1 U7694 ( .A1(n7743), .A2(n5888), .ZN(n5891) );
  OR2_X1 U7695 ( .A1(n7743), .A2(n5888), .ZN(n5889) );
  AND2_X1 U7696 ( .A1(n5891), .A2(n5889), .ZN(n8690) );
  NAND2_X1 U7697 ( .A1(n5890), .A2(n8690), .ZN(n8696) );
  NAND2_X1 U7698 ( .A1(n8696), .A2(n5891), .ZN(n8714) );
  INV_X1 U7699 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8876) );
  INV_X1 U7700 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n6117) );
  MUX2_X1 U7701 ( .A(n8876), .B(n6117), .S(n5895), .Z(n5892) );
  XNOR2_X1 U7702 ( .A(n8720), .B(n5892), .ZN(n8713) );
  NAND2_X1 U7703 ( .A1(n8714), .A2(n8713), .ZN(n8712) );
  INV_X1 U7704 ( .A(n5892), .ZN(n5893) );
  OR2_X1 U7705 ( .A1(n8720), .A2(n5893), .ZN(n5894) );
  NAND2_X1 U7706 ( .A1(n8712), .A2(n5894), .ZN(n5897) );
  INV_X1 U7707 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8945) );
  MUX2_X1 U7708 ( .A(n8865), .B(n8945), .S(n5895), .Z(n5896) );
  NAND2_X1 U7709 ( .A1(n5897), .A2(n5896), .ZN(n8737) );
  NOR2_X1 U7710 ( .A1(n5897), .A2(n5896), .ZN(n8739) );
  AOI21_X1 U7711 ( .B1(n7948), .B2(n8737), .A(n8739), .ZN(n5901) );
  MUX2_X1 U7712 ( .A(n5899), .B(n5898), .S(n6308), .Z(n5900) );
  XNOR2_X1 U7713 ( .A(n5901), .B(n5900), .ZN(n5910) );
  NAND2_X1 U7714 ( .A1(P2_U3893), .A2(n5804), .ZN(n8694) );
  NOR2_X1 U7715 ( .A1(n5895), .A2(P2_U3151), .ZN(n9090) );
  NAND2_X1 U7716 ( .A1(n5902), .A2(n9090), .ZN(n5903) );
  MUX2_X1 U7717 ( .A(n8614), .B(n5903), .S(n5804), .Z(n8721) );
  NOR2_X1 U7718 ( .A1(n8721), .A2(n8019), .ZN(n5908) );
  INV_X1 U7719 ( .A(n6500), .ZN(n5904) );
  NOR2_X1 U7720 ( .A1(n6492), .A2(n5904), .ZN(n5905) );
  NAND2_X1 U7721 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8467) );
  OAI21_X1 U7722 ( .B1(n7953), .B2(n5906), .A(n8467), .ZN(n5907) );
  INV_X1 U7723 ( .A(n5911), .ZN(n5912) );
  INV_X1 U7724 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5921) );
  OAI21_X1 U7725 ( .B1(n6784), .B2(n5915), .A(n6375), .ZN(n5916) );
  OAI22_X1 U7726 ( .A1(n8404), .A2(n9336), .B1(n6540), .B2(n9337), .ZN(n7295)
         );
  XNOR2_X1 U7727 ( .A(n5917), .B(n6784), .ZN(n9583) );
  OAI211_X1 U7728 ( .C1(n9908), .C2(n9598), .A(n9764), .B(n6379), .ZN(n9584)
         );
  NAND2_X1 U7729 ( .A1(n10073), .A2(n10064), .ZN(n9902) );
  XNOR2_X2 U7730 ( .A(n5925), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7731 ( .A1(n5926), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5934) );
  AND2_X4 U7732 ( .A1(n5927), .A2(n9084), .ZN(n5958) );
  INV_X1 U7733 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7733) );
  OR2_X1 U7734 ( .A1(n5957), .A2(n7733), .ZN(n5933) );
  OR2_X1 U7735 ( .A1(n5950), .A2(n5931), .ZN(n5932) );
  INV_X1 U7736 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7354) );
  INV_X1 U7737 ( .A(n7454), .ZN(n5935) );
  NAND2_X1 U7738 ( .A1(n5958), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5940) );
  INV_X1 U7739 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7461) );
  OR2_X1 U7740 ( .A1(n5957), .A2(n7461), .ZN(n5939) );
  OR2_X1 U7741 ( .A1(n5950), .A2(n5937), .ZN(n5938) );
  INV_X1 U7742 ( .A(SI_0_), .ZN(n5942) );
  INV_X1 U7743 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U7744 ( .B1(n4292), .B2(n5942), .A(n5941), .ZN(n5944) );
  AND2_X1 U7745 ( .A1(n5944), .A2(n5943), .ZN(n9100) );
  MUX2_X1 U7746 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9100), .S(n6316), .Z(n7530) );
  NAND2_X1 U7747 ( .A1(n7737), .A2(n7530), .ZN(n7730) );
  INV_X1 U7748 ( .A(n7730), .ZN(n5945) );
  NAND2_X1 U7749 ( .A1(n7732), .A2(n6837), .ZN(n7625) );
  NAND2_X1 U7750 ( .A1(n5958), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5947) );
  INV_X1 U7751 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7631) );
  OR2_X1 U7752 ( .A1(n5957), .A2(n7631), .ZN(n5946) );
  NAND2_X1 U7753 ( .A1(n5947), .A2(n5946), .ZN(n5948) );
  INV_X1 U7754 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7634) );
  OR2_X1 U7755 ( .A1(n6966), .A2(n7634), .ZN(n5951) );
  INV_X1 U7756 ( .A(n5953), .ZN(n7357) );
  OR2_X1 U7757 ( .A1(n6229), .A2(n7357), .ZN(n5954) );
  INV_X1 U7758 ( .A(n10118), .ZN(n7630) );
  NAND2_X1 U7759 ( .A1(n7625), .A2(n7627), .ZN(n5956) );
  NAND2_X1 U7760 ( .A1(n5956), .A2(n6843), .ZN(n7640) );
  OR2_X1 U7761 ( .A1(n5957), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5962) );
  INV_X1 U7762 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10158) );
  OR2_X1 U7763 ( .A1(n6969), .A2(n10158), .ZN(n5961) );
  INV_X1 U7764 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5959) );
  OR2_X1 U7765 ( .A1(n6097), .A2(n5959), .ZN(n5960) );
  AND4_X2 U7766 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n7629)
         );
  INV_X1 U7767 ( .A(n5964), .ZN(n7346) );
  OR2_X1 U7768 ( .A1(n7346), .A2(n6229), .ZN(n5966) );
  OR2_X1 U7769 ( .A1(n6976), .A2(n5072), .ZN(n5965) );
  OAI211_X1 U7770 ( .C1(n6316), .C2(n7345), .A(n5966), .B(n5965), .ZN(n7645)
         );
  INV_X1 U7771 ( .A(n7645), .ZN(n10121) );
  XNOR2_X1 U7772 ( .A(n7629), .B(n10121), .ZN(n7641) );
  NAND2_X1 U7773 ( .A1(n7640), .A2(n7641), .ZN(n5967) );
  NAND2_X1 U7774 ( .A1(n5967), .A2(n6850), .ZN(n10099) );
  NAND2_X1 U7775 ( .A1(n5958), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5975) );
  OR2_X1 U7776 ( .A1(n6966), .A2(n10106), .ZN(n5974) );
  INV_X2 U7777 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7778 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5970) );
  AND2_X1 U7779 ( .A1(n5980), .A2(n5970), .ZN(n10100) );
  OR2_X1 U7780 ( .A1(n5957), .A2(n10100), .ZN(n5973) );
  OR2_X1 U7781 ( .A1(n6969), .A2(n5971), .ZN(n5972) );
  NAND2_X1 U7782 ( .A1(n5988), .A2(n7347), .ZN(n5977) );
  OR2_X1 U7783 ( .A1(n6976), .A2(n7349), .ZN(n5976) );
  OAI211_X1 U7784 ( .C1(n6316), .C2(n7348), .A(n5977), .B(n5976), .ZN(n10124)
         );
  OR2_X1 U7785 ( .A1(n7533), .A2(n7654), .ZN(n6252) );
  NAND2_X1 U7786 ( .A1(n7533), .A2(n7654), .ZN(n6251) );
  NAND2_X1 U7787 ( .A1(n6252), .A2(n6251), .ZN(n10098) );
  NAND2_X1 U7788 ( .A1(n7533), .A2(n10124), .ZN(n6859) );
  NAND2_X1 U7789 ( .A1(n6211), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5986) );
  INV_X1 U7790 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5978) );
  OR2_X1 U7791 ( .A1(n6097), .A2(n5978), .ZN(n5985) );
  NAND2_X1 U7792 ( .A1(n5980), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5981) );
  AND2_X1 U7793 ( .A1(n5993), .A2(n5981), .ZN(n7801) );
  OR2_X1 U7794 ( .A1(n5957), .A2(n7801), .ZN(n5984) );
  INV_X1 U7795 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5982) );
  OR2_X1 U7796 ( .A1(n6969), .A2(n5982), .ZN(n5983) );
  NAND4_X1 U7797 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n10092)
         );
  AOI22_X1 U7798 ( .A1(n6127), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n4607), .B2(
        n5987), .ZN(n5990) );
  NAND2_X1 U7799 ( .A1(n7358), .A2(n5988), .ZN(n5989) );
  NAND2_X1 U7800 ( .A1(n5990), .A2(n5989), .ZN(n10129) );
  NOR2_X1 U7801 ( .A1(n10092), .A2(n7725), .ZN(n6858) );
  INV_X1 U7802 ( .A(n6858), .ZN(n5991) );
  NAND2_X1 U7803 ( .A1(n10092), .A2(n7725), .ZN(n6862) );
  NAND2_X1 U7804 ( .A1(n6211), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5999) );
  INV_X1 U7805 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5992) );
  OR2_X1 U7806 ( .A1(n6097), .A2(n5992), .ZN(n5998) );
  NAND2_X1 U7807 ( .A1(n5993), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5994) );
  AND2_X1 U7808 ( .A1(n6017), .A2(n5994), .ZN(n7788) );
  OR2_X1 U7809 ( .A1(n5957), .A2(n7788), .ZN(n5997) );
  OR2_X1 U7810 ( .A1(n6969), .A2(n5995), .ZN(n5996) );
  INV_X1 U7811 ( .A(n10079), .ZN(n7724) );
  NAND2_X1 U7812 ( .A1(n7369), .A2(n5988), .ZN(n6002) );
  AOI22_X1 U7813 ( .A1(n6127), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n4607), .B2(
        n6000), .ZN(n6001) );
  NAND2_X1 U7814 ( .A1(n7724), .A2(n7790), .ZN(n7989) );
  INV_X1 U7815 ( .A(n7790), .ZN(n10136) );
  NAND2_X1 U7816 ( .A1(n10136), .A2(n10079), .ZN(n6863) );
  NAND2_X1 U7817 ( .A1(n7989), .A2(n6863), .ZN(n7786) );
  NAND2_X1 U7818 ( .A1(n7378), .A2(n5988), .ZN(n6005) );
  AOI22_X1 U7819 ( .A1(n6127), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n4607), .B2(
        n7679), .ZN(n6004) );
  NAND2_X1 U7820 ( .A1(n6005), .A2(n6004), .ZN(n10150) );
  NAND2_X1 U7821 ( .A1(n5958), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6013) );
  OR2_X1 U7822 ( .A1(n6966), .A2(n7996), .ZN(n6012) );
  NAND2_X1 U7823 ( .A1(n6019), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6008) );
  AND2_X1 U7824 ( .A1(n6039), .A2(n6008), .ZN(n8105) );
  OR2_X1 U7825 ( .A1(n5957), .A2(n8105), .ZN(n6011) );
  OR2_X1 U7826 ( .A1(n6969), .A2(n6009), .ZN(n6010) );
  NAND2_X1 U7827 ( .A1(n10150), .A2(n8033), .ZN(n7006) );
  NAND2_X1 U7828 ( .A1(n7373), .A2(n5988), .ZN(n6016) );
  AOI22_X1 U7829 ( .A1(n6127), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n4607), .B2(
        n6014), .ZN(n6015) );
  NAND2_X1 U7830 ( .A1(n6016), .A2(n6015), .ZN(n10140) );
  NAND2_X1 U7831 ( .A1(n5958), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6023) );
  NAND2_X1 U7832 ( .A1(n6017), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6018) );
  AND2_X1 U7833 ( .A1(n6019), .A2(n6018), .ZN(n7873) );
  OR2_X1 U7834 ( .A1(n5957), .A2(n7873), .ZN(n6022) );
  OR2_X1 U7835 ( .A1(n6969), .A2(n7508), .ZN(n6021) );
  OR2_X1 U7836 ( .A1(n6966), .A2(n7510), .ZN(n6020) );
  NAND2_X1 U7837 ( .A1(n10140), .A2(n8102), .ZN(n6874) );
  AND3_X1 U7838 ( .A1(n7006), .A2(n6874), .A3(n7989), .ZN(n6024) );
  NAND2_X1 U7839 ( .A1(n7990), .A2(n6024), .ZN(n7969) );
  NAND2_X1 U7840 ( .A1(n7396), .A2(n5988), .ZN(n6026) );
  AOI22_X1 U7841 ( .A1(n6127), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n4607), .B2(
        n7777), .ZN(n6025) );
  NAND2_X1 U7842 ( .A1(n5958), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6033) );
  OR2_X1 U7843 ( .A1(n6966), .A2(n5779), .ZN(n6032) );
  NAND2_X1 U7844 ( .A1(n6028), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6029) );
  AND2_X1 U7845 ( .A1(n6051), .A2(n6029), .ZN(n8458) );
  OR2_X1 U7846 ( .A1(n5957), .A2(n8458), .ZN(n6031) );
  OR2_X1 U7847 ( .A1(n6969), .A2(n8214), .ZN(n6030) );
  OR2_X1 U7848 ( .A1(n10150), .A2(n8033), .ZN(n7007) );
  OR2_X1 U7849 ( .A1(n10140), .A2(n8102), .ZN(n7991) );
  NAND2_X1 U7850 ( .A1(n7007), .A2(n7991), .ZN(n6034) );
  NAND2_X1 U7851 ( .A1(n6034), .A2(n7006), .ZN(n7968) );
  NAND2_X1 U7852 ( .A1(n7393), .A2(n5988), .ZN(n6037) );
  AOI22_X1 U7853 ( .A1(n6127), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n4607), .B2(
        n6035), .ZN(n6036) );
  NAND2_X1 U7854 ( .A1(n6211), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6043) );
  INV_X1 U7855 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7856 ( .A1(n6097), .A2(n6038), .ZN(n6042) );
  XNOR2_X1 U7857 ( .A(n6039), .B(n10300), .ZN(n8034) );
  OR2_X1 U7858 ( .A1(n5957), .A2(n8034), .ZN(n6041) );
  OR2_X1 U7859 ( .A1(n6969), .A2(n7690), .ZN(n6040) );
  NAND4_X1 U7860 ( .A1(n6043), .A2(n6042), .A3(n6041), .A4(n6040), .ZN(n8610)
         );
  INV_X2 U7861 ( .A(n8610), .ZN(n8055) );
  NAND2_X1 U7862 ( .A1(n7969), .A2(n4982), .ZN(n6047) );
  INV_X1 U7863 ( .A(n7004), .ZN(n6044) );
  NAND2_X1 U7864 ( .A1(n8976), .A2(n8055), .ZN(n7005) );
  NAND2_X1 U7865 ( .A1(n8460), .A2(n8551), .ZN(n7003) );
  NAND2_X1 U7866 ( .A1(n6047), .A2(n6046), .ZN(n8076) );
  NAND2_X1 U7867 ( .A1(n7418), .A2(n5988), .ZN(n6050) );
  AOI22_X1 U7868 ( .A1(n6127), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6048), .B2(
        n4607), .ZN(n6049) );
  NAND2_X1 U7869 ( .A1(n6211), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6056) );
  INV_X1 U7870 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8080) );
  OR2_X1 U7871 ( .A1(n6097), .A2(n8080), .ZN(n6055) );
  NAND2_X1 U7872 ( .A1(n6051), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6052) );
  AND2_X1 U7873 ( .A1(n6062), .A2(n6052), .ZN(n8561) );
  OR2_X1 U7874 ( .A1(n5957), .A2(n8561), .ZN(n6054) );
  OR2_X1 U7875 ( .A1(n6969), .A2(n8088), .ZN(n6053) );
  OR2_X1 U7876 ( .A1(n8563), .A2(n8455), .ZN(n6884) );
  NAND2_X1 U7877 ( .A1(n8563), .A2(n8455), .ZN(n6885) );
  NAND2_X1 U7878 ( .A1(n6884), .A2(n6885), .ZN(n8075) );
  INV_X1 U7879 ( .A(n8075), .ZN(n8078) );
  INV_X1 U7880 ( .A(n6885), .ZN(n6057) );
  NAND2_X1 U7881 ( .A1(n7422), .A2(n5988), .ZN(n6059) );
  AOI22_X1 U7882 ( .A1(n7961), .A2(n4607), .B1(n6127), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7883 ( .A1(n5958), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6067) );
  OR2_X1 U7884 ( .A1(n6969), .A2(n8973), .ZN(n6066) );
  NAND2_X1 U7885 ( .A1(n6062), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6063) );
  AND2_X1 U7886 ( .A1(n6073), .A2(n6063), .ZN(n8196) );
  OR2_X1 U7887 ( .A1(n5957), .A2(n8196), .ZN(n6065) );
  OR2_X1 U7888 ( .A1(n6966), .A2(n5786), .ZN(n6064) );
  NAND4_X1 U7889 ( .A1(n6067), .A2(n6066), .A3(n6065), .A4(n6064), .ZN(n8607)
         );
  XNOR2_X1 U7890 ( .A(n8972), .B(n8607), .ZN(n8193) );
  INV_X1 U7891 ( .A(n8607), .ZN(n8557) );
  OR2_X1 U7892 ( .A1(n8972), .A2(n8557), .ZN(n6068) );
  NAND2_X1 U7893 ( .A1(n7541), .A2(n5988), .ZN(n6070) );
  AOI22_X1 U7894 ( .A1(n7543), .A2(n4607), .B1(n6127), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7895 ( .A1(n5958), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6078) );
  OR2_X1 U7896 ( .A1(n6966), .A2(n8323), .ZN(n6077) );
  NAND2_X1 U7897 ( .A1(n6073), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6074) );
  AND2_X1 U7898 ( .A1(n6083), .A2(n6074), .ZN(n8316) );
  OR2_X1 U7899 ( .A1(n5957), .A2(n8316), .ZN(n6076) );
  OR2_X1 U7900 ( .A1(n6969), .A2(n8966), .ZN(n6075) );
  NAND4_X1 U7901 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n8910)
         );
  INV_X1 U7902 ( .A(n8910), .ZN(n8442) );
  NAND2_X1 U7903 ( .A1(n9065), .A2(n8442), .ZN(n6079) );
  NAND2_X1 U7904 ( .A1(n7636), .A2(n5988), .ZN(n6082) );
  INV_X1 U7905 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7637) );
  OAI22_X1 U7906 ( .A1(n8663), .A2(n6316), .B1(n6976), .B2(n7637), .ZN(n6080)
         );
  INV_X1 U7907 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U7908 ( .A1(n6083), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7909 ( .A1(n6094), .A2(n6084), .ZN(n8912) );
  NAND2_X1 U7910 ( .A1(n6231), .A2(n8912), .ZN(n6089) );
  OR2_X1 U7911 ( .A1(n6966), .A2(n6085), .ZN(n6088) );
  INV_X1 U7912 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9058) );
  OR2_X1 U7913 ( .A1(n6097), .A2(n9058), .ZN(n6087) );
  OR2_X1 U7914 ( .A1(n6969), .A2(n8962), .ZN(n6086) );
  NAND4_X1 U7915 ( .A1(n6089), .A2(n6088), .A3(n6087), .A4(n6086), .ZN(n8606)
         );
  NAND2_X1 U7916 ( .A1(n9059), .A2(n8897), .ZN(n6900) );
  NAND2_X1 U7917 ( .A1(n8905), .A2(n6900), .ZN(n6090) );
  NAND2_X1 U7918 ( .A1(n6090), .A2(n6901), .ZN(n8890) );
  NAND2_X1 U7919 ( .A1(n7705), .A2(n5988), .ZN(n6093) );
  INV_X1 U7920 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7708) );
  OAI22_X1 U7921 ( .A1(n8678), .A2(n6316), .B1(n6976), .B2(n7708), .ZN(n6091)
         );
  INV_X1 U7922 ( .A(n6091), .ZN(n6092) );
  INV_X1 U7923 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U7924 ( .A1(n6094), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6095) );
  NAND2_X1 U7925 ( .A1(n6104), .A2(n6095), .ZN(n8899) );
  NAND2_X1 U7926 ( .A1(n8899), .A2(n6231), .ZN(n6101) );
  INV_X1 U7927 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6096) );
  OR2_X1 U7928 ( .A1(n6966), .A2(n6096), .ZN(n6099) );
  INV_X1 U7929 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9053) );
  OR2_X1 U7930 ( .A1(n6097), .A2(n9053), .ZN(n6098) );
  AND2_X1 U7931 ( .A1(n6099), .A2(n6098), .ZN(n6100) );
  OAI211_X1 U7932 ( .C1(n6969), .C2(n8959), .A(n6101), .B(n6100), .ZN(n8909)
         );
  INV_X1 U7933 ( .A(n8909), .ZN(n8510) );
  NAND2_X1 U7934 ( .A1(n8590), .A2(n8510), .ZN(n6910) );
  NAND2_X1 U7935 ( .A1(n7741), .A2(n5988), .ZN(n6103) );
  AOI22_X1 U7936 ( .A1(n7743), .A2(n4607), .B1(n6127), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7937 ( .A1(n6104), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7938 ( .A1(n6113), .A2(n6105), .ZN(n8887) );
  NAND2_X1 U7939 ( .A1(n8887), .A2(n6231), .ZN(n6107) );
  AOI22_X1 U7940 ( .A1(n6211), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n5958), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6106) );
  OAI211_X1 U7941 ( .C1(n6969), .C2(n8954), .A(n6107), .B(n6106), .ZN(n8870)
         );
  INV_X1 U7942 ( .A(n8870), .ZN(n8895) );
  OR2_X1 U7943 ( .A1(n9048), .A2(n8895), .ZN(n6912) );
  NAND2_X1 U7944 ( .A1(n9048), .A2(n8895), .ZN(n6905) );
  NAND2_X1 U7945 ( .A1(n6912), .A2(n6905), .ZN(n8883) );
  NAND2_X1 U7946 ( .A1(n7866), .A2(n5988), .ZN(n6110) );
  OAI22_X1 U7947 ( .A1(n8720), .A2(n6316), .B1(n6976), .B2(n10253), .ZN(n6108)
         );
  INV_X1 U7948 ( .A(n6108), .ZN(n6109) );
  NAND2_X1 U7949 ( .A1(n6113), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6114) );
  NAND2_X1 U7950 ( .A1(n6120), .A2(n6114), .ZN(n8873) );
  NAND2_X1 U7951 ( .A1(n8873), .A2(n6231), .ZN(n6116) );
  AOI22_X1 U7952 ( .A1(n6211), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n5958), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6115) );
  OAI211_X1 U7953 ( .C1(n6969), .C2(n6117), .A(n6116), .B(n6115), .ZN(n8885)
         );
  INV_X1 U7954 ( .A(n8885), .ZN(n8568) );
  NAND2_X1 U7955 ( .A1(n8948), .A2(n8568), .ZN(n6906) );
  NAND2_X1 U7956 ( .A1(n8859), .A2(n6906), .ZN(n8878) );
  NAND2_X1 U7957 ( .A1(n7924), .A2(n5988), .ZN(n6119) );
  AOI22_X1 U7958 ( .A1(n6127), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n4607), .B2(
        n8744), .ZN(n6118) );
  NAND2_X1 U7959 ( .A1(n6120), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7960 ( .A1(n6130), .A2(n6121), .ZN(n8866) );
  NAND2_X1 U7961 ( .A1(n8866), .A2(n6231), .ZN(n6126) );
  NAND2_X1 U7962 ( .A1(n6211), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U7963 ( .A1(n5958), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6122) );
  OAI211_X1 U7964 ( .C1(n8945), .C2(n6969), .A(n6123), .B(n6122), .ZN(n6124)
         );
  INV_X1 U7965 ( .A(n6124), .ZN(n6125) );
  OR2_X1 U7966 ( .A1(n9041), .A2(n8469), .ZN(n8858) );
  AND2_X1 U7967 ( .A1(n8858), .A2(n8859), .ZN(n7011) );
  NAND2_X1 U7968 ( .A1(n8018), .A2(n5988), .ZN(n6129) );
  AOI22_X1 U7969 ( .A1(n6127), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7028), .B2(
        n4607), .ZN(n6128) );
  NAND2_X1 U7970 ( .A1(n6130), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7971 ( .A1(n6138), .A2(n6131), .ZN(n8854) );
  INV_X1 U7972 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n6134) );
  NAND2_X1 U7973 ( .A1(n6211), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7974 ( .A1(n5958), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6132) );
  OAI211_X1 U7975 ( .C1(n6134), .C2(n6969), .A(n6133), .B(n6132), .ZN(n6135)
         );
  AOI21_X1 U7976 ( .B1(n8854), .B2(n6231), .A(n6135), .ZN(n8537) );
  NAND2_X1 U7977 ( .A1(n6447), .A2(n8537), .ZN(n6916) );
  NAND2_X1 U7978 ( .A1(n9041), .A2(n8469), .ZN(n8857) );
  AND2_X1 U7979 ( .A1(n6916), .A2(n8857), .ZN(n6835) );
  OR2_X1 U7980 ( .A1(n6447), .A2(n8537), .ZN(n6917) );
  NAND2_X1 U7981 ( .A1(n8186), .A2(n5988), .ZN(n6137) );
  OR2_X1 U7982 ( .A1(n6976), .A2(n8210), .ZN(n6136) );
  NAND2_X1 U7983 ( .A1(n6138), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7984 ( .A1(n6150), .A2(n6139), .ZN(n8840) );
  NAND2_X1 U7985 ( .A1(n8840), .A2(n6231), .ZN(n6144) );
  INV_X1 U7986 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U7987 ( .A1(n6211), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7988 ( .A1(n5958), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6140) );
  OAI211_X1 U7989 ( .C1(n8940), .C2(n6969), .A(n6141), .B(n6140), .ZN(n6142)
         );
  INV_X1 U7990 ( .A(n6142), .ZN(n6143) );
  OR2_X1 U7991 ( .A1(n6976), .A2(n10233), .ZN(n6146) );
  NAND2_X1 U7992 ( .A1(n6150), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6151) );
  NAND2_X1 U7993 ( .A1(n6166), .A2(n6151), .ZN(n8828) );
  INV_X1 U7994 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8937) );
  NAND2_X1 U7995 ( .A1(n6211), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7996 ( .A1(n5958), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7997 ( .C1(n8937), .C2(n6969), .A(n6153), .B(n6152), .ZN(n6154)
         );
  AOI21_X1 U7998 ( .B1(n8828), .B2(n6231), .A(n6154), .ZN(n6456) );
  INV_X1 U7999 ( .A(n6925), .ZN(n6929) );
  NAND2_X1 U8000 ( .A1(n6155), .A2(n5988), .ZN(n6157) );
  OR2_X1 U8001 ( .A1(n6976), .A2(n8347), .ZN(n6156) );
  INV_X1 U8002 ( .A(n6178), .ZN(n6179) );
  NAND2_X1 U8003 ( .A1(n6168), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U8004 ( .A1(n6179), .A2(n6158), .ZN(n8806) );
  NAND2_X1 U8005 ( .A1(n8806), .A2(n6231), .ZN(n6163) );
  INV_X1 U8006 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U8007 ( .A1(n6211), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U8008 ( .A1(n5958), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U8009 ( .C1(n8931), .C2(n6969), .A(n6160), .B(n6159), .ZN(n6161)
         );
  INV_X1 U8010 ( .A(n6161), .ZN(n6162) );
  OR2_X1 U8011 ( .A1(n9013), .A2(n8788), .ZN(n6950) );
  NAND2_X1 U8012 ( .A1(n8339), .A2(n5988), .ZN(n6165) );
  OR2_X1 U8013 ( .A1(n6976), .A2(n8344), .ZN(n6164) );
  NAND2_X1 U8014 ( .A1(n6166), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U8015 ( .A1(n6168), .A2(n6167), .ZN(n8815) );
  NAND2_X1 U8016 ( .A1(n8815), .A2(n6231), .ZN(n6173) );
  INV_X1 U8017 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8934) );
  NAND2_X1 U8018 ( .A1(n6211), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U8019 ( .A1(n5958), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6169) );
  OAI211_X1 U8020 ( .C1(n8934), .C2(n6969), .A(n6170), .B(n6169), .ZN(n6171)
         );
  INV_X1 U8021 ( .A(n6171), .ZN(n6172) );
  NAND2_X1 U8022 ( .A1(n6950), .A2(n8790), .ZN(n6932) );
  NAND2_X1 U8023 ( .A1(n9019), .A2(n8496), .ZN(n6283) );
  NAND2_X1 U8024 ( .A1(n6283), .A2(n8812), .ZN(n6174) );
  INV_X1 U8025 ( .A(n6283), .ZN(n8791) );
  AOI22_X1 U8026 ( .A1(n9013), .A2(n6174), .B1(n8791), .B2(n8788), .ZN(n6186)
         );
  NAND2_X1 U8027 ( .A1(n8372), .A2(n5988), .ZN(n6176) );
  OR2_X1 U8028 ( .A1(n6976), .A2(n8375), .ZN(n6175) );
  INV_X1 U8029 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U8030 ( .A1(n6179), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U8031 ( .A1(n6189), .A2(n6180), .ZN(n8789) );
  NAND2_X1 U8032 ( .A1(n8789), .A2(n6231), .ZN(n6185) );
  INV_X1 U8033 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U8034 ( .A1(n6211), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U8035 ( .A1(n5958), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6181) );
  OAI211_X1 U8036 ( .C1(n10222), .C2(n6969), .A(n6182), .B(n6181), .ZN(n6183)
         );
  INV_X1 U8037 ( .A(n6183), .ZN(n6184) );
  NAND2_X1 U8038 ( .A1(n9007), .A2(n8526), .ZN(n6995) );
  NAND2_X1 U8039 ( .A1(n8377), .A2(n5988), .ZN(n6188) );
  OR2_X1 U8040 ( .A1(n6976), .A2(n9098), .ZN(n6187) );
  NAND2_X1 U8041 ( .A1(n6189), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U8042 ( .A1(n6199), .A2(n6190), .ZN(n8779) );
  NAND2_X1 U8043 ( .A1(n8779), .A2(n6231), .ZN(n6195) );
  INV_X1 U8044 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U8045 ( .A1(n6211), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U8046 ( .A1(n5958), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6191) );
  OAI211_X1 U8047 ( .C1(n8925), .C2(n6969), .A(n6192), .B(n6191), .ZN(n6193)
         );
  INV_X1 U8048 ( .A(n6193), .ZN(n6194) );
  INV_X1 U8049 ( .A(n6938), .ZN(n6196) );
  NAND2_X1 U8050 ( .A1(n9001), .A2(n6469), .ZN(n6952) );
  NAND2_X1 U8051 ( .A1(n9094), .A2(n5988), .ZN(n6198) );
  OR2_X1 U8052 ( .A1(n6976), .A2(n9095), .ZN(n6197) );
  NAND2_X1 U8053 ( .A1(n6199), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U8054 ( .A1(n6209), .A2(n6200), .ZN(n8771) );
  INV_X1 U8055 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U8056 ( .A1(n6211), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6202) );
  NAND2_X1 U8057 ( .A1(n5958), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6201) );
  OAI211_X1 U8058 ( .C1(n8922), .C2(n6969), .A(n6202), .B(n6201), .ZN(n6203)
         );
  INV_X1 U8059 ( .A(n6203), .ZN(n6204) );
  NAND2_X1 U8060 ( .A1(n8995), .A2(n6502), .ZN(n6953) );
  NAND2_X1 U8061 ( .A1(n9089), .A2(n5988), .ZN(n6207) );
  OR2_X1 U8062 ( .A1(n6976), .A2(n6205), .ZN(n6206) );
  INV_X1 U8063 ( .A(n6209), .ZN(n6208) );
  INV_X1 U8064 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10199) );
  NAND2_X1 U8065 ( .A1(n6209), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U8066 ( .A1(n6220), .A2(n6210), .ZN(n8761) );
  NAND2_X1 U8067 ( .A1(n8761), .A2(n6231), .ZN(n6216) );
  INV_X1 U8068 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U8069 ( .A1(n5958), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U8070 ( .A1(n6211), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6212) );
  OAI211_X1 U8071 ( .C1(n6969), .C2(n8921), .A(n6213), .B(n6212), .ZN(n6214)
         );
  INV_X1 U8072 ( .A(n6214), .ZN(n6215) );
  NAND2_X1 U8073 ( .A1(n8989), .A2(n8584), .ZN(n6292) );
  INV_X1 U8074 ( .A(n6292), .ZN(n6955) );
  NAND2_X1 U8075 ( .A1(n8396), .A2(n5988), .ZN(n6219) );
  OR2_X1 U8076 ( .A1(n6976), .A2(n6217), .ZN(n6218) );
  NAND2_X1 U8077 ( .A1(n6220), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U8078 ( .A1(n6230), .A2(n6221), .ZN(n8476) );
  NAND2_X1 U8079 ( .A1(n8476), .A2(n6231), .ZN(n6227) );
  INV_X1 U8080 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U8081 ( .A1(n5926), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U8082 ( .A1(n5958), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6222) );
  OAI211_X1 U8083 ( .C1(n6966), .C2(n6224), .A(n6223), .B(n6222), .ZN(n6225)
         );
  INV_X1 U8084 ( .A(n6225), .ZN(n6226) );
  INV_X1 U8085 ( .A(n8759), .ZN(n6296) );
  NAND2_X1 U8086 ( .A1(n8480), .A2(n6296), .ZN(n6228) );
  INV_X1 U8087 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9085) );
  INV_X1 U8088 ( .A(n6958), .ZN(n6236) );
  NAND2_X1 U8089 ( .A1(n8380), .A2(n6231), .ZN(n6973) );
  INV_X1 U8090 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8381) );
  NAND2_X1 U8091 ( .A1(n5958), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6233) );
  NAND2_X1 U8092 ( .A1(n5926), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6232) );
  OAI211_X1 U8093 ( .C1(n8381), .C2(n6966), .A(n6233), .B(n6232), .ZN(n6234)
         );
  INV_X1 U8094 ( .A(n6234), .ZN(n6235) );
  NAND2_X1 U8095 ( .A1(n6973), .A2(n6235), .ZN(n8605) );
  INV_X1 U8096 ( .A(n8605), .ZN(n6956) );
  NAND2_X1 U8097 ( .A1(n6236), .A2(n6956), .ZN(n6987) );
  AOI21_X1 U8098 ( .B1(n7031), .B2(n8342), .A(n7028), .ZN(n6241) );
  AND2_X1 U8099 ( .A1(n10135), .A2(n6241), .ZN(n6243) );
  INV_X1 U8100 ( .A(n6384), .ZN(n6242) );
  INV_X1 U8101 ( .A(n7530), .ZN(n7478) );
  INV_X1 U8102 ( .A(n7454), .ZN(n10109) );
  NAND2_X1 U8103 ( .A1(n6245), .A2(n10109), .ZN(n6246) );
  NAND2_X1 U8104 ( .A1(n6247), .A2(n7630), .ZN(n6248) );
  NAND2_X1 U8105 ( .A1(n6249), .A2(n6248), .ZN(n7642) );
  AND2_X1 U8106 ( .A1(n7629), .A2(n10121), .ZN(n6250) );
  NAND2_X1 U8107 ( .A1(n10090), .A2(n6251), .ZN(n6253) );
  NAND2_X1 U8108 ( .A1(n6253), .A2(n6252), .ZN(n7795) );
  INV_X1 U8109 ( .A(n10092), .ZN(n7751) );
  NAND2_X1 U8110 ( .A1(n7751), .A2(n7725), .ZN(n6254) );
  NAND2_X1 U8111 ( .A1(n10092), .A2(n10129), .ZN(n6255) );
  INV_X1 U8112 ( .A(n8102), .ZN(n8612) );
  AND2_X1 U8113 ( .A1(n8612), .A2(n10140), .ZN(n6257) );
  OR2_X1 U8114 ( .A1(n8612), .A2(n10140), .ZN(n6256) );
  INV_X1 U8115 ( .A(n8033), .ZN(n10080) );
  AOI22_X1 U8116 ( .A1(n8976), .A2(n8610), .B1(n10150), .B2(n10080), .ZN(n6258) );
  NAND2_X1 U8117 ( .A1(n7974), .A2(n6258), .ZN(n6263) );
  INV_X1 U8118 ( .A(n8976), .ZN(n8039) );
  OAI21_X1 U8119 ( .B1(n10150), .B2(n10080), .A(n8610), .ZN(n6261) );
  NAND2_X1 U8120 ( .A1(n8055), .A2(n8033), .ZN(n6259) );
  NOR2_X1 U8121 ( .A1(n10150), .A2(n6259), .ZN(n6260) );
  AOI21_X1 U8122 ( .B1(n8039), .B2(n6261), .A(n6260), .ZN(n6262) );
  NAND2_X1 U8123 ( .A1(n6263), .A2(n6262), .ZN(n8053) );
  NAND2_X1 U8124 ( .A1(n8460), .A2(n8609), .ZN(n6264) );
  INV_X1 U8125 ( .A(n8455), .ZN(n8608) );
  NAND2_X1 U8126 ( .A1(n9065), .A2(n8910), .ZN(n6999) );
  NAND2_X1 U8127 ( .A1(n8314), .A2(n6999), .ZN(n6265) );
  OR2_X1 U8128 ( .A1(n9065), .A2(n8910), .ZN(n7000) );
  NAND2_X1 U8129 ( .A1(n6265), .A2(n7000), .ZN(n8907) );
  NAND2_X1 U8130 ( .A1(n9059), .A2(n8606), .ZN(n6266) );
  NAND2_X1 U8131 ( .A1(n8907), .A2(n6266), .ZN(n6268) );
  OR2_X1 U8132 ( .A1(n9059), .A2(n8606), .ZN(n6267) );
  NAND2_X1 U8133 ( .A1(n6268), .A2(n6267), .ZN(n8891) );
  NOR2_X1 U8134 ( .A1(n8590), .A2(n8909), .ZN(n6270) );
  NAND2_X1 U8135 ( .A1(n8590), .A2(n8909), .ZN(n6269) );
  NAND2_X1 U8136 ( .A1(n8948), .A2(n8885), .ZN(n6271) );
  AND2_X1 U8137 ( .A1(n9041), .A2(n8871), .ZN(n6274) );
  OR2_X1 U8138 ( .A1(n9041), .A2(n8871), .ZN(n6273) );
  INV_X1 U8139 ( .A(n8537), .ZN(n8863) );
  NAND2_X1 U8140 ( .A1(n6447), .A2(n8863), .ZN(n6276) );
  AND2_X1 U8141 ( .A1(n8835), .A2(n6276), .ZN(n6275) );
  INV_X1 U8142 ( .A(n6276), .ZN(n8834) );
  NOR2_X1 U8143 ( .A1(n8844), .A2(n8834), .ZN(n6279) );
  NOR2_X1 U8144 ( .A1(n6277), .A2(n8850), .ZN(n6278) );
  AOI21_X1 U8145 ( .B1(n8835), .B2(n6279), .A(n6278), .ZN(n8821) );
  INV_X1 U8146 ( .A(n6456), .ZN(n8837) );
  OR2_X1 U8147 ( .A1(n9025), .A2(n8837), .ZN(n6281) );
  NAND2_X1 U8148 ( .A1(n8790), .A2(n6283), .ZN(n8811) );
  OR2_X1 U8149 ( .A1(n9019), .A2(n8825), .ZN(n6284) );
  NAND2_X1 U8150 ( .A1(n9013), .A2(n8812), .ZN(n6286) );
  AND2_X1 U8151 ( .A1(n9007), .A2(n8803), .ZN(n6288) );
  NAND2_X1 U8152 ( .A1(n6938), .A2(n6952), .ZN(n8775) );
  OR2_X1 U8153 ( .A1(n9001), .A2(n8767), .ZN(n6289) );
  NAND2_X1 U8154 ( .A1(n8995), .A2(n8776), .ZN(n6291) );
  INV_X1 U8155 ( .A(n8758), .ZN(n6293) );
  NOR2_X1 U8156 ( .A1(n8989), .A2(n8768), .ZN(n7038) );
  INV_X1 U8157 ( .A(n7038), .ZN(n6295) );
  OAI211_X1 U8158 ( .C1(n8759), .C2(n8480), .A(n7016), .B(n6295), .ZN(n6307)
         );
  NAND2_X1 U8159 ( .A1(n8480), .A2(n8759), .ZN(n6298) );
  NAND3_X1 U8160 ( .A1(n8757), .A2(n6294), .A3(n6298), .ZN(n6306) );
  NAND2_X1 U8161 ( .A1(n6295), .A2(n8759), .ZN(n6297) );
  AOI22_X1 U8162 ( .A1(n7053), .A2(n6297), .B1(n7038), .B2(n6296), .ZN(n6303)
         );
  INV_X1 U8163 ( .A(n6298), .ZN(n6299) );
  NAND2_X1 U8164 ( .A1(n7016), .A2(n6299), .ZN(n6302) );
  OR2_X1 U8165 ( .A1(n8212), .A2(n6341), .ZN(n6301) );
  INV_X1 U8166 ( .A(n6342), .ZN(n6300) );
  OAI211_X1 U8167 ( .C1(n7016), .C2(n6303), .A(n6302), .B(n10096), .ZN(n6304)
         );
  INV_X1 U8168 ( .A(n6304), .ZN(n6305) );
  OAI211_X1 U8169 ( .C1(n8757), .C2(n6307), .A(n6306), .B(n6305), .ZN(n6319)
         );
  INV_X1 U8170 ( .A(n5804), .ZN(n7033) );
  NAND2_X1 U8171 ( .A1(n7033), .A2(n6308), .ZN(n6309) );
  INV_X1 U8172 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U8173 ( .A1(n5958), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6312) );
  INV_X1 U8174 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6310) );
  OR2_X1 U8175 ( .A1(n6966), .A2(n6310), .ZN(n6311) );
  OAI211_X1 U8176 ( .C1(n6313), .C2(n6969), .A(n6312), .B(n6311), .ZN(n6314)
         );
  INV_X1 U8177 ( .A(n6314), .ZN(n6315) );
  NAND2_X1 U8178 ( .A1(n6973), .A2(n6315), .ZN(n8604) );
  AND2_X1 U8179 ( .A1(n6316), .A2(P2_B_REG_SCAN_IN), .ZN(n6317) );
  NOR2_X1 U8180 ( .A1(n8896), .A2(n6317), .ZN(n8750) );
  AOI22_X1 U8181 ( .A1(n10093), .A2(n8759), .B1(n8604), .B2(n8750), .ZN(n6318)
         );
  INV_X1 U8182 ( .A(n10141), .ZN(n6321) );
  XNOR2_X1 U8183 ( .A(n6322), .B(P2_B_REG_SCAN_IN), .ZN(n6324) );
  NAND2_X1 U8184 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  INV_X1 U8185 ( .A(n6326), .ZN(n6327) );
  INV_X1 U8186 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U8187 ( .A1(n6327), .A2(n7368), .ZN(n6329) );
  INV_X1 U8188 ( .A(n7365), .ZN(n9096) );
  NAND2_X1 U8189 ( .A1(n6323), .A2(n9096), .ZN(n6328) );
  NAND2_X1 U8190 ( .A1(n6329), .A2(n6328), .ZN(n6358) );
  NAND2_X1 U8191 ( .A1(n6387), .A2(n6358), .ZN(n7305) );
  NOR2_X1 U8192 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .ZN(
        n6333) );
  NOR4_X1 U8193 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6332) );
  NOR4_X1 U8194 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6331) );
  NOR4_X1 U8195 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6330) );
  NAND4_X1 U8196 ( .A1(n6333), .A2(n6332), .A3(n6331), .A4(n6330), .ZN(n6339)
         );
  NOR4_X1 U8197 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6337) );
  NOR4_X1 U8198 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6336) );
  NOR4_X1 U8199 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6335) );
  NOR4_X1 U8200 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6334) );
  NAND4_X1 U8201 ( .A1(n6337), .A2(n6336), .A3(n6335), .A4(n6334), .ZN(n6338)
         );
  NOR2_X1 U8202 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  AND2_X1 U8203 ( .A1(n6980), .A2(n10135), .ZN(n6345) );
  NAND2_X1 U8204 ( .A1(n6341), .A2(n7031), .ZN(n6386) );
  INV_X1 U8205 ( .A(n6386), .ZN(n6343) );
  INV_X1 U8206 ( .A(n6489), .ZN(n6344) );
  NAND2_X1 U8207 ( .A1(n6345), .A2(n6344), .ZN(n6472) );
  NAND2_X1 U8208 ( .A1(n6472), .A2(n8778), .ZN(n6488) );
  NAND2_X1 U8209 ( .A1(n6485), .A2(n6488), .ZN(n6348) );
  OR2_X1 U8210 ( .A1(n6387), .A2(n6358), .ZN(n6355) );
  NOR2_X1 U8211 ( .A1(n6355), .A2(n6352), .ZN(n6486) );
  INV_X1 U8212 ( .A(n6495), .ZN(n7360) );
  NAND2_X1 U8213 ( .A1(n6486), .A2(n7360), .ZN(n6477) );
  INV_X1 U8214 ( .A(n6496), .ZN(n7525) );
  NOR2_X1 U8215 ( .A1(n7525), .A2(n6489), .ZN(n6346) );
  OR2_X1 U8216 ( .A1(n10152), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8217 ( .A1(n6236), .A2(n9066), .ZN(n6350) );
  NAND2_X1 U8218 ( .A1(n6351), .A2(n6350), .ZN(P2_U3456) );
  NOR2_X1 U8219 ( .A1(n6352), .A2(n6495), .ZN(n6353) );
  INV_X1 U8220 ( .A(n6354), .ZN(n7310) );
  AND2_X1 U8221 ( .A1(n6355), .A2(n6478), .ZN(n6362) );
  NAND2_X1 U8222 ( .A1(n7031), .A2(n8019), .ZN(n6356) );
  AOI21_X1 U8223 ( .B1(n6341), .B2(n6356), .A(n8342), .ZN(n6357) );
  OR2_X1 U8224 ( .A1(n6357), .A2(n6387), .ZN(n6361) );
  INV_X1 U8225 ( .A(n6357), .ZN(n6359) );
  NAND2_X1 U8226 ( .A1(n10164), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8227 ( .B1(n6365), .B2(n10164), .A(n4971), .ZN(P2_U3488) );
  NAND2_X1 U8228 ( .A1(n4777), .A2(n6366), .ZN(n6368) );
  NAND2_X1 U8229 ( .A1(n7060), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6367) );
  INV_X1 U8230 ( .A(n6371), .ZN(n6372) );
  INV_X1 U8231 ( .A(n6665), .ZN(n6789) );
  NAND2_X1 U8232 ( .A1(n6372), .A2(n6789), .ZN(n6374) );
  NAND2_X1 U8233 ( .A1(n6375), .A2(n6743), .ZN(n6376) );
  NAND2_X1 U8234 ( .A1(n6376), .A2(n6665), .ZN(n6378) );
  AOI22_X1 U8235 ( .A1(n9350), .A2(n9322), .B1(n9349), .B2(n9324), .ZN(n8412)
         );
  AOI21_X1 U8236 ( .B1(n8419), .B2(n6379), .A(n9784), .ZN(n6381) );
  AND2_X1 U8237 ( .A1(n6381), .A2(n6380), .ZN(n9573) );
  OR2_X1 U8238 ( .A1(n10070), .A2(n10298), .ZN(n6382) );
  OAI21_X1 U8239 ( .B1(n7061), .B2(n6383), .A(n4984), .ZN(P1_U3518) );
  OR2_X1 U8240 ( .A1(n6388), .A2(n6245), .ZN(n6389) );
  NAND2_X1 U8241 ( .A1(n6388), .A2(n6245), .ZN(n6393) );
  NAND2_X1 U8242 ( .A1(n6389), .A2(n6393), .ZN(n7449) );
  INV_X1 U8243 ( .A(n7449), .ZN(n6392) );
  OR2_X1 U8244 ( .A1(n6396), .A2(n7530), .ZN(n6390) );
  AND2_X1 U8245 ( .A1(n6390), .A2(n7730), .ZN(n7450) );
  NAND2_X1 U8246 ( .A1(n6392), .A2(n6391), .ZN(n7447) );
  NAND2_X1 U8247 ( .A1(n7447), .A2(n6393), .ZN(n7432) );
  XNOR2_X1 U8248 ( .A(n6396), .B(n10118), .ZN(n6394) );
  XNOR2_X1 U8249 ( .A(n6394), .B(n8615), .ZN(n7434) );
  NAND2_X1 U8250 ( .A1(n6394), .A2(n6247), .ZN(n6395) );
  NAND2_X1 U8251 ( .A1(n7433), .A2(n6395), .ZN(n7537) );
  INV_X1 U8252 ( .A(n7537), .ZN(n6398) );
  INV_X2 U8253 ( .A(n6396), .ZN(n6454) );
  XNOR2_X1 U8254 ( .A(n6471), .B(n7645), .ZN(n6402) );
  XNOR2_X1 U8255 ( .A(n6402), .B(n7629), .ZN(n7536) );
  INV_X1 U8256 ( .A(n7536), .ZN(n6397) );
  XNOR2_X1 U8257 ( .A(n6471), .B(n10124), .ZN(n6399) );
  NAND2_X1 U8258 ( .A1(n6399), .A2(n7533), .ZN(n7719) );
  INV_X1 U8259 ( .A(n6399), .ZN(n6400) );
  INV_X1 U8260 ( .A(n7533), .ZN(n8613) );
  NAND2_X1 U8261 ( .A1(n6400), .A2(n8613), .ZN(n6401) );
  AND2_X1 U8262 ( .A1(n7719), .A2(n6401), .ZN(n7651) );
  INV_X1 U8263 ( .A(n6402), .ZN(n6403) );
  INV_X1 U8264 ( .A(n7629), .ZN(n10094) );
  NAND2_X1 U8265 ( .A1(n6403), .A2(n10094), .ZN(n7648) );
  AND2_X1 U8266 ( .A1(n7651), .A2(n7648), .ZN(n6404) );
  XNOR2_X1 U8267 ( .A(n6471), .B(n10129), .ZN(n6405) );
  XNOR2_X1 U8268 ( .A(n6405), .B(n10092), .ZN(n7720) );
  NAND2_X1 U8269 ( .A1(n6405), .A2(n7751), .ZN(n6406) );
  XNOR2_X1 U8270 ( .A(n8473), .B(n7790), .ZN(n6407) );
  XNOR2_X1 U8271 ( .A(n6407), .B(n10079), .ZN(n7747) );
  NAND2_X1 U8272 ( .A1(n7748), .A2(n7747), .ZN(n7746) );
  INV_X1 U8273 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U8274 ( .A1(n6408), .A2(n10079), .ZN(n6409) );
  INV_X2 U8275 ( .A(n6454), .ZN(n8473) );
  XNOR2_X1 U8276 ( .A(n10140), .B(n8473), .ZN(n6411) );
  XNOR2_X1 U8277 ( .A(n6411), .B(n8102), .ZN(n7872) );
  NAND2_X1 U8278 ( .A1(n6411), .A2(n8102), .ZN(n6412) );
  XNOR2_X1 U8279 ( .A(n10150), .B(n8473), .ZN(n6413) );
  NAND2_X1 U8280 ( .A1(n6413), .A2(n8033), .ZN(n8107) );
  XNOR2_X1 U8281 ( .A(n8976), .B(n6454), .ZN(n8029) );
  NAND2_X1 U8282 ( .A1(n8029), .A2(n8610), .ZN(n8452) );
  INV_X1 U8283 ( .A(n6413), .ZN(n6414) );
  NAND2_X1 U8284 ( .A1(n6414), .A2(n10080), .ZN(n8109) );
  XNOR2_X1 U8285 ( .A(n8075), .B(n6454), .ZN(n8554) );
  XNOR2_X1 U8286 ( .A(n8460), .B(n8473), .ZN(n8552) );
  INV_X1 U8287 ( .A(n8029), .ZN(n6415) );
  AOI22_X1 U8288 ( .A1(n8552), .A2(n8551), .B1(n8055), .B2(n6415), .ZN(n6416)
         );
  NAND2_X1 U8289 ( .A1(n8473), .A2(n8609), .ZN(n6418) );
  OAI22_X1 U8290 ( .A1(n8460), .A2(n6418), .B1(n8455), .B2(n8473), .ZN(n6422)
         );
  NOR2_X1 U8291 ( .A1(n8473), .A2(n8551), .ZN(n6419) );
  AOI22_X1 U8292 ( .A1(n8460), .A2(n6419), .B1(n8608), .B2(n8473), .ZN(n6420)
         );
  NAND2_X1 U8293 ( .A1(n8075), .A2(n6420), .ZN(n6421) );
  OAI21_X1 U8294 ( .B1(n8075), .B2(n6422), .A(n6421), .ZN(n6423) );
  NAND2_X1 U8295 ( .A1(n6424), .A2(n6423), .ZN(n8094) );
  XNOR2_X1 U8296 ( .A(n8972), .B(n8473), .ZN(n6425) );
  XNOR2_X1 U8297 ( .A(n6425), .B(n8607), .ZN(n8093) );
  NAND2_X1 U8298 ( .A1(n8094), .A2(n8093), .ZN(n8092) );
  INV_X1 U8299 ( .A(n6425), .ZN(n6426) );
  NAND2_X1 U8300 ( .A1(n6426), .A2(n8607), .ZN(n6427) );
  NAND2_X1 U8301 ( .A1(n8092), .A2(n6427), .ZN(n8276) );
  XNOR2_X1 U8302 ( .A(n9065), .B(n8473), .ZN(n6428) );
  XNOR2_X1 U8303 ( .A(n6428), .B(n8910), .ZN(n8275) );
  NAND2_X1 U8304 ( .A1(n8276), .A2(n8275), .ZN(n8274) );
  INV_X1 U8305 ( .A(n6428), .ZN(n6429) );
  NAND2_X1 U8306 ( .A1(n6429), .A2(n8910), .ZN(n6430) );
  NAND2_X1 U8307 ( .A1(n8274), .A2(n6430), .ZN(n8439) );
  INV_X1 U8308 ( .A(n8439), .ZN(n6432) );
  XNOR2_X1 U8309 ( .A(n9059), .B(n6454), .ZN(n6433) );
  XNOR2_X1 U8310 ( .A(n6433), .B(n8606), .ZN(n8440) );
  INV_X1 U8311 ( .A(n8440), .ZN(n6431) );
  INV_X1 U8312 ( .A(n6433), .ZN(n6434) );
  NAND2_X1 U8313 ( .A1(n6434), .A2(n8897), .ZN(n6435) );
  XNOR2_X1 U8314 ( .A(n8590), .B(n8473), .ZN(n6436) );
  XNOR2_X1 U8315 ( .A(n6436), .B(n8909), .ZN(n8593) );
  INV_X1 U8316 ( .A(n6436), .ZN(n6437) );
  NAND2_X1 U8317 ( .A1(n6437), .A2(n8909), .ZN(n6438) );
  XNOR2_X1 U8318 ( .A(n9048), .B(n8473), .ZN(n6439) );
  XNOR2_X1 U8319 ( .A(n6439), .B(n8870), .ZN(n8507) );
  INV_X1 U8320 ( .A(n6439), .ZN(n6440) );
  NAND2_X1 U8321 ( .A1(n6440), .A2(n8870), .ZN(n6441) );
  XNOR2_X1 U8322 ( .A(n8948), .B(n6454), .ZN(n6443) );
  XNOR2_X1 U8323 ( .A(n6443), .B(n8885), .ZN(n8517) );
  INV_X1 U8324 ( .A(n8517), .ZN(n6442) );
  INV_X1 U8325 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8326 ( .A1(n6444), .A2(n8568), .ZN(n8570) );
  XNOR2_X1 U8327 ( .A(n9041), .B(n8473), .ZN(n6445) );
  XNOR2_X1 U8328 ( .A(n6445), .B(n8871), .ZN(n8569) );
  NAND2_X1 U8329 ( .A1(n6445), .A2(n8469), .ZN(n6446) );
  XNOR2_X1 U8330 ( .A(n6447), .B(n8473), .ZN(n6448) );
  XNOR2_X1 U8331 ( .A(n6448), .B(n8537), .ZN(n8463) );
  INV_X1 U8332 ( .A(n6448), .ZN(n6449) );
  NAND2_X1 U8333 ( .A1(n6449), .A2(n8863), .ZN(n6450) );
  XNOR2_X1 U8334 ( .A(n6277), .B(n8473), .ZN(n6452) );
  XNOR2_X1 U8335 ( .A(n6452), .B(n8850), .ZN(n8534) );
  NAND2_X1 U8336 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  XNOR2_X1 U8337 ( .A(n9025), .B(n6454), .ZN(n6455) );
  XNOR2_X1 U8338 ( .A(n6455), .B(n6456), .ZN(n8492) );
  INV_X1 U8339 ( .A(n6455), .ZN(n6457) );
  NAND2_X1 U8340 ( .A1(n6457), .A2(n6456), .ZN(n6458) );
  NAND2_X1 U8341 ( .A1(n6459), .A2(n6458), .ZN(n8542) );
  XNOR2_X1 U8342 ( .A(n9019), .B(n6471), .ZN(n6460) );
  XNOR2_X1 U8343 ( .A(n6460), .B(n8825), .ZN(n8543) );
  AND2_X1 U8344 ( .A1(n6460), .A2(n8496), .ZN(n6461) );
  XNOR2_X1 U8345 ( .A(n9007), .B(n8473), .ZN(n8527) );
  XNOR2_X1 U8346 ( .A(n9013), .B(n8473), .ZN(n6462) );
  OAI22_X1 U8347 ( .A1(n8527), .A2(n8526), .B1(n8788), .B2(n6462), .ZN(n6466)
         );
  OAI21_X1 U8348 ( .B1(n8523), .B2(n8812), .A(n8803), .ZN(n6463) );
  NOR3_X1 U8349 ( .A1(n8523), .A2(n8803), .A3(n8812), .ZN(n6464) );
  XNOR2_X1 U8350 ( .A(n9001), .B(n8473), .ZN(n6468) );
  XOR2_X1 U8351 ( .A(n8767), .B(n6468), .Z(n8500) );
  INV_X1 U8352 ( .A(n8500), .ZN(n6467) );
  XNOR2_X1 U8353 ( .A(n8995), .B(n8473), .ZN(n6470) );
  XNOR2_X1 U8354 ( .A(n6470), .B(n8776), .ZN(n8579) );
  XNOR2_X1 U8355 ( .A(n8989), .B(n6471), .ZN(n8485) );
  NOR2_X1 U8356 ( .A1(n8485), .A2(n8584), .ZN(n8481) );
  AOI21_X1 U8357 ( .B1(n8584), .B2(n8485), .A(n8481), .ZN(n6475) );
  NAND2_X1 U8358 ( .A1(n6476), .A2(n6475), .ZN(n8484) );
  NAND2_X1 U8359 ( .A1(n6485), .A2(n6489), .ZN(n6474) );
  OR2_X1 U8360 ( .A1(n6477), .A2(n6472), .ZN(n6473) );
  OAI211_X1 U8361 ( .C1(n6476), .C2(n6475), .A(n8484), .B(n8591), .ZN(n6508)
         );
  INV_X1 U8362 ( .A(n8989), .ZN(n6505) );
  OR2_X1 U8363 ( .A1(n6477), .A2(n10135), .ZN(n6479) );
  INV_X1 U8364 ( .A(n6485), .ZN(n6482) );
  OR2_X1 U8365 ( .A1(n6496), .A2(n6480), .ZN(n6481) );
  NOR2_X2 U8366 ( .A1(n6482), .A2(n6481), .ZN(n8595) );
  NOR2_X1 U8367 ( .A1(n6496), .A2(n6483), .ZN(n6484) );
  NAND2_X1 U8368 ( .A1(n6485), .A2(n6484), .ZN(n8597) );
  INV_X1 U8369 ( .A(n6486), .ZN(n6487) );
  NAND2_X1 U8370 ( .A1(n6488), .A2(n6487), .ZN(n6493) );
  NAND2_X1 U8371 ( .A1(n6497), .A2(n6489), .ZN(n6490) );
  NAND4_X1 U8372 ( .A1(n6493), .A2(n6492), .A3(n6491), .A4(n6490), .ZN(n6494)
         );
  NAND2_X1 U8373 ( .A1(n6494), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6499) );
  NOR2_X1 U8374 ( .A1(n6496), .A2(n6495), .ZN(n7034) );
  NAND2_X1 U8375 ( .A1(n7034), .A2(n6497), .ZN(n6498) );
  OR2_X1 U8376 ( .A1(n6500), .A2(P2_U3151), .ZN(n8345) );
  AOI22_X1 U8377 ( .A1(n8761), .A2(n8599), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n6501) );
  OAI21_X1 U8378 ( .B1(n6502), .B2(n8597), .A(n6501), .ZN(n6503) );
  AOI21_X1 U8379 ( .B1(n8595), .B2(n8759), .A(n6503), .ZN(n6504) );
  INV_X1 U8380 ( .A(n6506), .ZN(n6507) );
  INV_X1 U8381 ( .A(n6509), .ZN(n6519) );
  NAND2_X1 U8382 ( .A1(n6511), .A2(n6510), .ZN(n6513) );
  NAND2_X1 U8383 ( .A1(n6513), .A2(n6512), .ZN(n6514) );
  MUX2_X1 U8384 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7342), .Z(n6520) );
  XNOR2_X1 U8385 ( .A(n6520), .B(SI_30_), .ZN(n6521) );
  NAND2_X1 U8386 ( .A1(n8424), .A2(n5397), .ZN(n6517) );
  NAND2_X1 U8387 ( .A1(n5137), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n6516) );
  INV_X1 U8388 ( .A(n9567), .ZN(n6518) );
  NAND2_X1 U8389 ( .A1(n6519), .A2(n6518), .ZN(n6527) );
  MUX2_X1 U8390 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7342), .Z(n6524) );
  INV_X1 U8391 ( .A(SI_31_), .ZN(n6523) );
  XNOR2_X1 U8392 ( .A(n6524), .B(n6523), .ZN(n6525) );
  INV_X1 U8393 ( .A(n6529), .ZN(n6535) );
  INV_X1 U8394 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6533) );
  INV_X1 U8395 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6536) );
  OR2_X1 U8396 ( .A1(n6530), .A2(n6536), .ZN(n6532) );
  NAND2_X1 U8397 ( .A1(n5063), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6531) );
  OAI211_X1 U8398 ( .C1(n6534), .C2(n6533), .A(n6532), .B(n6531), .ZN(n9347)
         );
  NAND2_X1 U8399 ( .A1(n6535), .A2(n9347), .ZN(n9807) );
  MUX2_X1 U8400 ( .A(n8391), .B(n6536), .S(n7060), .Z(n6538) );
  NAND2_X1 U8401 ( .A1(n6687), .A2(n6366), .ZN(n6537) );
  NAND2_X1 U8402 ( .A1(n6538), .A2(n6537), .ZN(P1_U3553) );
  NOR2_X2 U8403 ( .A1(n7064), .A2(n9564), .ZN(n6679) );
  INV_X1 U8404 ( .A(n6786), .ZN(n6675) );
  OR2_X1 U8405 ( .A1(n9814), .A2(n6540), .ZN(n6542) );
  INV_X1 U8406 ( .A(n6740), .ZN(n6544) );
  NAND2_X1 U8407 ( .A1(n6544), .A2(n6802), .ZN(n6551) );
  OR2_X1 U8408 ( .A1(n7272), .A2(n6826), .ZN(n6547) );
  NOR2_X1 U8409 ( .A1(n6547), .A2(n8404), .ZN(n6546) );
  NAND2_X1 U8410 ( .A1(n7272), .A2(n6826), .ZN(n6666) );
  OAI21_X1 U8411 ( .B1(n5555), .B2(n6666), .A(n6668), .ZN(n6545) );
  OAI21_X1 U8412 ( .B1(n6546), .B2(n6668), .A(n6545), .ZN(n6550) );
  OAI22_X1 U8413 ( .A1(n6668), .A2(n6547), .B1(n8404), .B2(n6826), .ZN(n6548)
         );
  NAND2_X1 U8414 ( .A1(n9578), .A2(n6548), .ZN(n6549) );
  INV_X1 U8415 ( .A(n6551), .ZN(n6664) );
  NAND2_X1 U8416 ( .A1(n9354), .A2(n6826), .ZN(n6553) );
  OAI22_X1 U8417 ( .A1(n9922), .A2(n6553), .B1(n9119), .B2(n6679), .ZN(n6552)
         );
  INV_X1 U8418 ( .A(n6552), .ZN(n6556) );
  INV_X1 U8419 ( .A(n6553), .ZN(n6554) );
  NAND2_X1 U8420 ( .A1(n9353), .A2(n6554), .ZN(n6555) );
  OAI22_X1 U8421 ( .A1(n6556), .A2(n9920), .B1(n9922), .B2(n6555), .ZN(n6557)
         );
  AOI21_X1 U8422 ( .B1(n6732), .B2(n6826), .A(n6557), .ZN(n6663) );
  INV_X1 U8423 ( .A(n9847), .ZN(n9716) );
  NAND3_X1 U8424 ( .A1(n9672), .A2(n9716), .A3(n6630), .ZN(n6558) );
  OAI21_X1 U8425 ( .B1(n9313), .B2(n6679), .A(n6558), .ZN(n6560) );
  NAND2_X1 U8426 ( .A1(n6560), .A2(n6559), .ZN(n6562) );
  NAND3_X1 U8427 ( .A1(n9672), .A2(n6679), .A3(n6630), .ZN(n6561) );
  NAND2_X1 U8428 ( .A1(n6562), .A2(n6561), .ZN(n6624) );
  NAND2_X1 U8429 ( .A1(n7840), .A2(n6696), .ZN(n6563) );
  NAND3_X1 U8430 ( .A1(n6563), .A2(n6759), .A3(n7817), .ZN(n6564) );
  NAND3_X1 U8431 ( .A1(n6564), .A2(n6700), .A3(n6703), .ZN(n6565) );
  NAND3_X1 U8432 ( .A1(n6565), .A2(n8154), .A3(n6569), .ZN(n6566) );
  NAND2_X1 U8433 ( .A1(n6566), .A2(n8155), .ZN(n6574) );
  INV_X1 U8434 ( .A(n7817), .ZN(n6567) );
  OAI211_X1 U8435 ( .C1(n7840), .C2(n6567), .A(n6759), .B(n6696), .ZN(n6571)
         );
  NAND2_X1 U8436 ( .A1(n6569), .A2(n6568), .ZN(n6704) );
  INV_X1 U8437 ( .A(n6704), .ZN(n6570) );
  NAND2_X1 U8438 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  INV_X1 U8439 ( .A(n8241), .ZN(n6575) );
  NAND2_X1 U8440 ( .A1(n6577), .A2(n6576), .ZN(n6579) );
  NAND2_X1 U8441 ( .A1(n8158), .A2(n6765), .ZN(n6578) );
  MUX2_X1 U8442 ( .A(n6579), .B(n6578), .S(n6826), .Z(n6580) );
  INV_X1 U8443 ( .A(n6580), .ZN(n6581) );
  NAND2_X1 U8444 ( .A1(n6582), .A2(n6581), .ZN(n6586) );
  MUX2_X1 U8445 ( .A(n6583), .B(n6764), .S(n6679), .Z(n6584) );
  INV_X1 U8446 ( .A(n6584), .ZN(n6585) );
  NAND2_X1 U8447 ( .A1(n6586), .A2(n6585), .ZN(n6593) );
  NAND2_X1 U8448 ( .A1(n6593), .A2(n6587), .ZN(n6588) );
  NAND2_X1 U8449 ( .A1(n6588), .A2(n6594), .ZN(n6589) );
  NAND3_X1 U8450 ( .A1(n6590), .A2(n6712), .A3(n8283), .ZN(n6591) );
  NAND2_X1 U8451 ( .A1(n6593), .A2(n6592), .ZN(n6595) );
  NAND2_X1 U8452 ( .A1(n8283), .A2(n6594), .ZN(n6709) );
  AOI21_X1 U8453 ( .B1(n6595), .B2(n6710), .A(n6709), .ZN(n6598) );
  NAND2_X1 U8454 ( .A1(n6597), .A2(n6596), .ZN(n6714) );
  OAI21_X1 U8455 ( .B1(n6598), .B2(n6714), .A(n6712), .ZN(n6599) );
  AND2_X1 U8456 ( .A1(n6614), .A2(n6611), .ZN(n6723) );
  INV_X1 U8457 ( .A(n6723), .ZN(n6602) );
  NAND3_X1 U8458 ( .A1(n6773), .A2(n6826), .A3(n6716), .ZN(n6601) );
  NAND3_X1 U8459 ( .A1(n6772), .A2(n6679), .A3(n6713), .ZN(n6600) );
  OAI22_X1 U8460 ( .A1(n6602), .A2(n6601), .B1(n6692), .B2(n6600), .ZN(n6603)
         );
  NAND2_X1 U8461 ( .A1(n6604), .A2(n6603), .ZN(n6620) );
  NAND2_X1 U8462 ( .A1(n6716), .A2(n9338), .ZN(n6608) );
  OAI21_X1 U8463 ( .B1(n6716), .B2(n9338), .A(n9967), .ZN(n6605) );
  NAND4_X1 U8464 ( .A1(n9752), .A2(n6679), .A3(n6608), .A4(n6605), .ZN(n6606)
         );
  OAI21_X1 U8465 ( .B1(n6611), .B2(n6826), .A(n6606), .ZN(n6607) );
  NAND2_X1 U8466 ( .A1(n6607), .A2(n6691), .ZN(n6616) );
  AOI21_X1 U8467 ( .B1(n6713), .B2(n9363), .A(n6679), .ZN(n6610) );
  INV_X1 U8468 ( .A(n9967), .ZN(n7182) );
  OAI21_X1 U8469 ( .B1(n6608), .B2(n6713), .A(n7182), .ZN(n6609) );
  NAND3_X1 U8470 ( .A1(n6611), .A2(n6610), .A3(n6609), .ZN(n6612) );
  NAND2_X1 U8471 ( .A1(n6614), .A2(n6612), .ZN(n6613) );
  OAI21_X1 U8472 ( .B1(n6614), .B2(n6679), .A(n6613), .ZN(n6615) );
  OAI211_X1 U8473 ( .C1(n6617), .C2(n6679), .A(n6616), .B(n6615), .ZN(n6618)
         );
  INV_X1 U8474 ( .A(n6618), .ZN(n6619) );
  NAND2_X1 U8475 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NAND2_X1 U8476 ( .A1(n6621), .A2(n9738), .ZN(n6626) );
  AND2_X1 U8477 ( .A1(n6629), .A2(n9721), .ZN(n6721) );
  NAND2_X1 U8478 ( .A1(n6626), .A2(n6721), .ZN(n6622) );
  NAND4_X1 U8479 ( .A1(n6622), .A2(n6679), .A3(n6690), .A4(n6628), .ZN(n6623)
         );
  NAND2_X1 U8480 ( .A1(n6624), .A2(n6623), .ZN(n6638) );
  NAND2_X1 U8481 ( .A1(n6625), .A2(n6679), .ZN(n6637) );
  INV_X1 U8482 ( .A(n6626), .ZN(n6633) );
  AND2_X1 U8483 ( .A1(n6628), .A2(n6627), .ZN(n6726) );
  INV_X1 U8484 ( .A(n6726), .ZN(n6632) );
  NAND2_X1 U8485 ( .A1(n6630), .A2(n6629), .ZN(n6724) );
  INV_X1 U8486 ( .A(n6724), .ZN(n6631) );
  OAI211_X1 U8487 ( .C1(n6633), .C2(n6632), .A(n6631), .B(n6826), .ZN(n6634)
         );
  NAND2_X1 U8488 ( .A1(n6635), .A2(n6634), .ZN(n6636) );
  NOR2_X1 U8489 ( .A1(n6733), .A2(n6679), .ZN(n6640) );
  OAI22_X1 U8490 ( .A1(n6641), .A2(n6640), .B1(n6679), .B2(n6639), .ZN(n6651)
         );
  NAND2_X1 U8491 ( .A1(n6642), .A2(n9637), .ZN(n6728) );
  INV_X1 U8492 ( .A(n6728), .ZN(n6649) );
  NAND2_X1 U8493 ( .A1(n9920), .A2(n9353), .ZN(n6643) );
  NAND2_X1 U8494 ( .A1(n6644), .A2(n6643), .ZN(n6648) );
  AND2_X1 U8495 ( .A1(n6727), .A2(n6645), .ZN(n6739) );
  INV_X1 U8496 ( .A(n6739), .ZN(n6646) );
  NAND2_X1 U8497 ( .A1(n6646), .A2(n6826), .ZN(n6647) );
  OAI211_X1 U8498 ( .C1(n6649), .C2(n6826), .A(n6648), .B(n6647), .ZN(n6650)
         );
  AND2_X1 U8499 ( .A1(n9292), .A2(n6679), .ZN(n6652) );
  NAND2_X1 U8500 ( .A1(n9922), .A2(n6652), .ZN(n6655) );
  OAI21_X1 U8501 ( .B1(n6826), .B2(n9353), .A(n6655), .ZN(n6653) );
  NAND2_X1 U8502 ( .A1(n6653), .A2(n9920), .ZN(n6654) );
  OAI21_X1 U8503 ( .B1(n6655), .B2(n9353), .A(n6654), .ZN(n6657) );
  INV_X1 U8504 ( .A(n6732), .ZN(n6656) );
  OAI21_X1 U8505 ( .B1(n6658), .B2(n6657), .A(n6656), .ZN(n6662) );
  NAND2_X1 U8506 ( .A1(n6668), .A2(n9350), .ZN(n6659) );
  NAND2_X1 U8507 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  INV_X1 U8508 ( .A(n6666), .ZN(n6667) );
  NAND2_X1 U8509 ( .A1(n6668), .A2(n6667), .ZN(n6670) );
  NAND2_X1 U8510 ( .A1(n8404), .A2(n6826), .ZN(n6669) );
  NAND2_X1 U8511 ( .A1(n6670), .A2(n6669), .ZN(n6671) );
  NAND2_X1 U8512 ( .A1(n8419), .A2(n6671), .ZN(n6672) );
  MUX2_X1 U8513 ( .A(n6748), .B(n6809), .S(n6679), .Z(n6676) );
  INV_X1 U8514 ( .A(n6750), .ZN(n9348) );
  AND2_X1 U8515 ( .A1(n6687), .A2(n9348), .ZN(n6677) );
  NAND2_X1 U8516 ( .A1(n6678), .A2(n6677), .ZN(n6684) );
  INV_X1 U8517 ( .A(n9347), .ZN(n6686) );
  OR2_X1 U8518 ( .A1(n6750), .A2(n6686), .ZN(n6813) );
  AND2_X1 U8519 ( .A1(n6791), .A2(n6813), .ZN(n6681) );
  NAND2_X1 U8520 ( .A1(n6682), .A2(n6681), .ZN(n6683) );
  NAND2_X1 U8521 ( .A1(n6684), .A2(n6683), .ZN(n6830) );
  INV_X1 U8522 ( .A(n6830), .ZN(n6689) );
  INV_X1 U8523 ( .A(n6685), .ZN(n6687) );
  INV_X1 U8524 ( .A(n6827), .ZN(n6688) );
  INV_X1 U8525 ( .A(n6690), .ZN(n6735) );
  INV_X1 U8526 ( .A(n6691), .ZN(n6722) );
  INV_X1 U8527 ( .A(n6692), .ZN(n6719) );
  AOI21_X1 U8528 ( .B1(n6693), .B2(n7715), .A(n8301), .ZN(n6694) );
  OAI21_X1 U8529 ( .B1(n7073), .B2(n4293), .A(n6694), .ZN(n6695) );
  INV_X1 U8530 ( .A(n6695), .ZN(n6698) );
  OAI211_X1 U8531 ( .C1(n6699), .C2(n6698), .A(n6697), .B(n6696), .ZN(n6702)
         );
  INV_X1 U8532 ( .A(n6700), .ZN(n6701) );
  AOI21_X1 U8533 ( .B1(n6702), .B2(n7817), .A(n6701), .ZN(n6705) );
  OAI21_X1 U8534 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(n6706) );
  AND2_X1 U8535 ( .A1(n6706), .A2(n8154), .ZN(n6708) );
  OAI21_X1 U8536 ( .B1(n6708), .B2(n6768), .A(n6707), .ZN(n6711) );
  AOI21_X1 U8537 ( .B1(n6711), .B2(n6710), .A(n6709), .ZN(n6715) );
  OAI211_X1 U8538 ( .C1(n6715), .C2(n6714), .A(n6713), .B(n6712), .ZN(n6717)
         );
  NAND3_X1 U8539 ( .A1(n6717), .A2(n6773), .A3(n6716), .ZN(n6718) );
  NAND3_X1 U8540 ( .A1(n6719), .A2(n6772), .A3(n6718), .ZN(n6720) );
  OAI211_X1 U8541 ( .C1(n6723), .C2(n6722), .A(n6721), .B(n6720), .ZN(n6725)
         );
  AOI21_X1 U8542 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6734) );
  NAND2_X1 U8543 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  NAND2_X1 U8544 ( .A1(n6729), .A2(n9606), .ZN(n6730) );
  AND2_X1 U8545 ( .A1(n6730), .A2(n6738), .ZN(n6731) );
  NOR2_X2 U8546 ( .A1(n6732), .A2(n6731), .ZN(n6800) );
  OAI211_X1 U8547 ( .C1(n6735), .C2(n6734), .A(n6800), .B(n6733), .ZN(n6736)
         );
  NAND2_X1 U8548 ( .A1(n6736), .A2(n6802), .ZN(n6746) );
  NAND3_X1 U8549 ( .A1(n6739), .A2(n6738), .A3(n6737), .ZN(n6741) );
  AOI21_X1 U8550 ( .B1(n6800), .B2(n6741), .A(n6740), .ZN(n6745) );
  INV_X1 U8551 ( .A(n6807), .ZN(n6744) );
  OAI211_X1 U8552 ( .C1(n6745), .C2(n6744), .A(n6743), .B(n6742), .ZN(n6805)
         );
  AOI21_X1 U8553 ( .B1(n6807), .B2(n6746), .A(n6805), .ZN(n6749) );
  NAND2_X1 U8554 ( .A1(n6748), .A2(n6747), .ZN(n6810) );
  NAND2_X1 U8555 ( .A1(n9567), .A2(n6750), .ZN(n6788) );
  OAI211_X1 U8556 ( .C1(n6749), .C2(n6810), .A(n6809), .B(n6788), .ZN(n6751)
         );
  OR2_X1 U8557 ( .A1(n9567), .A2(n6750), .ZN(n6787) );
  AOI21_X1 U8558 ( .B1(n6751), .B2(n6787), .A(n6754), .ZN(n6752) );
  NOR2_X1 U8559 ( .A1(n6752), .A2(n6827), .ZN(n6753) );
  MUX2_X1 U8560 ( .A(n7065), .B(n7063), .S(n6753), .Z(n6821) );
  INV_X1 U8561 ( .A(n6754), .ZN(n6791) );
  INV_X1 U8562 ( .A(n6755), .ZN(n6756) );
  INV_X1 U8563 ( .A(n9753), .ZN(n9763) );
  INV_X1 U8564 ( .A(n8285), .ZN(n6771) );
  XNOR2_X1 U8565 ( .A(n6693), .B(n7836), .ZN(n9798) );
  NAND4_X1 U8566 ( .A1(n6759), .A2(n6758), .A3(n9798), .A4(n8301), .ZN(n6763)
         );
  XNOR2_X1 U8567 ( .A(n9374), .B(n7813), .ZN(n7832) );
  NAND2_X1 U8568 ( .A1(n6760), .A2(n7832), .ZN(n6762) );
  NOR3_X1 U8569 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n6767) );
  INV_X1 U8570 ( .A(n6764), .ZN(n6766) );
  NAND4_X1 U8571 ( .A1(n6767), .A2(n6766), .A3(n8154), .A4(n6765), .ZN(n6769)
         );
  NOR3_X1 U8572 ( .A1(n6769), .A2(n8000), .A3(n6768), .ZN(n6770) );
  NAND4_X1 U8573 ( .A1(n5654), .A2(n8071), .A3(n6771), .A4(n6770), .ZN(n6774)
         );
  NAND2_X1 U8574 ( .A1(n6773), .A2(n6772), .ZN(n8358) );
  NOR2_X1 U8575 ( .A1(n6774), .A2(n8358), .ZN(n6775) );
  NAND4_X1 U8576 ( .A1(n9738), .A2(n9776), .A3(n9763), .A4(n6775), .ZN(n6776)
         );
  NOR2_X1 U8577 ( .A1(n9723), .A2(n6776), .ZN(n6777) );
  AND2_X1 U8578 ( .A1(n9705), .A2(n6777), .ZN(n6780) );
  NAND2_X1 U8579 ( .A1(n6779), .A2(n6778), .ZN(n9692) );
  NAND4_X1 U8580 ( .A1(n9674), .A2(n9652), .A3(n6780), .A4(n9692), .ZN(n6781)
         );
  OR2_X1 U8581 ( .A1(n6781), .A2(n9642), .ZN(n6782) );
  NOR2_X1 U8582 ( .A1(n9625), .A2(n6782), .ZN(n6783) );
  NAND4_X1 U8583 ( .A1(n6784), .A2(n9607), .A3(n6783), .A4(n5666), .ZN(n6785)
         );
  NOR2_X1 U8584 ( .A1(n7444), .A2(n9564), .ZN(n6792) );
  INV_X1 U8585 ( .A(n7068), .ZN(n9796) );
  INV_X1 U8586 ( .A(n9801), .ZN(n6797) );
  NAND2_X1 U8587 ( .A1(n9796), .A2(n6797), .ZN(n6798) );
  NOR2_X1 U8588 ( .A1(n7445), .A2(n6798), .ZN(n7291) );
  NOR2_X1 U8589 ( .A1(n5674), .A2(n10002), .ZN(n9388) );
  OAI21_X1 U8590 ( .B1(n7444), .B2(n7064), .A(P1_B_REG_SCAN_IN), .ZN(n6799) );
  AOI21_X1 U8591 ( .B1(n7291), .B2(n9388), .A(n6799), .ZN(n6820) );
  INV_X1 U8592 ( .A(n6820), .ZN(n6819) );
  INV_X1 U8593 ( .A(n7444), .ZN(n8336) );
  OAI21_X1 U8594 ( .B1(n9564), .B2(n8188), .A(n8336), .ZN(n6818) );
  INV_X1 U8595 ( .A(n6800), .ZN(n6804) );
  OAI21_X1 U8596 ( .B1(n6804), .B2(n6803), .A(n6802), .ZN(n6806) );
  AOI21_X1 U8597 ( .B1(n6807), .B2(n6806), .A(n6805), .ZN(n6811) );
  NAND2_X1 U8598 ( .A1(n9567), .A2(n6813), .ZN(n6808) );
  OAI211_X1 U8599 ( .C1(n6811), .C2(n6810), .A(n6809), .B(n6808), .ZN(n6812)
         );
  OAI21_X1 U8600 ( .B1(n6813), .B2(n9567), .A(n6812), .ZN(n6814) );
  AOI211_X1 U8601 ( .C1(n6814), .C2(n6791), .A(n6827), .B(n7287), .ZN(n6816)
         );
  NOR4_X1 U8602 ( .A1(n6816), .A2(n6815), .A3(n6820), .A4(n8188), .ZN(n6817)
         );
  AOI21_X1 U8603 ( .B1(n6819), .B2(n6818), .A(n6817), .ZN(n6823) );
  NAND2_X1 U8604 ( .A1(n6823), .A2(n6822), .ZN(n6833) );
  NOR3_X1 U8605 ( .A1(n7444), .A2(n7064), .A3(n6824), .ZN(n6825) );
  OAI21_X1 U8606 ( .B1(n6791), .B2(n9564), .A(n6825), .ZN(n6828) );
  AOI21_X1 U8607 ( .B1(n6830), .B2(n6688), .A(n6829), .ZN(n6831) );
  NAND3_X1 U8608 ( .A1(n6834), .A2(n6833), .A3(n6832), .ZN(P1_U3242) );
  NAND2_X1 U8609 ( .A1(n9013), .A2(n8788), .ZN(n8793) );
  AND2_X1 U8610 ( .A1(n6995), .A2(n8793), .ZN(n6936) );
  INV_X1 U8611 ( .A(n6835), .ZN(n6909) );
  OR2_X1 U8612 ( .A1(n7737), .A2(n7530), .ZN(n7001) );
  NAND3_X1 U8613 ( .A1(n6838), .A2(n7730), .A3(n6837), .ZN(n6836) );
  MUX2_X1 U8614 ( .A(n6837), .B(n6836), .S(n6980), .Z(n6841) );
  NAND3_X1 U8615 ( .A1(n6841), .A2(n6840), .A3(n7627), .ZN(n6848) );
  OR2_X1 U8616 ( .A1(n7629), .A2(n7645), .ZN(n6857) );
  NAND2_X1 U8617 ( .A1(n6857), .A2(n6842), .ZN(n6845) );
  NAND2_X1 U8618 ( .A1(n6843), .A2(n6850), .ZN(n6844) );
  MUX2_X1 U8619 ( .A(n6845), .B(n6844), .S(n6980), .Z(n6846) );
  INV_X1 U8620 ( .A(n6846), .ZN(n6847) );
  NAND2_X1 U8621 ( .A1(n6848), .A2(n6847), .ZN(n6849) );
  NAND2_X1 U8622 ( .A1(n6849), .A2(n10098), .ZN(n6861) );
  INV_X1 U8623 ( .A(n6850), .ZN(n6853) );
  OAI21_X1 U8624 ( .B1(n7533), .B2(n10124), .A(n6862), .ZN(n6851) );
  INV_X1 U8625 ( .A(n6851), .ZN(n6852) );
  OAI21_X1 U8626 ( .B1(n6861), .B2(n6853), .A(n6852), .ZN(n6856) );
  INV_X1 U8627 ( .A(n7989), .ZN(n6864) );
  NOR2_X1 U8628 ( .A1(n6864), .A2(n6858), .ZN(n6855) );
  INV_X1 U8629 ( .A(n6863), .ZN(n6854) );
  AOI21_X1 U8630 ( .B1(n6856), .B2(n6855), .A(n6854), .ZN(n6868) );
  INV_X1 U8631 ( .A(n6857), .ZN(n6860) );
  OAI211_X1 U8632 ( .C1(n6861), .C2(n6860), .A(n5991), .B(n6859), .ZN(n6866)
         );
  AND2_X1 U8633 ( .A1(n6863), .A2(n6862), .ZN(n6865) );
  AOI21_X1 U8634 ( .B1(n6866), .B2(n6865), .A(n6864), .ZN(n6867) );
  NAND2_X1 U8635 ( .A1(n8050), .A2(n7007), .ZN(n6870) );
  AOI21_X1 U8636 ( .B1(n7005), .B2(n7006), .A(n6988), .ZN(n6869) );
  NAND2_X1 U8637 ( .A1(n7991), .A2(n6874), .ZN(n10075) );
  NOR2_X1 U8638 ( .A1(n6873), .A2(n10075), .ZN(n6871) );
  NAND2_X1 U8639 ( .A1(n6872), .A2(n6871), .ZN(n6883) );
  INV_X1 U8640 ( .A(n6873), .ZN(n6877) );
  NAND2_X1 U8641 ( .A1(n7006), .A2(n6874), .ZN(n6876) );
  NAND2_X1 U8642 ( .A1(n7003), .A2(n7005), .ZN(n6875) );
  AOI21_X1 U8643 ( .B1(n6877), .B2(n6876), .A(n6875), .ZN(n6881) );
  INV_X1 U8644 ( .A(n7005), .ZN(n6878) );
  OAI211_X1 U8645 ( .C1(n6878), .C2(n7968), .A(n7004), .B(n8050), .ZN(n6879)
         );
  INV_X1 U8646 ( .A(n6879), .ZN(n6880) );
  NAND2_X1 U8647 ( .A1(n6883), .A2(n6882), .ZN(n6888) );
  MUX2_X1 U8648 ( .A(n7004), .B(n7003), .S(n6980), .Z(n6886) );
  AND3_X1 U8649 ( .A1(n6886), .A2(n6885), .A3(n6884), .ZN(n6887) );
  NAND3_X1 U8650 ( .A1(n6888), .A2(n6887), .A3(n8193), .ZN(n6896) );
  OR2_X1 U8651 ( .A1(n8455), .A2(n6988), .ZN(n6890) );
  NAND3_X1 U8652 ( .A1(n8563), .A2(n6988), .A3(n8455), .ZN(n6889) );
  OAI21_X1 U8653 ( .B1(n8563), .B2(n6890), .A(n6889), .ZN(n6894) );
  NAND3_X1 U8654 ( .A1(n8972), .A2(n8557), .A3(n6988), .ZN(n6892) );
  OR3_X1 U8655 ( .A1(n8972), .A2(n6988), .A3(n8557), .ZN(n6891) );
  NAND2_X1 U8656 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  AOI21_X1 U8657 ( .B1(n8193), .B2(n6894), .A(n6893), .ZN(n6895) );
  NAND2_X1 U8658 ( .A1(n6896), .A2(n6895), .ZN(n6899) );
  INV_X1 U8659 ( .A(n7000), .ZN(n6898) );
  MUX2_X1 U8660 ( .A(n8910), .B(n9065), .S(n6988), .Z(n6897) );
  MUX2_X1 U8661 ( .A(n6901), .B(n6900), .S(n6980), .Z(n6902) );
  NAND3_X1 U8662 ( .A1(n6911), .A2(n6903), .A3(n6912), .ZN(n6904) );
  NAND2_X1 U8663 ( .A1(n8857), .A2(n6906), .ZN(n6998) );
  NAND2_X1 U8664 ( .A1(n6998), .A2(n6988), .ZN(n6907) );
  NAND3_X1 U8665 ( .A1(n6915), .A2(n8846), .A3(n8858), .ZN(n6908) );
  MUX2_X1 U8666 ( .A(n6909), .B(n6908), .S(n6988), .Z(n6923) );
  NAND2_X1 U8667 ( .A1(n6911), .A2(n6910), .ZN(n6913) );
  NAND3_X1 U8668 ( .A1(n6913), .A2(n6980), .A3(n6912), .ZN(n6914) );
  AOI21_X1 U8669 ( .B1(n6915), .B2(n6914), .A(n4613), .ZN(n6922) );
  AND2_X1 U8670 ( .A1(n6924), .A2(n6916), .ZN(n6920) );
  INV_X1 U8671 ( .A(n6917), .ZN(n6918) );
  NOR2_X1 U8672 ( .A1(n8835), .A2(n6918), .ZN(n6919) );
  MUX2_X1 U8673 ( .A(n6920), .B(n6919), .S(n6980), .Z(n6921) );
  NAND2_X1 U8674 ( .A1(n6925), .A2(n6924), .ZN(n6926) );
  AOI21_X1 U8675 ( .B1(n6928), .B2(n6927), .A(n6980), .ZN(n6931) );
  AOI21_X1 U8676 ( .B1(n6988), .B2(n6929), .A(n8811), .ZN(n6930) );
  MUX2_X1 U8677 ( .A(n6932), .B(n8791), .S(n6980), .Z(n6933) );
  INV_X1 U8678 ( .A(n6933), .ZN(n6934) );
  NAND4_X1 U8679 ( .A1(n6942), .A2(n6988), .A3(n6996), .A4(n6938), .ZN(n6935)
         );
  NAND2_X1 U8680 ( .A1(n6955), .A2(n6980), .ZN(n6940) );
  NAND3_X1 U8681 ( .A1(n6942), .A2(n6980), .A3(n6938), .ZN(n6939) );
  OAI211_X1 U8682 ( .C1(n6988), .C2(n6953), .A(n6940), .B(n6939), .ZN(n6947)
         );
  INV_X1 U8683 ( .A(n6952), .ZN(n6941) );
  INV_X1 U8684 ( .A(n6942), .ZN(n6943) );
  INV_X1 U8685 ( .A(n6949), .ZN(n6951) );
  NAND4_X1 U8686 ( .A1(n6953), .A2(n6980), .A3(n6952), .A4(n6995), .ZN(n6954)
         );
  NAND2_X1 U8687 ( .A1(n6956), .A2(n6988), .ZN(n6957) );
  MUX2_X1 U8688 ( .A(n8759), .B(n8480), .S(n6980), .Z(n6974) );
  INV_X1 U8689 ( .A(n6974), .ZN(n6961) );
  NAND2_X1 U8690 ( .A1(n9981), .A2(n5988), .ZN(n6964) );
  INV_X1 U8691 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9078) );
  OR2_X1 U8692 ( .A1(n6976), .A2(n9078), .ZN(n6963) );
  INV_X1 U8693 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6970) );
  NAND2_X1 U8694 ( .A1(n5958), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6968) );
  INV_X1 U8695 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n6965) );
  OR2_X1 U8696 ( .A1(n6966), .A2(n6965), .ZN(n6967) );
  OAI211_X1 U8697 ( .C1(n6970), .C2(n6969), .A(n6968), .B(n6967), .ZN(n6971)
         );
  INV_X1 U8698 ( .A(n6971), .ZN(n6972) );
  OAI21_X1 U8699 ( .B1(n6991), .B2(n8480), .A(n7023), .ZN(n6985) );
  NAND2_X1 U8700 ( .A1(n6975), .A2(n6974), .ZN(n6989) );
  INV_X1 U8701 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8425) );
  NOR2_X1 U8702 ( .A1(n6976), .A2(n8425), .ZN(n6977) );
  NAND2_X1 U8703 ( .A1(n8986), .A2(n8604), .ZN(n7024) );
  NAND3_X1 U8704 ( .A1(n6989), .A2(n7024), .A3(n7020), .ZN(n6984) );
  INV_X1 U8705 ( .A(n7023), .ZN(n6982) );
  INV_X1 U8706 ( .A(n8986), .ZN(n6979) );
  INV_X1 U8707 ( .A(n8604), .ZN(n6978) );
  AND2_X1 U8708 ( .A1(n6979), .A2(n6978), .ZN(n6986) );
  OAI21_X1 U8709 ( .B1(n6986), .B2(n6980), .A(n7024), .ZN(n6981) );
  INV_X1 U8710 ( .A(n6986), .ZN(n7017) );
  NAND2_X1 U8711 ( .A1(n7017), .A2(n6987), .ZN(n7019) );
  NOR2_X1 U8712 ( .A1(n7019), .A2(n6988), .ZN(n6990) );
  OAI211_X1 U8713 ( .C1(n6991), .C2(n8759), .A(n6990), .B(n6989), .ZN(n6992)
         );
  INV_X1 U8714 ( .A(n8345), .ZN(n7030) );
  AND2_X1 U8715 ( .A1(n7030), .A2(n8212), .ZN(n6994) );
  INV_X1 U8716 ( .A(n8775), .ZN(n8781) );
  INV_X1 U8717 ( .A(n8793), .ZN(n6997) );
  INV_X1 U8718 ( .A(n6998), .ZN(n7012) );
  INV_X1 U8719 ( .A(n8906), .ZN(n8908) );
  NAND2_X1 U8720 ( .A1(n7000), .A2(n6999), .ZN(n8319) );
  NAND2_X1 U8721 ( .A1(n7001), .A2(n7730), .ZN(n7524) );
  XNOR2_X1 U8722 ( .A(n10092), .B(n7725), .ZN(n7796) );
  NAND2_X1 U8723 ( .A1(n7004), .A2(n7003), .ZN(n8054) );
  NAND2_X1 U8724 ( .A1(n8050), .A2(n7005), .ZN(n7971) );
  NAND2_X1 U8725 ( .A1(n7007), .A2(n7006), .ZN(n7993) );
  NAND4_X1 U8726 ( .A1(n8319), .A2(n8078), .A3(n7008), .A4(n8193), .ZN(n7009)
         );
  NOR4_X1 U8727 ( .A1(n8883), .A2(n4657), .A3(n8908), .A4(n7009), .ZN(n7010)
         );
  NAND4_X1 U8728 ( .A1(n8846), .A2(n7012), .A3(n7011), .A4(n7010), .ZN(n7013)
         );
  NOR4_X1 U8729 ( .A1(n8823), .A2(n8811), .A3(n8835), .A4(n7013), .ZN(n7014)
         );
  NAND4_X1 U8730 ( .A1(n8781), .A2(n8795), .A3(n8802), .A4(n7014), .ZN(n7015)
         );
  XNOR2_X1 U8731 ( .A(n8480), .B(n8759), .ZN(n7047) );
  NAND2_X1 U8732 ( .A1(n7027), .A2(n7026), .ZN(n7029) );
  NAND3_X1 U8733 ( .A1(n7034), .A2(n7033), .A3(n5895), .ZN(n7035) );
  OAI211_X1 U8734 ( .C1(n7036), .C2(n8345), .A(n7035), .B(P2_B_REG_SCAN_IN), 
        .ZN(n7037) );
  INV_X1 U8735 ( .A(n7041), .ZN(n7039) );
  NAND2_X1 U8736 ( .A1(n7039), .A2(n7047), .ZN(n7043) );
  INV_X1 U8737 ( .A(n7047), .ZN(n7040) );
  AOI21_X1 U8738 ( .B1(n7041), .B2(n7040), .A(n8894), .ZN(n7042) );
  NAND2_X1 U8739 ( .A1(n7043), .A2(n7042), .ZN(n7045) );
  AOI22_X1 U8740 ( .A1(n8768), .A2(n10093), .B1(n8605), .B2(n10091), .ZN(n7044) );
  NAND2_X1 U8741 ( .A1(n7045), .A2(n7044), .ZN(n7309) );
  MUX2_X1 U8742 ( .A(n7309), .B(P2_REG0_REG_28__SCAN_IN), .S(n10154), .Z(n7046) );
  INV_X1 U8743 ( .A(n7046), .ZN(n7051) );
  XNOR2_X1 U8744 ( .A(n7048), .B(n7047), .ZN(n7312) );
  OAI22_X1 U8745 ( .A1(n7312), .A2(n9074), .B1(n7053), .B2(n9055), .ZN(n7049)
         );
  INV_X1 U8746 ( .A(n7049), .ZN(n7050) );
  NAND2_X1 U8747 ( .A1(n7051), .A2(n7050), .ZN(P2_U3455) );
  MUX2_X1 U8748 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n7309), .S(n10166), .Z(n7052) );
  INV_X1 U8749 ( .A(n7052), .ZN(n7056) );
  OAI22_X1 U8750 ( .A1(n7312), .A2(n8975), .B1(n7053), .B2(n8961), .ZN(n7054)
         );
  INV_X1 U8751 ( .A(n7054), .ZN(n7055) );
  NAND2_X1 U8752 ( .A1(n7056), .A2(n7055), .ZN(P2_U3487) );
  INV_X1 U8753 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7057) );
  OAI21_X1 U8754 ( .B1(n7061), .B2(n7060), .A(n7059), .ZN(P1_U3550) );
  NAND2_X1 U8755 ( .A1(n7063), .A2(n7062), .ZN(n7935) );
  NAND2_X1 U8756 ( .A1(n7068), .A2(n9801), .ZN(n7069) );
  OR2_X4 U8757 ( .A1(n7069), .A2(n7070), .ZN(n7270) );
  OR2_X2 U8758 ( .A1(n7070), .A2(n9801), .ZN(n7273) );
  OAI22_X1 U8759 ( .A1(n7110), .A2(n7715), .B1(n7071), .B2(n7273), .ZN(n7072)
         );
  AOI21_X1 U8760 ( .B1(n7070), .B2(P1_REG1_REG_0__SCAN_IN), .A(n7072), .ZN(
        n7713) );
  AOI222_X1 U8761 ( .A1(n6693), .A2(n7260), .B1(n7096), .B2(n7836), .C1(n7070), 
        .C2(P1_IR_REG_0__SCAN_IN), .ZN(n7714) );
  OAI22_X1 U8762 ( .A1(n7713), .A2(n7714), .B1(n7270), .B2(n7072), .ZN(n7758)
         );
  NAND2_X1 U8763 ( .A1(n7096), .A2(n9375), .ZN(n7074) );
  INV_X2 U8764 ( .A(n7270), .ZN(n8401) );
  XNOR2_X1 U8765 ( .A(n7075), .B(n8401), .ZN(n7079) );
  OR2_X1 U8766 ( .A1(n8403), .A2(n7073), .ZN(n7077) );
  NAND2_X1 U8767 ( .A1(n7096), .A2(n4293), .ZN(n7076) );
  AND2_X1 U8768 ( .A1(n7077), .A2(n7076), .ZN(n7078) );
  OAI21_X1 U8769 ( .B1(n7079), .B2(n7078), .A(n7080), .ZN(n7759) );
  INV_X1 U8770 ( .A(n7080), .ZN(n7808) );
  NAND2_X1 U8771 ( .A1(n8398), .A2(n7813), .ZN(n7082) );
  NAND2_X1 U8772 ( .A1(n7096), .A2(n9374), .ZN(n7081) );
  NAND2_X1 U8773 ( .A1(n7082), .A2(n7081), .ZN(n7083) );
  XNOR2_X1 U8774 ( .A(n7083), .B(n8401), .ZN(n7087) );
  INV_X1 U8775 ( .A(n9374), .ZN(n7084) );
  OR2_X1 U8776 ( .A1(n8403), .A2(n7084), .ZN(n7086) );
  NAND2_X1 U8777 ( .A1(n8406), .A2(n7813), .ZN(n7085) );
  AND2_X1 U8778 ( .A1(n7086), .A2(n7085), .ZN(n7088) );
  NAND2_X1 U8779 ( .A1(n7087), .A2(n7088), .ZN(n7092) );
  INV_X1 U8780 ( .A(n7087), .ZN(n7090) );
  INV_X1 U8781 ( .A(n7088), .ZN(n7089) );
  NAND2_X1 U8782 ( .A1(n7090), .A2(n7089), .ZN(n7091) );
  AND2_X1 U8783 ( .A1(n7092), .A2(n7091), .ZN(n7807) );
  OAI21_X2 U8784 ( .B1(n7809), .B2(n7808), .A(n7807), .ZN(n7806) );
  NAND2_X1 U8785 ( .A1(n7806), .A2(n7092), .ZN(n9137) );
  OAI22_X1 U8786 ( .A1(n8403), .A2(n7812), .B1(n7862), .B2(n7273), .ZN(n7102)
         );
  INV_X1 U8787 ( .A(n7862), .ZN(n10330) );
  NAND2_X1 U8788 ( .A1(n7246), .A2(n10330), .ZN(n7094) );
  NAND2_X1 U8789 ( .A1(n8406), .A2(n5084), .ZN(n7093) );
  NAND2_X1 U8790 ( .A1(n7094), .A2(n7093), .ZN(n7095) );
  XNOR2_X1 U8791 ( .A(n7095), .B(n7270), .ZN(n7101) );
  XOR2_X1 U8792 ( .A(n7102), .B(n7101), .Z(n9138) );
  NAND2_X1 U8793 ( .A1(n9137), .A2(n9138), .ZN(n9136) );
  AOI22_X1 U8794 ( .A1(n8398), .A2(n8044), .B1(n7204), .B2(n9373), .ZN(n7097)
         );
  XNOR2_X1 U8795 ( .A(n7097), .B(n7270), .ZN(n7108) );
  INV_X1 U8796 ( .A(n9373), .ZN(n7098) );
  OR2_X1 U8797 ( .A1(n8403), .A2(n7098), .ZN(n7100) );
  NAND2_X1 U8798 ( .A1(n7204), .A2(n8044), .ZN(n7099) );
  NAND2_X1 U8799 ( .A1(n7100), .A2(n7099), .ZN(n7106) );
  XNOR2_X1 U8800 ( .A(n7108), .B(n7106), .ZN(n7918) );
  INV_X1 U8801 ( .A(n7101), .ZN(n7104) );
  INV_X1 U8802 ( .A(n7102), .ZN(n7103) );
  NAND2_X1 U8803 ( .A1(n7104), .A2(n7103), .ZN(n7916) );
  INV_X1 U8804 ( .A(n7106), .ZN(n7107) );
  OR2_X1 U8805 ( .A1(n7108), .A2(n7107), .ZN(n7109) );
  OAI22_X1 U8806 ( .A1(n7110), .A2(n10057), .B1(n7111), .B2(n7273), .ZN(n7112)
         );
  XNOR2_X1 U8807 ( .A(n7112), .B(n7270), .ZN(n7113) );
  INV_X1 U8808 ( .A(n10057), .ZN(n8206) );
  AOI22_X1 U8809 ( .A1(n7260), .A2(n9372), .B1(n7204), .B2(n8206), .ZN(n8200)
         );
  NAND2_X1 U8810 ( .A1(n7246), .A2(n8219), .ZN(n7115) );
  NAND2_X1 U8811 ( .A1(n7204), .A2(n9371), .ZN(n7114) );
  NAND2_X1 U8812 ( .A1(n7115), .A2(n7114), .ZN(n7116) );
  XNOR2_X1 U8813 ( .A(n7116), .B(n7270), .ZN(n7121) );
  INV_X1 U8814 ( .A(n9371), .ZN(n7117) );
  OR2_X1 U8815 ( .A1(n8403), .A2(n7117), .ZN(n7119) );
  NAND2_X1 U8816 ( .A1(n7204), .A2(n8219), .ZN(n7118) );
  NAND2_X1 U8817 ( .A1(n7119), .A2(n7118), .ZN(n7120) );
  NOR2_X1 U8818 ( .A1(n7121), .A2(n7120), .ZN(n7122) );
  AOI21_X1 U8819 ( .B1(n7121), .B2(n7120), .A(n7122), .ZN(n8228) );
  NAND2_X1 U8820 ( .A1(n4284), .A2(n8228), .ZN(n8227) );
  INV_X1 U8821 ( .A(n7122), .ZN(n7123) );
  NAND2_X1 U8822 ( .A1(n8227), .A2(n7123), .ZN(n8328) );
  NAND2_X1 U8823 ( .A1(n7246), .A2(n10063), .ZN(n7125) );
  NAND2_X1 U8824 ( .A1(n7204), .A2(n9370), .ZN(n7124) );
  NAND2_X1 U8825 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  XNOR2_X1 U8826 ( .A(n7126), .B(n8401), .ZN(n7130) );
  INV_X1 U8827 ( .A(n9370), .ZN(n7127) );
  OR2_X1 U8828 ( .A1(n8403), .A2(n7127), .ZN(n7129) );
  NAND2_X1 U8829 ( .A1(n7204), .A2(n10063), .ZN(n7128) );
  AND2_X1 U8830 ( .A1(n7129), .A2(n7128), .ZN(n7131) );
  AND2_X1 U8831 ( .A1(n7130), .A2(n7131), .ZN(n8324) );
  INV_X1 U8832 ( .A(n7130), .ZN(n7133) );
  INV_X1 U8833 ( .A(n7131), .ZN(n7132) );
  NAND2_X1 U8834 ( .A1(n7133), .A2(n7132), .ZN(n8325) );
  OR2_X1 U8835 ( .A1(n8403), .A2(n7134), .ZN(n7136) );
  NAND2_X1 U8836 ( .A1(n7204), .A2(n9172), .ZN(n7135) );
  NAND2_X1 U8837 ( .A1(n7136), .A2(n7135), .ZN(n7144) );
  INV_X1 U8838 ( .A(n7144), .ZN(n9167) );
  NAND2_X1 U8839 ( .A1(n8398), .A2(n9172), .ZN(n7138) );
  NAND2_X1 U8840 ( .A1(n7204), .A2(n9369), .ZN(n7137) );
  NAND2_X1 U8841 ( .A1(n7138), .A2(n7137), .ZN(n7139) );
  XNOR2_X1 U8842 ( .A(n7139), .B(n7270), .ZN(n9251) );
  INV_X1 U8843 ( .A(n9251), .ZN(n9165) );
  NAND2_X1 U8844 ( .A1(n7246), .A2(n4435), .ZN(n7141) );
  NAND2_X1 U8845 ( .A1(n7204), .A2(n9368), .ZN(n7140) );
  NAND2_X1 U8846 ( .A1(n7141), .A2(n7140), .ZN(n7142) );
  XNOR2_X1 U8847 ( .A(n7142), .B(n8401), .ZN(n7147) );
  INV_X1 U8848 ( .A(n7147), .ZN(n9249) );
  NAND2_X1 U8849 ( .A1(n9249), .A2(n9248), .ZN(n9247) );
  OAI21_X1 U8850 ( .B1(n9167), .B2(n9165), .A(n9247), .ZN(n7149) );
  OAI21_X1 U8851 ( .B1(n9251), .B2(n7144), .A(n9248), .ZN(n7146) );
  NOR3_X1 U8852 ( .A1(n9251), .A2(n9248), .A3(n7144), .ZN(n7145) );
  AOI21_X1 U8853 ( .B1(n7147), .B2(n7146), .A(n7145), .ZN(n7148) );
  NAND2_X1 U8854 ( .A1(n9133), .A2(n7246), .ZN(n7151) );
  NAND2_X1 U8855 ( .A1(n7204), .A2(n9367), .ZN(n7150) );
  NAND2_X1 U8856 ( .A1(n7151), .A2(n7150), .ZN(n7152) );
  XNOR2_X1 U8857 ( .A(n7152), .B(n7270), .ZN(n9124) );
  NAND2_X1 U8858 ( .A1(n9133), .A2(n8406), .ZN(n7155) );
  OR2_X1 U8859 ( .A1(n8403), .A2(n7153), .ZN(n7154) );
  NAND2_X1 U8860 ( .A1(n7155), .A2(n7154), .ZN(n9128) );
  NOR2_X1 U8861 ( .A1(n9124), .A2(n9128), .ZN(n7163) );
  NAND2_X1 U8862 ( .A1(n9885), .A2(n7246), .ZN(n7157) );
  NAND2_X1 U8863 ( .A1(n7204), .A2(n9366), .ZN(n7156) );
  NAND2_X1 U8864 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  XNOR2_X1 U8865 ( .A(n7158), .B(n8401), .ZN(n7161) );
  NOR2_X1 U8866 ( .A1(n8403), .A2(n8288), .ZN(n7159) );
  AOI21_X1 U8867 ( .B1(n9885), .B2(n8406), .A(n7159), .ZN(n7160) );
  NAND2_X1 U8868 ( .A1(n7161), .A2(n7160), .ZN(n9194) );
  OAI21_X1 U8869 ( .B1(n7161), .B2(n7160), .A(n9194), .ZN(n9297) );
  AOI21_X1 U8870 ( .B1(n9124), .B2(n9128), .A(n9297), .ZN(n7162) );
  NAND2_X1 U8871 ( .A1(n8354), .A2(n7246), .ZN(n7165) );
  NAND2_X1 U8872 ( .A1(n7204), .A2(n9365), .ZN(n7164) );
  NAND2_X1 U8873 ( .A1(n7165), .A2(n7164), .ZN(n7166) );
  XNOR2_X1 U8874 ( .A(n7166), .B(n8401), .ZN(n7169) );
  NOR2_X1 U8875 ( .A1(n8403), .A2(n8304), .ZN(n7167) );
  AOI21_X1 U8876 ( .B1(n8354), .B2(n8406), .A(n7167), .ZN(n7168) );
  NAND2_X1 U8877 ( .A1(n7169), .A2(n7168), .ZN(n9274) );
  OR2_X1 U8878 ( .A1(n7169), .A2(n7168), .ZN(n7170) );
  AND2_X1 U8879 ( .A1(n9274), .A2(n7170), .ZN(n9195) );
  NAND2_X1 U8880 ( .A1(n7171), .A2(n9195), .ZN(n9196) );
  NAND2_X1 U8881 ( .A1(n9196), .A2(n9274), .ZN(n7179) );
  NAND2_X1 U8882 ( .A1(n9880), .A2(n7246), .ZN(n7173) );
  NAND2_X1 U8883 ( .A1(n7204), .A2(n9364), .ZN(n7172) );
  NAND2_X1 U8884 ( .A1(n7173), .A2(n7172), .ZN(n7174) );
  XNOR2_X1 U8885 ( .A(n7174), .B(n8401), .ZN(n7177) );
  NOR2_X1 U8886 ( .A1(n8403), .A2(n8287), .ZN(n7175) );
  AOI21_X1 U8887 ( .B1(n9880), .B2(n8406), .A(n7175), .ZN(n7176) );
  NAND2_X1 U8888 ( .A1(n7177), .A2(n7176), .ZN(n7180) );
  OR2_X1 U8889 ( .A1(n7177), .A2(n7176), .ZN(n7178) );
  AND2_X1 U8890 ( .A1(n7180), .A2(n7178), .ZN(n9275) );
  NAND2_X1 U8891 ( .A1(n7179), .A2(n9275), .ZN(n9278) );
  NAND2_X1 U8892 ( .A1(n9278), .A2(n7180), .ZN(n7183) );
  OAI22_X1 U8893 ( .A1(n7182), .A2(n7110), .B1(n9338), .B2(n7273), .ZN(n7181)
         );
  XOR2_X1 U8894 ( .A(n7270), .B(n7181), .Z(n7184) );
  OAI22_X1 U8895 ( .A1(n7182), .A2(n7273), .B1(n9338), .B2(n8403), .ZN(n9104)
         );
  NAND2_X1 U8896 ( .A1(n9843), .A2(n7246), .ZN(n7186) );
  NAND2_X1 U8897 ( .A1(n9357), .A2(n8406), .ZN(n7185) );
  NAND2_X1 U8898 ( .A1(n7186), .A2(n7185), .ZN(n7187) );
  XNOR2_X1 U8899 ( .A(n7187), .B(n7270), .ZN(n7198) );
  NAND2_X1 U8900 ( .A1(n9843), .A2(n8406), .ZN(n7189) );
  NAND2_X1 U8901 ( .A1(n9357), .A2(n7260), .ZN(n7188) );
  NAND2_X1 U8902 ( .A1(n7189), .A2(n7188), .ZN(n7197) );
  NAND2_X1 U8903 ( .A1(n7198), .A2(n7197), .ZN(n7219) );
  AOI22_X1 U8904 ( .A1(n9852), .A2(n7246), .B1(n7204), .B2(n9359), .ZN(n7190)
         );
  XNOR2_X1 U8905 ( .A(n7190), .B(n7270), .ZN(n9177) );
  AOI22_X1 U8906 ( .A1(n9852), .A2(n8406), .B1(n7260), .B2(n9359), .ZN(n9178)
         );
  NOR2_X1 U8907 ( .A1(n9313), .A2(n8403), .ZN(n7191) );
  AOI21_X1 U8908 ( .B1(n9847), .B2(n8406), .A(n7191), .ZN(n7225) );
  AOI21_X1 U8909 ( .B1(n9177), .B2(n9178), .A(n7225), .ZN(n7196) );
  NAND2_X1 U8910 ( .A1(n9847), .A2(n8398), .ZN(n7193) );
  NAND2_X1 U8911 ( .A1(n7204), .A2(n9358), .ZN(n7192) );
  NAND2_X1 U8912 ( .A1(n7193), .A2(n7192), .ZN(n7194) );
  XNOR2_X1 U8913 ( .A(n7194), .B(n7270), .ZN(n9155) );
  NAND3_X1 U8914 ( .A1(n7225), .A2(n9177), .A3(n9178), .ZN(n7195) );
  OAI21_X1 U8915 ( .B1(n7196), .B2(n9155), .A(n7195), .ZN(n7199) );
  NOR2_X1 U8916 ( .A1(n7198), .A2(n7197), .ZN(n9184) );
  NAND2_X1 U8917 ( .A1(n9870), .A2(n8398), .ZN(n7201) );
  NAND2_X1 U8918 ( .A1(n8406), .A2(n9362), .ZN(n7200) );
  NAND2_X1 U8919 ( .A1(n7201), .A2(n7200), .ZN(n7202) );
  XNOR2_X1 U8920 ( .A(n7202), .B(n8401), .ZN(n9146) );
  AOI22_X1 U8921 ( .A1(n9870), .A2(n8406), .B1(n7260), .B2(n9362), .ZN(n7220)
         );
  NAND2_X1 U8922 ( .A1(n9146), .A2(n7220), .ZN(n7213) );
  NOR2_X1 U8923 ( .A1(n8403), .A2(n9312), .ZN(n7203) );
  AOI21_X1 U8924 ( .B1(n9951), .B2(n8406), .A(n7203), .ZN(n7222) );
  NAND2_X1 U8925 ( .A1(n9951), .A2(n7246), .ZN(n7206) );
  NAND2_X1 U8926 ( .A1(n7204), .A2(n9360), .ZN(n7205) );
  NAND2_X1 U8927 ( .A1(n7206), .A2(n7205), .ZN(n7207) );
  XNOR2_X1 U8928 ( .A(n7207), .B(n7270), .ZN(n7224) );
  XOR2_X1 U8929 ( .A(n7222), .B(n7224), .Z(n9227) );
  NAND2_X1 U8930 ( .A1(n9861), .A2(n7246), .ZN(n7209) );
  NAND2_X1 U8931 ( .A1(n8406), .A2(n9361), .ZN(n7208) );
  NAND2_X1 U8932 ( .A1(n7209), .A2(n7208), .ZN(n7210) );
  XNOR2_X1 U8933 ( .A(n7210), .B(n7270), .ZN(n9218) );
  NAND2_X1 U8934 ( .A1(n9861), .A2(n8406), .ZN(n7212) );
  OR2_X1 U8935 ( .A1(n8403), .A2(n9335), .ZN(n7211) );
  NAND2_X1 U8936 ( .A1(n7212), .A2(n7211), .ZN(n9217) );
  NOR2_X1 U8937 ( .A1(n9218), .A2(n9217), .ZN(n9228) );
  NOR2_X1 U8938 ( .A1(n9227), .A2(n9228), .ZN(n7221) );
  NAND2_X1 U8939 ( .A1(n7218), .A2(n8398), .ZN(n7215) );
  NAND2_X1 U8940 ( .A1(n9356), .A2(n8406), .ZN(n7214) );
  AND2_X1 U8941 ( .A1(n9356), .A2(n7260), .ZN(n7217) );
  AOI21_X1 U8942 ( .B1(n7218), .B2(n8406), .A(n7217), .ZN(n7233) );
  XNOR2_X1 U8943 ( .A(n7235), .B(n7233), .ZN(n9185) );
  INV_X1 U8944 ( .A(n7219), .ZN(n9183) );
  INV_X1 U8945 ( .A(n9146), .ZN(n9145) );
  INV_X1 U8946 ( .A(n7220), .ZN(n9334) );
  AOI21_X1 U8947 ( .B1(n9145), .B2(n9334), .A(n9148), .ZN(n7227) );
  INV_X1 U8948 ( .A(n7221), .ZN(n9150) );
  INV_X1 U8949 ( .A(n9177), .ZN(n9153) );
  INV_X1 U8950 ( .A(n9178), .ZN(n9310) );
  INV_X1 U8951 ( .A(n7222), .ZN(n7223) );
  AOI21_X1 U8952 ( .B1(n9153), .B2(n9310), .A(n9152), .ZN(n7226) );
  INV_X1 U8953 ( .A(n7225), .ZN(n9154) );
  NAND2_X1 U8954 ( .A1(n9155), .A2(n9154), .ZN(n9265) );
  OAI211_X1 U8955 ( .C1(n7227), .C2(n9150), .A(n7226), .B(n9265), .ZN(n7229)
         );
  OAI21_X1 U8956 ( .B1(n9183), .B2(n7229), .A(n7228), .ZN(n7230) );
  INV_X1 U8957 ( .A(n7233), .ZN(n7234) );
  NAND2_X1 U8958 ( .A1(n9186), .A2(n7236), .ZN(n7239) );
  OAI22_X1 U8959 ( .A1(n9931), .A2(n7110), .B1(n9118), .B2(n7273), .ZN(n7237)
         );
  XOR2_X1 U8960 ( .A(n7270), .B(n7237), .Z(n7238) );
  OAI22_X1 U8961 ( .A1(n9931), .A2(n7273), .B1(n9118), .B2(n8403), .ZN(n9290)
         );
  NAND2_X1 U8962 ( .A1(n9922), .A2(n8398), .ZN(n7241) );
  NAND2_X1 U8963 ( .A1(n9354), .A2(n7204), .ZN(n7240) );
  NAND2_X1 U8964 ( .A1(n7241), .A2(n7240), .ZN(n7242) );
  XNOR2_X1 U8965 ( .A(n7242), .B(n8401), .ZN(n7245) );
  NOR2_X1 U8966 ( .A1(n9292), .A2(n8403), .ZN(n7243) );
  AOI21_X1 U8967 ( .B1(n9922), .B2(n8406), .A(n7243), .ZN(n7244) );
  OR2_X1 U8968 ( .A1(n7245), .A2(n7244), .ZN(n9114) );
  NAND2_X1 U8969 ( .A1(n7245), .A2(n7244), .ZN(n9116) );
  NAND2_X1 U8970 ( .A1(n9112), .A2(n9116), .ZN(n9236) );
  NAND2_X1 U8971 ( .A1(n9920), .A2(n7246), .ZN(n7248) );
  NAND2_X1 U8972 ( .A1(n9353), .A2(n8406), .ZN(n7247) );
  NAND2_X1 U8973 ( .A1(n7248), .A2(n7247), .ZN(n7249) );
  XNOR2_X1 U8974 ( .A(n7249), .B(n7270), .ZN(n7252) );
  AOI22_X1 U8975 ( .A1(n9920), .A2(n8406), .B1(n7260), .B2(n9353), .ZN(n7250)
         );
  XNOR2_X1 U8976 ( .A(n7252), .B(n7250), .ZN(n9237) );
  INV_X1 U8977 ( .A(n7250), .ZN(n7251) );
  OR2_X1 U8978 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  OAI22_X1 U8979 ( .A1(n9913), .A2(n7273), .B1(n7254), .B2(n8403), .ZN(n7258)
         );
  NAND2_X1 U8980 ( .A1(n9211), .A2(n8398), .ZN(n7256) );
  NAND2_X1 U8981 ( .A1(n9352), .A2(n7204), .ZN(n7255) );
  NAND2_X1 U8982 ( .A1(n7256), .A2(n7255), .ZN(n7257) );
  XNOR2_X1 U8983 ( .A(n7257), .B(n7270), .ZN(n7259) );
  XOR2_X1 U8984 ( .A(n7258), .B(n7259), .Z(n9206) );
  INV_X1 U8985 ( .A(n9318), .ZN(n7266) );
  AND2_X1 U8986 ( .A1(n9351), .A2(n7260), .ZN(n7261) );
  AOI21_X1 U8987 ( .B1(n9814), .B2(n8406), .A(n7261), .ZN(n7267) );
  NAND2_X1 U8988 ( .A1(n9814), .A2(n8398), .ZN(n7263) );
  NAND2_X1 U8989 ( .A1(n9351), .A2(n7204), .ZN(n7262) );
  NAND2_X1 U8990 ( .A1(n7263), .A2(n7262), .ZN(n7264) );
  XNOR2_X1 U8991 ( .A(n7264), .B(n7270), .ZN(n7269) );
  XOR2_X1 U8992 ( .A(n7267), .B(n7269), .Z(n9319) );
  INV_X1 U8993 ( .A(n9319), .ZN(n7265) );
  INV_X1 U8994 ( .A(n7267), .ZN(n7268) );
  NAND2_X1 U8995 ( .A1(n7269), .A2(n7268), .ZN(n7276) );
  NAND2_X1 U8996 ( .A1(n9320), .A2(n7276), .ZN(n7275) );
  OAI22_X1 U8997 ( .A1(n9908), .A2(n7110), .B1(n7272), .B2(n7273), .ZN(n7271)
         );
  XNOR2_X1 U8998 ( .A(n7271), .B(n7270), .ZN(n8411) );
  OAI22_X1 U8999 ( .A1(n9908), .A2(n7273), .B1(n7272), .B2(n8403), .ZN(n8410)
         );
  XNOR2_X1 U9000 ( .A(n8411), .B(n8410), .ZN(n7274) );
  INV_X1 U9001 ( .A(n7274), .ZN(n7277) );
  AND2_X1 U9002 ( .A1(n7277), .A2(n7276), .ZN(n7278) );
  INV_X1 U9003 ( .A(n7279), .ZN(n7329) );
  NAND3_X1 U9004 ( .A1(n7329), .A2(n7327), .A3(n7280), .ZN(n7298) );
  INV_X1 U9005 ( .A(n10064), .ZN(n10056) );
  NAND3_X1 U9006 ( .A1(n7296), .A2(n7287), .A3(n10056), .ZN(n7281) );
  NAND2_X1 U9007 ( .A1(n7296), .A2(n7332), .ZN(n7283) );
  OR2_X1 U9008 ( .A1(n7298), .A2(n7283), .ZN(n7286) );
  NAND2_X1 U9009 ( .A1(n7298), .A2(n10056), .ZN(n7288) );
  MUX2_X1 U9010 ( .A(n7065), .B(n7288), .S(n7287), .Z(n7289) );
  NAND2_X1 U9011 ( .A1(n7289), .A2(n7067), .ZN(n7712) );
  NAND2_X1 U9012 ( .A1(n7712), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7294) );
  AND2_X1 U9013 ( .A1(n7332), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7290) );
  OR2_X1 U9014 ( .A1(n7291), .A2(n7290), .ZN(n7292) );
  NAND2_X1 U9015 ( .A1(n7298), .A2(n7292), .ZN(n7709) );
  AND2_X1 U9016 ( .A1(n7709), .A2(n7444), .ZN(n7293) );
  INV_X1 U9017 ( .A(n7295), .ZN(n7300) );
  NAND2_X1 U9018 ( .A1(n7296), .A2(n7065), .ZN(n7297) );
  OAI22_X1 U9019 ( .A1(n7300), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7299), .ZN(n7301) );
  AOI21_X1 U9020 ( .B1(n9585), .B2(n9328), .A(n7301), .ZN(n7302) );
  INV_X1 U9021 ( .A(n7304), .ZN(n7307) );
  NAND3_X1 U9022 ( .A1(n7307), .A2(n7306), .A3(n7305), .ZN(n7313) );
  INV_X2 U9023 ( .A(n10107), .ZN(n7308) );
  NAND2_X1 U9024 ( .A1(n7309), .A2(n7308), .ZN(n7317) );
  OR2_X1 U9025 ( .A1(n7310), .A2(n6341), .ZN(n7794) );
  AND2_X1 U9026 ( .A1(n8059), .A2(n7794), .ZN(n7311) );
  AOI22_X1 U9027 ( .A1(n8480), .A2(n10101), .B1(n10102), .B2(n8476), .ZN(n7315) );
  NAND2_X1 U9028 ( .A1(n10107), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U9029 ( .A1(n7317), .A2(n4964), .ZN(P2_U3205) );
  INV_X1 U9030 ( .A(n7318), .ZN(n7319) );
  OR2_X1 U9031 ( .A1(n6760), .A2(n7319), .ZN(n7830) );
  NAND2_X1 U9032 ( .A1(n6760), .A2(n7319), .ZN(n7320) );
  NAND2_X1 U9033 ( .A1(n7830), .A2(n7320), .ZN(n7882) );
  INV_X1 U9034 ( .A(n7882), .ZN(n7338) );
  OAI21_X1 U9035 ( .B1(n7322), .B2(n6760), .A(n7321), .ZN(n7325) );
  NAND2_X1 U9036 ( .A1(n9322), .A2(n6693), .ZN(n7324) );
  NAND2_X1 U9037 ( .A1(n9324), .A2(n9374), .ZN(n7323) );
  NAND2_X1 U9038 ( .A1(n7324), .A2(n7323), .ZN(n7760) );
  AOI21_X1 U9039 ( .B1(n7325), .B2(n9778), .A(n7760), .ZN(n7326) );
  OAI21_X1 U9040 ( .B1(n7338), .B2(n8264), .A(n7326), .ZN(n7880) );
  INV_X1 U9041 ( .A(n7327), .ZN(n7330) );
  NAND3_X1 U9042 ( .A1(n7330), .A2(n7329), .A3(n7328), .ZN(n7331) );
  INV_X2 U9043 ( .A(n10337), .ZN(n10344) );
  MUX2_X1 U9044 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n7880), .S(n10344), .Z(n7341)
         );
  OAI22_X1 U9045 ( .A1(n9715), .A2(n7334), .B1(n9780), .B2(n7333), .ZN(n7340)
         );
  INV_X1 U9046 ( .A(n7935), .ZN(n7335) );
  NAND2_X1 U9047 ( .A1(n10344), .A2(n7335), .ZN(n8271) );
  XNOR2_X1 U9048 ( .A(n4293), .B(n7836), .ZN(n7336) );
  NOR2_X1 U9049 ( .A1(n9784), .A2(n7336), .ZN(n7881) );
  INV_X1 U9050 ( .A(n7881), .ZN(n7337) );
  OAI22_X1 U9051 ( .A1(n7338), .A2(n8271), .B1(n10341), .B2(n7337), .ZN(n7339)
         );
  OR3_X1 U9052 ( .A1(n7341), .A2(n7340), .A3(n7339), .ZN(P1_U3292) );
  NOR2_X1 U9053 ( .A1(n7342), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9988) );
  AOI22_X1 U9054 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n9988), .B1(n9409), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n7343) );
  OAI21_X1 U9055 ( .B1(n7346), .B2(n9994), .A(n7343), .ZN(P1_U3352) );
  INV_X2 U9056 ( .A(n9091), .ZN(n9097) );
  NOR2_X1 U9057 ( .A1(n7342), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9082) );
  OAI222_X1 U9058 ( .A1(n9097), .A2(n5072), .B1(n9093), .B2(n7346), .C1(
        P2_U3151), .C2(n7345), .ZN(P2_U3292) );
  INV_X1 U9059 ( .A(n7347), .ZN(n7351) );
  OAI222_X1 U9060 ( .A1(n9097), .A2(n7349), .B1(n9093), .B2(n7351), .C1(
        P2_U3151), .C2(n7348), .ZN(P2_U3291) );
  INV_X2 U9061 ( .A(n9988), .ZN(n9995) );
  OAI222_X1 U9062 ( .A1(n9995), .A2(n7350), .B1(n9994), .B2(n7357), .C1(
        P1_U3086), .C2(n4594), .ZN(P1_U3353) );
  INV_X1 U9063 ( .A(n9422), .ZN(n7562) );
  OAI222_X1 U9064 ( .A1(n9995), .A2(n7352), .B1(n9994), .B2(n7351), .C1(
        P1_U3086), .C2(n7562), .ZN(P1_U3351) );
  INV_X1 U9065 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7353) );
  OAI222_X1 U9066 ( .A1(n9995), .A2(n7353), .B1(n9994), .B2(n7355), .C1(
        P1_U3086), .C2(n7557), .ZN(P1_U3354) );
  OAI222_X1 U9067 ( .A1(n7587), .A2(P2_U3151), .B1(n9093), .B2(n7355), .C1(
        n7354), .C2(n9097), .ZN(P2_U3294) );
  INV_X1 U9068 ( .A(n7358), .ZN(n7359) );
  OAI222_X1 U9069 ( .A1(n9097), .A2(n5119), .B1(n9093), .B2(n7359), .C1(
        P2_U3151), .C2(n7503), .ZN(P2_U3290) );
  INV_X1 U9070 ( .A(n9436), .ZN(n7563) );
  OAI222_X1 U9071 ( .A1(n9995), .A2(n5117), .B1(n9994), .B2(n7359), .C1(
        P1_U3086), .C2(n7563), .ZN(P1_U3350) );
  NAND2_X1 U9072 ( .A1(n6326), .A2(n7360), .ZN(n7381) );
  INV_X1 U9073 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7363) );
  NOR3_X1 U9074 ( .A1(n7364), .A2(n7365), .A3(n7361), .ZN(n7362) );
  AOI21_X1 U9075 ( .B1(n7381), .B2(n7363), .A(n7362), .ZN(P2_U3376) );
  NOR3_X1 U9076 ( .A1(n7366), .A2(n7365), .A3(n7364), .ZN(n7367) );
  AOI21_X1 U9077 ( .B1(n7381), .B2(n7368), .A(n7367), .ZN(P2_U3377) );
  INV_X1 U9078 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7370) );
  INV_X1 U9079 ( .A(n7369), .ZN(n7371) );
  OAI222_X1 U9080 ( .A1(n9097), .A2(n7370), .B1(n9093), .B2(n7371), .C1(
        P2_U3151), .C2(n7614), .ZN(P2_U3289) );
  INV_X1 U9081 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n7372) );
  INV_X1 U9082 ( .A(n9449), .ZN(n7565) );
  OAI222_X1 U9083 ( .A1(n9995), .A2(n7372), .B1(n9994), .B2(n7371), .C1(
        P1_U3086), .C2(n7565), .ZN(P1_U3349) );
  INV_X1 U9084 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7374) );
  INV_X1 U9085 ( .A(n7373), .ZN(n7375) );
  INV_X1 U9086 ( .A(n9462), .ZN(n7568) );
  OAI222_X1 U9087 ( .A1(n9995), .A2(n7374), .B1(n9994), .B2(n7375), .C1(
        P1_U3086), .C2(n7568), .ZN(P1_U3348) );
  INV_X1 U9088 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7376) );
  OAI222_X1 U9089 ( .A1(n9097), .A2(n7376), .B1(n9093), .B2(n7375), .C1(
        P2_U3151), .C2(n4742), .ZN(P2_U3288) );
  INV_X1 U9090 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U9091 ( .A1(n4673), .A2(P2_U3893), .ZN(n7377) );
  OAI21_X1 U9092 ( .B1(P2_U3893), .B2(n10230), .A(n7377), .ZN(P2_U3491) );
  INV_X1 U9093 ( .A(n7378), .ZN(n7379) );
  INV_X1 U9094 ( .A(n9475), .ZN(n7569) );
  OAI222_X1 U9095 ( .A1(n9995), .A2(n10190), .B1(n9994), .B2(n7379), .C1(
        P1_U3086), .C2(n7569), .ZN(P1_U3347) );
  OAI222_X1 U9096 ( .A1(n9097), .A2(n7380), .B1(n9093), .B2(n7379), .C1(
        P2_U3151), .C2(n5771), .ZN(P2_U3287) );
  INV_X1 U9097 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n7382) );
  NOR2_X1 U9098 ( .A1(n7400), .A2(n7382), .ZN(P2_U3247) );
  INV_X1 U9099 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n7383) );
  NOR2_X1 U9100 ( .A1(n7400), .A2(n7383), .ZN(P2_U3255) );
  INV_X1 U9101 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n7384) );
  NOR2_X1 U9102 ( .A1(n7400), .A2(n7384), .ZN(P2_U3250) );
  INV_X1 U9103 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n7385) );
  NOR2_X1 U9104 ( .A1(n7400), .A2(n7385), .ZN(P2_U3254) );
  INV_X1 U9105 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n7386) );
  NOR2_X1 U9106 ( .A1(n7400), .A2(n7386), .ZN(P2_U3253) );
  INV_X1 U9107 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n7387) );
  NOR2_X1 U9108 ( .A1(n7400), .A2(n7387), .ZN(P2_U3256) );
  INV_X1 U9109 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n7388) );
  NOR2_X1 U9110 ( .A1(n7400), .A2(n7388), .ZN(P2_U3257) );
  INV_X1 U9111 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n7389) );
  NOR2_X1 U9112 ( .A1(n7400), .A2(n7389), .ZN(P2_U3248) );
  INV_X1 U9113 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7390) );
  NOR2_X1 U9114 ( .A1(n7400), .A2(n7390), .ZN(P2_U3251) );
  INV_X1 U9115 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n7391) );
  NOR2_X1 U9116 ( .A1(n7400), .A2(n7391), .ZN(P2_U3252) );
  INV_X1 U9117 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n7392) );
  NOR2_X1 U9118 ( .A1(n7400), .A2(n7392), .ZN(P2_U3246) );
  INV_X1 U9119 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10243) );
  NOR2_X1 U9120 ( .A1(n7400), .A2(n10243), .ZN(P2_U3249) );
  INV_X1 U9121 ( .A(n7393), .ZN(n7395) );
  INV_X1 U9122 ( .A(n7556), .ZN(n7594) );
  OAI222_X1 U9123 ( .A1(n9994), .A2(n7395), .B1(n7594), .B2(P1_U3086), .C1(
        n7394), .C2(n9995), .ZN(P1_U3346) );
  OAI222_X1 U9124 ( .A1(n9097), .A2(n10289), .B1(n9093), .B2(n7395), .C1(n7699), .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U9125 ( .A(n7396), .ZN(n7399) );
  INV_X1 U9126 ( .A(n9494), .ZN(n7596) );
  OAI222_X1 U9127 ( .A1(n9994), .A2(n7399), .B1(n7596), .B2(P1_U3086), .C1(
        n7397), .C2(n9995), .ZN(P1_U3345) );
  OAI222_X1 U9128 ( .A1(n9097), .A2(n10261), .B1(n9093), .B2(n7399), .C1(n7398), .C2(P2_U3151), .ZN(P2_U3285) );
  INV_X1 U9129 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n7401) );
  NOR2_X1 U9130 ( .A1(n7400), .A2(n7401), .ZN(P2_U3238) );
  INV_X1 U9131 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n7402) );
  NOR2_X1 U9132 ( .A1(n7400), .A2(n7402), .ZN(P2_U3239) );
  INV_X1 U9133 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n7403) );
  NOR2_X1 U9134 ( .A1(n7400), .A2(n7403), .ZN(P2_U3241) );
  INV_X1 U9135 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U9136 ( .A1(n7400), .A2(n10271), .ZN(P2_U3243) );
  INV_X1 U9137 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n7404) );
  NOR2_X1 U9138 ( .A1(n7400), .A2(n7404), .ZN(P2_U3237) );
  INV_X1 U9139 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n7405) );
  NOR2_X1 U9140 ( .A1(n7400), .A2(n7405), .ZN(P2_U3259) );
  INV_X1 U9141 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n7406) );
  NOR2_X1 U9142 ( .A1(n7400), .A2(n7406), .ZN(P2_U3245) );
  INV_X1 U9143 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n7407) );
  NOR2_X1 U9144 ( .A1(n7400), .A2(n7407), .ZN(P2_U3261) );
  INV_X1 U9145 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n7408) );
  NOR2_X1 U9146 ( .A1(n7400), .A2(n7408), .ZN(P2_U3262) );
  INV_X1 U9147 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n7409) );
  NOR2_X1 U9148 ( .A1(n7400), .A2(n7409), .ZN(P2_U3263) );
  INV_X1 U9149 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7410) );
  NOR2_X1 U9150 ( .A1(n7400), .A2(n7410), .ZN(P2_U3242) );
  INV_X1 U9151 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n7411) );
  NOR2_X1 U9152 ( .A1(n7400), .A2(n7411), .ZN(P2_U3234) );
  INV_X1 U9153 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n7412) );
  NOR2_X1 U9154 ( .A1(n7400), .A2(n7412), .ZN(P2_U3235) );
  INV_X1 U9155 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n7413) );
  NOR2_X1 U9156 ( .A1(n7400), .A2(n7413), .ZN(P2_U3244) );
  INV_X1 U9157 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n7414) );
  NOR2_X1 U9158 ( .A1(n7400), .A2(n7414), .ZN(P2_U3240) );
  INV_X1 U9159 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n7415) );
  NOR2_X1 U9160 ( .A1(n7400), .A2(n7415), .ZN(P2_U3258) );
  INV_X1 U9161 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n7416) );
  NOR2_X1 U9162 ( .A1(n7400), .A2(n7416), .ZN(P2_U3236) );
  INV_X1 U9163 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n7417) );
  NOR2_X1 U9164 ( .A1(n7400), .A2(n7417), .ZN(P2_U3260) );
  INV_X1 U9165 ( .A(n7418), .ZN(n7420) );
  OAI222_X1 U9166 ( .A1(n9097), .A2(n7419), .B1(n9093), .B2(n7420), .C1(
        P2_U3151), .C2(n7910), .ZN(P2_U3284) );
  INV_X1 U9167 ( .A(n9508), .ZN(n7597) );
  OAI222_X1 U9168 ( .A1(n9995), .A2(n7421), .B1(n9994), .B2(n7420), .C1(
        P1_U3086), .C2(n7597), .ZN(P1_U3344) );
  INV_X1 U9169 ( .A(n7422), .ZN(n7425) );
  OAI222_X1 U9170 ( .A1(n9994), .A2(n7425), .B1(n7665), .B2(P1_U3086), .C1(
        n7423), .C2(n9995), .ZN(P1_U3343) );
  OAI222_X1 U9171 ( .A1(n9097), .A2(n7426), .B1(n9093), .B2(n7425), .C1(n7424), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  NAND2_X1 U9172 ( .A1(n10052), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7428) );
  OAI21_X1 U9173 ( .B1(n10052), .B2(n7429), .A(n7428), .ZN(P1_U3439) );
  AND2_X1 U9174 ( .A1(n7431), .A2(n7430), .ZN(n7451) );
  OAI21_X1 U9175 ( .B1(n7434), .B2(n7432), .A(n7433), .ZN(n7435) );
  NAND2_X1 U9176 ( .A1(n7435), .A2(n8591), .ZN(n7438) );
  OAI22_X1 U9177 ( .A1(n8583), .A2(n7629), .B1(n6245), .B2(n8597), .ZN(n7436)
         );
  AOI21_X1 U9178 ( .B1(n10118), .B2(n8586), .A(n7436), .ZN(n7437) );
  OAI211_X1 U9179 ( .C1(n7451), .C2(n7631), .A(n7438), .B(n7437), .ZN(P2_U3177) );
  OAI22_X1 U9180 ( .A1(n8602), .A2(n7478), .B1(n8583), .B2(n6245), .ZN(n7439)
         );
  AOI21_X1 U9181 ( .B1(n7524), .B2(n8591), .A(n7439), .ZN(n7440) );
  OAI21_X1 U9182 ( .B1(n7451), .B2(n7461), .A(n7440), .ZN(P2_U3172) );
  AOI21_X1 U9183 ( .B1(n7443), .B2(n7442), .A(n7441), .ZN(n7552) );
  INV_X1 U9184 ( .A(n7552), .ZN(n7446) );
  NAND2_X1 U9185 ( .A1(n7445), .A2(n7444), .ZN(n7553) );
  NOR2_X1 U9186 ( .A1(n10004), .A2(n9390), .ZN(P1_U3085) );
  INV_X1 U9187 ( .A(n7447), .ZN(n7448) );
  AOI21_X1 U9188 ( .B1(n7450), .B2(n7449), .A(n7448), .ZN(n7456) );
  OAI22_X1 U9189 ( .A1(n8583), .A2(n6247), .B1(n7737), .B2(n8597), .ZN(n7453)
         );
  NOR2_X1 U9190 ( .A1(n7451), .A2(n7733), .ZN(n7452) );
  AOI211_X1 U9191 ( .C1(n7454), .C2(n8586), .A(n7453), .B(n7452), .ZN(n7455)
         );
  OAI21_X1 U9192 ( .B1(n8588), .B2(n7456), .A(n7455), .ZN(P2_U3162) );
  INV_X1 U9193 ( .A(n8694), .ZN(n8740) );
  OAI21_X1 U9194 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n7457), .A(n7577), .ZN(n7458) );
  OAI21_X1 U9195 ( .B1(n7459), .B2(n8740), .A(n7458), .ZN(n7460) );
  OAI21_X1 U9196 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n7461), .A(n7460), .ZN(n7462) );
  AOI21_X1 U9197 ( .B1(n8736), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7462), .ZN(
        n7463) );
  OAI21_X1 U9198 ( .B1(n4624), .B2(n8721), .A(n7463), .ZN(P2_U3182) );
  INV_X1 U9199 ( .A(n8626), .ZN(n7464) );
  AOI21_X1 U9200 ( .B1(n7466), .B2(n7465), .A(n7464), .ZN(n7476) );
  XNOR2_X1 U9201 ( .A(n7467), .B(n7644), .ZN(n7472) );
  NOR2_X1 U9202 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5969), .ZN(n7535) );
  XOR2_X1 U9203 ( .A(n7468), .B(P2_REG1_REG_3__SCAN_IN), .Z(n7470) );
  INV_X1 U9204 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n7469) );
  OAI22_X1 U9205 ( .A1(n8748), .A2(n7470), .B1(n7953), .B2(n7469), .ZN(n7471)
         );
  AOI211_X1 U9206 ( .C1(n8701), .C2(n7472), .A(n7535), .B(n7471), .ZN(n7475)
         );
  INV_X1 U9207 ( .A(n8721), .ZN(n8742) );
  NAND2_X1 U9208 ( .A1(n8742), .A2(n7473), .ZN(n7474) );
  OAI211_X1 U9209 ( .C1(n7476), .C2(n8694), .A(n7475), .B(n7474), .ZN(P2_U3185) );
  INV_X1 U9210 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n7480) );
  OAI21_X1 U9211 ( .B1(n10139), .B2(n10096), .A(n7524), .ZN(n7477) );
  OR2_X1 U9212 ( .A1(n6245), .A2(n8896), .ZN(n7527) );
  OAI211_X1 U9213 ( .C1(n10135), .C2(n7478), .A(n7477), .B(n7527), .ZN(n8980)
         );
  NAND2_X1 U9214 ( .A1(n10152), .A2(n8980), .ZN(n7479) );
  OAI21_X1 U9215 ( .B1(n10152), .B2(n7480), .A(n7479), .ZN(P2_U3390) );
  XOR2_X1 U9216 ( .A(n7481), .B(n7482), .Z(n7494) );
  OAI21_X1 U9217 ( .B1(n7485), .B2(n7484), .A(n7483), .ZN(n7486) );
  AOI22_X1 U9218 ( .A1(n8736), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8723), .B2(
        n7486), .ZN(n7491) );
  XNOR2_X1 U9219 ( .A(n7487), .B(n7488), .ZN(n7489) );
  AOI22_X1 U9220 ( .A1(n8701), .A2(n7489), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7490) );
  OAI211_X1 U9221 ( .C1(n7492), .C2(n8721), .A(n7491), .B(n7490), .ZN(n7493)
         );
  AOI21_X1 U9222 ( .B1(n8740), .B2(n7494), .A(n7493), .ZN(n7495) );
  INV_X1 U9223 ( .A(n7495), .ZN(P2_U3184) );
  XNOR2_X1 U9224 ( .A(n7497), .B(n7496), .ZN(n7507) );
  XNOR2_X1 U9225 ( .A(n7498), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7505) );
  XNOR2_X1 U9226 ( .A(n7499), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n7500) );
  NAND2_X1 U9227 ( .A1(n7500), .A2(n8701), .ZN(n7502) );
  AND2_X1 U9228 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7727) );
  AOI21_X1 U9229 ( .B1(n8736), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n7727), .ZN(
        n7501) );
  OAI211_X1 U9230 ( .C1(n8721), .C2(n7503), .A(n7502), .B(n7501), .ZN(n7504)
         );
  AOI21_X1 U9231 ( .B1(n8723), .B2(n7505), .A(n7504), .ZN(n7506) );
  OAI21_X1 U9232 ( .B1(n8694), .B2(n7507), .A(n7506), .ZN(P2_U3187) );
  XNOR2_X1 U9233 ( .A(n7509), .B(n7508), .ZN(n7523) );
  XNOR2_X1 U9234 ( .A(n7511), .B(n7510), .ZN(n7521) );
  INV_X1 U9235 ( .A(n7512), .ZN(n7607) );
  INV_X1 U9236 ( .A(n7513), .ZN(n7515) );
  NOR3_X1 U9237 ( .A1(n7607), .A2(n7515), .A3(n7514), .ZN(n7517) );
  INV_X1 U9238 ( .A(n7677), .ZN(n7516) );
  OAI21_X1 U9239 ( .B1(n7517), .B2(n7516), .A(n8740), .ZN(n7519) );
  AND2_X1 U9240 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7874) );
  AOI21_X1 U9241 ( .B1(n8736), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n7874), .ZN(
        n7518) );
  OAI211_X1 U9242 ( .C1(n8721), .C2(n4742), .A(n7519), .B(n7518), .ZN(n7520)
         );
  AOI21_X1 U9243 ( .B1(n7521), .B2(n8701), .A(n7520), .ZN(n7522) );
  OAI21_X1 U9244 ( .B1(n7523), .B2(n8748), .A(n7522), .ZN(P2_U3189) );
  INV_X1 U9245 ( .A(n7524), .ZN(n7526) );
  NOR3_X1 U9246 ( .A1(n7526), .A2(n7525), .A3(n10151), .ZN(n7529) );
  INV_X1 U9247 ( .A(n7527), .ZN(n7528) );
  OAI21_X1 U9248 ( .B1(n7529), .B2(n7528), .A(n7308), .ZN(n7532) );
  AOI22_X1 U9249 ( .A1(n10101), .A2(n7530), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10102), .ZN(n7531) );
  OAI211_X1 U9250 ( .C1(n5937), .C2(n7308), .A(n7532), .B(n7531), .ZN(P2_U3233) );
  OAI22_X1 U9251 ( .A1(n8602), .A2(n10121), .B1(n8583), .B2(n7533), .ZN(n7534)
         );
  AOI211_X1 U9252 ( .C1(n8580), .C2(n8615), .A(n7535), .B(n7534), .ZN(n7540)
         );
  AOI21_X1 U9253 ( .B1(n7537), .B2(n7536), .A(n8588), .ZN(n7538) );
  NAND2_X1 U9254 ( .A1(n7538), .A2(n7649), .ZN(n7539) );
  OAI211_X1 U9255 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8560), .A(n7540), .B(
        n7539), .ZN(P2_U3158) );
  INV_X1 U9256 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7542) );
  INV_X1 U9257 ( .A(n7541), .ZN(n7544) );
  INV_X1 U9258 ( .A(n9525), .ZN(n9513) );
  OAI222_X1 U9259 ( .A1(n9995), .A2(n7542), .B1(n9994), .B2(n7544), .C1(
        P1_U3086), .C2(n9513), .ZN(P1_U3342) );
  INV_X1 U9260 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7545) );
  OAI222_X1 U9261 ( .A1(n9097), .A2(n7545), .B1(n9093), .B2(n7544), .C1(
        P2_U3151), .C2(n4731), .ZN(P2_U3282) );
  XNOR2_X1 U9262 ( .A(n7556), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n7551) );
  INV_X1 U9263 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8247) );
  INV_X1 U9264 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n8217) );
  INV_X1 U9265 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n8042) );
  INV_X1 U9266 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8171) );
  MUX2_X1 U9267 ( .A(n5016), .B(P1_REG2_REG_1__SCAN_IN), .S(n7557), .Z(n9377)
         );
  AND2_X1 U9268 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9387) );
  NAND2_X1 U9269 ( .A1(n9377), .A2(n9387), .ZN(n9376) );
  NAND2_X1 U9270 ( .A1(n9381), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U9271 ( .A1(n9376), .A2(n7546), .ZN(n9401) );
  NAND2_X1 U9272 ( .A1(n9402), .A2(n9401), .ZN(n9400) );
  NAND2_X1 U9273 ( .A1(n9396), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7547) );
  INV_X1 U9274 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10334) );
  MUX2_X1 U9275 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10334), .S(n9409), .Z(n9415)
         );
  NAND2_X1 U9276 ( .A1(n9409), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7548) );
  XNOR2_X1 U9277 ( .A(n9422), .B(n8042), .ZN(n9425) );
  OAI21_X1 U9278 ( .B1(n7562), .B2(n8042), .A(n9423), .ZN(n9441) );
  XNOR2_X1 U9279 ( .A(n7563), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9442) );
  NAND2_X1 U9280 ( .A1(n9441), .A2(n9442), .ZN(n9440) );
  OAI21_X1 U9281 ( .B1(n7549), .B2(n7563), .A(n9440), .ZN(n9454) );
  XNOR2_X1 U9282 ( .A(n7565), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n9455) );
  NAND2_X1 U9283 ( .A1(n9454), .A2(n9455), .ZN(n9453) );
  OAI21_X1 U9284 ( .B1(n8217), .B2(n7565), .A(n9453), .ZN(n9467) );
  MUX2_X1 U9285 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n8247), .S(n9462), .Z(n9468)
         );
  NAND2_X1 U9286 ( .A1(n9467), .A2(n9468), .ZN(n9466) );
  OAI21_X1 U9287 ( .B1(n7568), .B2(n8247), .A(n9466), .ZN(n9477) );
  XNOR2_X1 U9288 ( .A(n7569), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n9478) );
  NAND2_X1 U9289 ( .A1(n9477), .A2(n9478), .ZN(n9476) );
  OAI21_X1 U9290 ( .B1(n8265), .B2(n7569), .A(n9476), .ZN(n7550) );
  AOI21_X1 U9291 ( .B1(n7551), .B2(n7550), .A(n7588), .ZN(n7576) );
  NAND2_X1 U9292 ( .A1(n7553), .A2(n7552), .ZN(n10006) );
  INV_X1 U9293 ( .A(n9388), .ZN(n7554) );
  AND2_X1 U9294 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9258) );
  NOR2_X1 U9295 ( .A1(n10043), .A2(n7594), .ZN(n7555) );
  AOI211_X1 U9296 ( .C1(n10004), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9258), .B(
        n7555), .ZN(n7575) );
  XNOR2_X1 U9297 ( .A(n7556), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7571) );
  INV_X1 U9298 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n9900) );
  INV_X1 U9299 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7567) );
  INV_X1 U9300 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n7566) );
  INV_X1 U9301 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7564) );
  INV_X1 U9302 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7561) );
  MUX2_X1 U9303 ( .A(n5015), .B(P1_REG1_REG_1__SCAN_IN), .S(n7557), .Z(n9380)
         );
  AND2_X1 U9304 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9379) );
  NAND2_X1 U9305 ( .A1(n9380), .A2(n9379), .ZN(n9378) );
  NAND2_X1 U9306 ( .A1(n9381), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7558) );
  NAND2_X1 U9307 ( .A1(n9378), .A2(n7558), .ZN(n9398) );
  NAND2_X1 U9308 ( .A1(n9399), .A2(n9398), .ZN(n9397) );
  NAND2_X1 U9309 ( .A1(n9396), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7559) );
  NAND2_X1 U9310 ( .A1(n9397), .A2(n7559), .ZN(n9411) );
  MUX2_X1 U9311 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5066), .S(n9409), .Z(n9412)
         );
  NAND2_X1 U9312 ( .A1(n9411), .A2(n9412), .ZN(n9410) );
  NAND2_X1 U9313 ( .A1(n9409), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n7560) );
  NAND2_X1 U9314 ( .A1(n9410), .A2(n7560), .ZN(n9427) );
  XNOR2_X1 U9315 ( .A(n9422), .B(n7561), .ZN(n9428) );
  NAND2_X1 U9316 ( .A1(n9427), .A2(n9428), .ZN(n9426) );
  OAI21_X1 U9317 ( .B1(n7562), .B2(n7561), .A(n9426), .ZN(n9438) );
  XOR2_X1 U9318 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9436), .Z(n9439) );
  XOR2_X1 U9319 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n9449), .Z(n9452) );
  NAND2_X1 U9320 ( .A1(n9451), .A2(n9452), .ZN(n9450) );
  MUX2_X1 U9321 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n7567), .S(n9462), .Z(n9465)
         );
  OAI21_X1 U9322 ( .B1(n7568), .B2(n7567), .A(n9463), .ZN(n9480) );
  XNOR2_X1 U9323 ( .A(n9475), .B(n9900), .ZN(n9481) );
  NAND2_X1 U9324 ( .A1(n9480), .A2(n9481), .ZN(n9479) );
  OAI21_X1 U9325 ( .B1(n9900), .B2(n7569), .A(n9479), .ZN(n7570) );
  NOR2_X1 U9326 ( .A1(n7570), .A2(n7571), .ZN(n7593) );
  AOI21_X1 U9327 ( .B1(n7571), .B2(n7570), .A(n7593), .ZN(n7573) );
  INV_X1 U9328 ( .A(n10002), .ZN(n7572) );
  OR2_X1 U9329 ( .A1(n7573), .A2(n10022), .ZN(n7574) );
  OAI211_X1 U9330 ( .C1(n7576), .C2(n10034), .A(n7575), .B(n7574), .ZN(
        P1_U3252) );
  XOR2_X1 U9331 ( .A(n7578), .B(n7577), .Z(n7585) );
  XOR2_X1 U9332 ( .A(n7579), .B(P2_REG1_REG_1__SCAN_IN), .Z(n7580) );
  INV_X1 U9333 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8114) );
  OAI22_X1 U9334 ( .A1(n8748), .A2(n7580), .B1(n8114), .B2(n7953), .ZN(n7584)
         );
  XNOR2_X1 U9335 ( .A(n7581), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n7582) );
  OAI22_X1 U9336 ( .A1(n8734), .A2(n7582), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7733), .ZN(n7583) );
  AOI211_X1 U9337 ( .C1(n8740), .C2(n7585), .A(n7584), .B(n7583), .ZN(n7586)
         );
  OAI21_X1 U9338 ( .B1(n7587), .B2(n8721), .A(n7586), .ZN(P2_U3183) );
  MUX2_X1 U9339 ( .A(n8294), .B(P1_REG2_REG_12__SCAN_IN), .S(n7592), .Z(n7591)
         );
  INV_X1 U9340 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8067) );
  AOI21_X1 U9341 ( .B1(n8164), .B2(n7594), .A(n7588), .ZN(n9490) );
  XNOR2_X1 U9342 ( .A(n7596), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U9343 ( .A1(n9490), .A2(n9489), .ZN(n9488) );
  OAI21_X1 U9344 ( .B1(n7596), .B2(n7589), .A(n9488), .ZN(n9504) );
  MUX2_X1 U9345 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n8067), .S(n9508), .Z(n9503)
         );
  NAND2_X1 U9346 ( .A1(n9504), .A2(n9503), .ZN(n9502) );
  OAI21_X1 U9347 ( .B1(n8067), .B2(n7597), .A(n9502), .ZN(n7590) );
  AOI21_X1 U9348 ( .B1(n7591), .B2(n7590), .A(n7658), .ZN(n7606) );
  XNOR2_X1 U9349 ( .A(n7592), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7600) );
  INV_X1 U9350 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7595) );
  XOR2_X1 U9351 ( .A(n9494), .B(P1_REG1_REG_10__SCAN_IN), .Z(n9486) );
  NAND2_X1 U9352 ( .A1(n9487), .A2(n9486), .ZN(n9485) );
  OAI21_X1 U9353 ( .B1(n7596), .B2(n7595), .A(n9485), .ZN(n9500) );
  XOR2_X1 U9354 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9508), .Z(n9499) );
  NOR2_X1 U9355 ( .A1(n7599), .A2(n7600), .ZN(n7664) );
  AOI21_X1 U9356 ( .B1(n7600), .B2(n7599), .A(n7664), .ZN(n7601) );
  OR2_X1 U9357 ( .A1(n7601), .A2(n10022), .ZN(n7605) );
  NOR2_X1 U9358 ( .A1(n7602), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9200) );
  NOR2_X1 U9359 ( .A1(n10043), .A2(n7665), .ZN(n7603) );
  AOI211_X1 U9360 ( .C1(n10004), .C2(P1_ADDR_REG_12__SCAN_IN), .A(n9200), .B(
        n7603), .ZN(n7604) );
  OAI211_X1 U9361 ( .C1(n7606), .C2(n10034), .A(n7605), .B(n7604), .ZN(
        P1_U3255) );
  AOI21_X1 U9362 ( .B1(n7609), .B2(n7608), .A(n7607), .ZN(n7623) );
  OAI21_X1 U9363 ( .B1(n7612), .B2(n7611), .A(n4287), .ZN(n7621) );
  NAND2_X1 U9364 ( .A1(n8736), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9365 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7749) );
  OAI211_X1 U9366 ( .C1(n8721), .C2(n7614), .A(n7613), .B(n7749), .ZN(n7620)
         );
  AOI21_X1 U9367 ( .B1(n7617), .B2(n7616), .A(n7615), .ZN(n7618) );
  NOR2_X1 U9368 ( .A1(n7618), .A2(n8734), .ZN(n7619) );
  AOI211_X1 U9369 ( .C1(n8723), .C2(n7621), .A(n7620), .B(n7619), .ZN(n7622)
         );
  OAI21_X1 U9370 ( .B1(n7623), .B2(n8694), .A(n7622), .ZN(P2_U3188) );
  XNOR2_X1 U9371 ( .A(n7625), .B(n7624), .ZN(n10115) );
  XNOR2_X1 U9372 ( .A(n7626), .B(n7627), .ZN(n7628) );
  OAI222_X1 U9373 ( .A1(n8896), .A2(n7629), .B1(n8898), .B2(n6245), .C1(n8894), 
        .C2(n7628), .ZN(n10116) );
  OAI22_X1 U9374 ( .A1(n8874), .A2(n7631), .B1(n7630), .B2(n8778), .ZN(n7632)
         );
  NOR2_X1 U9375 ( .A1(n10116), .A2(n7632), .ZN(n7633) );
  MUX2_X1 U9376 ( .A(n7634), .B(n7633), .S(n7308), .Z(n7635) );
  OAI21_X1 U9377 ( .B1(n8917), .B2(n10115), .A(n7635), .ZN(P2_U3231) );
  INV_X1 U9378 ( .A(n7636), .ZN(n7638) );
  OAI222_X1 U9379 ( .A1(n9097), .A2(n7637), .B1(n9093), .B2(n7638), .C1(
        P2_U3151), .C2(n8663), .ZN(P2_U3281) );
  INV_X1 U9380 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7639) );
  INV_X1 U9381 ( .A(n9527), .ZN(n10015) );
  OAI222_X1 U9382 ( .A1(n9995), .A2(n7639), .B1(n9994), .B2(n7638), .C1(
        P1_U3086), .C2(n10015), .ZN(P1_U3341) );
  XOR2_X1 U9383 ( .A(n7640), .B(n7641), .Z(n10119) );
  XOR2_X1 U9384 ( .A(n7642), .B(n7641), .Z(n7643) );
  AOI222_X1 U9385 ( .A1(n10096), .A2(n7643), .B1(n8613), .B2(n10091), .C1(
        n8615), .C2(n10093), .ZN(n10120) );
  MUX2_X1 U9386 ( .A(n7644), .B(n10120), .S(n7308), .Z(n7647) );
  AOI22_X1 U9387 ( .A1(n10101), .A2(n7645), .B1(n5969), .B2(n10102), .ZN(n7646) );
  OAI211_X1 U9388 ( .C1(n10119), .C2(n8917), .A(n7647), .B(n7646), .ZN(
        P2_U3230) );
  AND2_X1 U9389 ( .A1(n7649), .A2(n7648), .ZN(n7652) );
  OAI21_X1 U9390 ( .B1(n7652), .B2(n7651), .A(n7650), .ZN(n7653) );
  NAND2_X1 U9391 ( .A1(n7653), .A2(n8591), .ZN(n7657) );
  AND2_X1 U9392 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8623) );
  OAI22_X1 U9393 ( .A1(n8602), .A2(n7654), .B1(n8583), .B2(n7751), .ZN(n7655)
         );
  AOI211_X1 U9394 ( .C1(n8580), .C2(n10094), .A(n8623), .B(n7655), .ZN(n7656)
         );
  OAI211_X1 U9395 ( .C1(n10100), .C2(n8560), .A(n7657), .B(n7656), .ZN(
        P2_U3170) );
  INV_X1 U9396 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7659) );
  MUX2_X1 U9397 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n7659), .S(n9525), .Z(n7660)
         );
  OAI21_X1 U9398 ( .B1(n7661), .B2(n7660), .A(n9501), .ZN(n7670) );
  NOR2_X1 U9399 ( .A1(n10313), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9283) );
  INV_X1 U9400 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7662) );
  NOR2_X1 U9401 ( .A1(n10050), .A2(n7662), .ZN(n7663) );
  AOI211_X1 U9402 ( .C1(n10030), .C2(n9525), .A(n9283), .B(n7663), .ZN(n7669)
         );
  XOR2_X1 U9403 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9525), .Z(n7666) );
  NAND2_X1 U9404 ( .A1(n7667), .A2(n7666), .ZN(n9512) );
  OAI211_X1 U9405 ( .C1(n7667), .C2(n7666), .A(n9512), .B(n10037), .ZN(n7668)
         );
  OAI211_X1 U9406 ( .C1(n7670), .C2(n9524), .A(n7669), .B(n7668), .ZN(P1_U3256) );
  OAI21_X1 U9407 ( .B1(n7673), .B2(n7672), .A(n7671), .ZN(n7683) );
  INV_X1 U9408 ( .A(n7674), .ZN(n7675) );
  NAND3_X1 U9409 ( .A1(n7677), .A2(n7676), .A3(n7675), .ZN(n7678) );
  AOI21_X1 U9410 ( .B1(n7696), .B2(n7678), .A(n8694), .ZN(n7682) );
  INV_X1 U9411 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U9412 ( .A1(n8742), .A2(n7679), .ZN(n7680) );
  NAND2_X1 U9413 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n8101) );
  OAI211_X1 U9414 ( .C1(n8127), .C2(n7953), .A(n7680), .B(n8101), .ZN(n7681)
         );
  AOI211_X1 U9415 ( .C1(n7683), .C2(n8701), .A(n7682), .B(n7681), .ZN(n7689)
         );
  OAI21_X1 U9416 ( .B1(n7686), .B2(n7685), .A(n7684), .ZN(n7687) );
  NAND2_X1 U9417 ( .A1(n7687), .A2(n8723), .ZN(n7688) );
  NAND2_X1 U9418 ( .A1(n7689), .A2(n7688), .ZN(P2_U3190) );
  XNOR2_X1 U9419 ( .A(n7691), .B(n7690), .ZN(n7704) );
  XNOR2_X1 U9420 ( .A(n7692), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n7702) );
  INV_X1 U9421 ( .A(n7693), .ZN(n7694) );
  NAND3_X1 U9422 ( .A1(n7696), .A2(n7695), .A3(n7694), .ZN(n7697) );
  AOI21_X1 U9423 ( .B1(n7773), .B2(n7697), .A(n8694), .ZN(n7701) );
  NAND2_X1 U9424 ( .A1(n8736), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7698) );
  NAND2_X1 U9425 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8032) );
  OAI211_X1 U9426 ( .C1(n8721), .C2(n7699), .A(n7698), .B(n8032), .ZN(n7700)
         );
  AOI211_X1 U9427 ( .C1(n7702), .C2(n8701), .A(n7701), .B(n7700), .ZN(n7703)
         );
  OAI21_X1 U9428 ( .B1(n7704), .B2(n8748), .A(n7703), .ZN(P2_U3191) );
  INV_X1 U9429 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7706) );
  INV_X1 U9430 ( .A(n7705), .ZN(n7707) );
  INV_X1 U9431 ( .A(n10029), .ZN(n9528) );
  OAI222_X1 U9432 ( .A1(n9995), .A2(n7706), .B1(n9994), .B2(n7707), .C1(
        P1_U3086), .C2(n9528), .ZN(P1_U3340) );
  OAI222_X1 U9433 ( .A1(n9097), .A2(n7708), .B1(n9093), .B2(n7707), .C1(
        P2_U3151), .C2(n8678), .ZN(P2_U3280) );
  INV_X1 U9434 ( .A(n7709), .ZN(n7711) );
  NOR3_X1 U9435 ( .A1(n7712), .A2(n7711), .A3(n7710), .ZN(n7816) );
  XOR2_X1 U9436 ( .A(n7714), .B(n7713), .Z(n9392) );
  NAND2_X1 U9437 ( .A1(n9375), .A2(n9324), .ZN(n9794) );
  OAI22_X1 U9438 ( .A1(n9331), .A2(n7715), .B1(n9326), .B2(n9794), .ZN(n7716)
         );
  AOI21_X1 U9439 ( .B1(n9392), .B2(n9302), .A(n7716), .ZN(n7717) );
  OAI21_X1 U9440 ( .B1(n7816), .B2(n7718), .A(n7717), .ZN(P1_U3232) );
  INV_X1 U9441 ( .A(n7650), .ZN(n7722) );
  INV_X1 U9442 ( .A(n7719), .ZN(n7721) );
  NOR3_X1 U9443 ( .A1(n7722), .A2(n7721), .A3(n7720), .ZN(n7723) );
  OAI21_X1 U9444 ( .B1(n7723), .B2(n4378), .A(n8591), .ZN(n7729) );
  OAI22_X1 U9445 ( .A1(n8602), .A2(n7725), .B1(n8583), .B2(n7724), .ZN(n7726)
         );
  AOI211_X1 U9446 ( .C1(n8580), .C2(n8613), .A(n7727), .B(n7726), .ZN(n7728)
         );
  OAI211_X1 U9447 ( .C1(n7801), .C2(n8560), .A(n7729), .B(n7728), .ZN(P2_U3167) );
  NAND2_X1 U9448 ( .A1(n6244), .A2(n7730), .ZN(n7731) );
  NAND2_X1 U9449 ( .A1(n7732), .A2(n7731), .ZN(n10112) );
  OAI22_X1 U9450 ( .A1(n8901), .A2(n10109), .B1(n7733), .B2(n8874), .ZN(n7739)
         );
  XNOR2_X1 U9451 ( .A(n7735), .B(n7734), .ZN(n7736) );
  OAI222_X1 U9452 ( .A1(n8896), .A2(n6247), .B1(n8898), .B2(n7737), .C1(n8894), 
        .C2(n7736), .ZN(n10110) );
  MUX2_X1 U9453 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n10110), .S(n7308), .Z(n7738)
         );
  AOI211_X1 U9454 ( .C1(n10104), .C2(n10112), .A(n7739), .B(n7738), .ZN(n7740)
         );
  INV_X1 U9455 ( .A(n7740), .ZN(P2_U3232) );
  INV_X1 U9456 ( .A(n7741), .ZN(n7744) );
  INV_X1 U9457 ( .A(n9540), .ZN(n9523) );
  OAI222_X1 U9458 ( .A1(n9994), .A2(n7744), .B1(n9523), .B2(P1_U3086), .C1(
        n7742), .C2(n9995), .ZN(P1_U3339) );
  OAI222_X1 U9459 ( .A1(n9097), .A2(n7745), .B1(P2_U3151), .B2(n4631), .C1(
        n7744), .C2(n9093), .ZN(P2_U3279) );
  OAI211_X1 U9460 ( .C1(n7748), .C2(n7747), .A(n7746), .B(n8591), .ZN(n7754)
         );
  NAND2_X1 U9461 ( .A1(n8595), .A2(n8612), .ZN(n7750) );
  OAI211_X1 U9462 ( .C1(n8597), .C2(n7751), .A(n7750), .B(n7749), .ZN(n7752)
         );
  AOI21_X1 U9463 ( .B1(n7790), .B2(n8586), .A(n7752), .ZN(n7753) );
  OAI211_X1 U9464 ( .C1(n7788), .C2(n8560), .A(n7754), .B(n7753), .ZN(P2_U3179) );
  INV_X1 U9465 ( .A(n9798), .ZN(n9803) );
  OAI21_X1 U9466 ( .B1(n10061), .B2(n9778), .A(n9803), .ZN(n7756) );
  NAND2_X1 U9467 ( .A1(n9797), .A2(n7836), .ZN(n9795) );
  AND2_X1 U9468 ( .A1(n9794), .A2(n9795), .ZN(n7755) );
  AND2_X1 U9469 ( .A1(n7756), .A2(n7755), .ZN(n10054) );
  NAND2_X1 U9470 ( .A1(n7060), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7757) );
  OAI21_X1 U9471 ( .B1(n7060), .B2(n10054), .A(n7757), .ZN(P1_U3522) );
  AOI21_X1 U9472 ( .B1(n7758), .B2(n7759), .A(n7809), .ZN(n7764) );
  AOI22_X1 U9473 ( .A1(n9343), .A2(n4293), .B1(n9339), .B2(n7760), .ZN(n7763)
         );
  INV_X1 U9474 ( .A(n7816), .ZN(n7761) );
  NAND2_X1 U9475 ( .A1(n7761), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7762) );
  OAI211_X1 U9476 ( .C1(n7764), .C2(n9345), .A(n7763), .B(n7762), .ZN(P1_U3222) );
  INV_X1 U9477 ( .A(n7765), .ZN(n7766) );
  AOI21_X1 U9478 ( .B1(n7768), .B2(n7767), .A(n7766), .ZN(n7783) );
  INV_X1 U9479 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U9480 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8454) );
  OAI21_X1 U9481 ( .B1(n7953), .B2(n7769), .A(n8454), .ZN(n7776) );
  INV_X1 U9482 ( .A(n7770), .ZN(n7771) );
  NAND3_X1 U9483 ( .A1(n7773), .A2(n7772), .A3(n7771), .ZN(n7774) );
  AOI21_X1 U9484 ( .B1(n7907), .B2(n7774), .A(n8694), .ZN(n7775) );
  AOI211_X1 U9485 ( .C1(n8742), .C2(n7777), .A(n7776), .B(n7775), .ZN(n7782)
         );
  XNOR2_X1 U9486 ( .A(n7779), .B(n7778), .ZN(n7780) );
  NAND2_X1 U9487 ( .A1(n7780), .A2(n8723), .ZN(n7781) );
  OAI211_X1 U9488 ( .C1(n7783), .C2(n8734), .A(n7782), .B(n7781), .ZN(P2_U3192) );
  XOR2_X1 U9489 ( .A(n7786), .B(n7784), .Z(n10133) );
  XOR2_X1 U9490 ( .A(n7785), .B(n7786), .Z(n7787) );
  AOI222_X1 U9491 ( .A1(n10096), .A2(n7787), .B1(n8612), .B2(n10091), .C1(
        n10092), .C2(n10093), .ZN(n10134) );
  MUX2_X1 U9492 ( .A(n10286), .B(n10134), .S(n7308), .Z(n7792) );
  INV_X1 U9493 ( .A(n7788), .ZN(n7789) );
  AOI22_X1 U9494 ( .A1(n10101), .A2(n7790), .B1(n10102), .B2(n7789), .ZN(n7791) );
  OAI211_X1 U9495 ( .C1(n10133), .C2(n8917), .A(n7792), .B(n7791), .ZN(
        P2_U3227) );
  XOR2_X1 U9496 ( .A(n7796), .B(n7793), .Z(n10130) );
  INV_X1 U9497 ( .A(n10130), .ZN(n7805) );
  OR2_X1 U9498 ( .A1(n10107), .A2(n7794), .ZN(n10086) );
  INV_X1 U9499 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7800) );
  INV_X1 U9500 ( .A(n8059), .ZN(n10113) );
  XNOR2_X1 U9501 ( .A(n7795), .B(n7796), .ZN(n7798) );
  AOI22_X1 U9502 ( .A1(n8613), .A2(n10093), .B1(n10091), .B2(n10079), .ZN(
        n7797) );
  OAI21_X1 U9503 ( .B1(n7798), .B2(n8894), .A(n7797), .ZN(n7799) );
  AOI21_X1 U9504 ( .B1(n10130), .B2(n10113), .A(n7799), .ZN(n10132) );
  MUX2_X1 U9505 ( .A(n7800), .B(n10132), .S(n7308), .Z(n7804) );
  INV_X1 U9506 ( .A(n7801), .ZN(n7802) );
  AOI22_X1 U9507 ( .A1(n10101), .A2(n10129), .B1(n10102), .B2(n7802), .ZN(
        n7803) );
  OAI211_X1 U9508 ( .C1(n7805), .C2(n10086), .A(n7804), .B(n7803), .ZN(
        P2_U3228) );
  INV_X1 U9509 ( .A(n7806), .ZN(n7811) );
  NOR3_X1 U9510 ( .A1(n7809), .A2(n7808), .A3(n7807), .ZN(n7810) );
  OAI21_X1 U9511 ( .B1(n7811), .B2(n7810), .A(n9302), .ZN(n7815) );
  OAI22_X1 U9512 ( .A1(n7812), .A2(n9336), .B1(n9337), .B2(n7073), .ZN(n7834)
         );
  AOI22_X1 U9513 ( .A1(n9343), .A2(n7813), .B1(n9339), .B2(n7834), .ZN(n7814)
         );
  OAI211_X1 U9514 ( .C1(n7816), .C2(n9393), .A(n7815), .B(n7814), .ZN(P1_U3237) );
  NAND3_X1 U9515 ( .A1(n7818), .A2(n7817), .A3(n7825), .ZN(n7819) );
  AND2_X1 U9516 ( .A1(n7820), .A2(n7819), .ZN(n7821) );
  AOI22_X1 U9517 ( .A1(n9324), .A2(n9372), .B1(n9322), .B2(n5084), .ZN(n7920)
         );
  OAI21_X1 U9518 ( .B1(n7821), .B2(n9757), .A(n7920), .ZN(n8040) );
  NAND2_X1 U9519 ( .A1(n7846), .A2(n8044), .ZN(n7822) );
  NAND2_X1 U9520 ( .A1(n7822), .A2(n9764), .ZN(n7823) );
  NOR2_X1 U9521 ( .A1(n7939), .A2(n7823), .ZN(n8045) );
  NOR2_X1 U9522 ( .A1(n8040), .A2(n8045), .ZN(n7857) );
  AND2_X1 U9523 ( .A1(n7825), .A2(n7824), .ZN(n7932) );
  NOR2_X1 U9524 ( .A1(n7824), .A2(n7825), .ZN(n7826) );
  OR2_X1 U9525 ( .A1(n7932), .A2(n7826), .ZN(n8046) );
  OAI22_X1 U9526 ( .A1(n9902), .A2(n7854), .B1(n10073), .B2(n7561), .ZN(n7827)
         );
  AOI21_X1 U9527 ( .B1(n9858), .B2(n8046), .A(n7827), .ZN(n7828) );
  OAI21_X1 U9528 ( .B1(n7857), .B2(n7060), .A(n7828), .ZN(P1_U3526) );
  INV_X1 U9529 ( .A(n10061), .ZN(n9889) );
  NAND2_X1 U9530 ( .A1(n7073), .A2(n7334), .ZN(n7829) );
  NAND2_X1 U9531 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  XNOR2_X1 U9532 ( .A(n7831), .B(n7832), .ZN(n8179) );
  XNOR2_X1 U9533 ( .A(n7833), .B(n7832), .ZN(n7835) );
  AOI21_X1 U9534 ( .B1(n7835), .B2(n9778), .A(n7834), .ZN(n8175) );
  NOR2_X1 U9535 ( .A1(n4293), .A2(n7836), .ZN(n7837) );
  OAI211_X1 U9536 ( .C1(n8172), .C2(n7837), .A(n9764), .B(n7845), .ZN(n8170)
         );
  OAI211_X1 U9537 ( .C1(n9889), .C2(n8179), .A(n8175), .B(n8170), .ZN(n7860)
         );
  OAI22_X1 U9538 ( .A1(n9902), .A2(n8172), .B1(n10073), .B2(n5021), .ZN(n7838)
         );
  AOI21_X1 U9539 ( .B1(n10073), .B2(n7860), .A(n7838), .ZN(n7839) );
  INV_X1 U9540 ( .A(n7839), .ZN(P1_U3524) );
  XNOR2_X1 U9541 ( .A(n7840), .B(n7849), .ZN(n7844) );
  NAND2_X1 U9542 ( .A1(n9322), .A2(n9374), .ZN(n7842) );
  NAND2_X1 U9543 ( .A1(n9324), .A2(n9373), .ZN(n7841) );
  NAND2_X1 U9544 ( .A1(n7842), .A2(n7841), .ZN(n9140) );
  INV_X1 U9545 ( .A(n9140), .ZN(n7843) );
  OAI21_X1 U9546 ( .B1(n7844), .B2(n9757), .A(n7843), .ZN(n10343) );
  OAI211_X1 U9547 ( .C1(n5683), .C2(n7862), .A(n9764), .B(n7846), .ZN(n10340)
         );
  INV_X1 U9548 ( .A(n10340), .ZN(n7847) );
  NOR2_X1 U9549 ( .A1(n10343), .A2(n7847), .ZN(n7865) );
  OR2_X1 U9550 ( .A1(n7850), .A2(n7849), .ZN(n7851) );
  NAND2_X1 U9551 ( .A1(n7848), .A2(n7851), .ZN(n10332) );
  OAI22_X1 U9552 ( .A1(n9902), .A2(n7862), .B1(n10073), .B2(n5066), .ZN(n7852)
         );
  AOI21_X1 U9553 ( .B1(n9858), .B2(n10332), .A(n7852), .ZN(n7853) );
  OAI21_X1 U9554 ( .B1(n7865), .B2(n7060), .A(n7853), .ZN(P1_U3525) );
  OAI22_X1 U9555 ( .A1(n9978), .A2(n7854), .B1(n10070), .B2(n5086), .ZN(n7855)
         );
  AOI21_X1 U9556 ( .B1(n9952), .B2(n8046), .A(n7855), .ZN(n7856) );
  OAI21_X1 U9557 ( .B1(n7857), .B2(n6383), .A(n7856), .ZN(P1_U3465) );
  INV_X1 U9558 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7858) );
  OAI22_X1 U9559 ( .A1(n9978), .A2(n8172), .B1(n10070), .B2(n7858), .ZN(n7859)
         );
  AOI21_X1 U9560 ( .B1(n10070), .B2(n7860), .A(n7859), .ZN(n7861) );
  INV_X1 U9561 ( .A(n7861), .ZN(P1_U3459) );
  OAI22_X1 U9562 ( .A1(n9978), .A2(n7862), .B1(n10070), .B2(n5064), .ZN(n7863)
         );
  AOI21_X1 U9563 ( .B1(n9952), .B2(n10332), .A(n7863), .ZN(n7864) );
  OAI21_X1 U9564 ( .B1(n7865), .B2(n6383), .A(n7864), .ZN(P1_U3462) );
  INV_X1 U9565 ( .A(n7866), .ZN(n7867) );
  OAI222_X1 U9566 ( .A1(n9097), .A2(n10253), .B1(n9093), .B2(n7867), .C1(
        P2_U3151), .C2(n8720), .ZN(P2_U3278) );
  INV_X1 U9567 ( .A(n9553), .ZN(n9549) );
  OAI222_X1 U9568 ( .A1(n9995), .A2(n7868), .B1(n9994), .B2(n7867), .C1(
        P1_U3086), .C2(n9549), .ZN(P1_U3338) );
  INV_X1 U9569 ( .A(n7869), .ZN(n7870) );
  AOI21_X1 U9570 ( .B1(n7872), .B2(n7871), .A(n7870), .ZN(n7879) );
  INV_X1 U9571 ( .A(n7873), .ZN(n10088) );
  NAND2_X1 U9572 ( .A1(n8599), .A2(n10088), .ZN(n7876) );
  AOI21_X1 U9573 ( .B1(n8580), .B2(n10079), .A(n7874), .ZN(n7875) );
  OAI211_X1 U9574 ( .C1(n8033), .C2(n8583), .A(n7876), .B(n7875), .ZN(n7877)
         );
  AOI21_X1 U9575 ( .B1(n10140), .B2(n8586), .A(n7877), .ZN(n7878) );
  OAI21_X1 U9576 ( .B1(n7879), .B2(n8588), .A(n7878), .ZN(P2_U3153) );
  INV_X1 U9577 ( .A(n10067), .ZN(n9899) );
  AOI211_X1 U9578 ( .C1(n9899), .C2(n7882), .A(n7881), .B(n7880), .ZN(n7885)
         );
  AOI22_X1 U9579 ( .A1(n6366), .A2(n4293), .B1(n7060), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n7883) );
  OAI21_X1 U9580 ( .B1(n7885), .B2(n7060), .A(n7883), .ZN(P1_U3523) );
  AOI22_X1 U9581 ( .A1(n5687), .A2(n4293), .B1(n6383), .B2(
        P1_REG0_REG_1__SCAN_IN), .ZN(n7884) );
  OAI21_X1 U9582 ( .B1(n7885), .B2(n6383), .A(n7884), .ZN(P1_U3456) );
  INV_X1 U9583 ( .A(n7896), .ZN(n7887) );
  XNOR2_X1 U9584 ( .A(n8157), .B(n7887), .ZN(n7890) );
  NAND2_X1 U9585 ( .A1(n9324), .A2(n9370), .ZN(n7889) );
  NAND2_X1 U9586 ( .A1(n9322), .A2(n9372), .ZN(n7888) );
  NAND2_X1 U9587 ( .A1(n7889), .A2(n7888), .ZN(n8232) );
  AOI21_X1 U9588 ( .B1(n7890), .B2(n9778), .A(n8232), .ZN(n8226) );
  AOI21_X1 U9589 ( .B1(n7938), .B2(n8219), .A(n9784), .ZN(n7891) );
  NAND2_X1 U9590 ( .A1(n7891), .A2(n8248), .ZN(n8223) );
  AND2_X1 U9591 ( .A1(n8226), .A2(n8223), .ZN(n7901) );
  INV_X1 U9592 ( .A(n7892), .ZN(n7893) );
  NAND2_X1 U9593 ( .A1(n7894), .A2(n7893), .ZN(n7895) );
  XNOR2_X1 U9594 ( .A(n7896), .B(n7895), .ZN(n8220) );
  OAI22_X1 U9595 ( .A1(n9902), .A2(n8235), .B1(n10073), .B2(n7566), .ZN(n7897)
         );
  AOI21_X1 U9596 ( .B1(n9858), .B2(n8220), .A(n7897), .ZN(n7898) );
  OAI21_X1 U9597 ( .B1(n7901), .B2(n7060), .A(n7898), .ZN(P1_U3528) );
  OAI22_X1 U9598 ( .A1(n9978), .A2(n8235), .B1(n10070), .B2(n5132), .ZN(n7899)
         );
  AOI21_X1 U9599 ( .B1(n9952), .B2(n8220), .A(n7899), .ZN(n7900) );
  OAI21_X1 U9600 ( .B1(n7901), .B2(n6383), .A(n7900), .ZN(P1_U3471) );
  XNOR2_X1 U9601 ( .A(n7902), .B(n8083), .ZN(n7915) );
  XNOR2_X1 U9602 ( .A(n7903), .B(n8088), .ZN(n7913) );
  INV_X1 U9603 ( .A(n7904), .ZN(n7905) );
  NAND3_X1 U9604 ( .A1(n7907), .A2(n7906), .A3(n7905), .ZN(n7908) );
  AOI21_X1 U9605 ( .B1(n7957), .B2(n7908), .A(n8694), .ZN(n7912) );
  NAND2_X1 U9606 ( .A1(n8736), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n7909) );
  NAND2_X1 U9607 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8556) );
  OAI211_X1 U9608 ( .C1(n8721), .C2(n7910), .A(n7909), .B(n8556), .ZN(n7911)
         );
  AOI211_X1 U9609 ( .C1(n7913), .C2(n8723), .A(n7912), .B(n7911), .ZN(n7914)
         );
  OAI21_X1 U9610 ( .B1(n7915), .B2(n8734), .A(n7914), .ZN(P2_U3193) );
  AND2_X1 U9611 ( .A1(n9136), .A2(n7916), .ZN(n7919) );
  OAI211_X1 U9612 ( .C1(n7919), .C2(n7918), .A(n9302), .B(n7917), .ZN(n7923)
         );
  NAND2_X1 U9613 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9419) );
  OAI21_X1 U9614 ( .B1(n9326), .B2(n7920), .A(n9419), .ZN(n7921) );
  AOI21_X1 U9615 ( .B1(n9343), .B2(n8044), .A(n7921), .ZN(n7922) );
  OAI211_X1 U9616 ( .C1(n9341), .C2(n8041), .A(n7923), .B(n7922), .ZN(P1_U3230) );
  INV_X1 U9617 ( .A(n7924), .ZN(n7947) );
  INV_X1 U9618 ( .A(n9557), .ZN(n10042) );
  OAI222_X1 U9619 ( .A1(n9994), .A2(n7947), .B1(n10042), .B2(P1_U3086), .C1(
        n10314), .C2(n9995), .ZN(P1_U3337) );
  OAI21_X1 U9620 ( .B1(n7933), .B2(n7926), .A(n7925), .ZN(n7927) );
  NAND2_X1 U9621 ( .A1(n7927), .A2(n9778), .ZN(n7930) );
  NAND2_X1 U9622 ( .A1(n9322), .A2(n9373), .ZN(n7929) );
  NAND2_X1 U9623 ( .A1(n9324), .A2(n9371), .ZN(n7928) );
  AND2_X1 U9624 ( .A1(n7929), .A2(n7928), .ZN(n8204) );
  NAND2_X1 U9625 ( .A1(n7930), .A2(n8204), .ZN(n10058) );
  INV_X1 U9626 ( .A(n10058), .ZN(n7945) );
  NOR2_X1 U9627 ( .A1(n7932), .A2(n7931), .ZN(n7934) );
  XNOR2_X1 U9628 ( .A(n7934), .B(n7933), .ZN(n10060) );
  NAND2_X1 U9629 ( .A1(n8264), .A2(n7935), .ZN(n7936) );
  OAI211_X1 U9630 ( .C1(n7939), .C2(n10057), .A(n7938), .B(n9764), .ZN(n10055)
         );
  INV_X1 U9631 ( .A(n8209), .ZN(n7940) );
  INV_X1 U9632 ( .A(n9780), .ZN(n10336) );
  AOI22_X1 U9633 ( .A1(n10337), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7940), .B2(
        n10336), .ZN(n7942) );
  NAND2_X1 U9634 ( .A1(n10331), .A2(n8206), .ZN(n7941) );
  OAI211_X1 U9635 ( .C1(n10341), .C2(n10055), .A(n7942), .B(n7941), .ZN(n7943)
         );
  AOI21_X1 U9636 ( .B1(n10060), .B2(n10333), .A(n7943), .ZN(n7944) );
  OAI21_X1 U9637 ( .B1(n7945), .B2(n9712), .A(n7944), .ZN(P1_U3288) );
  OAI222_X1 U9638 ( .A1(P2_U3151), .A2(n7948), .B1(n9093), .B2(n7947), .C1(
        n7946), .C2(n9097), .ZN(P2_U3277) );
  AOI21_X1 U9639 ( .B1(n7951), .B2(n7950), .A(n7949), .ZN(n7967) );
  INV_X1 U9640 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U9641 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8095) );
  OAI21_X1 U9642 ( .B1(n7953), .B2(n7952), .A(n8095), .ZN(n7960) );
  INV_X1 U9643 ( .A(n7954), .ZN(n7955) );
  NAND3_X1 U9644 ( .A1(n7957), .A2(n7956), .A3(n7955), .ZN(n7958) );
  AOI21_X1 U9645 ( .B1(n8640), .B2(n7958), .A(n8694), .ZN(n7959) );
  AOI211_X1 U9646 ( .C1(n8742), .C2(n7961), .A(n7960), .B(n7959), .ZN(n7966)
         );
  XNOR2_X1 U9647 ( .A(n7963), .B(n7962), .ZN(n7964) );
  NAND2_X1 U9648 ( .A1(n7964), .A2(n8723), .ZN(n7965) );
  OAI211_X1 U9649 ( .C1(n7967), .C2(n8734), .A(n7966), .B(n7965), .ZN(P2_U3194) );
  NAND2_X1 U9650 ( .A1(n7969), .A2(n7968), .ZN(n7972) );
  INV_X1 U9651 ( .A(n7972), .ZN(n7970) );
  NAND2_X1 U9652 ( .A1(n7970), .A2(n7971), .ZN(n7973) );
  INV_X1 U9653 ( .A(n7971), .ZN(n7978) );
  NAND2_X1 U9654 ( .A1(n7972), .A2(n7978), .ZN(n8051) );
  NAND2_X1 U9655 ( .A1(n7975), .A2(n8033), .ZN(n7976) );
  NAND2_X1 U9656 ( .A1(n7976), .A2(n10150), .ZN(n7977) );
  OAI21_X1 U9657 ( .B1(n8033), .B2(n7975), .A(n7977), .ZN(n7979) );
  XNOR2_X1 U9658 ( .A(n7979), .B(n7978), .ZN(n7980) );
  NAND2_X1 U9659 ( .A1(n7980), .A2(n10096), .ZN(n7984) );
  OAI22_X1 U9660 ( .A1(n8033), .A2(n8898), .B1(n8551), .B2(n8896), .ZN(n7981)
         );
  AOI21_X1 U9661 ( .B1(n7982), .B2(n10113), .A(n7981), .ZN(n7983) );
  AND2_X1 U9662 ( .A1(n7984), .A2(n7983), .ZN(n8978) );
  MUX2_X1 U9663 ( .A(n7985), .B(n8978), .S(n7308), .Z(n7988) );
  INV_X1 U9664 ( .A(n8034), .ZN(n7986) );
  AOI22_X1 U9665 ( .A1(n10101), .A2(n8976), .B1(n7986), .B2(n10102), .ZN(n7987) );
  OAI211_X1 U9666 ( .C1(n8979), .C2(n10086), .A(n7988), .B(n7987), .ZN(
        P2_U3224) );
  NAND2_X1 U9667 ( .A1(n10074), .A2(n4401), .ZN(n10078) );
  NAND2_X1 U9668 ( .A1(n10078), .A2(n7991), .ZN(n7992) );
  XOR2_X1 U9669 ( .A(n7993), .B(n7992), .Z(n10147) );
  XOR2_X1 U9670 ( .A(n7975), .B(n7993), .Z(n7994) );
  OAI222_X1 U9671 ( .A1(n8896), .A2(n8055), .B1(n8898), .B2(n8102), .C1(n8894), 
        .C2(n7994), .ZN(n10148) );
  INV_X1 U9672 ( .A(n10148), .ZN(n7995) );
  MUX2_X1 U9673 ( .A(n7996), .B(n7995), .S(n7308), .Z(n7999) );
  INV_X1 U9674 ( .A(n8105), .ZN(n7997) );
  AOI22_X1 U9675 ( .A1(n10101), .A2(n10150), .B1(n10102), .B2(n7997), .ZN(
        n7998) );
  OAI211_X1 U9676 ( .C1(n10147), .C2(n8917), .A(n7999), .B(n7998), .ZN(
        P2_U3225) );
  OR2_X1 U9677 ( .A1(n8001), .A2(n8000), .ZN(n8002) );
  NAND2_X1 U9678 ( .A1(n8003), .A2(n8002), .ZN(n8024) );
  INV_X1 U9679 ( .A(n8024), .ZN(n8017) );
  OAI21_X1 U9680 ( .B1(n8006), .B2(n8005), .A(n8004), .ZN(n8007) );
  NAND2_X1 U9681 ( .A1(n8007), .A2(n9778), .ZN(n8008) );
  AOI22_X1 U9682 ( .A1(n9322), .A2(n9368), .B1(n9366), .B2(n9324), .ZN(n9129)
         );
  NAND2_X1 U9683 ( .A1(n8008), .A2(n9129), .ZN(n8021) );
  NAND2_X1 U9684 ( .A1(n8021), .A2(n7937), .ZN(n8016) );
  INV_X1 U9685 ( .A(n8066), .ZN(n8010) );
  AOI211_X1 U9686 ( .C1(n9133), .C2(n8009), .A(n9784), .B(n8010), .ZN(n8020)
         );
  INV_X1 U9687 ( .A(n9133), .ZN(n8013) );
  INV_X1 U9688 ( .A(n9130), .ZN(n8011) );
  AOI22_X1 U9689 ( .A1(n10337), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n8011), .B2(
        n10336), .ZN(n8012) );
  OAI21_X1 U9690 ( .B1(n8013), .B2(n9715), .A(n8012), .ZN(n8014) );
  AOI21_X1 U9691 ( .B1(n8020), .B2(n9788), .A(n8014), .ZN(n8015) );
  OAI211_X1 U9692 ( .C1(n8017), .C2(n9793), .A(n8016), .B(n8015), .ZN(P1_U3283) );
  INV_X1 U9693 ( .A(n8018), .ZN(n8388) );
  OAI222_X1 U9694 ( .A1(n9097), .A2(n10259), .B1(n9093), .B2(n8388), .C1(
        P2_U3151), .C2(n8019), .ZN(P2_U3276) );
  NOR2_X1 U9695 ( .A1(n8021), .A2(n8020), .ZN(n8027) );
  AOI22_X1 U9696 ( .A1(n6366), .A2(n9133), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n7060), .ZN(n8023) );
  NAND2_X1 U9697 ( .A1(n8024), .A2(n9858), .ZN(n8022) );
  OAI211_X1 U9698 ( .C1(n8027), .C2(n7060), .A(n8023), .B(n8022), .ZN(P1_U3532) );
  AOI22_X1 U9699 ( .A1(n5687), .A2(n9133), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n6383), .ZN(n8026) );
  NAND2_X1 U9700 ( .A1(n8024), .A2(n9952), .ZN(n8025) );
  OAI211_X1 U9701 ( .C1(n8027), .C2(n6383), .A(n8026), .B(n8025), .ZN(P1_U3483) );
  NAND2_X1 U9702 ( .A1(n8028), .A2(n8109), .ZN(n8031) );
  XNOR2_X1 U9703 ( .A(n8029), .B(n8055), .ZN(n8030) );
  NAND2_X1 U9704 ( .A1(n8031), .A2(n8030), .ZN(n8453) );
  OAI211_X1 U9705 ( .C1(n8031), .C2(n8030), .A(n8453), .B(n8591), .ZN(n8038)
         );
  OAI21_X1 U9706 ( .B1(n8597), .B2(n8033), .A(n8032), .ZN(n8036) );
  NOR2_X1 U9707 ( .A1(n8560), .A2(n8034), .ZN(n8035) );
  AOI211_X1 U9708 ( .C1(n8595), .C2(n8609), .A(n8036), .B(n8035), .ZN(n8037)
         );
  OAI211_X1 U9709 ( .C1(n8039), .C2(n8602), .A(n8038), .B(n8037), .ZN(P2_U3171) );
  INV_X1 U9710 ( .A(n8040), .ZN(n8049) );
  OAI22_X1 U9711 ( .A1(n10344), .A2(n8042), .B1(n8041), .B2(n9780), .ZN(n8043)
         );
  AOI21_X1 U9712 ( .B1(n10331), .B2(n8044), .A(n8043), .ZN(n8048) );
  AOI22_X1 U9713 ( .A1(n10333), .A2(n8046), .B1(n9788), .B2(n8045), .ZN(n8047)
         );
  OAI211_X1 U9714 ( .C1(n8049), .C2(n10337), .A(n8048), .B(n8047), .ZN(
        P1_U3289) );
  NAND2_X1 U9715 ( .A1(n8051), .A2(n8050), .ZN(n8052) );
  XOR2_X1 U9716 ( .A(n8054), .B(n8052), .Z(n8185) );
  INV_X1 U9717 ( .A(n8185), .ZN(n8060) );
  XNOR2_X1 U9718 ( .A(n8053), .B(n8054), .ZN(n8057) );
  OAI22_X1 U9719 ( .A1(n8055), .A2(n8898), .B1(n8455), .B2(n8896), .ZN(n8056)
         );
  AOI21_X1 U9720 ( .B1(n8057), .B2(n10096), .A(n8056), .ZN(n8058) );
  OAI21_X1 U9721 ( .B1(n8185), .B2(n8059), .A(n8058), .ZN(n8180) );
  AOI21_X1 U9722 ( .B1(n10141), .B2(n8060), .A(n8180), .ZN(n8213) );
  AOI22_X1 U9723 ( .A1(n9066), .A2(n8460), .B1(n10154), .B2(
        P2_REG0_REG_10__SCAN_IN), .ZN(n8061) );
  OAI21_X1 U9724 ( .B1(n8213), .B2(n10154), .A(n8061), .ZN(P2_U3420) );
  OAI21_X1 U9725 ( .B1(n8071), .B2(n8062), .A(n8284), .ZN(n8065) );
  NAND2_X1 U9726 ( .A1(n9367), .A2(n9322), .ZN(n8064) );
  NAND2_X1 U9727 ( .A1(n9365), .A2(n9324), .ZN(n8063) );
  NAND2_X1 U9728 ( .A1(n8064), .A2(n8063), .ZN(n9307) );
  AOI21_X1 U9729 ( .B1(n8065), .B2(n9778), .A(n9307), .ZN(n9887) );
  AOI211_X1 U9730 ( .C1(n9885), .C2(n8066), .A(n9784), .B(n8291), .ZN(n9884)
         );
  NOR2_X1 U9731 ( .A1(n9715), .A2(n4771), .ZN(n8069) );
  OAI22_X1 U9732 ( .A1(n10344), .A2(n8067), .B1(n9305), .B2(n9780), .ZN(n8068)
         );
  AOI211_X1 U9733 ( .C1(n9884), .C2(n9788), .A(n8069), .B(n8068), .ZN(n8074)
         );
  XNOR2_X1 U9734 ( .A(n8070), .B(n8071), .ZN(n9888) );
  INV_X1 U9735 ( .A(n9888), .ZN(n8072) );
  NAND2_X1 U9736 ( .A1(n8072), .A2(n10333), .ZN(n8073) );
  OAI211_X1 U9737 ( .C1(n9887), .C2(n10337), .A(n8074), .B(n8073), .ZN(
        P1_U3282) );
  XNOR2_X1 U9738 ( .A(n8076), .B(n8075), .ZN(n8091) );
  XNOR2_X1 U9739 ( .A(n8077), .B(n8078), .ZN(n8079) );
  AOI222_X1 U9740 ( .A1(n10096), .A2(n8079), .B1(n8607), .B2(n10091), .C1(
        n8609), .C2(n10093), .ZN(n8087) );
  MUX2_X1 U9741 ( .A(n8080), .B(n8087), .S(n10152), .Z(n8082) );
  NAND2_X1 U9742 ( .A1(n8563), .A2(n9066), .ZN(n8081) );
  OAI211_X1 U9743 ( .C1(n8091), .C2(n9074), .A(n8082), .B(n8081), .ZN(P2_U3423) );
  MUX2_X1 U9744 ( .A(n8083), .B(n8087), .S(n7308), .Z(n8086) );
  INV_X1 U9745 ( .A(n8561), .ZN(n8084) );
  AOI22_X1 U9746 ( .A1(n8563), .A2(n10101), .B1(n10102), .B2(n8084), .ZN(n8085) );
  OAI211_X1 U9747 ( .C1(n8091), .C2(n8917), .A(n8086), .B(n8085), .ZN(P2_U3222) );
  MUX2_X1 U9748 ( .A(n8088), .B(n8087), .S(n10166), .Z(n8090) );
  NAND2_X1 U9749 ( .A1(n8563), .A2(n8967), .ZN(n8089) );
  OAI211_X1 U9750 ( .C1(n8975), .C2(n8091), .A(n8090), .B(n8089), .ZN(P2_U3470) );
  INV_X1 U9751 ( .A(n8972), .ZN(n8100) );
  OAI211_X1 U9752 ( .C1(n8094), .C2(n8093), .A(n8092), .B(n8591), .ZN(n8099)
         );
  OAI21_X1 U9753 ( .B1(n8583), .B2(n8442), .A(n8095), .ZN(n8097) );
  NOR2_X1 U9754 ( .A1(n8560), .A2(n8196), .ZN(n8096) );
  AOI211_X1 U9755 ( .C1(n8580), .C2(n8608), .A(n8097), .B(n8096), .ZN(n8098)
         );
  OAI211_X1 U9756 ( .C1(n8100), .C2(n8602), .A(n8099), .B(n8098), .ZN(P2_U3164) );
  OAI21_X1 U9757 ( .B1(n8597), .B2(n8102), .A(n8101), .ZN(n8103) );
  AOI21_X1 U9758 ( .B1(n8595), .B2(n8610), .A(n8103), .ZN(n8104) );
  OAI21_X1 U9759 ( .B1(n8105), .B2(n8560), .A(n8104), .ZN(n8112) );
  INV_X1 U9760 ( .A(n8028), .ZN(n8110) );
  AOI21_X1 U9761 ( .B1(n8107), .B2(n8109), .A(n8106), .ZN(n8108) );
  AOI211_X1 U9762 ( .C1(n8110), .C2(n8109), .A(n8588), .B(n8108), .ZN(n8111)
         );
  AOI211_X1 U9763 ( .C1(n10150), .C2(n8586), .A(n8112), .B(n8111), .ZN(n8113)
         );
  INV_X1 U9764 ( .A(n8113), .ZN(P2_U3161) );
  NOR2_X1 U9765 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n8147) );
  NOR2_X1 U9766 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8145) );
  NOR2_X1 U9767 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n8143) );
  NOR2_X1 U9768 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8141) );
  NOR2_X1 U9769 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8139) );
  NOR2_X1 U9770 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8137) );
  NOR2_X1 U9771 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8135) );
  NOR2_X1 U9772 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8133) );
  NOR2_X1 U9773 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8131) );
  NOR2_X1 U9774 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8129) );
  NOR2_X1 U9775 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8126) );
  NOR2_X1 U9776 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8124) );
  NOR2_X1 U9777 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8122) );
  NOR2_X1 U9778 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8120) );
  NAND2_X1 U9779 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n8118) );
  XOR2_X1 U9780 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10360) );
  NAND2_X1 U9781 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8116) );
  XOR2_X1 U9782 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10358) );
  AOI21_X1 U9783 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10167) );
  NAND3_X1 U9784 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10169) );
  OAI21_X1 U9785 ( .B1(n10167), .B2(n8114), .A(n10169), .ZN(n10357) );
  NAND2_X1 U9786 ( .A1(n10358), .A2(n10357), .ZN(n8115) );
  NAND2_X1 U9787 ( .A1(n8116), .A2(n8115), .ZN(n10359) );
  NAND2_X1 U9788 ( .A1(n10360), .A2(n10359), .ZN(n8117) );
  NAND2_X1 U9789 ( .A1(n8118), .A2(n8117), .ZN(n10362) );
  XNOR2_X1 U9790 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10361) );
  NOR2_X1 U9791 ( .A1(n10362), .A2(n10361), .ZN(n8119) );
  NOR2_X1 U9792 ( .A1(n8120), .A2(n8119), .ZN(n10350) );
  XNOR2_X1 U9793 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n10349) );
  NOR2_X1 U9794 ( .A1(n10350), .A2(n10349), .ZN(n8121) );
  NOR2_X1 U9795 ( .A1(n8122), .A2(n8121), .ZN(n10348) );
  XNOR2_X1 U9796 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10347) );
  NOR2_X1 U9797 ( .A1(n10348), .A2(n10347), .ZN(n8123) );
  NOR2_X1 U9798 ( .A1(n8124), .A2(n8123), .ZN(n10354) );
  XNOR2_X1 U9799 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10353) );
  NOR2_X1 U9800 ( .A1(n10354), .A2(n10353), .ZN(n8125) );
  NOR2_X1 U9801 ( .A1(n8126), .A2(n8125), .ZN(n10356) );
  INV_X1 U9802 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9473) );
  AOI22_X1 U9803 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9473), .B1(
        P1_ADDR_REG_8__SCAN_IN), .B2(n8127), .ZN(n10355) );
  NOR2_X1 U9804 ( .A1(n10356), .A2(n10355), .ZN(n8128) );
  XNOR2_X1 U9805 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n10351) );
  NOR2_X1 U9806 ( .A1(n10352), .A2(n10351), .ZN(n8130) );
  XNOR2_X1 U9807 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10188) );
  NOR2_X1 U9808 ( .A1(n10189), .A2(n10188), .ZN(n8132) );
  XNOR2_X1 U9809 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10186) );
  NOR2_X1 U9810 ( .A1(n10187), .A2(n10186), .ZN(n8134) );
  XNOR2_X1 U9811 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10184) );
  NOR2_X1 U9812 ( .A1(n10185), .A2(n10184), .ZN(n8136) );
  XNOR2_X1 U9813 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10182) );
  NOR2_X1 U9814 ( .A1(n10183), .A2(n10182), .ZN(n8138) );
  XNOR2_X1 U9815 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10180) );
  NOR2_X1 U9816 ( .A1(n10181), .A2(n10180), .ZN(n8140) );
  NOR2_X1 U9817 ( .A1(n8141), .A2(n8140), .ZN(n10179) );
  XNOR2_X1 U9818 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10178) );
  NOR2_X1 U9819 ( .A1(n10179), .A2(n10178), .ZN(n8142) );
  NOR2_X1 U9820 ( .A1(n8143), .A2(n8142), .ZN(n10177) );
  XNOR2_X1 U9821 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10176) );
  NOR2_X1 U9822 ( .A1(n10177), .A2(n10176), .ZN(n8144) );
  NOR2_X1 U9823 ( .A1(n8145), .A2(n8144), .ZN(n10175) );
  XNOR2_X1 U9824 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10174) );
  NOR2_X1 U9825 ( .A1(n10175), .A2(n10174), .ZN(n8146) );
  NOR2_X1 U9826 ( .A1(n8147), .A2(n8146), .ZN(n8148) );
  AND2_X1 U9827 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8148), .ZN(n10171) );
  NOR2_X1 U9828 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10171), .ZN(n8149) );
  NOR2_X1 U9829 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n8148), .ZN(n10172) );
  NOR2_X1 U9830 ( .A1(n8149), .A2(n10172), .ZN(n8151) );
  XNOR2_X1 U9831 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8150) );
  XNOR2_X1 U9832 ( .A(n8151), .B(n8150), .ZN(ADD_1068_U4) );
  OAI21_X1 U9833 ( .B1(n8153), .B2(n8159), .A(n8152), .ZN(n9892) );
  INV_X1 U9834 ( .A(n9892), .ZN(n8169) );
  INV_X1 U9835 ( .A(n8154), .ZN(n8156) );
  OAI21_X1 U9836 ( .B1(n8157), .B2(n8156), .A(n8155), .ZN(n8240) );
  NOR2_X1 U9837 ( .A1(n8240), .A2(n8241), .ZN(n8260) );
  OAI21_X1 U9838 ( .B1(n8260), .B2(n8259), .A(n8258), .ZN(n8257) );
  NAND2_X1 U9839 ( .A1(n8257), .A2(n8158), .ZN(n8160) );
  XNOR2_X1 U9840 ( .A(n8160), .B(n8159), .ZN(n8161) );
  NAND2_X1 U9841 ( .A1(n9369), .A2(n9322), .ZN(n9256) );
  OAI21_X1 U9842 ( .B1(n8161), .B2(n9757), .A(n9256), .ZN(n9890) );
  NAND2_X1 U9843 ( .A1(n9890), .A2(n7937), .ZN(n8168) );
  OAI211_X1 U9844 ( .C1(n9974), .C2(n8162), .A(n8009), .B(n9764), .ZN(n8163)
         );
  NAND2_X1 U9845 ( .A1(n9367), .A2(n9324), .ZN(n9255) );
  NAND2_X1 U9846 ( .A1(n8163), .A2(n9255), .ZN(n9891) );
  NOR2_X1 U9847 ( .A1(n9715), .A2(n9974), .ZN(n8166) );
  OAI22_X1 U9848 ( .A1(n10344), .A2(n8164), .B1(n9262), .B2(n9780), .ZN(n8165)
         );
  AOI211_X1 U9849 ( .C1(n9891), .C2(n9788), .A(n8166), .B(n8165), .ZN(n8167)
         );
  OAI211_X1 U9850 ( .C1(n8169), .C2(n9793), .A(n8168), .B(n8167), .ZN(P1_U3284) );
  INV_X1 U9851 ( .A(n8170), .ZN(n8174) );
  OAI22_X1 U9852 ( .A1(n9715), .A2(n8172), .B1(n8171), .B2(n10344), .ZN(n8173)
         );
  AOI21_X1 U9853 ( .B1(n9788), .B2(n8174), .A(n8173), .ZN(n8178) );
  OAI21_X1 U9854 ( .B1(n9393), .B2(n9780), .A(n8175), .ZN(n8176) );
  NAND2_X1 U9855 ( .A1(n8176), .A2(n7937), .ZN(n8177) );
  OAI211_X1 U9856 ( .C1(n8179), .C2(n9793), .A(n8178), .B(n8177), .ZN(P1_U3291) );
  INV_X1 U9857 ( .A(n8180), .ZN(n8181) );
  MUX2_X1 U9858 ( .A(n5779), .B(n8181), .S(n7308), .Z(n8184) );
  INV_X1 U9859 ( .A(n8458), .ZN(n8182) );
  AOI22_X1 U9860 ( .A1(n8460), .A2(n10101), .B1(n10102), .B2(n8182), .ZN(n8183) );
  OAI211_X1 U9861 ( .C1(n8185), .C2(n10086), .A(n8184), .B(n8183), .ZN(
        P2_U3223) );
  INV_X1 U9862 ( .A(n8186), .ZN(n8211) );
  OAI222_X1 U9863 ( .A1(n9994), .A2(n8211), .B1(n8188), .B2(P1_U3086), .C1(
        n8187), .C2(n9995), .ZN(P1_U3335) );
  OR2_X1 U9864 ( .A1(n8189), .A2(n8193), .ZN(n8190) );
  NAND2_X1 U9865 ( .A1(n8191), .A2(n8190), .ZN(n9075) );
  XOR2_X1 U9866 ( .A(n8193), .B(n8192), .Z(n8194) );
  OAI222_X1 U9867 ( .A1(n8896), .A2(n8442), .B1(n8898), .B2(n8455), .C1(n8894), 
        .C2(n8194), .ZN(n8971) );
  NAND2_X1 U9868 ( .A1(n8971), .A2(n7308), .ZN(n8199) );
  NAND2_X1 U9869 ( .A1(n10107), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8195) );
  OAI21_X1 U9870 ( .B1(n8196), .B2(n8874), .A(n8195), .ZN(n8197) );
  AOI21_X1 U9871 ( .B1(n8972), .B2(n10101), .A(n8197), .ZN(n8198) );
  OAI211_X1 U9872 ( .C1(n9075), .C2(n8917), .A(n8199), .B(n8198), .ZN(P2_U3221) );
  NOR2_X1 U9873 ( .A1(n4379), .A2(n4307), .ZN(n8201) );
  XNOR2_X1 U9874 ( .A(n8201), .B(n8200), .ZN(n8202) );
  NAND2_X1 U9875 ( .A1(n8202), .A2(n9302), .ZN(n8208) );
  OAI22_X1 U9876 ( .A1(n9326), .A2(n8204), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8203), .ZN(n8205) );
  AOI21_X1 U9877 ( .B1(n9343), .B2(n8206), .A(n8205), .ZN(n8207) );
  OAI211_X1 U9878 ( .C1(n9341), .C2(n8209), .A(n8208), .B(n8207), .ZN(P1_U3227) );
  OAI222_X1 U9879 ( .A1(P2_U3151), .A2(n8212), .B1(n9093), .B2(n8211), .C1(
        n8210), .C2(n9097), .ZN(P2_U3275) );
  INV_X1 U9880 ( .A(n8460), .ZN(n8216) );
  MUX2_X1 U9881 ( .A(n8214), .B(n8213), .S(n10166), .Z(n8215) );
  OAI21_X1 U9882 ( .B1(n8216), .B2(n8961), .A(n8215), .ZN(P2_U3469) );
  OAI22_X1 U9883 ( .A1(n10344), .A2(n8217), .B1(n8229), .B2(n9780), .ZN(n8218)
         );
  AOI21_X1 U9884 ( .B1(n10331), .B2(n8219), .A(n8218), .ZN(n8222) );
  NAND2_X1 U9885 ( .A1(n8220), .A2(n10333), .ZN(n8221) );
  OAI211_X1 U9886 ( .C1(n8223), .C2(n10341), .A(n8222), .B(n8221), .ZN(n8224)
         );
  INV_X1 U9887 ( .A(n8224), .ZN(n8225) );
  OAI21_X1 U9888 ( .B1(n8226), .B2(n9712), .A(n8225), .ZN(P1_U3287) );
  OAI21_X1 U9889 ( .B1(n8228), .B2(n4284), .A(n8227), .ZN(n8237) );
  INV_X1 U9890 ( .A(n8229), .ZN(n8230) );
  NAND2_X1 U9891 ( .A1(n9328), .A2(n8230), .ZN(n8234) );
  NAND2_X1 U9892 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9446) );
  INV_X1 U9893 ( .A(n9446), .ZN(n8231) );
  AOI21_X1 U9894 ( .B1(n9339), .B2(n8232), .A(n8231), .ZN(n8233) );
  OAI211_X1 U9895 ( .C1(n8235), .C2(n9331), .A(n8234), .B(n8233), .ZN(n8236)
         );
  AOI21_X1 U9896 ( .B1(n8237), .B2(n9302), .A(n8236), .ZN(n8238) );
  INV_X1 U9897 ( .A(n8238), .ZN(P1_U3239) );
  OAI21_X1 U9898 ( .B1(n8239), .B2(n8241), .A(n8255), .ZN(n8245) );
  INV_X1 U9899 ( .A(n8245), .ZN(n10068) );
  INV_X1 U9900 ( .A(n8264), .ZN(n8246) );
  AOI22_X1 U9901 ( .A1(n9369), .A2(n9324), .B1(n9322), .B2(n9371), .ZN(n8330)
         );
  INV_X1 U9902 ( .A(n8330), .ZN(n8244) );
  AOI21_X1 U9903 ( .B1(n8241), .B2(n8240), .A(n8260), .ZN(n8242) );
  NOR2_X1 U9904 ( .A1(n8242), .A2(n9757), .ZN(n8243) );
  AOI211_X1 U9905 ( .C1(n8246), .C2(n8245), .A(n8244), .B(n8243), .ZN(n10066)
         );
  MUX2_X1 U9906 ( .A(n8247), .B(n10066), .S(n10344), .Z(n8252) );
  AOI211_X1 U9907 ( .C1(n10063), .C2(n8248), .A(n9784), .B(n8267), .ZN(n10062)
         );
  OAI22_X1 U9908 ( .A1(n9715), .A2(n8249), .B1(n8331), .B2(n9780), .ZN(n8250)
         );
  AOI21_X1 U9909 ( .B1(n10062), .B2(n9788), .A(n8250), .ZN(n8251) );
  OAI211_X1 U9910 ( .C1(n10068), .C2(n8271), .A(n8252), .B(n8251), .ZN(
        P1_U3286) );
  INV_X1 U9911 ( .A(n8253), .ZN(n8254) );
  NAND2_X1 U9912 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  XNOR2_X1 U9913 ( .A(n8258), .B(n8256), .ZN(n9895) );
  INV_X1 U9914 ( .A(n8257), .ZN(n8262) );
  NOR3_X1 U9915 ( .A1(n8260), .A2(n8259), .A3(n8258), .ZN(n8261) );
  OAI21_X1 U9916 ( .B1(n8262), .B2(n8261), .A(n9778), .ZN(n8263) );
  AOI22_X1 U9917 ( .A1(n9368), .A2(n9324), .B1(n9322), .B2(n9370), .ZN(n9170)
         );
  OAI211_X1 U9918 ( .C1(n9895), .C2(n8264), .A(n8263), .B(n9170), .ZN(n9896)
         );
  OAI22_X1 U9919 ( .A1(n10344), .A2(n8265), .B1(n9175), .B2(n9780), .ZN(n8266)
         );
  AOI21_X1 U9920 ( .B1(n10331), .B2(n9172), .A(n8266), .ZN(n8270) );
  OAI21_X1 U9921 ( .B1(n8267), .B2(n9979), .A(n9764), .ZN(n8268) );
  NOR2_X1 U9922 ( .A1(n8268), .A2(n8162), .ZN(n9897) );
  NAND2_X1 U9923 ( .A1(n9897), .A2(n9788), .ZN(n8269) );
  OAI211_X1 U9924 ( .C1(n9895), .C2(n8271), .A(n8270), .B(n8269), .ZN(n8272)
         );
  AOI21_X1 U9925 ( .B1(n9896), .B2(n7937), .A(n8272), .ZN(n8273) );
  INV_X1 U9926 ( .A(n8273), .ZN(P1_U3285) );
  INV_X1 U9927 ( .A(n9065), .ZN(n8317) );
  OAI211_X1 U9928 ( .C1(n8276), .C2(n8275), .A(n8274), .B(n8591), .ZN(n8280)
         );
  NAND2_X1 U9929 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8642) );
  OAI21_X1 U9930 ( .B1(n8583), .B2(n8897), .A(n8642), .ZN(n8278) );
  NOR2_X1 U9931 ( .A1(n8560), .A2(n8316), .ZN(n8277) );
  AOI211_X1 U9932 ( .C1(n8580), .C2(n8607), .A(n8278), .B(n8277), .ZN(n8279)
         );
  OAI211_X1 U9933 ( .C1(n8317), .C2(n8602), .A(n8280), .B(n8279), .ZN(P2_U3174) );
  OAI21_X1 U9934 ( .B1(n8282), .B2(n8285), .A(n8281), .ZN(n8355) );
  INV_X1 U9935 ( .A(n8355), .ZN(n8299) );
  NAND2_X1 U9936 ( .A1(n8284), .A2(n8283), .ZN(n8286) );
  XNOR2_X1 U9937 ( .A(n8286), .B(n8285), .ZN(n8290) );
  OAI22_X1 U9938 ( .A1(n8288), .A2(n9337), .B1(n9336), .B2(n8287), .ZN(n9201)
         );
  INV_X1 U9939 ( .A(n9201), .ZN(n8289) );
  OAI21_X1 U9940 ( .B1(n8290), .B2(n9757), .A(n8289), .ZN(n8349) );
  NAND2_X1 U9941 ( .A1(n8349), .A2(n7937), .ZN(n8298) );
  INV_X1 U9942 ( .A(n8291), .ZN(n8293) );
  AOI211_X1 U9943 ( .C1(n8354), .C2(n8293), .A(n9784), .B(n8292), .ZN(n8348)
         );
  NOR2_X1 U9944 ( .A1(n9204), .A2(n9715), .ZN(n8296) );
  OAI22_X1 U9945 ( .A1(n10344), .A2(n8294), .B1(n9198), .B2(n9780), .ZN(n8295)
         );
  AOI211_X1 U9946 ( .C1(n8348), .C2(n9788), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI211_X1 U9947 ( .C1(n8299), .C2(n9793), .A(n8298), .B(n8297), .ZN(P1_U3281) );
  INV_X1 U9948 ( .A(n6145), .ZN(n8426) );
  OAI222_X1 U9949 ( .A1(n9994), .A2(n8426), .B1(n8301), .B2(P1_U3086), .C1(
        n8300), .C2(n9995), .ZN(P1_U3334) );
  OAI21_X1 U9950 ( .B1(n8303), .B2(n5654), .A(n8302), .ZN(n8305) );
  OAI22_X1 U9951 ( .A1(n8304), .A2(n9337), .B1(n9336), .B2(n9338), .ZN(n9284)
         );
  AOI21_X1 U9952 ( .B1(n8305), .B2(n9778), .A(n9284), .ZN(n9882) );
  INV_X1 U9953 ( .A(n8292), .ZN(n8306) );
  AOI211_X1 U9954 ( .C1(n9880), .C2(n8306), .A(n9784), .B(n4767), .ZN(n9879)
         );
  NOR2_X1 U9955 ( .A1(n9287), .A2(n9715), .ZN(n8308) );
  OAI22_X1 U9956 ( .A1(n10344), .A2(n7659), .B1(n9281), .B2(n9780), .ZN(n8307)
         );
  AOI211_X1 U9957 ( .C1(n9879), .C2(n9788), .A(n8308), .B(n8307), .ZN(n8313)
         );
  OAI21_X1 U9958 ( .B1(n8311), .B2(n8310), .A(n8309), .ZN(n9878) );
  NAND2_X1 U9959 ( .A1(n9878), .A2(n10333), .ZN(n8312) );
  OAI211_X1 U9960 ( .C1(n9882), .C2(n10337), .A(n8313), .B(n8312), .ZN(
        P1_U3280) );
  XNOR2_X1 U9961 ( .A(n8314), .B(n8319), .ZN(n8315) );
  OAI222_X1 U9962 ( .A1(n8898), .A2(n8557), .B1(n8896), .B2(n8897), .C1(n8315), 
        .C2(n8894), .ZN(n8965) );
  OAI22_X1 U9963 ( .A1(n8317), .A2(n8778), .B1(n8316), .B2(n8874), .ZN(n8318)
         );
  OAI21_X1 U9964 ( .B1(n8965), .B2(n8318), .A(n7308), .ZN(n8322) );
  XOR2_X1 U9965 ( .A(n8320), .B(n8319), .Z(n9068) );
  NAND2_X1 U9966 ( .A1(n9068), .A2(n10104), .ZN(n8321) );
  OAI211_X1 U9967 ( .C1(n7308), .C2(n8323), .A(n8322), .B(n8321), .ZN(P2_U3220) );
  INV_X1 U9968 ( .A(n8324), .ZN(n8326) );
  NAND2_X1 U9969 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  XNOR2_X1 U9970 ( .A(n8328), .B(n8327), .ZN(n8335) );
  OAI22_X1 U9971 ( .A1(n9326), .A2(n8330), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8329), .ZN(n8333) );
  NOR2_X1 U9972 ( .A1(n9341), .A2(n8331), .ZN(n8332) );
  AOI211_X1 U9973 ( .C1(n10063), .C2(n9343), .A(n8333), .B(n8332), .ZN(n8334)
         );
  OAI21_X1 U9974 ( .B1(n8335), .B2(n9345), .A(n8334), .ZN(P1_U3213) );
  INV_X1 U9975 ( .A(n6155), .ZN(n8338) );
  AOI21_X1 U9976 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9988), .A(n8336), .ZN(
        n8337) );
  OAI21_X1 U9977 ( .B1(n8338), .B2(n9994), .A(n8337), .ZN(P1_U3332) );
  INV_X1 U9978 ( .A(n8339), .ZN(n8343) );
  OAI222_X1 U9979 ( .A1(n9995), .A2(n8341), .B1(n9994), .B2(n8343), .C1(
        P1_U3086), .C2(n8340), .ZN(P1_U3333) );
  OAI222_X1 U9980 ( .A1(n9097), .A2(n8344), .B1(n9093), .B2(n8343), .C1(
        P2_U3151), .C2(n8342), .ZN(P2_U3273) );
  NAND2_X1 U9981 ( .A1(n6155), .A2(n9082), .ZN(n8346) );
  OAI211_X1 U9982 ( .C1(n8347), .C2(n9097), .A(n8346), .B(n8345), .ZN(P2_U3272) );
  INV_X1 U9983 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8350) );
  NOR2_X1 U9984 ( .A1(n8349), .A2(n8348), .ZN(n8353) );
  MUX2_X1 U9985 ( .A(n8350), .B(n8353), .S(n10070), .Z(n8352) );
  AOI22_X1 U9986 ( .A1(n8355), .A2(n9952), .B1(n5687), .B2(n8354), .ZN(n8351)
         );
  NAND2_X1 U9987 ( .A1(n8352), .A2(n8351), .ZN(P1_U3489) );
  MUX2_X1 U9988 ( .A(n10196), .B(n8353), .S(n10073), .Z(n8357) );
  AOI22_X1 U9989 ( .A1(n8355), .A2(n9858), .B1(n6366), .B2(n8354), .ZN(n8356)
         );
  NAND2_X1 U9990 ( .A1(n8357), .A2(n8356), .ZN(P1_U3534) );
  INV_X1 U9991 ( .A(n8358), .ZN(n8362) );
  XNOR2_X1 U9992 ( .A(n8359), .B(n8362), .ZN(n8361) );
  AOI22_X1 U9993 ( .A1(n9364), .A2(n9322), .B1(n9324), .B2(n9362), .ZN(n9106)
         );
  INV_X1 U9994 ( .A(n9106), .ZN(n8360) );
  AOI21_X1 U9995 ( .B1(n8361), .B2(n9778), .A(n8360), .ZN(n9874) );
  XNOR2_X1 U9996 ( .A(n8363), .B(n8362), .ZN(n9875) );
  INV_X1 U9997 ( .A(n9875), .ZN(n8370) );
  AOI21_X1 U9998 ( .B1(n8364), .B2(n9967), .A(n9784), .ZN(n8366) );
  NAND2_X1 U9999 ( .A1(n8366), .A2(n9785), .ZN(n9873) );
  OAI22_X1 U10000 ( .A1(n10344), .A2(n10255), .B1(n9107), .B2(n9780), .ZN(
        n8367) );
  AOI21_X1 U10001 ( .B1(n9967), .B2(n10331), .A(n8367), .ZN(n8368) );
  OAI21_X1 U10002 ( .B1(n9873), .B2(n10341), .A(n8368), .ZN(n8369) );
  AOI21_X1 U10003 ( .B1(n8370), .B2(n10333), .A(n8369), .ZN(n8371) );
  OAI21_X1 U10004 ( .B1(n9712), .B2(n9874), .A(n8371), .ZN(P1_U3279) );
  INV_X1 U10005 ( .A(n8372), .ZN(n8376) );
  OAI222_X1 U10006 ( .A1(n9994), .A2(n8376), .B1(P1_U3086), .B2(n8374), .C1(
        n8373), .C2(n9995), .ZN(P1_U3331) );
  OAI222_X1 U10007 ( .A1(n6322), .A2(P2_U3151), .B1(n9093), .B2(n8376), .C1(
        n8375), .C2(n9097), .ZN(P2_U3271) );
  INV_X1 U10008 ( .A(n8377), .ZN(n9099) );
  OAI222_X1 U10009 ( .A1(n9994), .A2(n9099), .B1(P1_U3086), .B2(n8378), .C1(
        n10191), .C2(n9995), .ZN(P1_U3330) );
  NAND2_X1 U10010 ( .A1(n8379), .A2(n7308), .ZN(n8384) );
  NAND2_X1 U10011 ( .A1(n8380), .A2(n10102), .ZN(n8752) );
  OAI21_X1 U10012 ( .B1(n7308), .B2(n8381), .A(n8752), .ZN(n8382) );
  AOI21_X1 U10013 ( .B1(n6236), .B2(n10101), .A(n8382), .ZN(n8383) );
  OAI211_X1 U10014 ( .C1(n8385), .C2(n10086), .A(n8384), .B(n8383), .ZN(
        P2_U3204) );
  INV_X1 U10015 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8387) );
  OAI222_X1 U10016 ( .A1(n9994), .A2(n8386), .B1(n4999), .B2(P1_U3086), .C1(
        n8387), .C2(n9995), .ZN(P1_U3326) );
  OAI222_X1 U10017 ( .A1(n9995), .A2(n8389), .B1(n9994), .B2(n8388), .C1(
        P1_U3086), .C2(n9564), .ZN(P1_U3336) );
  INV_X1 U10018 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n8390) );
  MUX2_X2 U10019 ( .A(n8391), .B(n8390), .S(n6383), .Z(n8392) );
  OAI21_X1 U10020 ( .B1(n6685), .B2(n9978), .A(n8392), .ZN(P1_U3521) );
  NOR2_X1 U10021 ( .A1(n10337), .A2(n9807), .ZN(n9569) );
  NOR2_X1 U10022 ( .A1(n6685), .A2(n9715), .ZN(n8393) );
  AOI211_X1 U10023 ( .C1(n9712), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9569), .B(
        n8393), .ZN(n8394) );
  OAI21_X1 U10024 ( .B1(n8395), .B2(n10341), .A(n8394), .ZN(P1_U3263) );
  INV_X1 U10025 ( .A(n8396), .ZN(n9088) );
  OAI222_X1 U10026 ( .A1(n9994), .A2(n9088), .B1(n5674), .B2(P1_U3086), .C1(
        n8397), .C2(n9995), .ZN(P1_U3327) );
  NAND2_X1 U10027 ( .A1(n8419), .A2(n8398), .ZN(n8400) );
  NAND2_X1 U10028 ( .A1(n5555), .A2(n8406), .ZN(n8399) );
  NAND2_X1 U10029 ( .A1(n8400), .A2(n8399), .ZN(n8402) );
  XNOR2_X1 U10030 ( .A(n8402), .B(n8401), .ZN(n8408) );
  NOR2_X1 U10031 ( .A1(n8404), .A2(n8403), .ZN(n8405) );
  AOI21_X1 U10032 ( .B1(n8419), .B2(n8406), .A(n8405), .ZN(n8407) );
  XNOR2_X1 U10033 ( .A(n8408), .B(n8407), .ZN(n8416) );
  INV_X1 U10034 ( .A(n8416), .ZN(n8409) );
  NAND2_X1 U10035 ( .A1(n8409), .A2(n9302), .ZN(n8423) );
  OR2_X1 U10036 ( .A1(n8411), .A2(n8410), .ZN(n8415) );
  NAND4_X1 U10037 ( .A1(n8422), .A2(n9302), .A3(n8416), .A4(n8415), .ZN(n8421)
         );
  INV_X1 U10038 ( .A(n8412), .ZN(n8413) );
  AOI22_X1 U10039 ( .A1(n8413), .A2(n9339), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8414) );
  OAI21_X1 U10040 ( .B1(n9341), .B2(n9574), .A(n8414), .ZN(n8418) );
  NOR3_X1 U10041 ( .A1(n8416), .A2(n9345), .A3(n8415), .ZN(n8417) );
  AOI211_X1 U10042 ( .C1(n9343), .C2(n8419), .A(n8418), .B(n8417), .ZN(n8420)
         );
  OAI211_X1 U10043 ( .C1(n8423), .C2(n8422), .A(n8421), .B(n8420), .ZN(
        P1_U3220) );
  INV_X1 U10044 ( .A(n8424), .ZN(n9990) );
  OAI222_X1 U10045 ( .A1(n9097), .A2(n8425), .B1(n9093), .B2(n9990), .C1(
        P2_U3151), .C2(n5927), .ZN(P2_U3265) );
  OAI222_X1 U10046 ( .A1(n9097), .A2(n10233), .B1(n9093), .B2(n8426), .C1(
        n6341), .C2(P2_U3151), .ZN(P2_U3274) );
  INV_X1 U10047 ( .A(n8427), .ZN(n8435) );
  NOR2_X1 U10048 ( .A1(n8428), .A2(n10341), .ZN(n8434) );
  INV_X1 U10049 ( .A(n8429), .ZN(n8430) );
  AOI22_X1 U10050 ( .A1(n8430), .A2(n10336), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n10337), .ZN(n8431) );
  OAI21_X1 U10051 ( .B1(n8432), .B2(n9715), .A(n8431), .ZN(n8433) );
  INV_X1 U10052 ( .A(n8437), .ZN(n8438) );
  AOI21_X1 U10053 ( .B1(n8440), .B2(n8439), .A(n8438), .ZN(n8446) );
  NAND2_X1 U10054 ( .A1(n8595), .A2(n8909), .ZN(n8441) );
  NAND2_X1 U10055 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8661) );
  OAI211_X1 U10056 ( .C1(n8597), .C2(n8442), .A(n8441), .B(n8661), .ZN(n8443)
         );
  AOI21_X1 U10057 ( .B1(n8912), .B2(n8599), .A(n8443), .ZN(n8445) );
  NAND2_X1 U10058 ( .A1(n9059), .A2(n8586), .ZN(n8444) );
  OAI211_X1 U10059 ( .C1(n8446), .C2(n8588), .A(n8445), .B(n8444), .ZN(
        P2_U3155) );
  XNOR2_X1 U10060 ( .A(n8525), .B(n8788), .ZN(n8451) );
  AOI22_X1 U10061 ( .A1(n8825), .A2(n8580), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8448) );
  NAND2_X1 U10062 ( .A1(n8806), .A2(n8599), .ZN(n8447) );
  OAI211_X1 U10063 ( .C1(n8526), .C2(n8583), .A(n8448), .B(n8447), .ZN(n8449)
         );
  AOI21_X1 U10064 ( .B1(n9013), .B2(n8586), .A(n8449), .ZN(n8450) );
  OAI21_X1 U10065 ( .B1(n8451), .B2(n8588), .A(n8450), .ZN(P2_U3156) );
  NAND2_X1 U10066 ( .A1(n8453), .A2(n8452), .ZN(n8549) );
  XNOR2_X1 U10067 ( .A(n8549), .B(n8551), .ZN(n8553) );
  XOR2_X1 U10068 ( .A(n8552), .B(n8553), .Z(n8462) );
  OAI21_X1 U10069 ( .B1(n8583), .B2(n8455), .A(n8454), .ZN(n8456) );
  AOI21_X1 U10070 ( .B1(n8580), .B2(n8610), .A(n8456), .ZN(n8457) );
  OAI21_X1 U10071 ( .B1(n8458), .B2(n8560), .A(n8457), .ZN(n8459) );
  AOI21_X1 U10072 ( .B1(n8460), .B2(n8586), .A(n8459), .ZN(n8461) );
  OAI21_X1 U10073 ( .B1(n8462), .B2(n8588), .A(n8461), .ZN(P2_U3157) );
  INV_X1 U10074 ( .A(n6447), .ZN(n9035) );
  AOI21_X1 U10075 ( .B1(n8464), .B2(n8463), .A(n8588), .ZN(n8466) );
  NAND2_X1 U10076 ( .A1(n8466), .A2(n8465), .ZN(n8472) );
  NAND2_X1 U10077 ( .A1(n8850), .A2(n8595), .ZN(n8468) );
  OAI211_X1 U10078 ( .C1(n8469), .C2(n8597), .A(n8468), .B(n8467), .ZN(n8470)
         );
  AOI21_X1 U10079 ( .B1(n8854), .B2(n8599), .A(n8470), .ZN(n8471) );
  OAI211_X1 U10080 ( .C1(n9035), .C2(n8602), .A(n8472), .B(n8471), .ZN(
        P2_U3159) );
  INV_X1 U10081 ( .A(n8484), .ZN(n8475) );
  XNOR2_X1 U10082 ( .A(n8759), .B(n8473), .ZN(n8474) );
  XNOR2_X1 U10083 ( .A(n8480), .B(n8474), .ZN(n8482) );
  INV_X1 U10084 ( .A(n8482), .ZN(n8487) );
  NAND3_X1 U10085 ( .A1(n8475), .A2(n8487), .A3(n8591), .ZN(n8491) );
  NAND2_X1 U10086 ( .A1(n8605), .A2(n8595), .ZN(n8478) );
  AOI22_X1 U10087 ( .A1(n8476), .A2(n8599), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8477) );
  OAI211_X1 U10088 ( .C1(n8584), .C2(n8597), .A(n8478), .B(n8477), .ZN(n8479)
         );
  AOI21_X1 U10089 ( .B1(n8480), .B2(n8586), .A(n8479), .ZN(n8490) );
  INV_X1 U10090 ( .A(n8481), .ZN(n8483) );
  NAND4_X1 U10091 ( .A1(n8484), .A2(n8591), .A3(n8483), .A4(n8482), .ZN(n8489)
         );
  INV_X1 U10092 ( .A(n8485), .ZN(n8486) );
  NAND4_X1 U10093 ( .A1(n8487), .A2(n8486), .A3(n8768), .A4(n8591), .ZN(n8488)
         );
  NAND4_X1 U10094 ( .A1(n8491), .A2(n8490), .A3(n8489), .A4(n8488), .ZN(
        P2_U3160) );
  XOR2_X1 U10095 ( .A(n8493), .B(n8492), .Z(n8499) );
  AOI22_X1 U10096 ( .A1(n8850), .A2(n8580), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8495) );
  NAND2_X1 U10097 ( .A1(n8828), .A2(n8599), .ZN(n8494) );
  OAI211_X1 U10098 ( .C1(n8496), .C2(n8583), .A(n8495), .B(n8494), .ZN(n8497)
         );
  AOI21_X1 U10099 ( .B1(n9025), .B2(n8586), .A(n8497), .ZN(n8498) );
  OAI21_X1 U10100 ( .B1(n8499), .B2(n8588), .A(n8498), .ZN(P2_U3163) );
  XOR2_X1 U10101 ( .A(n8500), .B(n4311), .Z(n8505) );
  NAND2_X1 U10102 ( .A1(n8776), .A2(n8595), .ZN(n8502) );
  AOI22_X1 U10103 ( .A1(n8779), .A2(n8599), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8501) );
  OAI211_X1 U10104 ( .C1(n8526), .C2(n8597), .A(n8502), .B(n8501), .ZN(n8503)
         );
  AOI21_X1 U10105 ( .B1(n9001), .B2(n8586), .A(n8503), .ZN(n8504) );
  OAI21_X1 U10106 ( .B1(n8505), .B2(n8588), .A(n8504), .ZN(P2_U3165) );
  INV_X1 U10107 ( .A(n9048), .ZN(n8514) );
  OAI211_X1 U10108 ( .C1(n8508), .C2(n8507), .A(n8506), .B(n8591), .ZN(n8513)
         );
  NAND2_X1 U10109 ( .A1(n8595), .A2(n8885), .ZN(n8509) );
  NAND2_X1 U10110 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8697) );
  OAI211_X1 U10111 ( .C1(n8597), .C2(n8510), .A(n8509), .B(n8697), .ZN(n8511)
         );
  AOI21_X1 U10112 ( .B1(n8887), .B2(n8599), .A(n8511), .ZN(n8512) );
  OAI211_X1 U10113 ( .C1(n8514), .C2(n8602), .A(n8513), .B(n8512), .ZN(
        P2_U3166) );
  INV_X1 U10114 ( .A(n8572), .ZN(n8515) );
  AOI21_X1 U10115 ( .B1(n8517), .B2(n8516), .A(n8515), .ZN(n8522) );
  NAND2_X1 U10116 ( .A1(n8595), .A2(n8871), .ZN(n8518) );
  NAND2_X1 U10117 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8718) );
  OAI211_X1 U10118 ( .C1(n8597), .C2(n8895), .A(n8518), .B(n8718), .ZN(n8519)
         );
  AOI21_X1 U10119 ( .B1(n8873), .B2(n8599), .A(n8519), .ZN(n8521) );
  NAND2_X1 U10120 ( .A1(n8948), .A2(n8586), .ZN(n8520) );
  OAI211_X1 U10121 ( .C1(n8522), .C2(n8588), .A(n8521), .B(n8520), .ZN(
        P2_U3168) );
  XNOR2_X1 U10122 ( .A(n8527), .B(n8526), .ZN(n8528) );
  AOI22_X1 U10123 ( .A1(n8812), .A2(n8580), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8530) );
  NAND2_X1 U10124 ( .A1(n8789), .A2(n8599), .ZN(n8529) );
  OAI211_X1 U10125 ( .C1(n6469), .C2(n8583), .A(n8530), .B(n8529), .ZN(n8531)
         );
  AOI21_X1 U10126 ( .B1(n9007), .B2(n8586), .A(n8531), .ZN(n8532) );
  INV_X1 U10127 ( .A(n6277), .ZN(n8541) );
  OAI21_X1 U10128 ( .B1(n4366), .B2(n8534), .A(n8533), .ZN(n8535) );
  NAND2_X1 U10129 ( .A1(n8535), .A2(n8591), .ZN(n8540) );
  AOI22_X1 U10130 ( .A1(n8837), .A2(n8595), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8536) );
  OAI21_X1 U10131 ( .B1(n8537), .B2(n8597), .A(n8536), .ZN(n8538) );
  AOI21_X1 U10132 ( .B1(n8840), .B2(n8599), .A(n8538), .ZN(n8539) );
  OAI211_X1 U10133 ( .C1(n8541), .C2(n8602), .A(n8540), .B(n8539), .ZN(
        P2_U3173) );
  XOR2_X1 U10134 ( .A(n8543), .B(n8542), .Z(n8548) );
  AOI22_X1 U10135 ( .A1(n8837), .A2(n8580), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8545) );
  NAND2_X1 U10136 ( .A1(n8815), .A2(n8599), .ZN(n8544) );
  OAI211_X1 U10137 ( .C1(n8788), .C2(n8583), .A(n8545), .B(n8544), .ZN(n8546)
         );
  AOI21_X1 U10138 ( .B1(n9019), .B2(n8586), .A(n8546), .ZN(n8547) );
  OAI21_X1 U10139 ( .B1(n8548), .B2(n8588), .A(n8547), .ZN(P2_U3175) );
  INV_X1 U10140 ( .A(n8549), .ZN(n8550) );
  AOI22_X1 U10141 ( .A1(n8553), .A2(n8552), .B1(n8551), .B2(n8550), .ZN(n8555)
         );
  XNOR2_X1 U10142 ( .A(n8555), .B(n8554), .ZN(n8565) );
  OAI21_X1 U10143 ( .B1(n8583), .B2(n8557), .A(n8556), .ZN(n8558) );
  AOI21_X1 U10144 ( .B1(n8580), .B2(n8609), .A(n8558), .ZN(n8559) );
  OAI21_X1 U10145 ( .B1(n8561), .B2(n8560), .A(n8559), .ZN(n8562) );
  AOI21_X1 U10146 ( .B1(n8563), .B2(n8586), .A(n8562), .ZN(n8564) );
  OAI21_X1 U10147 ( .B1(n8565), .B2(n8588), .A(n8564), .ZN(P2_U3176) );
  AND2_X1 U10148 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8735) );
  AOI21_X1 U10149 ( .B1(n8863), .B2(n8595), .A(n8735), .ZN(n8567) );
  NAND2_X1 U10150 ( .A1(n8599), .A2(n8866), .ZN(n8566) );
  OAI211_X1 U10151 ( .C1(n8568), .C2(n8597), .A(n8567), .B(n8566), .ZN(n8576)
         );
  INV_X1 U10152 ( .A(n8569), .ZN(n8571) );
  NAND3_X1 U10153 ( .A1(n8572), .A2(n8571), .A3(n8570), .ZN(n8573) );
  AOI21_X1 U10154 ( .B1(n8574), .B2(n8573), .A(n8588), .ZN(n8575) );
  AOI211_X1 U10155 ( .C1(n9041), .C2(n8586), .A(n8576), .B(n8575), .ZN(n8577)
         );
  INV_X1 U10156 ( .A(n8577), .ZN(P2_U3178) );
  XOR2_X1 U10157 ( .A(n8579), .B(n8578), .Z(n8589) );
  AOI22_X1 U10158 ( .A1(n8771), .A2(n8599), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8582) );
  NAND2_X1 U10159 ( .A1(n8767), .A2(n8580), .ZN(n8581) );
  OAI211_X1 U10160 ( .C1(n8584), .C2(n8583), .A(n8582), .B(n8581), .ZN(n8585)
         );
  AOI21_X1 U10161 ( .B1(n8995), .B2(n8586), .A(n8585), .ZN(n8587) );
  OAI21_X1 U10162 ( .B1(n8589), .B2(n8588), .A(n8587), .ZN(P2_U3180) );
  OAI211_X1 U10163 ( .C1(n8594), .C2(n8593), .A(n8592), .B(n8591), .ZN(n8601)
         );
  NAND2_X1 U10164 ( .A1(n8595), .A2(n8870), .ZN(n8596) );
  NAND2_X1 U10165 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8676) );
  OAI211_X1 U10166 ( .C1(n8597), .C2(n8897), .A(n8596), .B(n8676), .ZN(n8598)
         );
  AOI21_X1 U10167 ( .B1(n8899), .B2(n8599), .A(n8598), .ZN(n8600) );
  OAI211_X1 U10168 ( .C1(n9056), .C2(n8602), .A(n8601), .B(n8600), .ZN(
        P2_U3181) );
  INV_X1 U10169 ( .A(n8603), .ZN(n8751) );
  MUX2_X1 U10170 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8751), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10171 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8604), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10172 ( .A(n8605), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8614), .Z(
        P2_U3520) );
  MUX2_X1 U10173 ( .A(n8759), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8614), .Z(
        P2_U3519) );
  MUX2_X1 U10174 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8768), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10175 ( .A(n8776), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8614), .Z(
        P2_U3517) );
  INV_X1 U10176 ( .A(n8614), .ZN(n8611) );
  MUX2_X1 U10177 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8767), .S(n8611), .Z(
        P2_U3516) );
  MUX2_X1 U10178 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8803), .S(n8611), .Z(
        P2_U3515) );
  MUX2_X1 U10179 ( .A(n8812), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8614), .Z(
        P2_U3514) );
  MUX2_X1 U10180 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8825), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10181 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8837), .S(n8611), .Z(
        P2_U3512) );
  MUX2_X1 U10182 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8850), .S(n8611), .Z(
        P2_U3511) );
  MUX2_X1 U10183 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8863), .S(n8611), .Z(
        P2_U3510) );
  MUX2_X1 U10184 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8871), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10185 ( .A(n8885), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8614), .Z(
        P2_U3508) );
  MUX2_X1 U10186 ( .A(n8870), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8614), .Z(
        P2_U3507) );
  MUX2_X1 U10187 ( .A(n8909), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8614), .Z(
        P2_U3506) );
  MUX2_X1 U10188 ( .A(n8606), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8614), .Z(
        P2_U3505) );
  MUX2_X1 U10189 ( .A(n8910), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8614), .Z(
        P2_U3504) );
  MUX2_X1 U10190 ( .A(n8607), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8614), .Z(
        P2_U3503) );
  MUX2_X1 U10191 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8608), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10192 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8609), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10193 ( .A(n8610), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8614), .Z(
        P2_U3500) );
  MUX2_X1 U10194 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n10080), .S(n8611), .Z(
        P2_U3499) );
  MUX2_X1 U10195 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8612), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10196 ( .A(n10079), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8614), .Z(
        P2_U3497) );
  MUX2_X1 U10197 ( .A(n10092), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8614), .Z(
        P2_U3496) );
  MUX2_X1 U10198 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8613), .S(P2_U3893), .Z(
        P2_U3495) );
  MUX2_X1 U10199 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n10094), .S(P2_U3893), .Z(
        P2_U3494) );
  MUX2_X1 U10200 ( .A(n8615), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8614), .Z(
        P2_U3493) );
  MUX2_X1 U10201 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5936), .S(P2_U3893), .Z(
        P2_U3492) );
  OAI21_X1 U10202 ( .B1(n8618), .B2(n8617), .A(n8616), .ZN(n8619) );
  AOI22_X1 U10203 ( .A1(n8736), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n8701), .B2(
        n8619), .ZN(n8634) );
  OAI21_X1 U10204 ( .B1(n8622), .B2(n8621), .A(n8620), .ZN(n8624) );
  AOI21_X1 U10205 ( .B1(n8723), .B2(n8624), .A(n8623), .ZN(n8633) );
  AND2_X1 U10206 ( .A1(n8626), .A2(n8625), .ZN(n8629) );
  OAI211_X1 U10207 ( .C1(n8629), .C2(n8628), .A(n8740), .B(n8627), .ZN(n8632)
         );
  NAND2_X1 U10208 ( .A1(n8742), .A2(n8630), .ZN(n8631) );
  NAND4_X1 U10209 ( .A1(n8634), .A2(n8633), .A3(n8632), .A4(n8631), .ZN(
        P2_U3186) );
  XNOR2_X1 U10210 ( .A(n8635), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n8648) );
  XNOR2_X1 U10211 ( .A(n8636), .B(n8966), .ZN(n8646) );
  INV_X1 U10212 ( .A(n8637), .ZN(n8638) );
  NAND3_X1 U10213 ( .A1(n8640), .A2(n8639), .A3(n8638), .ZN(n8641) );
  AOI21_X1 U10214 ( .B1(n8659), .B2(n8641), .A(n8694), .ZN(n8645) );
  NAND2_X1 U10215 ( .A1(n8736), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n8643) );
  OAI211_X1 U10216 ( .C1(n8721), .C2(n4731), .A(n8643), .B(n8642), .ZN(n8644)
         );
  AOI211_X1 U10217 ( .C1(n8646), .C2(n8723), .A(n8645), .B(n8644), .ZN(n8647)
         );
  OAI21_X1 U10218 ( .B1(n8648), .B2(n8734), .A(n8647), .ZN(P2_U3195) );
  OAI21_X1 U10219 ( .B1(n8651), .B2(n8650), .A(n8649), .ZN(n8652) );
  NAND2_X1 U10220 ( .A1(n8652), .A2(n8701), .ZN(n8668) );
  OAI21_X1 U10221 ( .B1(n8655), .B2(n8654), .A(n8653), .ZN(n8666) );
  INV_X1 U10222 ( .A(n8656), .ZN(n8657) );
  NAND3_X1 U10223 ( .A1(n8659), .A2(n8658), .A3(n8657), .ZN(n8660) );
  AOI21_X1 U10224 ( .B1(n8674), .B2(n8660), .A(n8694), .ZN(n8665) );
  NAND2_X1 U10225 ( .A1(n8736), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8662) );
  OAI211_X1 U10226 ( .C1(n8721), .C2(n8663), .A(n8662), .B(n8661), .ZN(n8664)
         );
  AOI211_X1 U10227 ( .C1(n8666), .C2(n8723), .A(n8665), .B(n8664), .ZN(n8667)
         );
  NAND2_X1 U10228 ( .A1(n8668), .A2(n8667), .ZN(P2_U3196) );
  OAI21_X1 U10229 ( .B1(n8670), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8669), .ZN(
        n8681) );
  INV_X1 U10230 ( .A(n8671), .ZN(n8672) );
  NAND3_X1 U10231 ( .A1(n8674), .A2(n8673), .A3(n8672), .ZN(n8675) );
  AOI21_X1 U10232 ( .B1(n8693), .B2(n8675), .A(n8694), .ZN(n8680) );
  NAND2_X1 U10233 ( .A1(n8736), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8677) );
  OAI211_X1 U10234 ( .C1(n8721), .C2(n8678), .A(n8677), .B(n8676), .ZN(n8679)
         );
  AOI211_X1 U10235 ( .C1(n8681), .C2(n8701), .A(n8680), .B(n8679), .ZN(n8686)
         );
  OAI21_X1 U10236 ( .B1(n8683), .B2(P2_REG1_REG_15__SCAN_IN), .A(n8682), .ZN(
        n8684) );
  NAND2_X1 U10237 ( .A1(n8684), .A2(n8723), .ZN(n8685) );
  NAND2_X1 U10238 ( .A1(n8686), .A2(n8685), .ZN(P2_U3197) );
  OAI21_X1 U10239 ( .B1(n8689), .B2(n8688), .A(n8687), .ZN(n8702) );
  INV_X1 U10240 ( .A(n8690), .ZN(n8691) );
  NAND3_X1 U10241 ( .A1(n8693), .A2(n8692), .A3(n8691), .ZN(n8695) );
  AOI21_X1 U10242 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n8700) );
  NAND2_X1 U10243 ( .A1(n8736), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8698) );
  OAI211_X1 U10244 ( .C1(n4631), .C2(n8721), .A(n8698), .B(n8697), .ZN(n8699)
         );
  AOI211_X1 U10245 ( .C1(n8702), .C2(n8701), .A(n8700), .B(n8699), .ZN(n8708)
         );
  OAI21_X1 U10246 ( .B1(n8705), .B2(n8704), .A(n8703), .ZN(n8706) );
  NAND2_X1 U10247 ( .A1(n8706), .A2(n8723), .ZN(n8707) );
  NAND2_X1 U10248 ( .A1(n8708), .A2(n8707), .ZN(P2_U3198) );
  INV_X1 U10249 ( .A(n8709), .ZN(n8711) );
  INV_X1 U10250 ( .A(n8732), .ZN(n8710) );
  AOI21_X1 U10251 ( .B1(n8711), .B2(n8876), .A(n8710), .ZN(n8727) );
  OAI21_X1 U10252 ( .B1(n8714), .B2(n8713), .A(n8712), .ZN(n8715) );
  NAND2_X1 U10253 ( .A1(n8715), .A2(n8740), .ZN(n8726) );
  OAI21_X1 U10254 ( .B1(n8717), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8716), .ZN(
        n8724) );
  NAND2_X1 U10255 ( .A1(n8736), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8719) );
  OAI211_X1 U10256 ( .C1(n8721), .C2(n8720), .A(n8719), .B(n8718), .ZN(n8722)
         );
  AOI21_X1 U10257 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8725) );
  OAI211_X1 U10258 ( .C1(n8727), .C2(n8734), .A(n8726), .B(n8725), .ZN(
        P2_U3199) );
  XOR2_X1 U10259 ( .A(n8729), .B(n8728), .Z(n8749) );
  INV_X1 U10260 ( .A(n8737), .ZN(n8738) );
  INV_X1 U10261 ( .A(n8743), .ZN(n8741) );
  NAND2_X1 U10262 ( .A1(n8741), .A2(n8740), .ZN(n8746) );
  AOI21_X1 U10263 ( .B1(n8743), .B2(P2_U3893), .A(n8742), .ZN(n8745) );
  NAND2_X1 U10264 ( .A1(n8751), .A2(n8750), .ZN(n8981) );
  OAI21_X1 U10265 ( .B1(n8981), .B2(n10107), .A(n8752), .ZN(n8754) );
  AOI21_X1 U10266 ( .B1(P2_REG2_REG_31__SCAN_IN), .B2(n10107), .A(n8754), .ZN(
        n8753) );
  OAI21_X1 U10267 ( .B1(n8983), .B2(n8901), .A(n8753), .ZN(P2_U3202) );
  AOI21_X1 U10268 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(n10107), .A(n8754), .ZN(
        n8755) );
  OAI21_X1 U10269 ( .B1(n8986), .B2(n8901), .A(n8755), .ZN(P2_U3203) );
  XNOR2_X1 U10270 ( .A(n8756), .B(n8758), .ZN(n8992) );
  INV_X1 U10271 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8760) );
  MUX2_X1 U10272 ( .A(n8760), .B(n8987), .S(n7308), .Z(n8763) );
  AOI22_X1 U10273 ( .A1(n8989), .A2(n10101), .B1(n10102), .B2(n8761), .ZN(
        n8762) );
  OAI211_X1 U10274 ( .C1(n8992), .C2(n8917), .A(n8763), .B(n8762), .ZN(
        P2_U3206) );
  XNOR2_X1 U10275 ( .A(n8764), .B(n8766), .ZN(n8998) );
  INV_X1 U10276 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8770) );
  XNOR2_X1 U10277 ( .A(n8765), .B(n8766), .ZN(n8769) );
  AOI222_X1 U10278 ( .A1(n10096), .A2(n8769), .B1(n8768), .B2(n10091), .C1(
        n8767), .C2(n10093), .ZN(n8993) );
  MUX2_X1 U10279 ( .A(n8770), .B(n8993), .S(n7308), .Z(n8773) );
  AOI22_X1 U10280 ( .A1(n8995), .A2(n10101), .B1(n10102), .B2(n8771), .ZN(
        n8772) );
  OAI211_X1 U10281 ( .C1(n8998), .C2(n8917), .A(n8773), .B(n8772), .ZN(
        P2_U3207) );
  XNOR2_X1 U10282 ( .A(n8774), .B(n8775), .ZN(n8777) );
  AOI222_X1 U10283 ( .A1(n10096), .A2(n8777), .B1(n8803), .B2(n10093), .C1(
        n8776), .C2(n10091), .ZN(n8999) );
  INV_X1 U10284 ( .A(n8778), .ZN(n8913) );
  AOI22_X1 U10285 ( .A1(n9001), .A2(n8913), .B1(n10102), .B2(n8779), .ZN(n8780) );
  AND2_X1 U10286 ( .A1(n8999), .A2(n8780), .ZN(n8785) );
  XNOR2_X1 U10287 ( .A(n8782), .B(n8781), .ZN(n9004) );
  INV_X1 U10288 ( .A(n9004), .ZN(n8783) );
  AOI22_X1 U10289 ( .A1(n8783), .A2(n10104), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10107), .ZN(n8784) );
  OAI21_X1 U10290 ( .B1(n8785), .B2(n10107), .A(n8784), .ZN(P2_U3208) );
  XOR2_X1 U10291 ( .A(n8786), .B(n8795), .Z(n8787) );
  OAI222_X1 U10292 ( .A1(n8898), .A2(n8788), .B1(n8896), .B2(n6469), .C1(n8787), .C2(n8894), .ZN(n8928) );
  AOI21_X1 U10293 ( .B1(n8913), .B2(n9007), .A(n8928), .ZN(n8799) );
  AOI22_X1 U10294 ( .A1(n8789), .A2(n10102), .B1(n10107), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8798) );
  INV_X1 U10295 ( .A(n8809), .ZN(n8792) );
  OAI21_X1 U10296 ( .B1(n8792), .B2(n8791), .A(n8790), .ZN(n8800) );
  OAI21_X1 U10297 ( .B1(n8800), .B2(n8794), .A(n8793), .ZN(n8796) );
  XNOR2_X1 U10298 ( .A(n8796), .B(n8795), .ZN(n9008) );
  NAND2_X1 U10299 ( .A1(n9008), .A2(n10104), .ZN(n8797) );
  OAI211_X1 U10300 ( .C1(n8799), .C2(n10107), .A(n8798), .B(n8797), .ZN(
        P2_U3209) );
  XNOR2_X1 U10301 ( .A(n8800), .B(n8802), .ZN(n9016) );
  INV_X1 U10302 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8805) );
  XOR2_X1 U10303 ( .A(n8801), .B(n8802), .Z(n8804) );
  AOI222_X1 U10304 ( .A1(n10096), .A2(n8804), .B1(n8825), .B2(n10093), .C1(
        n8803), .C2(n10091), .ZN(n9011) );
  MUX2_X1 U10305 ( .A(n8805), .B(n9011), .S(n7308), .Z(n8808) );
  AOI22_X1 U10306 ( .A1(n9013), .A2(n10101), .B1(n10102), .B2(n8806), .ZN(
        n8807) );
  OAI211_X1 U10307 ( .C1(n9016), .C2(n8917), .A(n8808), .B(n8807), .ZN(
        P2_U3210) );
  XNOR2_X1 U10308 ( .A(n8809), .B(n8811), .ZN(n9020) );
  INV_X1 U10309 ( .A(n9020), .ZN(n8818) );
  INV_X1 U10310 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8814) );
  XNOR2_X1 U10311 ( .A(n8810), .B(n8811), .ZN(n8813) );
  AOI222_X1 U10312 ( .A1(n10096), .A2(n8813), .B1(n8812), .B2(n10091), .C1(
        n8837), .C2(n10093), .ZN(n9017) );
  MUX2_X1 U10313 ( .A(n8814), .B(n9017), .S(n7308), .Z(n8817) );
  AOI22_X1 U10314 ( .A1(n9019), .A2(n10101), .B1(n10102), .B2(n8815), .ZN(
        n8816) );
  OAI211_X1 U10315 ( .C1(n8818), .C2(n8917), .A(n8817), .B(n8816), .ZN(
        P2_U3211) );
  XNOR2_X1 U10316 ( .A(n8820), .B(n8819), .ZN(n9026) );
  INV_X1 U10317 ( .A(n9026), .ZN(n8831) );
  INV_X1 U10318 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8827) );
  NAND2_X1 U10319 ( .A1(n8822), .A2(n8821), .ZN(n8824) );
  XNOR2_X1 U10320 ( .A(n8824), .B(n8823), .ZN(n8826) );
  AOI222_X1 U10321 ( .A1(n10096), .A2(n8826), .B1(n8850), .B2(n10093), .C1(
        n8825), .C2(n10091), .ZN(n9023) );
  MUX2_X1 U10322 ( .A(n8827), .B(n9023), .S(n7308), .Z(n8830) );
  AOI22_X1 U10323 ( .A1(n9025), .A2(n10101), .B1(n10102), .B2(n8828), .ZN(
        n8829) );
  OAI211_X1 U10324 ( .C1(n8831), .C2(n8917), .A(n8830), .B(n8829), .ZN(
        P2_U3212) );
  XOR2_X1 U10325 ( .A(n8832), .B(n8835), .Z(n9033) );
  INV_X1 U10326 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8839) );
  NOR2_X1 U10327 ( .A1(n8833), .A2(n8846), .ZN(n8849) );
  NOR2_X1 U10328 ( .A1(n8849), .A2(n8834), .ZN(n8836) );
  XNOR2_X1 U10329 ( .A(n8836), .B(n8835), .ZN(n8838) );
  AOI222_X1 U10330 ( .A1(n10096), .A2(n8838), .B1(n8837), .B2(n10091), .C1(
        n8863), .C2(n10093), .ZN(n9029) );
  MUX2_X1 U10331 ( .A(n8839), .B(n9029), .S(n7308), .Z(n8842) );
  AOI22_X1 U10332 ( .A1(n6277), .A2(n10101), .B1(n10102), .B2(n8840), .ZN(
        n8841) );
  OAI211_X1 U10333 ( .C1(n9033), .C2(n8917), .A(n8842), .B(n8841), .ZN(
        P2_U3213) );
  NAND2_X1 U10334 ( .A1(n8843), .A2(n8857), .ZN(n8845) );
  XNOR2_X1 U10335 ( .A(n8845), .B(n8844), .ZN(n9036) );
  NAND2_X1 U10336 ( .A1(n8833), .A2(n8846), .ZN(n8847) );
  NAND2_X1 U10337 ( .A1(n8847), .A2(n10096), .ZN(n8848) );
  OR2_X1 U10338 ( .A1(n8849), .A2(n8848), .ZN(n8852) );
  AOI22_X1 U10339 ( .A1(n8850), .A2(n10091), .B1(n10093), .B2(n8871), .ZN(
        n8851) );
  NAND2_X1 U10340 ( .A1(n8852), .A2(n8851), .ZN(n9034) );
  MUX2_X1 U10341 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9034), .S(n7308), .Z(n8853) );
  INV_X1 U10342 ( .A(n8853), .ZN(n8856) );
  AOI22_X1 U10343 ( .A1(n6447), .A2(n10101), .B1(n10102), .B2(n8854), .ZN(
        n8855) );
  OAI211_X1 U10344 ( .C1(n9036), .C2(n8917), .A(n8856), .B(n8855), .ZN(
        P2_U3214) );
  NAND2_X1 U10345 ( .A1(n8858), .A2(n8857), .ZN(n8862) );
  NAND2_X1 U10346 ( .A1(n8950), .A2(n8859), .ZN(n8860) );
  XOR2_X1 U10347 ( .A(n8862), .B(n8860), .Z(n9044) );
  XOR2_X1 U10348 ( .A(n8862), .B(n8861), .Z(n8864) );
  AOI222_X1 U10349 ( .A1(n10096), .A2(n8864), .B1(n8863), .B2(n10091), .C1(
        n8885), .C2(n10093), .ZN(n9039) );
  MUX2_X1 U10350 ( .A(n8865), .B(n9039), .S(n7308), .Z(n8868) );
  AOI22_X1 U10351 ( .A1(n9041), .A2(n10101), .B1(n10102), .B2(n8866), .ZN(
        n8867) );
  OAI211_X1 U10352 ( .C1(n9044), .C2(n8917), .A(n8868), .B(n8867), .ZN(
        P2_U3215) );
  XNOR2_X1 U10353 ( .A(n8869), .B(n4908), .ZN(n8872) );
  AOI222_X1 U10354 ( .A1(n10096), .A2(n8872), .B1(n8871), .B2(n10091), .C1(
        n8870), .C2(n10093), .ZN(n8952) );
  INV_X1 U10355 ( .A(n8873), .ZN(n8875) );
  OAI22_X1 U10356 ( .A1(n7308), .A2(n8876), .B1(n8875), .B2(n8874), .ZN(n8877)
         );
  AOI21_X1 U10357 ( .B1(n8948), .B2(n10101), .A(n8877), .ZN(n8881) );
  NAND2_X1 U10358 ( .A1(n8879), .A2(n8878), .ZN(n8949) );
  NAND3_X1 U10359 ( .A1(n8950), .A2(n10104), .A3(n8949), .ZN(n8880) );
  OAI211_X1 U10360 ( .C1(n8952), .C2(n10107), .A(n8881), .B(n8880), .ZN(
        P2_U3216) );
  XOR2_X1 U10361 ( .A(n8883), .B(n8882), .Z(n9051) );
  XOR2_X1 U10362 ( .A(n8884), .B(n8883), .Z(n8886) );
  AOI222_X1 U10363 ( .A1(n10096), .A2(n8886), .B1(n8909), .B2(n10093), .C1(
        n8885), .C2(n10091), .ZN(n9046) );
  MUX2_X1 U10364 ( .A(n10277), .B(n9046), .S(n7308), .Z(n8889) );
  AOI22_X1 U10365 ( .A1(n9048), .A2(n10101), .B1(n10102), .B2(n8887), .ZN(
        n8888) );
  OAI211_X1 U10366 ( .C1(n9051), .C2(n8917), .A(n8889), .B(n8888), .ZN(
        P2_U3217) );
  XNOR2_X1 U10367 ( .A(n8890), .B(n4657), .ZN(n8958) );
  INV_X1 U10368 ( .A(n8958), .ZN(n8904) );
  XNOR2_X1 U10369 ( .A(n8891), .B(n8892), .ZN(n8893) );
  OAI222_X1 U10370 ( .A1(n8898), .A2(n8897), .B1(n8896), .B2(n8895), .C1(n8894), .C2(n8893), .ZN(n8957) );
  AOI22_X1 U10371 ( .A1(n10107), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n10102), 
        .B2(n8899), .ZN(n8900) );
  OAI21_X1 U10372 ( .B1(n9056), .B2(n8901), .A(n8900), .ZN(n8902) );
  AOI21_X1 U10373 ( .B1(n8957), .B2(n7308), .A(n8902), .ZN(n8903) );
  OAI21_X1 U10374 ( .B1(n8904), .B2(n8917), .A(n8903), .ZN(P2_U3218) );
  XNOR2_X1 U10375 ( .A(n8905), .B(n8906), .ZN(n9062) );
  XNOR2_X1 U10376 ( .A(n8907), .B(n8908), .ZN(n8911) );
  AOI222_X1 U10377 ( .A1(n10096), .A2(n8911), .B1(n8910), .B2(n10093), .C1(
        n8909), .C2(n10091), .ZN(n9057) );
  AOI22_X1 U10378 ( .A1(n9059), .A2(n8913), .B1(n10102), .B2(n8912), .ZN(n8914) );
  AOI21_X1 U10379 ( .B1(n9057), .B2(n8914), .A(n10107), .ZN(n8915) );
  AOI21_X1 U10380 ( .B1(n10107), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8915), .ZN(
        n8916) );
  OAI21_X1 U10381 ( .B1(n9062), .B2(n8917), .A(n8916), .ZN(P2_U3219) );
  NOR2_X1 U10382 ( .A1(n8981), .A2(n10164), .ZN(n8919) );
  AOI21_X1 U10383 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10164), .A(n8919), .ZN(
        n8918) );
  OAI21_X1 U10384 ( .B1(n8983), .B2(n8961), .A(n8918), .ZN(P2_U3490) );
  AOI21_X1 U10385 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10164), .A(n8919), .ZN(
        n8920) );
  OAI21_X1 U10386 ( .B1(n8986), .B2(n8961), .A(n8920), .ZN(P2_U3489) );
  MUX2_X1 U10387 ( .A(n8922), .B(n8993), .S(n10166), .Z(n8924) );
  NAND2_X1 U10388 ( .A1(n8995), .A2(n8967), .ZN(n8923) );
  OAI211_X1 U10389 ( .C1(n8975), .C2(n8998), .A(n8924), .B(n8923), .ZN(
        P2_U3485) );
  MUX2_X1 U10390 ( .A(n8925), .B(n8999), .S(n10166), .Z(n8927) );
  NAND2_X1 U10391 ( .A1(n9001), .A2(n8967), .ZN(n8926) );
  OAI211_X1 U10392 ( .C1(n9004), .C2(n8975), .A(n8927), .B(n8926), .ZN(
        P2_U3484) );
  INV_X1 U10393 ( .A(n8928), .ZN(n9005) );
  MUX2_X1 U10394 ( .A(n10222), .B(n9005), .S(n10166), .Z(n8930) );
  INV_X1 U10395 ( .A(n8975), .ZN(n8968) );
  AOI22_X1 U10396 ( .A1(n9008), .A2(n8968), .B1(n8967), .B2(n9007), .ZN(n8929)
         );
  NAND2_X1 U10397 ( .A1(n8930), .A2(n8929), .ZN(P2_U3483) );
  MUX2_X1 U10398 ( .A(n8931), .B(n9011), .S(n10166), .Z(n8933) );
  NAND2_X1 U10399 ( .A1(n9013), .A2(n8967), .ZN(n8932) );
  OAI211_X1 U10400 ( .C1(n9016), .C2(n8975), .A(n8933), .B(n8932), .ZN(
        P2_U3482) );
  MUX2_X1 U10401 ( .A(n8934), .B(n9017), .S(n10166), .Z(n8936) );
  AOI22_X1 U10402 ( .A1(n9020), .A2(n8968), .B1(n8967), .B2(n9019), .ZN(n8935)
         );
  NAND2_X1 U10403 ( .A1(n8936), .A2(n8935), .ZN(P2_U3481) );
  MUX2_X1 U10404 ( .A(n8937), .B(n9023), .S(n10166), .Z(n8939) );
  AOI22_X1 U10405 ( .A1(n9026), .A2(n8968), .B1(n8967), .B2(n9025), .ZN(n8938)
         );
  NAND2_X1 U10406 ( .A1(n8939), .A2(n8938), .ZN(P2_U3480) );
  MUX2_X1 U10407 ( .A(n8940), .B(n9029), .S(n10166), .Z(n8942) );
  NAND2_X1 U10408 ( .A1(n6277), .A2(n8967), .ZN(n8941) );
  OAI211_X1 U10409 ( .C1(n9033), .C2(n8975), .A(n8942), .B(n8941), .ZN(
        P2_U3479) );
  MUX2_X1 U10410 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9034), .S(n10166), .Z(
        n8944) );
  OAI22_X1 U10411 ( .A1(n9036), .A2(n8975), .B1(n9035), .B2(n8961), .ZN(n8943)
         );
  OR2_X1 U10412 ( .A1(n8944), .A2(n8943), .ZN(P2_U3478) );
  MUX2_X1 U10413 ( .A(n8945), .B(n9039), .S(n10166), .Z(n8947) );
  NAND2_X1 U10414 ( .A1(n9041), .A2(n8967), .ZN(n8946) );
  OAI211_X1 U10415 ( .C1(n9044), .C2(n8975), .A(n8947), .B(n8946), .ZN(
        P2_U3477) );
  INV_X1 U10416 ( .A(n8948), .ZN(n8953) );
  NAND3_X1 U10417 ( .A1(n8950), .A2(n10139), .A3(n8949), .ZN(n8951) );
  OAI211_X1 U10418 ( .C1(n8953), .C2(n10135), .A(n8952), .B(n8951), .ZN(n9045)
         );
  MUX2_X1 U10419 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9045), .S(n10166), .Z(
        P2_U3476) );
  MUX2_X1 U10420 ( .A(n8954), .B(n9046), .S(n10166), .Z(n8956) );
  NAND2_X1 U10421 ( .A1(n9048), .A2(n8967), .ZN(n8955) );
  OAI211_X1 U10422 ( .C1(n9051), .C2(n8975), .A(n8956), .B(n8955), .ZN(
        P2_U3475) );
  AOI21_X1 U10423 ( .B1(n10139), .B2(n8958), .A(n8957), .ZN(n9052) );
  MUX2_X1 U10424 ( .A(n8959), .B(n9052), .S(n10166), .Z(n8960) );
  OAI21_X1 U10425 ( .B1(n9056), .B2(n8961), .A(n8960), .ZN(P2_U3474) );
  MUX2_X1 U10426 ( .A(n8962), .B(n9057), .S(n10166), .Z(n8964) );
  NAND2_X1 U10427 ( .A1(n9059), .A2(n8967), .ZN(n8963) );
  OAI211_X1 U10428 ( .C1(n9062), .C2(n8975), .A(n8964), .B(n8963), .ZN(
        P2_U3473) );
  INV_X1 U10429 ( .A(n8965), .ZN(n9063) );
  MUX2_X1 U10430 ( .A(n8966), .B(n9063), .S(n10166), .Z(n8970) );
  AOI22_X1 U10431 ( .A1(n9068), .A2(n8968), .B1(n8967), .B2(n9065), .ZN(n8969)
         );
  NAND2_X1 U10432 ( .A1(n8970), .A2(n8969), .ZN(P2_U3472) );
  AOI21_X1 U10433 ( .B1(n10151), .B2(n8972), .A(n8971), .ZN(n9071) );
  MUX2_X1 U10434 ( .A(n8973), .B(n9071), .S(n10166), .Z(n8974) );
  OAI21_X1 U10435 ( .B1(n8975), .B2(n9075), .A(n8974), .ZN(P2_U3471) );
  NAND2_X1 U10436 ( .A1(n8976), .A2(n10151), .ZN(n8977) );
  OAI211_X1 U10437 ( .C1(n8979), .C2(n6321), .A(n8978), .B(n8977), .ZN(n9076)
         );
  MUX2_X1 U10438 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9076), .S(n10166), .Z(
        P2_U3468) );
  MUX2_X1 U10439 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8980), .S(n10166), .Z(
        P2_U3459) );
  NOR2_X1 U10440 ( .A1(n8981), .A2(n10154), .ZN(n8984) );
  AOI21_X1 U10441 ( .B1(n10154), .B2(P2_REG0_REG_31__SCAN_IN), .A(n8984), .ZN(
        n8982) );
  OAI21_X1 U10442 ( .B1(n8983), .B2(n9055), .A(n8982), .ZN(P2_U3458) );
  AOI21_X1 U10443 ( .B1(n10154), .B2(P2_REG0_REG_30__SCAN_IN), .A(n8984), .ZN(
        n8985) );
  OAI21_X1 U10444 ( .B1(n8986), .B2(n9055), .A(n8985), .ZN(P2_U3457) );
  INV_X1 U10445 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8988) );
  MUX2_X1 U10446 ( .A(n8988), .B(n8987), .S(n10152), .Z(n8991) );
  NAND2_X1 U10447 ( .A1(n8989), .A2(n9066), .ZN(n8990) );
  OAI211_X1 U10448 ( .C1(n8992), .C2(n9074), .A(n8991), .B(n8990), .ZN(
        P2_U3454) );
  INV_X1 U10449 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8994) );
  MUX2_X1 U10450 ( .A(n8994), .B(n8993), .S(n10152), .Z(n8997) );
  NAND2_X1 U10451 ( .A1(n8995), .A2(n9066), .ZN(n8996) );
  OAI211_X1 U10452 ( .C1(n8998), .C2(n9074), .A(n8997), .B(n8996), .ZN(
        P2_U3453) );
  INV_X1 U10453 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9000) );
  MUX2_X1 U10454 ( .A(n9000), .B(n8999), .S(n10152), .Z(n9003) );
  NAND2_X1 U10455 ( .A1(n9001), .A2(n9066), .ZN(n9002) );
  OAI211_X1 U10456 ( .C1(n9004), .C2(n9074), .A(n9003), .B(n9002), .ZN(
        P2_U3452) );
  INV_X1 U10457 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9006) );
  MUX2_X1 U10458 ( .A(n9006), .B(n9005), .S(n10152), .Z(n9010) );
  INV_X1 U10459 ( .A(n9074), .ZN(n9067) );
  AOI22_X1 U10460 ( .A1(n9008), .A2(n9067), .B1(n9066), .B2(n9007), .ZN(n9009)
         );
  NAND2_X1 U10461 ( .A1(n9010), .A2(n9009), .ZN(P2_U3451) );
  INV_X1 U10462 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9012) );
  MUX2_X1 U10463 ( .A(n9012), .B(n9011), .S(n10152), .Z(n9015) );
  NAND2_X1 U10464 ( .A1(n9013), .A2(n9066), .ZN(n9014) );
  OAI211_X1 U10465 ( .C1(n9016), .C2(n9074), .A(n9015), .B(n9014), .ZN(
        P2_U3450) );
  INV_X1 U10466 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9018) );
  MUX2_X1 U10467 ( .A(n9018), .B(n9017), .S(n10152), .Z(n9022) );
  AOI22_X1 U10468 ( .A1(n9020), .A2(n9067), .B1(n9066), .B2(n9019), .ZN(n9021)
         );
  NAND2_X1 U10469 ( .A1(n9022), .A2(n9021), .ZN(P2_U3449) );
  INV_X1 U10470 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9024) );
  MUX2_X1 U10471 ( .A(n9024), .B(n9023), .S(n10152), .Z(n9028) );
  AOI22_X1 U10472 ( .A1(n9026), .A2(n9067), .B1(n9066), .B2(n9025), .ZN(n9027)
         );
  NAND2_X1 U10473 ( .A1(n9028), .A2(n9027), .ZN(P2_U3448) );
  INV_X1 U10474 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9030) );
  MUX2_X1 U10475 ( .A(n9030), .B(n9029), .S(n10152), .Z(n9032) );
  NAND2_X1 U10476 ( .A1(n6277), .A2(n9066), .ZN(n9031) );
  OAI211_X1 U10477 ( .C1(n9033), .C2(n9074), .A(n9032), .B(n9031), .ZN(
        P2_U3447) );
  MUX2_X1 U10478 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9034), .S(n10152), .Z(
        n9038) );
  OAI22_X1 U10479 ( .A1(n9036), .A2(n9074), .B1(n9035), .B2(n9055), .ZN(n9037)
         );
  OR2_X1 U10480 ( .A1(n9038), .A2(n9037), .ZN(P2_U3446) );
  INV_X1 U10481 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9040) );
  MUX2_X1 U10482 ( .A(n9040), .B(n9039), .S(n10152), .Z(n9043) );
  NAND2_X1 U10483 ( .A1(n9041), .A2(n9066), .ZN(n9042) );
  OAI211_X1 U10484 ( .C1(n9044), .C2(n9074), .A(n9043), .B(n9042), .ZN(
        P2_U3444) );
  MUX2_X1 U10485 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9045), .S(n10152), .Z(
        P2_U3441) );
  INV_X1 U10486 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9047) );
  MUX2_X1 U10487 ( .A(n9047), .B(n9046), .S(n10152), .Z(n9050) );
  NAND2_X1 U10488 ( .A1(n9048), .A2(n9066), .ZN(n9049) );
  OAI211_X1 U10489 ( .C1(n9051), .C2(n9074), .A(n9050), .B(n9049), .ZN(
        P2_U3438) );
  MUX2_X1 U10490 ( .A(n9053), .B(n9052), .S(n10152), .Z(n9054) );
  OAI21_X1 U10491 ( .B1(n9056), .B2(n9055), .A(n9054), .ZN(P2_U3435) );
  MUX2_X1 U10492 ( .A(n9058), .B(n9057), .S(n10152), .Z(n9061) );
  NAND2_X1 U10493 ( .A1(n9059), .A2(n9066), .ZN(n9060) );
  OAI211_X1 U10494 ( .C1(n9062), .C2(n9074), .A(n9061), .B(n9060), .ZN(
        P2_U3432) );
  INV_X1 U10495 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9064) );
  MUX2_X1 U10496 ( .A(n9064), .B(n9063), .S(n10152), .Z(n9070) );
  AOI22_X1 U10497 ( .A1(n9068), .A2(n9067), .B1(n9066), .B2(n9065), .ZN(n9069)
         );
  NAND2_X1 U10498 ( .A1(n9070), .A2(n9069), .ZN(P2_U3429) );
  INV_X1 U10499 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9072) );
  MUX2_X1 U10500 ( .A(n9072), .B(n9071), .S(n10152), .Z(n9073) );
  OAI21_X1 U10501 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(P2_U3426) );
  MUX2_X1 U10502 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n9076), .S(n10152), .Z(
        P2_U3417) );
  NAND3_X1 U10503 ( .A1(n9077), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n9079) );
  OAI22_X1 U10504 ( .A1(n9080), .A2(n9079), .B1(n9078), .B2(n9097), .ZN(n9081)
         );
  AOI21_X1 U10505 ( .B1(n9981), .B2(n9082), .A(n9081), .ZN(n9083) );
  INV_X1 U10506 ( .A(n9083), .ZN(P2_U3264) );
  OAI222_X1 U10507 ( .A1(n9097), .A2(n9085), .B1(n9093), .B2(n8386), .C1(n9084), .C2(P2_U3151), .ZN(P2_U3266) );
  AOI21_X1 U10508 ( .B1(n9091), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n9086), .ZN(
        n9087) );
  OAI21_X1 U10509 ( .B1(n9088), .B2(n9093), .A(n9087), .ZN(P2_U3267) );
  INV_X1 U10510 ( .A(n9089), .ZN(n9993) );
  AOI21_X1 U10511 ( .B1(n9091), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n9090), .ZN(
        n9092) );
  OAI21_X1 U10512 ( .B1(n9993), .B2(n9093), .A(n9092), .ZN(P2_U3268) );
  INV_X1 U10513 ( .A(n9094), .ZN(n9998) );
  OAI222_X1 U10514 ( .A1(n9096), .A2(P2_U3151), .B1(n9093), .B2(n9998), .C1(
        n9095), .C2(n9097), .ZN(P2_U3269) );
  OAI222_X1 U10515 ( .A1(n6323), .A2(P2_U3151), .B1(n9093), .B2(n9099), .C1(
        n9098), .C2(n9097), .ZN(P2_U3270) );
  MUX2_X1 U10516 ( .A(n9100), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10517 ( .A1(n9102), .A2(n9101), .ZN(n9103) );
  XOR2_X1 U10518 ( .A(n9104), .B(n9103), .Z(n9111) );
  OAI22_X1 U10519 ( .A1(n9326), .A2(n9106), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9105), .ZN(n9109) );
  NOR2_X1 U10520 ( .A1(n9341), .A2(n9107), .ZN(n9108) );
  AOI211_X1 U10521 ( .C1(n9967), .C2(n9343), .A(n9109), .B(n9108), .ZN(n9110)
         );
  OAI21_X1 U10522 ( .B1(n9111), .B2(n9345), .A(n9110), .ZN(P1_U3215) );
  INV_X1 U10523 ( .A(n9112), .ZN(n9117) );
  AOI21_X1 U10524 ( .B1(n9114), .B2(n9116), .A(n9113), .ZN(n9115) );
  AOI21_X1 U10525 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9123) );
  OAI22_X1 U10526 ( .A1(n9119), .A2(n9336), .B1(n9118), .B2(n9337), .ZN(n9639)
         );
  AOI22_X1 U10527 ( .A1(n9639), .A2(n9339), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9120) );
  OAI21_X1 U10528 ( .B1(n9341), .B2(n9646), .A(n9120), .ZN(n9121) );
  AOI21_X1 U10529 ( .B1(n9922), .B2(n9343), .A(n9121), .ZN(n9122) );
  OAI21_X1 U10530 ( .B1(n9123), .B2(n9345), .A(n9122), .ZN(P1_U3216) );
  INV_X1 U10531 ( .A(n9124), .ZN(n9125) );
  NAND2_X1 U10532 ( .A1(n9126), .A2(n9125), .ZN(n9298) );
  OAI21_X1 U10533 ( .B1(n9126), .B2(n9125), .A(n9298), .ZN(n9127) );
  NOR2_X1 U10534 ( .A1(n9127), .A2(n9128), .ZN(n9301) );
  AOI21_X1 U10535 ( .B1(n9128), .B2(n9127), .A(n9301), .ZN(n9135) );
  NAND2_X1 U10536 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9491) );
  OAI21_X1 U10537 ( .B1(n9326), .B2(n9129), .A(n9491), .ZN(n9132) );
  NOR2_X1 U10538 ( .A1(n9341), .A2(n9130), .ZN(n9131) );
  AOI211_X1 U10539 ( .C1(n9133), .C2(n9343), .A(n9132), .B(n9131), .ZN(n9134)
         );
  OAI21_X1 U10540 ( .B1(n9135), .B2(n9345), .A(n9134), .ZN(P1_U3217) );
  OAI21_X1 U10541 ( .B1(n9138), .B2(n9137), .A(n9136), .ZN(n9139) );
  NAND2_X1 U10542 ( .A1(n9139), .A2(n9302), .ZN(n9143) );
  AOI22_X1 U10543 ( .A1(n9343), .A2(n10330), .B1(n9339), .B2(n9140), .ZN(n9142) );
  MUX2_X1 U10544 ( .A(n9341), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n9141) );
  NAND3_X1 U10545 ( .A1(n9143), .A2(n9142), .A3(n9141), .ZN(P1_U3218) );
  NOR2_X1 U10546 ( .A1(n9148), .A2(n9334), .ZN(n9151) );
  NAND2_X1 U10547 ( .A1(n9144), .A2(n9145), .ZN(n9214) );
  INV_X1 U10548 ( .A(n9144), .ZN(n9147) );
  NOR2_X1 U10549 ( .A1(n9215), .A2(n9148), .ZN(n9149) );
  XNOR2_X1 U10550 ( .A(n9179), .B(n9153), .ZN(n9311) );
  AOI22_X1 U10551 ( .A1(n9311), .A2(n9178), .B1(n9177), .B2(n9179), .ZN(n9158)
         );
  NOR2_X1 U10552 ( .A1(n9155), .A2(n9154), .ZN(n9176) );
  INV_X1 U10553 ( .A(n9265), .ZN(n9156) );
  NOR2_X1 U10554 ( .A1(n9176), .A2(n9156), .ZN(n9157) );
  XNOR2_X1 U10555 ( .A(n9158), .B(n9157), .ZN(n9163) );
  NOR2_X1 U10556 ( .A1(n9341), .A2(n9710), .ZN(n9161) );
  AOI22_X1 U10557 ( .A1(n9357), .A2(n9324), .B1(n9322), .B2(n9359), .ZN(n9707)
         );
  OAI22_X1 U10558 ( .A1(n9326), .A2(n9707), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9159), .ZN(n9160) );
  AOI211_X1 U10559 ( .C1(n9847), .C2(n9343), .A(n9161), .B(n9160), .ZN(n9162)
         );
  OAI21_X1 U10560 ( .B1(n9163), .B2(n9345), .A(n9162), .ZN(P1_U3219) );
  XNOR2_X1 U10561 ( .A(n9164), .B(n9165), .ZN(n9166) );
  NAND2_X1 U10562 ( .A1(n9166), .A2(n9167), .ZN(n9250) );
  OAI21_X1 U10563 ( .B1(n9167), .B2(n9166), .A(n9250), .ZN(n9168) );
  NAND2_X1 U10564 ( .A1(n9168), .A2(n9302), .ZN(n9174) );
  OAI22_X1 U10565 ( .A1(n9326), .A2(n9170), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9169), .ZN(n9171) );
  AOI21_X1 U10566 ( .B1(n9343), .B2(n9172), .A(n9171), .ZN(n9173) );
  OAI211_X1 U10567 ( .C1(n9341), .C2(n9175), .A(n9174), .B(n9173), .ZN(
        P1_U3221) );
  INV_X1 U10568 ( .A(n9179), .ZN(n9182) );
  INV_X1 U10569 ( .A(n9176), .ZN(n9181) );
  OAI211_X1 U10570 ( .C1(n9182), .C2(n9310), .A(n9181), .B(n9180), .ZN(n9266)
         );
  NOR2_X1 U10571 ( .A1(n9184), .A2(n9183), .ZN(n9264) );
  NAND3_X1 U10572 ( .A1(n9266), .A2(n9264), .A3(n9265), .ZN(n9263) );
  NOR2_X1 U10573 ( .A1(n9185), .A2(n9184), .ZN(n9188) );
  INV_X1 U10574 ( .A(n9186), .ZN(n9187) );
  AOI21_X1 U10575 ( .B1(n9263), .B2(n9188), .A(n9187), .ZN(n9193) );
  AND2_X1 U10576 ( .A1(n9357), .A2(n9322), .ZN(n9189) );
  AOI21_X1 U10577 ( .B1(n9355), .B2(n9324), .A(n9189), .ZN(n9675) );
  OAI22_X1 U10578 ( .A1(n9675), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10221), .ZN(n9191) );
  NOR2_X1 U10579 ( .A1(n9933), .A2(n9331), .ZN(n9190) );
  AOI211_X1 U10580 ( .C1(n9681), .C2(n9328), .A(n9191), .B(n9190), .ZN(n9192)
         );
  OAI21_X1 U10581 ( .B1(n9193), .B2(n9345), .A(n9192), .ZN(P1_U3223) );
  NOR3_X1 U10582 ( .A1(n4373), .A2(n4809), .A3(n9195), .ZN(n9197) );
  INV_X1 U10583 ( .A(n9196), .ZN(n9277) );
  OAI21_X1 U10584 ( .B1(n9197), .B2(n9277), .A(n9302), .ZN(n9203) );
  NOR2_X1 U10585 ( .A1(n9341), .A2(n9198), .ZN(n9199) );
  AOI211_X1 U10586 ( .C1(n9339), .C2(n9201), .A(n9200), .B(n9199), .ZN(n9202)
         );
  OAI211_X1 U10587 ( .C1(n9204), .C2(n9331), .A(n9203), .B(n9202), .ZN(
        P1_U3224) );
  XOR2_X1 U10588 ( .A(n9206), .B(n9205), .Z(n9213) );
  NAND2_X1 U10589 ( .A1(n9351), .A2(n9324), .ZN(n9208) );
  NAND2_X1 U10590 ( .A1(n9353), .A2(n9322), .ZN(n9207) );
  NAND2_X1 U10591 ( .A1(n9208), .A2(n9207), .ZN(n9610) );
  AOI22_X1 U10592 ( .A1(n9610), .A2(n9339), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3086), .ZN(n9209) );
  OAI21_X1 U10593 ( .B1(n9341), .B2(n9614), .A(n9209), .ZN(n9210) );
  AOI21_X1 U10594 ( .B1(n9211), .B2(n9343), .A(n9210), .ZN(n9212) );
  OAI21_X1 U10595 ( .B1(n9213), .B2(n9345), .A(n9212), .ZN(P1_U3225) );
  NAND2_X1 U10596 ( .A1(n9215), .A2(n9214), .ZN(n9333) );
  NOR2_X1 U10597 ( .A1(n9333), .A2(n9334), .ZN(n9332) );
  INV_X1 U10598 ( .A(n9215), .ZN(n9216) );
  NOR2_X1 U10599 ( .A1(n9332), .A2(n9216), .ZN(n9220) );
  XNOR2_X1 U10600 ( .A(n9218), .B(n9217), .ZN(n9219) );
  NOR2_X1 U10601 ( .A1(n9220), .A2(n9219), .ZN(n9229) );
  AOI21_X1 U10602 ( .B1(n9220), .B2(n9219), .A(n9229), .ZN(n9226) );
  OAI22_X1 U10603 ( .A1(n9221), .A2(n9337), .B1(n9336), .B2(n9312), .ZN(n9755)
         );
  NOR2_X1 U10604 ( .A1(n9222), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9521) );
  AOI21_X1 U10605 ( .B1(n9339), .B2(n9755), .A(n9521), .ZN(n9223) );
  OAI21_X1 U10606 ( .B1(n9341), .B2(n9759), .A(n9223), .ZN(n9224) );
  AOI21_X1 U10607 ( .B1(n9861), .B2(n9343), .A(n9224), .ZN(n9225) );
  OAI21_X1 U10608 ( .B1(n9226), .B2(n9345), .A(n9225), .ZN(P1_U3226) );
  OAI21_X1 U10609 ( .B1(n9229), .B2(n9228), .A(n9227), .ZN(n9230) );
  NAND3_X1 U10610 ( .A1(n9230), .A2(n9302), .A3(n4391), .ZN(n9234) );
  INV_X1 U10611 ( .A(n9744), .ZN(n9232) );
  AOI22_X1 U10612 ( .A1(n9361), .A2(n9322), .B1(n9324), .B2(n9359), .ZN(n9739)
         );
  NAND2_X1 U10613 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9541) );
  OAI21_X1 U10614 ( .B1(n9326), .B2(n9739), .A(n9541), .ZN(n9231) );
  AOI21_X1 U10615 ( .B1(n9328), .B2(n9232), .A(n9231), .ZN(n9233) );
  OAI211_X1 U10616 ( .C1(n9743), .C2(n9331), .A(n9234), .B(n9233), .ZN(
        P1_U3228) );
  INV_X1 U10617 ( .A(n9920), .ZN(n9246) );
  OAI21_X1 U10618 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9238) );
  NAND2_X1 U10619 ( .A1(n9238), .A2(n9302), .ZN(n9245) );
  NAND2_X1 U10620 ( .A1(n9352), .A2(n9324), .ZN(n9240) );
  NAND2_X1 U10621 ( .A1(n9354), .A2(n9322), .ZN(n9239) );
  NAND2_X1 U10622 ( .A1(n9240), .A2(n9239), .ZN(n9622) );
  INV_X1 U10623 ( .A(n9622), .ZN(n9242) );
  OAI22_X1 U10624 ( .A1(n9242), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9241), .ZN(n9243) );
  AOI21_X1 U10625 ( .B1(n9631), .B2(n9328), .A(n9243), .ZN(n9244) );
  OAI211_X1 U10626 ( .C1(n9246), .C2(n9331), .A(n9245), .B(n9244), .ZN(
        P1_U3229) );
  OAI21_X1 U10627 ( .B1(n9249), .B2(n9248), .A(n9247), .ZN(n9253) );
  OAI21_X1 U10628 ( .B1(n9251), .B2(n9164), .A(n9250), .ZN(n9252) );
  XOR2_X1 U10629 ( .A(n9253), .B(n9252), .Z(n9254) );
  NAND2_X1 U10630 ( .A1(n9254), .A2(n9302), .ZN(n9261) );
  AOI21_X1 U10631 ( .B1(n9256), .B2(n9255), .A(n9326), .ZN(n9257) );
  AOI211_X1 U10632 ( .C1(n4435), .C2(n9343), .A(n9258), .B(n9257), .ZN(n9260)
         );
  OAI211_X1 U10633 ( .C1(n9341), .C2(n9262), .A(n9261), .B(n9260), .ZN(
        P1_U3231) );
  INV_X1 U10634 ( .A(n9263), .ZN(n9268) );
  AOI21_X1 U10635 ( .B1(n9266), .B2(n9265), .A(n9264), .ZN(n9267) );
  INV_X1 U10636 ( .A(n9269), .ZN(n9697) );
  AOI22_X1 U10637 ( .A1(n9356), .A2(n9324), .B1(n9322), .B2(n9358), .ZN(n9694)
         );
  OAI22_X1 U10638 ( .A1(n9326), .A2(n9694), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9270), .ZN(n9271) );
  AOI21_X1 U10639 ( .B1(n9328), .B2(n9697), .A(n9271), .ZN(n9272) );
  OAI211_X1 U10640 ( .C1(n9700), .C2(n9331), .A(n9273), .B(n9272), .ZN(
        P1_U3233) );
  INV_X1 U10641 ( .A(n9274), .ZN(n9276) );
  NOR3_X1 U10642 ( .A1(n9277), .A2(n9276), .A3(n9275), .ZN(n9280) );
  INV_X1 U10643 ( .A(n9278), .ZN(n9279) );
  OAI21_X1 U10644 ( .B1(n9280), .B2(n9279), .A(n9302), .ZN(n9286) );
  NOR2_X1 U10645 ( .A1(n9341), .A2(n9281), .ZN(n9282) );
  AOI211_X1 U10646 ( .C1(n9339), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9285)
         );
  OAI211_X1 U10647 ( .C1(n9287), .C2(n9331), .A(n9286), .B(n9285), .ZN(
        P1_U3234) );
  NOR2_X1 U10648 ( .A1(n9289), .A2(n9290), .ZN(n9288) );
  AOI21_X1 U10649 ( .B1(n9290), .B2(n9289), .A(n9288), .ZN(n9296) );
  OAI22_X1 U10650 ( .A1(n9292), .A2(n9336), .B1(n9291), .B2(n9337), .ZN(n9658)
         );
  AOI22_X1 U10651 ( .A1(n9658), .A2(n9339), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9293) );
  OAI21_X1 U10652 ( .B1(n9341), .B2(n9663), .A(n9293), .ZN(n9294) );
  AOI21_X1 U10653 ( .B1(n9662), .B2(n9343), .A(n9294), .ZN(n9295) );
  OAI21_X1 U10654 ( .B1(n9296), .B2(n9345), .A(n9295), .ZN(P1_U3235) );
  INV_X1 U10655 ( .A(n9297), .ZN(n9300) );
  INV_X1 U10656 ( .A(n9298), .ZN(n9299) );
  NOR3_X1 U10657 ( .A1(n9301), .A2(n9300), .A3(n9299), .ZN(n9303) );
  OAI21_X1 U10658 ( .B1(n9303), .B2(n4373), .A(n9302), .ZN(n9309) );
  NOR2_X1 U10659 ( .A1(n9304), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9507) );
  NOR2_X1 U10660 ( .A1(n9341), .A2(n9305), .ZN(n9306) );
  AOI211_X1 U10661 ( .C1(n9339), .C2(n9307), .A(n9507), .B(n9306), .ZN(n9308)
         );
  OAI211_X1 U10662 ( .C1(n4771), .C2(n9331), .A(n9309), .B(n9308), .ZN(
        P1_U3236) );
  XNOR2_X1 U10663 ( .A(n9311), .B(n9310), .ZN(n9317) );
  OAI22_X1 U10664 ( .A1(n9313), .A2(n9336), .B1(n9337), .B2(n9312), .ZN(n9724)
         );
  AOI22_X1 U10665 ( .A1(n9339), .A2(n9724), .B1(P1_REG3_REG_18__SCAN_IN), .B2(
        P1_U3086), .ZN(n9314) );
  OAI21_X1 U10666 ( .B1(n9341), .B2(n9729), .A(n9314), .ZN(n9315) );
  AOI21_X1 U10667 ( .B1(n9852), .B2(n9343), .A(n9315), .ZN(n9316) );
  OAI21_X1 U10668 ( .B1(n9317), .B2(n9345), .A(n9316), .ZN(P1_U3238) );
  AOI21_X1 U10669 ( .B1(n9318), .B2(n9319), .A(n9345), .ZN(n9321) );
  NAND2_X1 U10670 ( .A1(n9321), .A2(n9320), .ZN(n9330) );
  AND2_X1 U10671 ( .A1(n9352), .A2(n9322), .ZN(n9323) );
  AOI21_X1 U10672 ( .B1(n9350), .B2(n9324), .A(n9323), .ZN(n9595) );
  OAI22_X1 U10673 ( .A1(n9595), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9325), .ZN(n9327) );
  AOI21_X1 U10674 ( .B1(n9599), .B2(n9328), .A(n9327), .ZN(n9329) );
  OAI211_X1 U10675 ( .C1(n9602), .C2(n9331), .A(n9330), .B(n9329), .ZN(
        P1_U3240) );
  AOI21_X1 U10676 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9346) );
  NAND2_X1 U10677 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10031)
         );
  OAI22_X1 U10678 ( .A1(n9338), .A2(n9337), .B1(n9336), .B2(n9335), .ZN(n9777)
         );
  NAND2_X1 U10679 ( .A1(n9339), .A2(n9777), .ZN(n9340) );
  OAI211_X1 U10680 ( .C1(n9341), .C2(n9781), .A(n10031), .B(n9340), .ZN(n9342)
         );
  AOI21_X1 U10681 ( .B1(n9870), .B2(n9343), .A(n9342), .ZN(n9344) );
  OAI21_X1 U10682 ( .B1(n9346), .B2(n9345), .A(n9344), .ZN(P1_U3241) );
  MUX2_X1 U10683 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n9347), .S(n9390), .Z(
        P1_U3585) );
  MUX2_X1 U10684 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9348), .S(n9390), .Z(
        P1_U3584) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9349), .S(n9390), .Z(
        P1_U3583) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n5555), .S(n9390), .Z(
        P1_U3582) );
  MUX2_X1 U10687 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9350), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10688 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9351), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9352), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9353), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9354), .S(n9390), .Z(
        P1_U3577) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9355), .S(n9390), .Z(
        P1_U3576) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9356), .S(n9390), .Z(
        P1_U3575) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9357), .S(n9390), .Z(
        P1_U3574) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9358), .S(n9390), .Z(
        P1_U3573) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9359), .S(n9390), .Z(
        P1_U3572) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9360), .S(n9390), .Z(
        P1_U3571) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9361), .S(n9390), .Z(
        P1_U3570) );
  MUX2_X1 U10699 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9362), .S(n9390), .Z(
        P1_U3569) );
  MUX2_X1 U10700 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9363), .S(n9390), .Z(
        P1_U3568) );
  MUX2_X1 U10701 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9364), .S(n9390), .Z(
        P1_U3567) );
  MUX2_X1 U10702 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9365), .S(n9390), .Z(
        P1_U3566) );
  MUX2_X1 U10703 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9366), .S(n9390), .Z(
        P1_U3565) );
  MUX2_X1 U10704 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9367), .S(n9390), .Z(
        P1_U3564) );
  MUX2_X1 U10705 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9368), .S(n9390), .Z(
        P1_U3563) );
  MUX2_X1 U10706 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9369), .S(n9390), .Z(
        P1_U3562) );
  MUX2_X1 U10707 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9370), .S(n9390), .Z(
        P1_U3561) );
  MUX2_X1 U10708 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9371), .S(n9390), .Z(
        P1_U3560) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9372), .S(n9390), .Z(
        P1_U3559) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9373), .S(n9390), .Z(
        P1_U3558) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n5084), .S(n9390), .Z(
        P1_U3557) );
  MUX2_X1 U10712 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9374), .S(n9390), .Z(
        P1_U3556) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9375), .S(n9390), .Z(
        P1_U3555) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n6693), .S(n9390), .Z(
        P1_U3554) );
  OAI211_X1 U10715 ( .C1(n9377), .C2(n9387), .A(n9501), .B(n9376), .ZN(n9385)
         );
  OAI211_X1 U10716 ( .C1(n9380), .C2(n9379), .A(n10037), .B(n9378), .ZN(n9384)
         );
  AOI22_X1 U10717 ( .A1(n10004), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9383) );
  NAND2_X1 U10718 ( .A1(n10030), .A2(n9381), .ZN(n9382) );
  NAND4_X1 U10719 ( .A1(n9385), .A2(n9384), .A3(n9383), .A4(n9382), .ZN(
        P1_U3244) );
  NAND2_X1 U10720 ( .A1(n9386), .A2(n10002), .ZN(n9391) );
  OAI21_X1 U10721 ( .B1(n10002), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9386), .ZN(
        n10000) );
  AOI22_X1 U10722 ( .A1(n4778), .A2(n10000), .B1(n9388), .B2(n9387), .ZN(n9389) );
  OAI211_X1 U10723 ( .C1(n9392), .C2(n9391), .A(n9390), .B(n9389), .ZN(n9432)
         );
  INV_X1 U10724 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9394) );
  OAI22_X1 U10725 ( .A1(n10050), .A2(n9394), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9393), .ZN(n9395) );
  AOI21_X1 U10726 ( .B1(n9396), .B2(n10030), .A(n9395), .ZN(n9405) );
  OAI211_X1 U10727 ( .C1(n9399), .C2(n9398), .A(n10037), .B(n9397), .ZN(n9404)
         );
  OAI211_X1 U10728 ( .C1(n9402), .C2(n9401), .A(n9501), .B(n9400), .ZN(n9403)
         );
  NAND4_X1 U10729 ( .A1(n9432), .A2(n9405), .A3(n9404), .A4(n9403), .ZN(
        P1_U3245) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U10731 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9406) );
  OAI21_X1 U10732 ( .B1(n10050), .B2(n9407), .A(n9406), .ZN(n9408) );
  AOI21_X1 U10733 ( .B1(n9409), .B2(n10030), .A(n9408), .ZN(n9418) );
  OAI211_X1 U10734 ( .C1(n9412), .C2(n9411), .A(n10037), .B(n9410), .ZN(n9417)
         );
  OAI211_X1 U10735 ( .C1(n9415), .C2(n9414), .A(n9501), .B(n9413), .ZN(n9416)
         );
  NAND3_X1 U10736 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(P1_U3246) );
  INV_X1 U10737 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9420) );
  OAI21_X1 U10738 ( .B1(n10050), .B2(n9420), .A(n9419), .ZN(n9421) );
  AOI21_X1 U10739 ( .B1(n9422), .B2(n10030), .A(n9421), .ZN(n9431) );
  OAI211_X1 U10740 ( .C1(n9425), .C2(n9424), .A(n9501), .B(n9423), .ZN(n9430)
         );
  OAI211_X1 U10741 ( .C1(n9428), .C2(n9427), .A(n10037), .B(n9426), .ZN(n9429)
         );
  NAND4_X1 U10742 ( .A1(n9432), .A2(n9431), .A3(n9430), .A4(n9429), .ZN(
        P1_U3247) );
  INV_X1 U10743 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9434) );
  NAND2_X1 U10744 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9433) );
  OAI21_X1 U10745 ( .B1(n10050), .B2(n9434), .A(n9433), .ZN(n9435) );
  AOI21_X1 U10746 ( .B1(n9436), .B2(n10030), .A(n9435), .ZN(n9445) );
  OAI211_X1 U10747 ( .C1(n9439), .C2(n9438), .A(n10037), .B(n9437), .ZN(n9444)
         );
  OAI211_X1 U10748 ( .C1(n9442), .C2(n9441), .A(n9501), .B(n9440), .ZN(n9443)
         );
  NAND3_X1 U10749 ( .A1(n9445), .A2(n9444), .A3(n9443), .ZN(P1_U3248) );
  INV_X1 U10750 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9447) );
  OAI21_X1 U10751 ( .B1(n10050), .B2(n9447), .A(n9446), .ZN(n9448) );
  AOI21_X1 U10752 ( .B1(n9449), .B2(n10030), .A(n9448), .ZN(n9458) );
  OAI211_X1 U10753 ( .C1(n9452), .C2(n9451), .A(n10037), .B(n9450), .ZN(n9457)
         );
  OAI211_X1 U10754 ( .C1(n9455), .C2(n9454), .A(n9501), .B(n9453), .ZN(n9456)
         );
  NAND3_X1 U10755 ( .A1(n9458), .A2(n9457), .A3(n9456), .ZN(P1_U3249) );
  INV_X1 U10756 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U10757 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9459) );
  OAI21_X1 U10758 ( .B1(n10050), .B2(n9460), .A(n9459), .ZN(n9461) );
  AOI21_X1 U10759 ( .B1(n9462), .B2(n10030), .A(n9461), .ZN(n9471) );
  OAI211_X1 U10760 ( .C1(n9465), .C2(n9464), .A(n10037), .B(n9463), .ZN(n9470)
         );
  OAI211_X1 U10761 ( .C1(n9468), .C2(n9467), .A(n9501), .B(n9466), .ZN(n9469)
         );
  NAND3_X1 U10762 ( .A1(n9471), .A2(n9470), .A3(n9469), .ZN(P1_U3250) );
  NAND2_X1 U10763 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n9472) );
  OAI21_X1 U10764 ( .B1(n10050), .B2(n9473), .A(n9472), .ZN(n9474) );
  AOI21_X1 U10765 ( .B1(n9475), .B2(n10030), .A(n9474), .ZN(n9484) );
  OAI211_X1 U10766 ( .C1(n9478), .C2(n9477), .A(n9501), .B(n9476), .ZN(n9483)
         );
  OAI211_X1 U10767 ( .C1(n9481), .C2(n9480), .A(n10037), .B(n9479), .ZN(n9482)
         );
  NAND3_X1 U10768 ( .A1(n9484), .A2(n9483), .A3(n9482), .ZN(P1_U3251) );
  OAI211_X1 U10769 ( .C1(n9487), .C2(n9486), .A(n9485), .B(n10037), .ZN(n9497)
         );
  OAI211_X1 U10770 ( .C1(n9490), .C2(n9489), .A(n9488), .B(n9501), .ZN(n9496)
         );
  INV_X1 U10771 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9492) );
  OAI21_X1 U10772 ( .B1(n10050), .B2(n9492), .A(n9491), .ZN(n9493) );
  AOI21_X1 U10773 ( .B1(n9494), .B2(n10030), .A(n9493), .ZN(n9495) );
  NAND3_X1 U10774 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(P1_U3253) );
  OAI211_X1 U10775 ( .C1(n9500), .C2(n9499), .A(n9498), .B(n10037), .ZN(n9511)
         );
  OAI211_X1 U10776 ( .C1(n9504), .C2(n9503), .A(n9502), .B(n9501), .ZN(n9510)
         );
  INV_X1 U10777 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9505) );
  NOR2_X1 U10778 ( .A1(n10050), .A2(n9505), .ZN(n9506) );
  AOI211_X1 U10779 ( .C1(n10030), .C2(n9508), .A(n9507), .B(n9506), .ZN(n9509)
         );
  NAND3_X1 U10780 ( .A1(n9511), .A2(n9510), .A3(n9509), .ZN(P1_U3254) );
  OAI21_X1 U10781 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n10013) );
  XOR2_X1 U10782 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9527), .Z(n10012) );
  NAND2_X1 U10783 ( .A1(n10013), .A2(n10012), .ZN(n10011) );
  OAI21_X1 U10784 ( .B1(n9515), .B2(n10015), .A(n10011), .ZN(n9517) );
  AND2_X1 U10785 ( .A1(n9517), .A2(n10029), .ZN(n9518) );
  INV_X1 U10786 ( .A(n9518), .ZN(n9516) );
  OAI21_X1 U10787 ( .B1(n10029), .B2(n9517), .A(n9516), .ZN(n10023) );
  INV_X1 U10788 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10024) );
  NOR2_X1 U10789 ( .A1(n10023), .A2(n10024), .ZN(n10021) );
  AOI22_X1 U10790 ( .A1(n9540), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9865), .B2(
        n9523), .ZN(n9519) );
  OAI21_X1 U10791 ( .B1(n9520), .B2(n9519), .A(n9539), .ZN(n9536) );
  AOI21_X1 U10792 ( .B1(n10004), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n9521), .ZN(
        n9522) );
  OAI21_X1 U10793 ( .B1(n9523), .B2(n10043), .A(n9522), .ZN(n9535) );
  INV_X1 U10794 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n10255) );
  NOR2_X1 U10795 ( .A1(n9527), .A2(n10255), .ZN(n9526) );
  AOI21_X1 U10796 ( .B1(n9527), .B2(n10255), .A(n9526), .ZN(n10010) );
  NOR2_X1 U10797 ( .A1(n10009), .A2(n10010), .ZN(n10008) );
  NOR2_X1 U10798 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  NAND2_X1 U10799 ( .A1(n9540), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9531) );
  OAI21_X1 U10800 ( .B1(n9540), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9531), .ZN(
        n9532) );
  NOR2_X1 U10801 ( .A1(n9533), .A2(n9532), .ZN(n9538) );
  AOI211_X1 U10802 ( .C1(n9533), .C2(n9532), .A(n9538), .B(n10034), .ZN(n9534)
         );
  AOI211_X1 U10803 ( .C1(n10037), .C2(n9536), .A(n9535), .B(n9534), .ZN(n9537)
         );
  INV_X1 U10804 ( .A(n9537), .ZN(P1_U3259) );
  XNOR2_X1 U10805 ( .A(n9553), .B(n9745), .ZN(n9547) );
  XOR2_X1 U10806 ( .A(n9547), .B(n9548), .Z(n9546) );
  OAI21_X1 U10807 ( .B1(n9540), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9539), .ZN(
        n9556) );
  XNOR2_X1 U10808 ( .A(n9553), .B(n9857), .ZN(n9555) );
  XNOR2_X1 U10809 ( .A(n9556), .B(n9555), .ZN(n9544) );
  NAND2_X1 U10810 ( .A1(n10004), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n9542) );
  OAI211_X1 U10811 ( .C1(n10043), .C2(n9549), .A(n9542), .B(n9541), .ZN(n9543)
         );
  AOI21_X1 U10812 ( .B1(n9544), .B2(n10037), .A(n9543), .ZN(n9545) );
  OAI21_X1 U10813 ( .B1(n9546), .B2(n10034), .A(n9545), .ZN(P1_U3260) );
  NAND2_X1 U10814 ( .A1(n9549), .A2(n9745), .ZN(n9550) );
  NAND2_X1 U10815 ( .A1(n9557), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9551) );
  OAI21_X1 U10816 ( .B1(n9557), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9551), .ZN(
        n10035) );
  INV_X1 U10817 ( .A(n9563), .ZN(n9561) );
  NOR2_X1 U10818 ( .A1(n9553), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n9554) );
  AOI21_X1 U10819 ( .B1(n9556), .B2(n9555), .A(n9554), .ZN(n10040) );
  OR2_X1 U10820 ( .A1(n9557), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9558) );
  NAND2_X1 U10821 ( .A1(n9557), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9559) );
  AND2_X1 U10822 ( .A1(n9558), .A2(n9559), .ZN(n10039) );
  NAND2_X1 U10823 ( .A1(n10040), .A2(n10039), .ZN(n10038) );
  NAND2_X1 U10824 ( .A1(n10038), .A2(n9559), .ZN(n9560) );
  XNOR2_X1 U10825 ( .A(n9560), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9562) );
  NAND2_X1 U10826 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9565) );
  XNOR2_X1 U10827 ( .A(n6509), .B(n9567), .ZN(n9568) );
  NAND2_X1 U10828 ( .A1(n9809), .A2(n9788), .ZN(n9571) );
  AOI21_X1 U10829 ( .B1(n9712), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9569), .ZN(
        n9570) );
  OAI211_X1 U10830 ( .C1(n6518), .C2(n9715), .A(n9571), .B(n9570), .ZN(
        P1_U3264) );
  INV_X1 U10831 ( .A(n9572), .ZN(n9582) );
  NAND2_X1 U10832 ( .A1(n9573), .A2(n9788), .ZN(n9577) );
  INV_X1 U10833 ( .A(n9574), .ZN(n9575) );
  AOI22_X1 U10834 ( .A1(n9575), .A2(n10336), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10337), .ZN(n9576) );
  OAI211_X1 U10835 ( .C1(n9578), .C2(n9715), .A(n9577), .B(n9576), .ZN(n9579)
         );
  OAI21_X1 U10836 ( .B1(n9582), .B2(n9793), .A(n9581), .ZN(P1_U3265) );
  NAND2_X1 U10837 ( .A1(n9583), .A2(n10333), .ZN(n9589) );
  AOI22_X1 U10838 ( .A1(n9585), .A2(n10336), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10337), .ZN(n9586) );
  OAI21_X1 U10839 ( .B1(n9908), .B2(n9715), .A(n9586), .ZN(n9587) );
  AOI21_X1 U10840 ( .B1(n5918), .B2(n9788), .A(n9587), .ZN(n9588) );
  OAI211_X1 U10841 ( .C1(n9590), .C2(n10337), .A(n9589), .B(n9588), .ZN(
        P1_U3266) );
  XNOR2_X1 U10842 ( .A(n9591), .B(n5666), .ZN(n9912) );
  XNOR2_X1 U10843 ( .A(n9592), .B(n9593), .ZN(n9594) );
  NAND2_X1 U10844 ( .A1(n9594), .A2(n9778), .ZN(n9596) );
  INV_X1 U10845 ( .A(n9597), .ZN(n9613) );
  AOI211_X1 U10846 ( .C1(n9814), .C2(n9613), .A(n9784), .B(n9598), .ZN(n9813)
         );
  NAND2_X1 U10847 ( .A1(n9813), .A2(n9788), .ZN(n9601) );
  AOI22_X1 U10848 ( .A1(n9599), .A2(n10336), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10337), .ZN(n9600) );
  OAI211_X1 U10849 ( .C1(n9602), .C2(n9715), .A(n9601), .B(n9600), .ZN(n9603)
         );
  AOI21_X1 U10850 ( .B1(n9812), .B2(n10344), .A(n9603), .ZN(n9604) );
  OAI21_X1 U10851 ( .B1(n9912), .B2(n9793), .A(n9604), .ZN(P1_U3267) );
  XNOR2_X1 U10852 ( .A(n9605), .B(n9607), .ZN(n9914) );
  NOR2_X1 U10853 ( .A1(n9607), .A2(n4945), .ZN(n9608) );
  AOI21_X1 U10854 ( .B1(n9609), .B2(n9608), .A(n9757), .ZN(n9611) );
  AOI21_X1 U10855 ( .B1(n9612), .B2(n9611), .A(n9610), .ZN(n9818) );
  INV_X1 U10856 ( .A(n9818), .ZN(n9619) );
  OAI211_X1 U10857 ( .C1(n9913), .C2(n9628), .A(n9613), .B(n9764), .ZN(n9817)
         );
  NOR2_X1 U10858 ( .A1(n9817), .A2(n10341), .ZN(n9618) );
  INV_X1 U10859 ( .A(n9614), .ZN(n9615) );
  AOI22_X1 U10860 ( .A1(n9615), .A2(n10336), .B1(n10337), .B2(
        P1_REG2_REG_25__SCAN_IN), .ZN(n9616) );
  OAI21_X1 U10861 ( .B1(n9913), .B2(n9715), .A(n9616), .ZN(n9617) );
  AOI211_X1 U10862 ( .C1(n9619), .C2(n10344), .A(n9618), .B(n9617), .ZN(n9620)
         );
  OAI21_X1 U10863 ( .B1(n9914), .B2(n9793), .A(n9620), .ZN(P1_U3268) );
  XNOR2_X1 U10864 ( .A(n9621), .B(n5665), .ZN(n9623) );
  AOI21_X1 U10865 ( .B1(n9623), .B2(n9778), .A(n9622), .ZN(n9823) );
  OR2_X1 U10866 ( .A1(n9626), .A2(n9625), .ZN(n9627) );
  NAND2_X1 U10867 ( .A1(n9624), .A2(n9627), .ZN(n9821) );
  INV_X1 U10868 ( .A(n9628), .ZN(n9630) );
  AOI21_X1 U10869 ( .B1(n9644), .B2(n9920), .A(n9784), .ZN(n9629) );
  NAND2_X1 U10870 ( .A1(n9630), .A2(n9629), .ZN(n9822) );
  AOI22_X1 U10871 ( .A1(n10337), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n9631), 
        .B2(n10336), .ZN(n9633) );
  NAND2_X1 U10872 ( .A1(n9920), .A2(n10331), .ZN(n9632) );
  OAI211_X1 U10873 ( .C1(n9822), .C2(n10341), .A(n9633), .B(n9632), .ZN(n9634)
         );
  AOI21_X1 U10874 ( .B1(n9821), .B2(n10333), .A(n9634), .ZN(n9635) );
  OAI21_X1 U10875 ( .B1(n10337), .B2(n9823), .A(n9635), .ZN(P1_U3269) );
  NAND2_X1 U10876 ( .A1(n9654), .A2(n9637), .ZN(n9638) );
  XNOR2_X1 U10877 ( .A(n9642), .B(n9638), .ZN(n9640) );
  AOI21_X1 U10878 ( .B1(n9640), .B2(n9778), .A(n9639), .ZN(n9828) );
  OAI21_X1 U10879 ( .B1(n9643), .B2(n9642), .A(n9641), .ZN(n9923) );
  AOI21_X1 U10880 ( .B1(n9660), .B2(n9922), .A(n9784), .ZN(n9645) );
  NAND2_X1 U10881 ( .A1(n9645), .A2(n9644), .ZN(n9827) );
  INV_X1 U10882 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9647) );
  OAI22_X1 U10883 ( .A1(n10344), .A2(n9647), .B1(n9646), .B2(n9780), .ZN(n9648) );
  AOI21_X1 U10884 ( .B1(n9922), .B2(n10331), .A(n9648), .ZN(n9649) );
  OAI21_X1 U10885 ( .B1(n9827), .B2(n10341), .A(n9649), .ZN(n9650) );
  AOI21_X1 U10886 ( .B1(n9923), .B2(n10333), .A(n9650), .ZN(n9651) );
  OAI21_X1 U10887 ( .B1(n9712), .B2(n9828), .A(n9651), .ZN(P1_U3270) );
  XNOR2_X1 U10888 ( .A(n9653), .B(n9652), .ZN(n9834) );
  INV_X1 U10889 ( .A(n9834), .ZN(n9669) );
  INV_X1 U10890 ( .A(n9654), .ZN(n9655) );
  AOI211_X1 U10891 ( .C1(n9657), .C2(n9656), .A(n9757), .B(n9655), .ZN(n9659)
         );
  OR2_X1 U10892 ( .A1(n9659), .A2(n9658), .ZN(n9832) );
  NAND2_X1 U10893 ( .A1(n9832), .A2(n7937), .ZN(n9668) );
  INV_X1 U10894 ( .A(n9660), .ZN(n9661) );
  AOI211_X1 U10895 ( .C1(n9662), .C2(n4326), .A(n9784), .B(n9661), .ZN(n9833)
         );
  NOR2_X1 U10896 ( .A1(n9931), .A2(n9715), .ZN(n9666) );
  OAI22_X1 U10897 ( .A1(n10344), .A2(n9664), .B1(n9663), .B2(n9780), .ZN(n9665) );
  AOI211_X1 U10898 ( .C1(n9833), .C2(n9788), .A(n9666), .B(n9665), .ZN(n9667)
         );
  OAI211_X1 U10899 ( .C1(n9669), .C2(n9793), .A(n9668), .B(n9667), .ZN(
        P1_U3271) );
  XNOR2_X1 U10900 ( .A(n9670), .B(n9674), .ZN(n9934) );
  INV_X1 U10901 ( .A(n9671), .ZN(n9693) );
  NAND2_X1 U10902 ( .A1(n9693), .A2(n9692), .ZN(n9691) );
  NAND2_X1 U10903 ( .A1(n9691), .A2(n9672), .ZN(n9673) );
  XOR2_X1 U10904 ( .A(n9674), .B(n9673), .Z(n9677) );
  INV_X1 U10905 ( .A(n9675), .ZN(n9676) );
  AOI21_X1 U10906 ( .B1(n9677), .B2(n9778), .A(n9676), .ZN(n9838) );
  INV_X1 U10907 ( .A(n9838), .ZN(n9685) );
  INV_X1 U10908 ( .A(n9678), .ZN(n9679) );
  NAND2_X1 U10909 ( .A1(n9679), .A2(n7218), .ZN(n9680) );
  NAND3_X1 U10910 ( .A1(n4326), .A2(n9680), .A3(n9764), .ZN(n9837) );
  AOI22_X1 U10911 ( .A1(n10337), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9681), 
        .B2(n10336), .ZN(n9683) );
  NAND2_X1 U10912 ( .A1(n7218), .A2(n10331), .ZN(n9682) );
  OAI211_X1 U10913 ( .C1(n9837), .C2(n10341), .A(n9683), .B(n9682), .ZN(n9684)
         );
  AOI21_X1 U10914 ( .B1(n9685), .B2(n10344), .A(n9684), .ZN(n9686) );
  OAI21_X1 U10915 ( .B1(n9793), .B2(n9934), .A(n9686), .ZN(P1_U3272) );
  NAND2_X1 U10916 ( .A1(n9703), .A2(n9687), .ZN(n9689) );
  NAND2_X1 U10917 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  XOR2_X1 U10918 ( .A(n9692), .B(n9690), .Z(n9940) );
  OAI211_X1 U10919 ( .C1(n9693), .C2(n9692), .A(n9691), .B(n9778), .ZN(n9695)
         );
  NAND2_X1 U10920 ( .A1(n9695), .A2(n9694), .ZN(n9841) );
  INV_X1 U10921 ( .A(n9709), .ZN(n9696) );
  AOI211_X1 U10922 ( .C1(n9843), .C2(n9696), .A(n9784), .B(n9678), .ZN(n9842)
         );
  NAND2_X1 U10923 ( .A1(n9842), .A2(n9788), .ZN(n9699) );
  AOI22_X1 U10924 ( .A1(n10337), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9697), 
        .B2(n10336), .ZN(n9698) );
  OAI211_X1 U10925 ( .C1(n9700), .C2(n9715), .A(n9699), .B(n9698), .ZN(n9701)
         );
  AOI21_X1 U10926 ( .B1(n9841), .B2(n10344), .A(n9701), .ZN(n9702) );
  OAI21_X1 U10927 ( .B1(n9940), .B2(n9793), .A(n9702), .ZN(P1_U3273) );
  XOR2_X1 U10928 ( .A(n9705), .B(n9703), .Z(n9944) );
  XOR2_X1 U10929 ( .A(n9706), .B(n9705), .Z(n9708) );
  OAI21_X1 U10930 ( .B1(n9708), .B2(n9757), .A(n9707), .ZN(n9845) );
  AOI211_X1 U10931 ( .C1(n9847), .C2(n9727), .A(n9784), .B(n9709), .ZN(n9846)
         );
  NAND2_X1 U10932 ( .A1(n9846), .A2(n9788), .ZN(n9714) );
  INV_X1 U10933 ( .A(n9710), .ZN(n9711) );
  AOI22_X1 U10934 ( .A1(n9712), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9711), .B2(
        n10336), .ZN(n9713) );
  OAI211_X1 U10935 ( .C1(n9716), .C2(n9715), .A(n9714), .B(n9713), .ZN(n9717)
         );
  AOI21_X1 U10936 ( .B1(n9845), .B2(n10344), .A(n9717), .ZN(n9718) );
  OAI21_X1 U10937 ( .B1(n9793), .B2(n9944), .A(n9718), .ZN(P1_U3274) );
  XOR2_X1 U10938 ( .A(n9719), .B(n9723), .Z(n9948) );
  NAND2_X1 U10939 ( .A1(n9720), .A2(n9721), .ZN(n9722) );
  XOR2_X1 U10940 ( .A(n9723), .B(n9722), .Z(n9726) );
  INV_X1 U10941 ( .A(n9724), .ZN(n9725) );
  OAI21_X1 U10942 ( .B1(n9726), .B2(n9757), .A(n9725), .ZN(n9850) );
  AOI21_X1 U10943 ( .B1(n9742), .B2(n9852), .A(n9784), .ZN(n9728) );
  AND2_X1 U10944 ( .A1(n9728), .A2(n9727), .ZN(n9851) );
  NAND2_X1 U10945 ( .A1(n9851), .A2(n9788), .ZN(n9733) );
  OAI22_X1 U10946 ( .A1(n10344), .A2(n9730), .B1(n9729), .B2(n9780), .ZN(n9731) );
  AOI21_X1 U10947 ( .B1(n9852), .B2(n10331), .A(n9731), .ZN(n9732) );
  NAND2_X1 U10948 ( .A1(n9733), .A2(n9732), .ZN(n9734) );
  AOI21_X1 U10949 ( .B1(n9850), .B2(n7937), .A(n9734), .ZN(n9735) );
  OAI21_X1 U10950 ( .B1(n9948), .B2(n9793), .A(n9735), .ZN(P1_U3275) );
  XNOR2_X1 U10951 ( .A(n9736), .B(n9738), .ZN(n9953) );
  INV_X1 U10952 ( .A(n9953), .ZN(n9751) );
  OAI211_X1 U10953 ( .C1(n9738), .C2(n9737), .A(n9720), .B(n9778), .ZN(n9740)
         );
  AND2_X1 U10954 ( .A1(n9740), .A2(n9739), .ZN(n9856) );
  INV_X1 U10955 ( .A(n9856), .ZN(n9749) );
  OAI211_X1 U10956 ( .C1(n9767), .C2(n9743), .A(n9742), .B(n9764), .ZN(n9855)
         );
  OAI22_X1 U10957 ( .A1(n10344), .A2(n9745), .B1(n9744), .B2(n9780), .ZN(n9746) );
  AOI21_X1 U10958 ( .B1(n9951), .B2(n10331), .A(n9746), .ZN(n9747) );
  OAI21_X1 U10959 ( .B1(n9855), .B2(n10341), .A(n9747), .ZN(n9748) );
  AOI21_X1 U10960 ( .B1(n9749), .B2(n7937), .A(n9748), .ZN(n9750) );
  OAI21_X1 U10961 ( .B1(n9793), .B2(n9751), .A(n9750), .ZN(P1_U3276) );
  NAND2_X1 U10962 ( .A1(n9774), .A2(n9752), .ZN(n9754) );
  XNOR2_X1 U10963 ( .A(n9754), .B(n9753), .ZN(n9758) );
  INV_X1 U10964 ( .A(n9755), .ZN(n9756) );
  OAI21_X1 U10965 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9862) );
  NAND2_X1 U10966 ( .A1(n9862), .A2(n7937), .ZN(n9771) );
  OAI22_X1 U10967 ( .A1(n10344), .A2(n9760), .B1(n9759), .B2(n9780), .ZN(n9761) );
  AOI21_X1 U10968 ( .B1(n9861), .B2(n10331), .A(n9761), .ZN(n9770) );
  XNOR2_X1 U10969 ( .A(n9762), .B(n9763), .ZN(n9864) );
  NAND2_X1 U10970 ( .A1(n9864), .A2(n10333), .ZN(n9769) );
  NAND2_X1 U10971 ( .A1(n9787), .A2(n9861), .ZN(n9765) );
  NAND2_X1 U10972 ( .A1(n9765), .A2(n9764), .ZN(n9766) );
  NOR2_X1 U10973 ( .A1(n9767), .A2(n9766), .ZN(n9863) );
  NAND2_X1 U10974 ( .A1(n9863), .A2(n9788), .ZN(n9768) );
  NAND4_X1 U10975 ( .A1(n9771), .A2(n9770), .A3(n9769), .A4(n9768), .ZN(
        P1_U3277) );
  XNOR2_X1 U10976 ( .A(n9772), .B(n9776), .ZN(n9964) );
  OAI21_X1 U10977 ( .B1(n9776), .B2(n9775), .A(n9774), .ZN(n9779) );
  AOI21_X1 U10978 ( .B1(n9779), .B2(n9778), .A(n9777), .ZN(n9867) );
  OAI22_X1 U10979 ( .A1(n10344), .A2(n9782), .B1(n9781), .B2(n9780), .ZN(n9783) );
  AOI21_X1 U10980 ( .B1(n9870), .B2(n10331), .A(n9783), .ZN(n9790) );
  AOI21_X1 U10981 ( .B1(n9785), .B2(n9870), .A(n9784), .ZN(n9786) );
  AND2_X1 U10982 ( .A1(n9787), .A2(n9786), .ZN(n9869) );
  NAND2_X1 U10983 ( .A1(n9869), .A2(n9788), .ZN(n9789) );
  OAI211_X1 U10984 ( .C1(n9867), .C2(n10337), .A(n9790), .B(n9789), .ZN(n9791)
         );
  INV_X1 U10985 ( .A(n9791), .ZN(n9792) );
  OAI21_X1 U10986 ( .B1(n9964), .B2(n9793), .A(n9792), .ZN(P1_U3278) );
  OAI21_X1 U10987 ( .B1(n7063), .B2(n9795), .A(n9794), .ZN(n9800) );
  NOR3_X1 U10988 ( .A1(n9798), .A2(n9797), .A3(n9796), .ZN(n9799) );
  AOI211_X1 U10989 ( .C1(n10336), .C2(P1_REG3_REG_0__SCAN_IN), .A(n9800), .B(
        n9799), .ZN(n9805) );
  NAND3_X1 U10990 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n9804) );
  NAND2_X1 U10991 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  MUX2_X1 U10992 ( .A(P1_REG2_REG_0__SCAN_IN), .B(n9806), .S(n10344), .Z(
        P1_U3293) );
  INV_X1 U10993 ( .A(n9807), .ZN(n9808) );
  NOR2_X1 U10994 ( .A1(n9809), .A2(n9808), .ZN(n9903) );
  MUX2_X1 U10995 ( .A(n9810), .B(n9903), .S(n10073), .Z(n9811) );
  OAI21_X1 U10996 ( .B1(n6518), .B2(n9902), .A(n9811), .ZN(P1_U3552) );
  INV_X1 U10997 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9815) );
  MUX2_X1 U10998 ( .A(n9815), .B(n9909), .S(n10073), .Z(n9816) );
  OAI22_X1 U10999 ( .A1(n9914), .A2(n9872), .B1(n9913), .B2(n9902), .ZN(n9820)
         );
  NAND2_X1 U11000 ( .A1(n9818), .A2(n9817), .ZN(n9915) );
  MUX2_X1 U11001 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9915), .S(n10073), .Z(
        n9819) );
  OR2_X1 U11002 ( .A1(n9820), .A2(n9819), .ZN(P1_U3547) );
  NAND2_X1 U11003 ( .A1(n9821), .A2(n10061), .ZN(n9824) );
  NAND3_X1 U11004 ( .A1(n9824), .A2(n9823), .A3(n9822), .ZN(n9918) );
  MUX2_X1 U11005 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9918), .S(n10073), .Z(
        n9825) );
  AOI21_X1 U11006 ( .B1(n6366), .B2(n9920), .A(n9825), .ZN(n9826) );
  INV_X1 U11007 ( .A(n9826), .ZN(P1_U3546) );
  AOI22_X1 U11008 ( .A1(n9923), .A2(n9858), .B1(n6366), .B2(n9922), .ZN(n9831)
         );
  INV_X1 U11009 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9829) );
  AND2_X1 U11010 ( .A1(n9828), .A2(n9827), .ZN(n9924) );
  MUX2_X1 U11011 ( .A(n9829), .B(n9924), .S(n10073), .Z(n9830) );
  NAND2_X1 U11012 ( .A1(n9831), .A2(n9830), .ZN(P1_U3545) );
  INV_X1 U11013 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9835) );
  AOI211_X1 U11014 ( .C1(n9834), .C2(n10061), .A(n9833), .B(n9832), .ZN(n9928)
         );
  MUX2_X1 U11015 ( .A(n9835), .B(n9928), .S(n10073), .Z(n9836) );
  OAI21_X1 U11016 ( .B1(n9931), .B2(n9902), .A(n9836), .ZN(P1_U3544) );
  NAND2_X1 U11017 ( .A1(n9838), .A2(n9837), .ZN(n9932) );
  MUX2_X1 U11018 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9932), .S(n10073), .Z(
        n9840) );
  OAI22_X1 U11019 ( .A1(n9934), .A2(n9872), .B1(n9933), .B2(n9902), .ZN(n9839)
         );
  OR2_X1 U11020 ( .A1(n9840), .A2(n9839), .ZN(P1_U3543) );
  INV_X1 U11021 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10258) );
  AOI211_X1 U11022 ( .C1(n10064), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9937)
         );
  MUX2_X1 U11023 ( .A(n10258), .B(n9937), .S(n10073), .Z(n9844) );
  OAI21_X1 U11024 ( .B1(n9940), .B2(n9872), .A(n9844), .ZN(P1_U3542) );
  INV_X1 U11025 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9848) );
  AOI211_X1 U11026 ( .C1(n10064), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9941)
         );
  MUX2_X1 U11027 ( .A(n9848), .B(n9941), .S(n10073), .Z(n9849) );
  OAI21_X1 U11028 ( .B1(n9872), .B2(n9944), .A(n9849), .ZN(P1_U3541) );
  INV_X1 U11029 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9853) );
  AOI211_X1 U11030 ( .C1(n10064), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9945)
         );
  MUX2_X1 U11031 ( .A(n9853), .B(n9945), .S(n10073), .Z(n9854) );
  OAI21_X1 U11032 ( .B1(n9948), .B2(n9872), .A(n9854), .ZN(P1_U3540) );
  AND2_X1 U11033 ( .A1(n9856), .A2(n9855), .ZN(n9950) );
  MUX2_X1 U11034 ( .A(n9950), .B(n9857), .S(n7060), .Z(n9860) );
  AOI22_X1 U11035 ( .A1(n9953), .A2(n9858), .B1(n6366), .B2(n9951), .ZN(n9859)
         );
  NAND2_X1 U11036 ( .A1(n9860), .A2(n9859), .ZN(P1_U3539) );
  INV_X1 U11037 ( .A(n9861), .ZN(n9959) );
  AOI211_X1 U11038 ( .C1(n9864), .C2(n10061), .A(n9863), .B(n9862), .ZN(n9956)
         );
  MUX2_X1 U11039 ( .A(n9865), .B(n9956), .S(n10073), .Z(n9866) );
  OAI21_X1 U11040 ( .B1(n9959), .B2(n9902), .A(n9866), .ZN(P1_U3538) );
  INV_X1 U11041 ( .A(n9867), .ZN(n9868) );
  AOI211_X1 U11042 ( .C1(n10064), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9960)
         );
  MUX2_X1 U11043 ( .A(n10024), .B(n9960), .S(n10073), .Z(n9871) );
  OAI21_X1 U11044 ( .B1(n9964), .B2(n9872), .A(n9871), .ZN(P1_U3537) );
  OAI211_X1 U11045 ( .C1(n9875), .C2(n9889), .A(n9874), .B(n9873), .ZN(n9965)
         );
  MUX2_X1 U11046 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9965), .S(n10073), .Z(
        n9876) );
  AOI21_X1 U11047 ( .B1(n6366), .B2(n9967), .A(n9876), .ZN(n9877) );
  INV_X1 U11048 ( .A(n9877), .ZN(P1_U3536) );
  INV_X1 U11049 ( .A(n9878), .ZN(n9883) );
  AOI21_X1 U11050 ( .B1(n10064), .B2(n9880), .A(n9879), .ZN(n9881) );
  OAI211_X1 U11051 ( .C1(n9883), .C2(n9889), .A(n9882), .B(n9881), .ZN(n9969)
         );
  MUX2_X1 U11052 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9969), .S(n10073), .Z(
        P1_U3535) );
  AOI21_X1 U11053 ( .B1(n10064), .B2(n9885), .A(n9884), .ZN(n9886) );
  OAI211_X1 U11054 ( .C1(n9889), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9970)
         );
  MUX2_X1 U11055 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9970), .S(n10073), .Z(
        P1_U3533) );
  AOI211_X1 U11056 ( .C1(n10061), .C2(n9892), .A(n9891), .B(n9890), .ZN(n9971)
         );
  MUX2_X1 U11057 ( .A(n9893), .B(n9971), .S(n10073), .Z(n9894) );
  OAI21_X1 U11058 ( .B1(n9974), .B2(n9902), .A(n9894), .ZN(P1_U3531) );
  INV_X1 U11059 ( .A(n9895), .ZN(n9898) );
  AOI211_X1 U11060 ( .C1(n9899), .C2(n9898), .A(n9897), .B(n9896), .ZN(n9975)
         );
  MUX2_X1 U11061 ( .A(n9900), .B(n9975), .S(n10073), .Z(n9901) );
  OAI21_X1 U11062 ( .B1(n9979), .B2(n9902), .A(n9901), .ZN(P1_U3530) );
  INV_X1 U11063 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9904) );
  MUX2_X1 U11064 ( .A(n9904), .B(n9903), .S(n10070), .Z(n9905) );
  OAI21_X1 U11065 ( .B1(n6518), .B2(n9978), .A(n9905), .ZN(P1_U3520) );
  INV_X1 U11066 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9910) );
  MUX2_X1 U11067 ( .A(n9910), .B(n9909), .S(n10070), .Z(n9911) );
  OAI22_X1 U11068 ( .A1(n9914), .A2(n9963), .B1(n9913), .B2(n9978), .ZN(n9917)
         );
  MUX2_X1 U11069 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9915), .S(n10070), .Z(
        n9916) );
  OR2_X1 U11070 ( .A1(n9917), .A2(n9916), .ZN(P1_U3515) );
  MUX2_X1 U11071 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9918), .S(n10070), .Z(
        n9919) );
  AOI21_X1 U11072 ( .B1(n5687), .B2(n9920), .A(n9919), .ZN(n9921) );
  INV_X1 U11073 ( .A(n9921), .ZN(P1_U3514) );
  AOI22_X1 U11074 ( .A1(n9923), .A2(n9952), .B1(n5687), .B2(n9922), .ZN(n9927)
         );
  MUX2_X1 U11075 ( .A(n9925), .B(n9924), .S(n10070), .Z(n9926) );
  NAND2_X1 U11076 ( .A1(n9927), .A2(n9926), .ZN(P1_U3513) );
  INV_X1 U11077 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9929) );
  MUX2_X1 U11078 ( .A(n9929), .B(n9928), .S(n10070), .Z(n9930) );
  OAI21_X1 U11079 ( .B1(n9931), .B2(n9978), .A(n9930), .ZN(P1_U3512) );
  MUX2_X1 U11080 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9932), .S(n10070), .Z(
        n9936) );
  OAI22_X1 U11081 ( .A1(n9934), .A2(n9963), .B1(n9933), .B2(n9978), .ZN(n9935)
         );
  OR2_X1 U11082 ( .A1(n9936), .A2(n9935), .ZN(P1_U3511) );
  MUX2_X1 U11083 ( .A(n9938), .B(n9937), .S(n10070), .Z(n9939) );
  OAI21_X1 U11084 ( .B1(n9940), .B2(n9963), .A(n9939), .ZN(P1_U3510) );
  MUX2_X1 U11085 ( .A(n9942), .B(n9941), .S(n10070), .Z(n9943) );
  OAI21_X1 U11086 ( .B1(n9944), .B2(n9963), .A(n9943), .ZN(P1_U3509) );
  INV_X1 U11087 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9946) );
  MUX2_X1 U11088 ( .A(n9946), .B(n9945), .S(n10070), .Z(n9947) );
  OAI21_X1 U11089 ( .B1(n9948), .B2(n9963), .A(n9947), .ZN(P1_U3507) );
  INV_X1 U11090 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9949) );
  MUX2_X1 U11091 ( .A(n9950), .B(n9949), .S(n6383), .Z(n9955) );
  AOI22_X1 U11092 ( .A1(n9953), .A2(n9952), .B1(n5687), .B2(n9951), .ZN(n9954)
         );
  NAND2_X1 U11093 ( .A1(n9955), .A2(n9954), .ZN(P1_U3504) );
  INV_X1 U11094 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9957) );
  MUX2_X1 U11095 ( .A(n9957), .B(n9956), .S(n10070), .Z(n9958) );
  OAI21_X1 U11096 ( .B1(n9959), .B2(n9978), .A(n9958), .ZN(P1_U3501) );
  MUX2_X1 U11097 ( .A(n9961), .B(n9960), .S(n10070), .Z(n9962) );
  OAI21_X1 U11098 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(P1_U3498) );
  MUX2_X1 U11099 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9965), .S(n10070), .Z(
        n9966) );
  AOI21_X1 U11100 ( .B1(n5687), .B2(n9967), .A(n9966), .ZN(n9968) );
  INV_X1 U11101 ( .A(n9968), .ZN(P1_U3495) );
  MUX2_X1 U11102 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9969), .S(n10070), .Z(
        P1_U3492) );
  MUX2_X1 U11103 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9970), .S(n10070), .Z(
        P1_U3486) );
  INV_X1 U11104 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9972) );
  MUX2_X1 U11105 ( .A(n9972), .B(n9971), .S(n10070), .Z(n9973) );
  OAI21_X1 U11106 ( .B1(n9974), .B2(n9978), .A(n9973), .ZN(P1_U3480) );
  MUX2_X1 U11107 ( .A(n9976), .B(n9975), .S(n10070), .Z(n9977) );
  OAI21_X1 U11108 ( .B1(n9979), .B2(n9978), .A(n9977), .ZN(P1_U3477) );
  MUX2_X1 U11109 ( .A(P1_D_REG_1__SCAN_IN), .B(n9980), .S(n10051), .Z(P1_U3440) );
  INV_X1 U11110 ( .A(n9981), .ZN(n9986) );
  NOR4_X1 U11111 ( .A1(n9982), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9983), .ZN(n9984) );
  AOI21_X1 U11112 ( .B1(n9988), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9984), .ZN(
        n9985) );
  OAI21_X1 U11113 ( .B1(n9986), .B2(n9994), .A(n9985), .ZN(P1_U3324) );
  AOI22_X1 U11114 ( .A1(n9987), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9988), .ZN(n9989) );
  OAI21_X1 U11115 ( .B1(n9990), .B2(n9994), .A(n9989), .ZN(P1_U3325) );
  OAI222_X1 U11116 ( .A1(n9994), .A2(n9993), .B1(n10002), .B2(P1_U3086), .C1(
        n9991), .C2(n9995), .ZN(P1_U3328) );
  OAI222_X1 U11117 ( .A1(n9994), .A2(n9998), .B1(P1_U3086), .B2(n9997), .C1(
        n9996), .C2(n9995), .ZN(P1_U3329) );
  MUX2_X1 U11118 ( .A(n9999), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11119 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11120 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI21_X1 U11121 ( .B1(n10002), .B2(n10001), .A(n10000), .ZN(n10003) );
  XNOR2_X1 U11122 ( .A(n10003), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11123 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10004), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10005) );
  OAI21_X1 U11124 ( .B1(n10007), .B2(n10006), .A(n10005), .ZN(P1_U3243) );
  INV_X1 U11125 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10020) );
  AOI211_X1 U11126 ( .C1(n10010), .C2(n10009), .A(n10034), .B(n10008), .ZN(
        n10017) );
  OAI211_X1 U11127 ( .C1(n10013), .C2(n10012), .A(n10011), .B(n10037), .ZN(
        n10014) );
  OAI21_X1 U11128 ( .B1(n10043), .B2(n10015), .A(n10014), .ZN(n10016) );
  NOR2_X1 U11129 ( .A1(n10017), .A2(n10016), .ZN(n10019) );
  NAND2_X1 U11130 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10018)
         );
  OAI211_X1 U11131 ( .C1(n10050), .C2(n10020), .A(n10019), .B(n10018), .ZN(
        P1_U3257) );
  INV_X1 U11132 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10033) );
  AOI211_X1 U11133 ( .C1(n10024), .C2(n10023), .A(n10022), .B(n10021), .ZN(
        n10028) );
  AOI211_X1 U11134 ( .C1(n10026), .C2(n9782), .A(n10025), .B(n10034), .ZN(
        n10027) );
  AOI211_X1 U11135 ( .C1(n10030), .C2(n10029), .A(n10028), .B(n10027), .ZN(
        n10032) );
  OAI211_X1 U11136 ( .C1(n10050), .C2(n10033), .A(n10032), .B(n10031), .ZN(
        P1_U3258) );
  INV_X1 U11137 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10049) );
  AOI21_X1 U11138 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10046) );
  OAI211_X1 U11139 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10041) );
  OAI21_X1 U11140 ( .B1(n10043), .B2(n10042), .A(n10041), .ZN(n10044) );
  AOI21_X1 U11141 ( .B1(n10046), .B2(n10045), .A(n10044), .ZN(n10048) );
  NAND2_X1 U11142 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3086), .ZN(n10047)
         );
  OAI211_X1 U11143 ( .C1(n10050), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        P1_U3261) );
  AND2_X1 U11144 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10052), .ZN(P1_U3294) );
  AND2_X1 U11145 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10052), .ZN(P1_U3295) );
  INV_X1 U11146 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10273) );
  NOR2_X1 U11147 ( .A1(n10051), .A2(n10273), .ZN(P1_U3296) );
  AND2_X1 U11148 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10052), .ZN(P1_U3297) );
  AND2_X1 U11149 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10052), .ZN(P1_U3298) );
  AND2_X1 U11150 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10052), .ZN(P1_U3299) );
  AND2_X1 U11151 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10052), .ZN(P1_U3300) );
  AND2_X1 U11152 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10052), .ZN(P1_U3301) );
  AND2_X1 U11153 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10052), .ZN(P1_U3302) );
  AND2_X1 U11154 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10052), .ZN(P1_U3303) );
  AND2_X1 U11155 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10052), .ZN(P1_U3304) );
  AND2_X1 U11156 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10052), .ZN(P1_U3305) );
  AND2_X1 U11157 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10052), .ZN(P1_U3306) );
  AND2_X1 U11158 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10052), .ZN(P1_U3307) );
  AND2_X1 U11159 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10052), .ZN(P1_U3308) );
  AND2_X1 U11160 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10052), .ZN(P1_U3309) );
  AND2_X1 U11161 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10052), .ZN(P1_U3310) );
  AND2_X1 U11162 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10052), .ZN(P1_U3311) );
  AND2_X1 U11163 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10052), .ZN(P1_U3312) );
  AND2_X1 U11164 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10052), .ZN(P1_U3313) );
  AND2_X1 U11165 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10052), .ZN(P1_U3314) );
  AND2_X1 U11166 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10052), .ZN(P1_U3315) );
  AND2_X1 U11167 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10052), .ZN(P1_U3316) );
  INV_X1 U11168 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U11169 ( .A1(n10051), .A2(n10218), .ZN(P1_U3317) );
  AND2_X1 U11170 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10052), .ZN(P1_U3318) );
  AND2_X1 U11171 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10052), .ZN(P1_U3319) );
  AND2_X1 U11172 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10052), .ZN(P1_U3320) );
  AND2_X1 U11173 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10052), .ZN(P1_U3321) );
  AND2_X1 U11174 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10052), .ZN(P1_U3322) );
  AND2_X1 U11175 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10052), .ZN(P1_U3323) );
  INV_X1 U11176 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10053) );
  AOI22_X1 U11177 ( .A1(n10070), .A2(n10054), .B1(n10053), .B2(n6383), .ZN(
        P1_U3453) );
  OAI21_X1 U11178 ( .B1(n10057), .B2(n10056), .A(n10055), .ZN(n10059) );
  AOI211_X1 U11179 ( .C1(n10061), .C2(n10060), .A(n10059), .B(n10058), .ZN(
        n10071) );
  AOI22_X1 U11180 ( .A1(n10070), .A2(n10071), .B1(n5103), .B2(n6383), .ZN(
        P1_U3468) );
  AOI21_X1 U11181 ( .B1(n10064), .B2(n10063), .A(n10062), .ZN(n10065) );
  OAI211_X1 U11182 ( .C1(n10068), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10069) );
  INV_X1 U11183 ( .A(n10069), .ZN(n10072) );
  AOI22_X1 U11184 ( .A1(n10070), .A2(n10072), .B1(n5156), .B2(n6383), .ZN(
        P1_U3474) );
  AOI22_X1 U11185 ( .A1(n10073), .A2(n10071), .B1(n7564), .B2(n7060), .ZN(
        P1_U3527) );
  AOI22_X1 U11186 ( .A1(n10073), .A2(n10072), .B1(n7567), .B2(n7060), .ZN(
        P1_U3529) );
  INV_X1 U11187 ( .A(n10074), .ZN(n10076) );
  NAND2_X1 U11188 ( .A1(n10076), .A2(n10075), .ZN(n10077) );
  NAND2_X1 U11189 ( .A1(n10142), .A2(n10113), .ZN(n10085) );
  AOI22_X1 U11190 ( .A1(n10080), .A2(n10091), .B1(n10093), .B2(n10079), .ZN(
        n10084) );
  XNOR2_X1 U11191 ( .A(n10081), .B(n4401), .ZN(n10082) );
  NAND2_X1 U11192 ( .A1(n10082), .A2(n10096), .ZN(n10083) );
  INV_X1 U11193 ( .A(n10086), .ZN(n10087) );
  AOI222_X1 U11194 ( .A1(n10088), .A2(n10102), .B1(n10142), .B2(n10087), .C1(
        n10140), .C2(n10101), .ZN(n10089) );
  OAI221_X1 U11195 ( .B1(n10107), .B2(n10144), .C1(n7308), .C2(n7510), .A(
        n10089), .ZN(P2_U3226) );
  XNOR2_X1 U11196 ( .A(n10090), .B(n10098), .ZN(n10095) );
  AOI222_X1 U11197 ( .A1(n10096), .A2(n10095), .B1(n10094), .B2(n10093), .C1(
        n10092), .C2(n10091), .ZN(n10127) );
  OAI21_X1 U11198 ( .B1(n10099), .B2(n10098), .A(n10097), .ZN(n10125) );
  INV_X1 U11199 ( .A(n10100), .ZN(n10103) );
  AOI222_X1 U11200 ( .A1(n10125), .A2(n10104), .B1(n10103), .B2(n10102), .C1(
        n10124), .C2(n10101), .ZN(n10105) );
  OAI221_X1 U11201 ( .B1(n10107), .B2(n10127), .C1(n7308), .C2(n10106), .A(
        n10105), .ZN(P2_U3229) );
  INV_X1 U11202 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10114) );
  NAND2_X1 U11203 ( .A1(n10112), .A2(n10141), .ZN(n10108) );
  OAI21_X1 U11204 ( .B1(n10109), .B2(n10135), .A(n10108), .ZN(n10111) );
  AOI211_X1 U11205 ( .C1(n10113), .C2(n10112), .A(n10111), .B(n10110), .ZN(
        n10156) );
  AOI22_X1 U11206 ( .A1(n10154), .A2(n10114), .B1(n10156), .B2(n10152), .ZN(
        P2_U3393) );
  INV_X1 U11207 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U11208 ( .A1(n10115), .A2(n10146), .ZN(n10117) );
  AOI211_X1 U11209 ( .C1(n10151), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        n10157) );
  AOI22_X1 U11210 ( .A1(n10154), .A2(n10217), .B1(n10157), .B2(n10152), .ZN(
        P2_U3396) );
  INV_X1 U11211 ( .A(n10119), .ZN(n10123) );
  OAI21_X1 U11212 ( .B1(n10121), .B2(n10135), .A(n10120), .ZN(n10122) );
  AOI21_X1 U11213 ( .B1(n10139), .B2(n10123), .A(n10122), .ZN(n10159) );
  AOI22_X1 U11214 ( .A1(n10154), .A2(n5959), .B1(n10159), .B2(n10152), .ZN(
        P2_U3399) );
  INV_X1 U11215 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10128) );
  AOI22_X1 U11216 ( .A1(n10125), .A2(n10139), .B1(n10151), .B2(n10124), .ZN(
        n10126) );
  AND2_X1 U11217 ( .A1(n10127), .A2(n10126), .ZN(n10160) );
  AOI22_X1 U11218 ( .A1(n10154), .A2(n10128), .B1(n10160), .B2(n10152), .ZN(
        P2_U3402) );
  AOI22_X1 U11219 ( .A1(n10130), .A2(n10141), .B1(n10151), .B2(n10129), .ZN(
        n10131) );
  AND2_X1 U11220 ( .A1(n10132), .A2(n10131), .ZN(n10161) );
  AOI22_X1 U11221 ( .A1(n10154), .A2(n5978), .B1(n10161), .B2(n10152), .ZN(
        P2_U3405) );
  INV_X1 U11222 ( .A(n10133), .ZN(n10138) );
  OAI21_X1 U11223 ( .B1(n10136), .B2(n10135), .A(n10134), .ZN(n10137) );
  AOI21_X1 U11224 ( .B1(n10139), .B2(n10138), .A(n10137), .ZN(n10162) );
  AOI22_X1 U11225 ( .A1(n10154), .A2(n5992), .B1(n10162), .B2(n10152), .ZN(
        P2_U3408) );
  INV_X1 U11226 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U11227 ( .A1(n10142), .A2(n10141), .B1(n10151), .B2(n10140), .ZN(
        n10143) );
  AOI22_X1 U11228 ( .A1(n10154), .A2(n10145), .B1(n10163), .B2(n10152), .ZN(
        P2_U3411) );
  INV_X1 U11229 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10153) );
  NOR2_X1 U11230 ( .A1(n10147), .A2(n10146), .ZN(n10149) );
  AOI211_X1 U11231 ( .C1(n10151), .C2(n10150), .A(n10149), .B(n10148), .ZN(
        n10165) );
  AOI22_X1 U11232 ( .A1(n10154), .A2(n10153), .B1(n10165), .B2(n10152), .ZN(
        P2_U3414) );
  INV_X1 U11233 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U11234 ( .A1(n10166), .A2(n10156), .B1(n10155), .B2(n10164), .ZN(
        P2_U3460) );
  AOI22_X1 U11235 ( .A1(n10166), .A2(n10157), .B1(n5806), .B2(n10164), .ZN(
        P2_U3461) );
  AOI22_X1 U11236 ( .A1(n10166), .A2(n10159), .B1(n10158), .B2(n10164), .ZN(
        P2_U3462) );
  AOI22_X1 U11237 ( .A1(n10166), .A2(n10160), .B1(n5971), .B2(n10164), .ZN(
        P2_U3463) );
  AOI22_X1 U11238 ( .A1(n10166), .A2(n10161), .B1(n5982), .B2(n10164), .ZN(
        P2_U3464) );
  AOI22_X1 U11239 ( .A1(n10166), .A2(n10162), .B1(n5995), .B2(n10164), .ZN(
        P2_U3465) );
  AOI22_X1 U11240 ( .A1(n10166), .A2(n10163), .B1(n7508), .B2(n10164), .ZN(
        P2_U3466) );
  AOI22_X1 U11241 ( .A1(n10166), .A2(n10165), .B1(n6009), .B2(n10164), .ZN(
        P2_U3467) );
  INV_X1 U11242 ( .A(n10167), .ZN(n10168) );
  NAND2_X1 U11243 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  XNOR2_X1 U11244 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10170), .ZN(ADD_1068_U5)
         );
  XOR2_X1 U11245 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  NOR2_X1 U11246 ( .A1(n10172), .A2(n10171), .ZN(n10173) );
  XOR2_X1 U11247 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10173), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11248 ( .A(n10175), .B(n10174), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11249 ( .A(n10177), .B(n10176), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11250 ( .A(n10179), .B(n10178), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11251 ( .A(n10181), .B(n10180), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11252 ( .A(n10183), .B(n10182), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11253 ( .A(n10185), .B(n10184), .ZN(ADD_1068_U61) );
  XNOR2_X1 U11254 ( .A(n10187), .B(n10186), .ZN(ADD_1068_U62) );
  XNOR2_X1 U11255 ( .A(n10189), .B(n10188), .ZN(ADD_1068_U63) );
  NAND4_X1 U11256 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(P2_REG2_REG_6__SCAN_IN), 
        .A3(P1_REG2_REG_30__SCAN_IN), .A4(n7508), .ZN(n10195) );
  INV_X1 U11257 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10291) );
  NAND4_X1 U11258 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(P2_REG2_REG_28__SCAN_IN), 
        .A3(n9664), .A4(n10291), .ZN(n10194) );
  NAND4_X1 U11259 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(SI_26_), .A3(
        P1_D_REG_29__SCAN_IN), .A4(n10274), .ZN(n10193) );
  NAND4_X1 U11260 ( .A1(n10191), .A2(n10190), .A3(n5103), .A4(
        P2_D_REG_22__SCAN_IN), .ZN(n10192) );
  NOR4_X1 U11261 ( .A1(n10195), .A2(n10194), .A3(n10193), .A4(n10192), .ZN(
        n10329) );
  NAND3_X1 U11262 ( .A1(P1_REG0_REG_29__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .A3(n10314), .ZN(n10215) );
  NOR3_X1 U11263 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .A3(n10298), .ZN(n10198) );
  NOR4_X1 U11264 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P1_REG1_REG_24__SCAN_IN), 
        .A3(P1_REG2_REG_20__SCAN_IN), .A4(n10196), .ZN(n10197) );
  NAND3_X1 U11265 ( .A1(n10199), .A2(n10198), .A3(n10197), .ZN(n10200) );
  NOR3_X1 U11266 ( .A1(n10200), .A2(SI_9_), .A3(P2_REG3_REG_9__SCAN_IN), .ZN(
        n10201) );
  NAND3_X1 U11267 ( .A1(n10201), .A2(P2_DATAO_REG_1__SCAN_IN), .A3(SI_16_), 
        .ZN(n10214) );
  NOR4_X1 U11268 ( .A1(P2_REG1_REG_24__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), 
        .A3(P1_REG3_REG_21__SCAN_IN), .A4(n10217), .ZN(n10212) );
  NAND4_X1 U11269 ( .A1(SI_29_), .A2(P1_IR_REG_2__SCAN_IN), .A3(
        P2_ADDR_REG_2__SCAN_IN), .A4(P1_ADDR_REG_1__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U11270 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .A3(P1_REG0_REG_20__SCAN_IN), .A4(n10230), .ZN(n10203) );
  NAND3_X1 U11271 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P1_DATAO_REG_21__SCAN_IN), 
        .A3(SI_31_), .ZN(n10202) );
  NOR4_X1 U11272 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(n10204), .A3(n10203), .A4(
        n10202), .ZN(n10211) );
  NOR4_X1 U11273 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), 
        .A3(P1_REG2_REG_14__SCAN_IN), .A4(n10258), .ZN(n10210) );
  NAND4_X1 U11274 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10256), .A3(n8381), 
        .A4(n10253), .ZN(n10208) );
  NAND4_X1 U11275 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_REG2_REG_18__SCAN_IN), 
        .A3(P1_IR_REG_30__SCAN_IN), .A4(P1_REG3_REG_22__SCAN_IN), .ZN(n10205)
         );
  OR3_X1 U11276 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), 
        .A3(n10205), .ZN(n10206) );
  NOR4_X1 U11277 ( .A1(n10208), .A2(P1_REG3_REG_4__SCAN_IN), .A3(n10207), .A4(
        n10206), .ZN(n10209) );
  NAND4_X1 U11278 ( .A1(n10212), .A2(n10211), .A3(n10210), .A4(n10209), .ZN(
        n10213) );
  NOR4_X1 U11279 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n10215), .A3(n10214), 
        .A4(n10213), .ZN(n10328) );
  AOI22_X1 U11280 ( .A1(n10218), .A2(keyinput58), .B1(n10217), .B2(keyinput53), 
        .ZN(n10216) );
  OAI221_X1 U11281 ( .B1(n10218), .B2(keyinput58), .C1(n10217), .C2(keyinput53), .A(n10216), .ZN(n10228) );
  AOI22_X1 U11282 ( .A1(n4985), .A2(keyinput59), .B1(n5572), .B2(keyinput26), 
        .ZN(n10219) );
  OAI221_X1 U11283 ( .B1(n4985), .B2(keyinput59), .C1(n5572), .C2(keyinput26), 
        .A(n10219), .ZN(n10227) );
  AOI22_X1 U11284 ( .A1(n10222), .A2(keyinput1), .B1(keyinput63), .B2(n10221), 
        .ZN(n10220) );
  OAI221_X1 U11285 ( .B1(n10222), .B2(keyinput1), .C1(n10221), .C2(keyinput63), 
        .A(n10220), .ZN(n10226) );
  XNOR2_X1 U11286 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput41), .ZN(n10224)
         );
  XNOR2_X1 U11287 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput12), .ZN(n10223) );
  NAND2_X1 U11288 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  NOR4_X1 U11289 ( .A1(n10228), .A2(n10227), .A3(n10226), .A4(n10225), .ZN(
        n10269) );
  INV_X1 U11290 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U11291 ( .A1(n10231), .A2(keyinput42), .B1(n10230), .B2(keyinput0), 
        .ZN(n10229) );
  OAI221_X1 U11292 ( .B1(n10231), .B2(keyinput42), .C1(n10230), .C2(keyinput0), 
        .A(n10229), .ZN(n10240) );
  AOI22_X1 U11293 ( .A1(n10233), .A2(keyinput36), .B1(keyinput60), .B2(n6523), 
        .ZN(n10232) );
  OAI221_X1 U11294 ( .B1(n10233), .B2(keyinput36), .C1(n6523), .C2(keyinput60), 
        .A(n10232), .ZN(n10239) );
  XNOR2_X1 U11295 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput47), .ZN(n10237)
         );
  XNOR2_X1 U11296 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput50), .ZN(n10236) );
  XNOR2_X1 U11297 ( .A(P2_REG2_REG_18__SCAN_IN), .B(keyinput24), .ZN(n10235)
         );
  XNOR2_X1 U11298 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput18), .ZN(n10234) );
  NAND4_X1 U11299 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10238) );
  NOR3_X1 U11300 ( .A1(n10240), .A2(n10239), .A3(n10238), .ZN(n10268) );
  INV_X1 U11301 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U11302 ( .A1(n10242), .A2(keyinput31), .B1(n8381), .B2(keyinput32), 
        .ZN(n10241) );
  OAI221_X1 U11303 ( .B1(n10242), .B2(keyinput31), .C1(n8381), .C2(keyinput32), 
        .A(n10241), .ZN(n10251) );
  XNOR2_X1 U11304 ( .A(keyinput34), .B(n4995), .ZN(n10250) );
  XNOR2_X1 U11305 ( .A(keyinput4), .B(n10243), .ZN(n10249) );
  XNOR2_X1 U11306 ( .A(P2_IR_REG_7__SCAN_IN), .B(keyinput2), .ZN(n10247) );
  XNOR2_X1 U11307 ( .A(P1_REG3_REG_22__SCAN_IN), .B(keyinput13), .ZN(n10246)
         );
  XNOR2_X1 U11308 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput33), .ZN(n10245) );
  XNOR2_X1 U11309 ( .A(P1_REG3_REG_4__SCAN_IN), .B(keyinput55), .ZN(n10244) );
  NAND4_X1 U11310 ( .A1(n10247), .A2(n10246), .A3(n10245), .A4(n10244), .ZN(
        n10248) );
  NOR4_X1 U11311 ( .A1(n10251), .A2(n10250), .A3(n10249), .A4(n10248), .ZN(
        n10267) );
  AOI22_X1 U11312 ( .A1(n10253), .A2(keyinput23), .B1(keyinput7), .B2(n9745), 
        .ZN(n10252) );
  OAI221_X1 U11313 ( .B1(n10253), .B2(keyinput23), .C1(n9745), .C2(keyinput7), 
        .A(n10252), .ZN(n10265) );
  AOI22_X1 U11314 ( .A1(n10256), .A2(keyinput61), .B1(keyinput45), .B2(n10255), 
        .ZN(n10254) );
  OAI221_X1 U11315 ( .B1(n10256), .B2(keyinput61), .C1(n10255), .C2(keyinput45), .A(n10254), .ZN(n10264) );
  AOI22_X1 U11316 ( .A1(n10259), .A2(keyinput37), .B1(keyinput46), .B2(n10258), 
        .ZN(n10257) );
  OAI221_X1 U11317 ( .B1(n10259), .B2(keyinput37), .C1(n10258), .C2(keyinput46), .A(n10257), .ZN(n10263) );
  AOI22_X1 U11318 ( .A1(n4997), .A2(keyinput52), .B1(n10261), .B2(keyinput21), 
        .ZN(n10260) );
  OAI221_X1 U11319 ( .B1(n4997), .B2(keyinput52), .C1(n10261), .C2(keyinput21), 
        .A(n10260), .ZN(n10262) );
  NOR4_X1 U11320 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10266) );
  NAND4_X1 U11321 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10327) );
  AOI22_X1 U11322 ( .A1(n5103), .A2(keyinput40), .B1(n10271), .B2(keyinput56), 
        .ZN(n10270) );
  OAI221_X1 U11323 ( .B1(n5103), .B2(keyinput40), .C1(n10271), .C2(keyinput56), 
        .A(n10270), .ZN(n10283) );
  AOI22_X1 U11324 ( .A1(n10274), .A2(keyinput19), .B1(n10273), .B2(keyinput9), 
        .ZN(n10272) );
  OAI221_X1 U11325 ( .B1(n10274), .B2(keyinput19), .C1(n10273), .C2(keyinput9), 
        .A(n10272), .ZN(n10282) );
  AOI22_X1 U11326 ( .A1(n10277), .A2(keyinput11), .B1(n10276), .B2(keyinput38), 
        .ZN(n10275) );
  OAI221_X1 U11327 ( .B1(n10277), .B2(keyinput11), .C1(n10276), .C2(keyinput38), .A(n10275), .ZN(n10281) );
  XNOR2_X1 U11328 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput3), .ZN(n10279) );
  XNOR2_X1 U11329 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput25), .ZN(n10278)
         );
  NAND2_X1 U11330 ( .A1(n10279), .A2(n10278), .ZN(n10280) );
  NOR4_X1 U11331 ( .A1(n10283), .A2(n10282), .A3(n10281), .A4(n10280), .ZN(
        n10325) );
  INV_X1 U11332 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10285) );
  AOI22_X1 U11333 ( .A1(n10286), .A2(keyinput14), .B1(keyinput6), .B2(n10285), 
        .ZN(n10284) );
  OAI221_X1 U11334 ( .B1(n10286), .B2(keyinput14), .C1(n10285), .C2(keyinput6), 
        .A(n10284), .ZN(n10295) );
  AOI22_X1 U11335 ( .A1(n5675), .A2(keyinput43), .B1(n7508), .B2(keyinput20), 
        .ZN(n10287) );
  OAI221_X1 U11336 ( .B1(n5675), .B2(keyinput43), .C1(n7508), .C2(keyinput20), 
        .A(n10287), .ZN(n10294) );
  AOI22_X1 U11337 ( .A1(n9664), .A2(keyinput44), .B1(n10289), .B2(keyinput62), 
        .ZN(n10288) );
  OAI221_X1 U11338 ( .B1(n9664), .B2(keyinput44), .C1(n10289), .C2(keyinput62), 
        .A(n10288), .ZN(n10293) );
  AOI22_X1 U11339 ( .A1(n10291), .A2(keyinput16), .B1(n6224), .B2(keyinput17), 
        .ZN(n10290) );
  OAI221_X1 U11340 ( .B1(n10291), .B2(keyinput16), .C1(n6224), .C2(keyinput17), 
        .A(n10290), .ZN(n10292) );
  NOR4_X1 U11341 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10324) );
  INV_X1 U11342 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11343 ( .A1(n10298), .A2(keyinput5), .B1(keyinput35), .B2(n10297), 
        .ZN(n10296) );
  OAI221_X1 U11344 ( .B1(n10298), .B2(keyinput5), .C1(n10297), .C2(keyinput35), 
        .A(n10296), .ZN(n10308) );
  AOI22_X1 U11345 ( .A1(n10301), .A2(keyinput57), .B1(n10300), .B2(keyinput22), 
        .ZN(n10299) );
  OAI221_X1 U11346 ( .B1(n10301), .B2(keyinput57), .C1(n10300), .C2(keyinput22), .A(n10299), .ZN(n10307) );
  XNOR2_X1 U11347 ( .A(SI_16_), .B(keyinput27), .ZN(n10305) );
  XNOR2_X1 U11348 ( .A(P1_REG3_REG_0__SCAN_IN), .B(keyinput10), .ZN(n10304) );
  XNOR2_X1 U11349 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput54), .ZN(n10303)
         );
  XNOR2_X1 U11350 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput48), .ZN(n10302)
         );
  NAND4_X1 U11351 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n10306) );
  NOR3_X1 U11352 ( .A1(n10308), .A2(n10307), .A3(n10306), .ZN(n10323) );
  INV_X1 U11353 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U11354 ( .A1(n10311), .A2(keyinput28), .B1(keyinput51), .B2(n10310), 
        .ZN(n10309) );
  OAI221_X1 U11355 ( .B1(n10311), .B2(keyinput28), .C1(n10310), .C2(keyinput51), .A(n10309), .ZN(n10321) );
  AOI22_X1 U11356 ( .A1(n10314), .A2(keyinput49), .B1(keyinput39), .B2(n10313), 
        .ZN(n10312) );
  OAI221_X1 U11357 ( .B1(n10314), .B2(keyinput49), .C1(n10313), .C2(keyinput39), .A(n10312), .ZN(n10320) );
  XNOR2_X1 U11358 ( .A(P1_REG1_REG_12__SCAN_IN), .B(keyinput30), .ZN(n10318)
         );
  XNOR2_X1 U11359 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput15), .ZN(n10317) );
  XNOR2_X1 U11360 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(keyinput29), .ZN(n10316)
         );
  XNOR2_X1 U11361 ( .A(P1_REG0_REG_29__SCAN_IN), .B(keyinput8), .ZN(n10315) );
  NAND4_X1 U11362 ( .A1(n10318), .A2(n10317), .A3(n10316), .A4(n10315), .ZN(
        n10319) );
  NOR3_X1 U11363 ( .A1(n10321), .A2(n10320), .A3(n10319), .ZN(n10322) );
  NAND4_X1 U11364 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10326) );
  AOI211_X1 U11365 ( .C1(n10329), .C2(n10328), .A(n10327), .B(n10326), .ZN(
        n10346) );
  AOI22_X1 U11366 ( .A1(n10333), .A2(n10332), .B1(n10331), .B2(n10330), .ZN(
        n10339) );
  INV_X1 U11367 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U11368 ( .A1(n10337), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10336), 
        .B2(n10335), .ZN(n10338) );
  OAI211_X1 U11369 ( .C1(n10341), .C2(n10340), .A(n10339), .B(n10338), .ZN(
        n10342) );
  AOI21_X1 U11370 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(n10345) );
  XNOR2_X1 U11371 ( .A(n10346), .B(n10345), .ZN(P1_U3290) );
  XNOR2_X1 U11372 ( .A(n10348), .B(n10347), .ZN(ADD_1068_U50) );
  XNOR2_X1 U11373 ( .A(n10350), .B(n10349), .ZN(ADD_1068_U51) );
  XNOR2_X1 U11374 ( .A(n10352), .B(n10351), .ZN(ADD_1068_U47) );
  XNOR2_X1 U11375 ( .A(n10354), .B(n10353), .ZN(ADD_1068_U49) );
  XNOR2_X1 U11376 ( .A(n10356), .B(n10355), .ZN(ADD_1068_U48) );
  XOR2_X1 U11377 ( .A(n10358), .B(n10357), .Z(ADD_1068_U54) );
  XOR2_X1 U11378 ( .A(n10360), .B(n10359), .Z(ADD_1068_U53) );
  XNOR2_X1 U11379 ( .A(n10362), .B(n10361), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4816 ( .A(n6801), .Z(n6803) );
  CLKBUF_X1 U4822 ( .A(n9636), .Z(n9654) );
  CLKBUF_X1 U6500 ( .A(n5640), .Z(n4293) );
  CLKBUF_X1 U6550 ( .A(n5642), .Z(n9374) );
endmodule

