

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676;

  AOI21_X1 U11010 ( .B1(n16168), .B2(n16419), .A(n16161), .ZN(n16427) );
  NAND2_X1 U11011 ( .A1(n9799), .A2(n9798), .ZN(n16196) );
  BUF_X1 U11012 ( .A(n10995), .Z(n14501) );
  NAND2_X1 U11013 ( .A1(n9628), .A2(n14236), .ZN(n20051) );
  NAND2_X1 U11014 ( .A1(n10300), .A2(n12426), .ZN(n16762) );
  INV_X1 U11015 ( .A(n18565), .ZN(n18659) );
  INV_X1 U11016 ( .A(n12428), .ZN(n12404) );
  CLKBUF_X2 U11017 ( .A(n12945), .Z(n12999) );
  INV_X1 U11018 ( .A(n12932), .ZN(n14731) );
  BUF_X2 U11019 ( .A(n12410), .Z(n15822) );
  INV_X1 U11020 ( .A(n14214), .ZN(n18992) );
  XNOR2_X1 U11021 ( .A(n11770), .B(n12400), .ZN(n16665) );
  INV_X1 U11022 ( .A(n17109), .ZN(n18141) );
  INV_X4 U11023 ( .A(n12183), .ZN(n12216) );
  INV_X2 U11024 ( .A(n18086), .ZN(n18132) );
  NAND2_X1 U11025 ( .A1(n10398), .A2(n10399), .ZN(n10128) );
  CLKBUF_X2 U11026 ( .A(n12165), .Z(n12295) );
  AND2_X2 U11027 ( .A1(n11790), .A2(n11656), .ZN(n11872) );
  AND2_X2 U11028 ( .A1(n11784), .A2(n11656), .ZN(n12160) );
  CLKBUF_X2 U11029 ( .A(n11797), .Z(n9581) );
  AND2_X2 U11030 ( .A1(n11972), .A2(n11656), .ZN(n11813) );
  AND2_X1 U11031 ( .A1(n10594), .A2(n10202), .ZN(n14039) );
  OR2_X1 U11032 ( .A1(n10568), .A2(n10567), .ZN(n10607) );
  INV_X1 U11033 ( .A(n10587), .ZN(n10609) );
  AND2_X1 U11034 ( .A1(n10491), .A2(n10490), .ZN(n10496) );
  NAND3_X1 U11035 ( .A1(n13925), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        n14583), .ZN(n10570) );
  AND2_X2 U11036 ( .A1(n10136), .A2(n10468), .ZN(n10626) );
  INV_X1 U11037 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10948) );
  CLKBUF_X1 U11038 ( .A(n18413), .Z(n9566) );
  NOR2_X1 U11039 ( .A1(n18380), .A2(n19442), .ZN(n18413) );
  CLKBUF_X1 U11040 ( .A(n20853), .Z(n9567) );
  NOR2_X1 U11041 ( .A1(n15135), .A2(n17244), .ZN(n20853) );
  INV_X1 U11042 ( .A(n11472), .ZN(n11555) );
  AND2_X2 U11043 ( .A1(n9923), .A2(n13925), .ZN(n10663) );
  NOR2_X1 U11044 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11606) );
  NAND2_X1 U11045 ( .A1(n13707), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10737) );
  NOR2_X2 U11046 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10097) );
  AND2_X1 U11047 ( .A1(n14597), .A2(n11656), .ZN(n12165) );
  NAND2_X2 U11048 ( .A1(n10737), .A2(n10736), .ZN(n10966) );
  XNOR2_X1 U11049 ( .A(n11732), .B(n11734), .ZN(n10162) );
  AND2_X1 U11050 ( .A1(n14167), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13177) );
  INV_X1 U11051 ( .A(n13423), .ZN(n17089) );
  NAND2_X1 U11052 ( .A1(n10599), .A2(n10587), .ZN(n13028) );
  NAND3_X1 U11053 ( .A1(n10274), .A2(n14039), .A3(n10601), .ZN(n13023) );
  INV_X1 U11054 ( .A(n13070), .ZN(n12887) );
  AND2_X1 U11055 ( .A1(n16203), .A2(n12740), .ZN(n16190) );
  NOR2_X1 U11056 ( .A1(n12412), .A2(n15822), .ZN(n9937) );
  NAND2_X1 U11057 ( .A1(n12402), .A2(n10164), .ZN(n20305) );
  INV_X2 U11058 ( .A(n9626), .ZN(n17057) );
  AND2_X1 U11059 ( .A1(n11461), .A2(n11460), .ZN(n11489) );
  CLKBUF_X3 U11060 ( .A(n10901), .Z(n15353) );
  INV_X1 U11061 ( .A(n15353), .ZN(n15333) );
  INV_X1 U11062 ( .A(n12969), .ZN(n12959) );
  MUX2_X1 U11063 ( .A(n13066), .B(n14623), .S(n9587), .Z(n14700) );
  NAND2_X1 U11064 ( .A1(n13663), .A2(n13674), .ZN(n9792) );
  OR2_X1 U11065 ( .A1(n15822), .A2(n10349), .ZN(n20089) );
  INV_X1 U11066 ( .A(n14217), .ZN(n17775) );
  AND2_X1 U11067 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14389) );
  NOR3_X1 U11068 ( .A1(n17117), .A2(n17653), .A3(n17633), .ZN(n18046) );
  INV_X1 U11069 ( .A(n9580), .ZN(n18035) );
  INV_X1 U11070 ( .A(n20677), .ZN(n13732) );
  INV_X1 U11071 ( .A(n20888), .ZN(n20876) );
  AOI21_X1 U11072 ( .B1(n14012), .B2(n14011), .A(n11779), .ZN(n14228) );
  OR2_X1 U11073 ( .A1(n16381), .A2(n9775), .ZN(n10118) );
  NOR2_X1 U11074 ( .A1(n16268), .A2(n16517), .ZN(n16253) );
  INV_X1 U11075 ( .A(n16720), .ZN(n20157) );
  INV_X1 U11076 ( .A(n17807), .ZN(n17712) );
  INV_X1 U11077 ( .A(n17791), .ZN(n17805) );
  AND2_X1 U11078 ( .A1(n9954), .A2(n9953), .ZN(n18120) );
  OR2_X1 U11079 ( .A1(n13731), .A2(n13710), .ZN(n20691) );
  INV_X2 U11080 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U11081 ( .A1(n14232), .A2(n14235), .ZN(n20582) );
  INV_X1 U11082 ( .A(n16665), .ZN(n15847) );
  INV_X1 U11083 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20581) );
  INV_X2 U11084 ( .A(n20619), .ZN(n20618) );
  INV_X2 U11085 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14167) );
  AND2_X1 U11086 ( .A1(n13614), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15135)
         );
  INV_X2 U11087 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11656) );
  AND4_X2 U11088 ( .A1(n9825), .A2(n10933), .A3(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A4(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9568) );
  XOR2_X1 U11089 ( .A(n16195), .B(n16194), .Z(n9569) );
  INV_X2 U11090 ( .A(n10885), .ZN(n10886) );
  INV_X2 U11091 ( .A(n10881), .ZN(n10885) );
  AND3_X1 U11092 ( .A1(n10086), .A2(n12528), .A3(n12527), .ZN(n12540) );
  NAND2_X2 U11094 ( .A1(n10586), .A2(n10790), .ZN(n10602) );
  NAND2_X4 U11095 ( .A1(n10456), .A2(n10496), .ZN(n10790) );
  OR2_X2 U11096 ( .A1(n14437), .A2(n10830), .ZN(n10832) );
  OAI21_X2 U11097 ( .B1(n15359), .B2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n15357), .ZN(n10083) );
  CLKBUF_X3 U11098 ( .A(n11591), .Z(n15359) );
  OAI21_X2 U11099 ( .B1(n13084), .B2(n13083), .A(n13082), .ZN(n13091) );
  NAND2_X2 U11100 ( .A1(n12636), .A2(n12637), .ZN(n12609) );
  AND2_X2 U11101 ( .A1(n15651), .A2(n16144), .ZN(n15638) );
  NAND3_X2 U11102 ( .A1(n10122), .A2(n12551), .A3(n12550), .ZN(n16340) );
  NAND2_X2 U11103 ( .A1(n14048), .A2(n12254), .ZN(n16083) );
  NAND2_X2 U11104 ( .A1(n14051), .A2(n14050), .ZN(n14048) );
  AND2_X2 U11105 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  NAND2_X2 U11106 ( .A1(n10267), .A2(n13333), .ZN(n13338) );
  NAND2_X2 U11107 ( .A1(n9946), .A2(n9945), .ZN(n19997) );
  NAND4_X2 U11108 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12590) );
  AND2_X1 U11109 ( .A1(n12556), .A2(n12102), .ZN(n9571) );
  AND2_X1 U11110 ( .A1(n12556), .A2(n12102), .ZN(n9572) );
  XNOR2_X2 U11111 ( .A(n13286), .B(n13285), .ZN(n18697) );
  NAND2_X2 U11112 ( .A1(n16922), .A2(n13269), .ZN(n13286) );
  AND2_X1 U11113 ( .A1(n9816), .A2(n9815), .ZN(n16370) );
  NAND2_X1 U11114 ( .A1(n16285), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16539) );
  INV_X1 U11115 ( .A(n16268), .ZN(n16285) );
  NAND2_X1 U11116 ( .A1(n9989), .A2(n9988), .ZN(n10212) );
  AND2_X1 U11117 ( .A1(n14785), .A2(n14784), .ZN(n14802) );
  CLKBUF_X1 U11118 ( .A(n16275), .Z(n16276) );
  OAI211_X1 U11119 ( .C1(n12617), .C2(n9782), .A(n12618), .B(n9781), .ZN(
        n16278) );
  NAND2_X1 U11120 ( .A1(n14468), .A2(n14469), .ZN(n14467) );
  AND4_X1 U11121 ( .A1(n15313), .A2(n15316), .A3(n10880), .A4(n15302), .ZN(
        n15304) );
  NAND2_X1 U11122 ( .A1(n14482), .A2(n10835), .ZN(n20775) );
  INV_X4 U11123 ( .A(n20691), .ZN(n20709) );
  CLKBUF_X1 U11124 ( .A(n13347), .Z(n18522) );
  AND2_X2 U11125 ( .A1(n12316), .A2(n9611), .ZN(n13977) );
  NAND2_X1 U11126 ( .A1(n12685), .A2(n12700), .ZN(n12619) );
  NAND2_X1 U11127 ( .A1(n10703), .A2(n20931), .ZN(n10279) );
  NAND2_X1 U11128 ( .A1(n20931), .A2(n10702), .ZN(n10709) );
  XNOR2_X1 U11129 ( .A(n11772), .B(n10128), .ZN(n12400) );
  NAND2_X1 U11130 ( .A1(n14388), .A2(n13768), .ZN(n18978) );
  NAND2_X1 U11131 ( .A1(n9839), .A2(n13248), .ZN(n13268) );
  AOI21_X1 U11132 ( .B1(n14207), .B2(n14206), .A(n19449), .ZN(n17005) );
  NOR2_X4 U11133 ( .A1(n13788), .A2(n12050), .ZN(n11723) );
  INV_X1 U11134 ( .A(n10618), .ZN(n13025) );
  BUF_X2 U11135 ( .A(n12215), .Z(n13640) );
  OR2_X1 U11136 ( .A1(n19004), .A2(n13480), .ZN(n13478) );
  NAND2_X1 U11137 ( .A1(n10970), .A2(n12932), .ZN(n13913) );
  AND2_X1 U11138 ( .A1(n11693), .A2(n11692), .ZN(n12154) );
  AND2_X1 U11139 ( .A1(n10616), .A2(n10916), .ZN(n10274) );
  INV_X1 U11140 ( .A(n14511), .ZN(n13707) );
  INV_X1 U11141 ( .A(n19019), .ZN(n18186) );
  INV_X4 U11142 ( .A(n19001), .ZN(n19570) );
  CLKBUF_X1 U11143 ( .A(n10790), .Z(n20838) );
  INV_X2 U11144 ( .A(n12178), .ZN(n12721) );
  NAND2_X2 U11145 ( .A1(n10607), .A2(n14511), .ZN(n12969) );
  CLKBUF_X2 U11146 ( .A(n10607), .Z(n20819) );
  CLKBUF_X2 U11147 ( .A(n10598), .Z(n20833) );
  INV_X2 U11148 ( .A(n11686), .ZN(n12178) );
  NAND4_X2 U11149 ( .A1(n13381), .A2(n13380), .A3(n13379), .A4(n13378), .ZN(
        n19001) );
  CLKBUF_X2 U11150 ( .A(n11713), .Z(n16735) );
  AND4_X1 U11151 ( .A1(n13176), .A2(n13175), .A3(n13174), .A4(n13173), .ZN(
        n9591) );
  INV_X1 U11152 ( .A(n11702), .ZN(n11699) );
  NAND4_X1 U11153 ( .A1(n10482), .A2(n10481), .A3(n10480), .A4(n10479), .ZN(
        n10598) );
  AND4_X1 U11154 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10481) );
  INV_X4 U11155 ( .A(n17112), .ZN(n18111) );
  CLKBUF_X2 U11156 ( .A(n9568), .Z(n11497) );
  BUF_X2 U11157 ( .A(n10663), .Z(n10651) );
  BUF_X2 U11158 ( .A(n11556), .Z(n11400) );
  INV_X2 U11159 ( .A(n9626), .ZN(n18056) );
  CLKBUF_X2 U11160 ( .A(n10627), .Z(n11551) );
  AND2_X1 U11161 ( .A1(n9579), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11797) );
  INV_X4 U11162 ( .A(n10448), .ZN(n9573) );
  CLKBUF_X2 U11163 ( .A(n10635), .Z(n11557) );
  AND2_X2 U11164 ( .A1(n10468), .A2(n10474), .ZN(n11556) );
  NAND2_X1 U11165 ( .A1(n10136), .A2(n14409), .ZN(n11465) );
  INV_X2 U11166 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n9587) );
  OAI22_X1 U11167 ( .A1(n9599), .A2(n9943), .B1(n9673), .B2(n9762), .ZN(n13694) );
  AND2_X1 U11168 ( .A1(n9792), .A2(n9791), .ZN(n16466) );
  NAND2_X1 U11169 ( .A1(n13584), .A2(n16196), .ZN(n16467) );
  NAND2_X1 U11170 ( .A1(n9799), .A2(n9593), .ZN(n16207) );
  NAND2_X1 U11171 ( .A1(n16141), .A2(n9617), .ZN(n16111) );
  OAI21_X1 U11172 ( .B1(n16141), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16123), .ZN(n16397) );
  AND2_X1 U11173 ( .A1(n10025), .A2(n10193), .ZN(n13680) );
  AND2_X1 U11174 ( .A1(n10103), .A2(n10101), .ZN(n15212) );
  AOI21_X1 U11175 ( .B1(n16382), .B2(n19962), .A(n10118), .ZN(n16383) );
  AND2_X1 U11176 ( .A1(n10194), .A2(n10192), .ZN(n14586) );
  XNOR2_X1 U11177 ( .A(n9759), .B(n9702), .ZN(n10064) );
  NAND2_X1 U11178 ( .A1(n9760), .A2(n16203), .ZN(n9759) );
  OAI21_X1 U11179 ( .B1(n10210), .B2(n10102), .A(n15353), .ZN(n10101) );
  INV_X1 U11180 ( .A(n10212), .ZN(n15237) );
  AND2_X1 U11181 ( .A1(n10096), .A2(n10094), .ZN(n15203) );
  NOR2_X1 U11182 ( .A1(n15210), .A2(n15211), .ZN(n10103) );
  NAND2_X1 U11183 ( .A1(n10012), .A2(n10011), .ZN(n16191) );
  AND2_X1 U11184 ( .A1(n9593), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9798) );
  OAI21_X1 U11185 ( .B1(n16241), .B2(n9590), .A(n10013), .ZN(n16205) );
  AND2_X1 U11186 ( .A1(n10301), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9934) );
  AOI21_X1 U11187 ( .B1(n13727), .B2(n13729), .A(n13728), .ZN(n15032) );
  AND2_X1 U11188 ( .A1(n10301), .A2(n10305), .ZN(n9593) );
  NOR2_X1 U11189 ( .A1(n13644), .A2(n13643), .ZN(n13647) );
  NOR2_X1 U11190 ( .A1(n10903), .A2(n10095), .ZN(n10094) );
  NOR2_X1 U11191 ( .A1(n15244), .A2(n10211), .ZN(n10096) );
  AOI21_X1 U11192 ( .B1(n14612), .B2(n16002), .A(n10425), .ZN(n14613) );
  NAND2_X1 U11193 ( .A1(n10037), .A2(n10394), .ZN(n10903) );
  AND2_X1 U11194 ( .A1(n13664), .A2(n12552), .ZN(n9826) );
  AND2_X1 U11195 ( .A1(n13580), .A2(n12526), .ZN(n13664) );
  AND2_X1 U11196 ( .A1(n13580), .A2(n16552), .ZN(n10301) );
  XNOR2_X1 U11197 ( .A(n13072), .B(n13071), .ZN(n14696) );
  AND2_X1 U11198 ( .A1(n9892), .A2(n9890), .ZN(n16331) );
  NAND2_X1 U11199 ( .A1(n9636), .A2(n9813), .ZN(n16248) );
  NAND2_X1 U11200 ( .A1(n12524), .A2(n9800), .ZN(n13580) );
  NAND2_X1 U11201 ( .A1(n13113), .A2(n12375), .ZN(n16360) );
  OAI21_X1 U11202 ( .B1(n15666), .B2(n15665), .A(n15664), .ZN(n16414) );
  XNOR2_X1 U11203 ( .A(n14539), .B(n14540), .ZN(n16392) );
  OR2_X1 U11204 ( .A1(n15625), .A2(n12374), .ZN(n12375) );
  AND2_X1 U11205 ( .A1(n15649), .A2(n9722), .ZN(n13681) );
  OR2_X1 U11206 ( .A1(n16833), .A2(n16834), .ZN(n20487) );
  NAND2_X1 U11207 ( .A1(n12670), .A2(n16275), .ZN(n9813) );
  AND2_X1 U11208 ( .A1(n18440), .A2(n18439), .ZN(n18441) );
  OR2_X1 U11209 ( .A1(n15625), .A2(n15624), .ZN(n16374) );
  AND2_X1 U11210 ( .A1(n10186), .A2(n10185), .ZN(n15869) );
  OR2_X1 U11211 ( .A1(n16635), .A2(n12546), .ZN(n12550) );
  OAI21_X1 U11212 ( .B1(n12768), .B2(n10213), .A(n10047), .ZN(n10046) );
  AOI21_X1 U11213 ( .B1(n10133), .B2(n10131), .A(n10130), .ZN(n10129) );
  AOI21_X1 U11214 ( .B1(n16278), .B2(n12682), .A(n12681), .ZN(n9772) );
  NAND2_X1 U11215 ( .A1(n9802), .A2(n12769), .ZN(n16315) );
  NAND2_X1 U11216 ( .A1(n12539), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16635) );
  NAND2_X1 U11217 ( .A1(n10017), .A2(n10183), .ZN(n10186) );
  AND2_X1 U11218 ( .A1(n17232), .A2(n10862), .ZN(n10205) );
  NAND2_X1 U11219 ( .A1(n16350), .A2(n12661), .ZN(n16628) );
  INV_X1 U11220 ( .A(n12542), .ZN(n9802) );
  AND2_X1 U11221 ( .A1(n12542), .A2(n12541), .ZN(n12547) );
  OAI21_X1 U11222 ( .B1(n10135), .B2(n10438), .A(n12749), .ZN(n10117) );
  XOR2_X1 U11223 ( .A(n12774), .B(n13085), .Z(n14692) );
  NAND2_X1 U11224 ( .A1(n12540), .A2(n12546), .ZN(n12542) );
  OR2_X1 U11225 ( .A1(n12540), .A2(n12546), .ZN(n12541) );
  OR2_X1 U11226 ( .A1(n16348), .A2(n12769), .ZN(n16350) );
  NAND2_X1 U11227 ( .A1(n10055), .A2(n10054), .ZN(n16876) );
  OAI21_X1 U11228 ( .B1(n11994), .B2(n15883), .A(n9697), .ZN(n10184) );
  AND2_X1 U11229 ( .A1(n13353), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9589) );
  NOR2_X1 U11230 ( .A1(n12773), .A2(n12772), .ZN(n13085) );
  AND2_X1 U11231 ( .A1(n15311), .A2(n15315), .ZN(n15285) );
  NAND2_X1 U11232 ( .A1(n11042), .A2(n11041), .ZN(n15100) );
  OAI211_X1 U11233 ( .C1(n9633), .C2(n10837), .A(n10199), .B(n10836), .ZN(
        n14468) );
  NAND2_X1 U11234 ( .A1(n14253), .A2(n10994), .ZN(n14450) );
  NOR2_X2 U11235 ( .A1(n20269), .A2(n16765), .ZN(n20378) );
  AND2_X1 U11236 ( .A1(n10271), .A2(n10269), .ZN(n10268) );
  AND2_X1 U11237 ( .A1(n18469), .A2(n13348), .ZN(n13349) );
  NOR2_X2 U11238 ( .A1(n20178), .A2(n20574), .ZN(n10443) );
  OR2_X1 U11239 ( .A1(n20049), .A2(n16765), .ZN(n16720) );
  OR2_X1 U11240 ( .A1(n12764), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16158) );
  NOR2_X2 U11241 ( .A1(n20574), .A2(n20049), .ZN(n20202) );
  NOR2_X2 U11242 ( .A1(n20178), .A2(n20308), .ZN(n20088) );
  AND2_X1 U11243 ( .A1(n12498), .A2(n12497), .ZN(n12614) );
  NAND2_X1 U11244 ( .A1(n16746), .A2(n16745), .ZN(n20269) );
  NAND2_X1 U11245 ( .A1(n10026), .A2(n9629), .ZN(n14369) );
  NOR2_X2 U11246 ( .A1(n20049), .A2(n20308), .ZN(n10452) );
  INV_X1 U11247 ( .A(n20582), .ZN(n16746) );
  NAND2_X1 U11248 ( .A1(n20582), .A2(n16745), .ZN(n20049) );
  NAND2_X1 U11249 ( .A1(n20582), .A2(n20601), .ZN(n20178) );
  INV_X1 U11250 ( .A(n18579), .ZN(n18559) );
  NAND2_X1 U11251 ( .A1(n21296), .A2(n21191), .ZN(n21401) );
  NAND2_X1 U11252 ( .A1(n21296), .A2(n21263), .ZN(n21335) );
  OAI21_X1 U11253 ( .B1(n19633), .B2(n12523), .A(n16481), .ZN(n16203) );
  NAND2_X1 U11254 ( .A1(n13347), .A2(n13342), .ZN(n18548) );
  AND2_X1 U11255 ( .A1(n13347), .A2(n9886), .ZN(n9885) );
  NAND2_X1 U11256 ( .A1(n10085), .A2(n10084), .ZN(n10788) );
  NOR2_X1 U11257 ( .A1(n12458), .A2(n12457), .ZN(n12466) );
  OR2_X1 U11258 ( .A1(n12442), .A2(n12443), .ZN(n10149) );
  AND2_X1 U11259 ( .A1(n19660), .A2(n12769), .ZN(n12731) );
  OR2_X1 U11260 ( .A1(n14233), .A2(n14234), .ZN(n14235) );
  OR2_X1 U11261 ( .A1(n20590), .A2(n19968), .ZN(n20574) );
  NAND2_X1 U11262 ( .A1(n13337), .A2(n10435), .ZN(n18568) );
  NAND2_X1 U11263 ( .A1(n20590), .A2(n19968), .ZN(n20246) );
  NOR2_X1 U11264 ( .A1(n20388), .A2(n12456), .ZN(n12457) );
  INV_X1 U11265 ( .A(n18432), .ZN(n18610) );
  OAI22_X1 U11266 ( .A1(n12414), .A2(n12515), .B1(n12502), .B2(n12413), .ZN(
        n12415) );
  OAI22_X1 U11267 ( .A1(n12421), .A2(n12516), .B1(n12501), .B2(n12420), .ZN(
        n12422) );
  AND2_X1 U11268 ( .A1(n12699), .A2(n12703), .ZN(n19660) );
  NAND2_X1 U11269 ( .A1(n20590), .A2(n16744), .ZN(n20308) );
  OR2_X1 U11270 ( .A1(n12419), .A2(n12412), .ZN(n12502) );
  INV_X1 U11271 ( .A(n18594), .ZN(n13337) );
  NAND2_X1 U11272 ( .A1(n9674), .A2(n12404), .ZN(n20388) );
  OR2_X1 U11273 ( .A1(n12419), .A2(n12417), .ZN(n12516) );
  OR2_X1 U11274 ( .A1(n12419), .A2(n12424), .ZN(n12515) );
  OAI21_X1 U11275 ( .B1(n16927), .B2(n18495), .A(n19180), .ZN(n18432) );
  OR2_X1 U11276 ( .A1(n12419), .A2(n12425), .ZN(n12501) );
  NAND2_X1 U11277 ( .A1(n10164), .A2(n9937), .ZN(n19973) );
  AND2_X1 U11278 ( .A1(n11761), .A2(n11780), .ZN(n14229) );
  OR2_X2 U11279 ( .A1(n12428), .A2(n12427), .ZN(n20216) );
  NAND2_X1 U11280 ( .A1(n13335), .A2(n9733), .ZN(n18594) );
  INV_X1 U11281 ( .A(n18672), .ZN(n13335) );
  NOR2_X2 U11282 ( .A1(n14031), .A2(n15135), .ZN(n13615) );
  NAND2_X1 U11283 ( .A1(n12698), .A2(n12721), .ZN(n13087) );
  NAND2_X1 U11284 ( .A1(n9876), .A2(n10753), .ZN(n14428) );
  NAND2_X1 U11285 ( .A1(n10976), .A2(n10979), .ZN(n14417) );
  OAI21_X2 U11286 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19567), .A(n17423), 
        .ZN(n18708) );
  NAND2_X1 U11287 ( .A1(n11736), .A2(n11735), .ZN(n12805) );
  NAND2_X1 U11288 ( .A1(n9986), .A2(n10694), .ZN(n10978) );
  NAND2_X1 U11289 ( .A1(n11769), .A2(n11768), .ZN(n16654) );
  AND2_X1 U11290 ( .A1(n13526), .A2(n13525), .ZN(n19409) );
  NOR2_X2 U11291 ( .A1(n19441), .A2(n13778), .ZN(n17807) );
  INV_X1 U11292 ( .A(n16652), .ZN(n13909) );
  AOI21_X1 U11293 ( .B1(n16665), .B2(n11776), .A(n11775), .ZN(n14011) );
  NAND2_X1 U11294 ( .A1(n10823), .A2(n9657), .ZN(n10695) );
  AND2_X1 U11295 ( .A1(n11762), .A2(n11767), .ZN(n16652) );
  NAND2_X1 U11296 ( .A1(n9818), .A2(n9853), .ZN(n20862) );
  NAND2_X1 U11297 ( .A1(n9925), .A2(n10659), .ZN(n10819) );
  AND2_X1 U11298 ( .A1(n14453), .A2(n14455), .ZN(n14454) );
  NOR2_X1 U11299 ( .A1(n15995), .A2(n14442), .ZN(n14453) );
  NAND2_X1 U11300 ( .A1(n13110), .A2(n13810), .ZN(n13163) );
  NOR2_X2 U11301 ( .A1(n19400), .A2(n18978), .ZN(n18882) );
  AND2_X1 U11302 ( .A1(n12785), .A2(n12784), .ZN(n15995) );
  AND2_X1 U11303 ( .A1(n12812), .A2(n12811), .ZN(n14376) );
  INV_X2 U11304 ( .A(n16002), .ZN(n9574) );
  AND2_X1 U11305 ( .A1(n12791), .A2(n12790), .ZN(n14442) );
  NAND2_X1 U11306 ( .A1(n16922), .A2(n9663), .ZN(n13287) );
  NAND2_X1 U11307 ( .A1(n11731), .A2(n11730), .ZN(n11734) );
  AOI21_X2 U11308 ( .B1(n16836), .B2(n14152), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n20397) );
  NAND2_X1 U11309 ( .A1(n10021), .A2(n10019), .ZN(n11772) );
  NAND2_X1 U11310 ( .A1(n11715), .A2(n11714), .ZN(n11763) );
  OR2_X2 U11311 ( .A1(n13330), .A2(n18302), .ZN(n18565) );
  NAND2_X1 U11312 ( .A1(n16920), .A2(n16919), .ZN(n16922) );
  AND2_X1 U11313 ( .A1(n11729), .A2(n11728), .ZN(n11732) );
  INV_X1 U11314 ( .A(n12783), .ZN(n12843) );
  NOR2_X1 U11315 ( .A1(n12238), .A2(n12237), .ZN(n15806) );
  NAND3_X1 U11316 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18180), .A3(n18159), .ZN(
        n18155) );
  NAND2_X1 U11317 ( .A1(n13094), .A2(n12134), .ZN(n9786) );
  AND2_X1 U11318 ( .A1(n14667), .A2(n9736), .ZN(n14675) );
  OR2_X1 U11319 ( .A1(n13305), .A2(n18305), .ZN(n13330) );
  NOR2_X1 U11320 ( .A1(n18424), .A2(n19570), .ZN(n18425) );
  OR2_X1 U11321 ( .A1(n13268), .A2(n13267), .ZN(n13269) );
  XNOR2_X1 U11322 ( .A(n13268), .B(n13266), .ZN(n16920) );
  AND2_X2 U11323 ( .A1(n17006), .A2(n17005), .ZN(n18180) );
  NAND2_X1 U11324 ( .A1(n17422), .A2(n14160), .ZN(n13770) );
  NAND2_X1 U11325 ( .A1(n14663), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14664) );
  AND2_X1 U11326 ( .A1(n9770), .A2(n9769), .ZN(n10399) );
  CLKBUF_X1 U11327 ( .A(n11724), .Z(n16694) );
  AND2_X1 U11328 ( .A1(n13132), .A2(n11709), .ZN(n10061) );
  INV_X1 U11329 ( .A(n17421), .ZN(n17413) );
  AND3_X1 U11330 ( .A1(n13025), .A2(n10603), .A3(n14140), .ZN(n12920) );
  NOR2_X1 U11331 ( .A1(n12645), .A2(n12649), .ZN(n12582) );
  NAND2_X1 U11332 ( .A1(n12577), .A2(n12576), .ZN(n12644) );
  NAND3_X1 U11333 ( .A1(n10292), .A2(n13127), .A3(n10293), .ZN(n16673) );
  NAND2_X1 U11334 ( .A1(n9810), .A2(n9809), .ZN(n13132) );
  OAI21_X1 U11335 ( .B1(n12373), .B2(n20509), .A(n12184), .ZN(n12200) );
  OR2_X1 U11336 ( .A1(n10320), .A2(n12591), .ZN(n10319) );
  OAI21_X1 U11337 ( .B1(n10618), .B2(n10584), .A(n13707), .ZN(n10597) );
  NAND3_X1 U11338 ( .A1(n10589), .A2(n10610), .A3(n13599), .ZN(n12904) );
  AND3_X1 U11339 ( .A1(n14205), .A2(n13475), .A3(n13483), .ZN(n14175) );
  CLKBUF_X1 U11340 ( .A(n12927), .Z(n14733) );
  OR2_X1 U11341 ( .A1(n12176), .A2(n12175), .ZN(n13893) );
  NAND2_X1 U11342 ( .A1(n12902), .A2(n10591), .ZN(n14576) );
  AND2_X1 U11343 ( .A1(n12927), .A2(n10595), .ZN(n13026) );
  AND2_X1 U11344 ( .A1(n11691), .A2(n11690), .ZN(n10292) );
  NOR2_X1 U11345 ( .A1(n12341), .A2(n12523), .ZN(n12310) );
  INV_X1 U11346 ( .A(n14137), .ZN(n21499) );
  AND2_X1 U11347 ( .A1(n10588), .A2(n10599), .ZN(n10610) );
  INV_X1 U11348 ( .A(n13474), .ZN(n19008) );
  CLKBUF_X1 U11349 ( .A(n12468), .Z(n12530) );
  NOR2_X2 U11350 ( .A1(n13460), .A2(n13459), .ZN(n14205) );
  AND2_X1 U11351 ( .A1(n12178), .A2(n11685), .ZN(n11693) );
  OAI211_X1 U11352 ( .C1(n9591), .C2(n9830), .A(n9829), .B(n9828), .ZN(n16936)
         );
  AND3_X2 U11353 ( .A1(n16735), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12445), 
        .ZN(n14368) );
  BUF_X2 U11354 ( .A(n12445), .Z(n15871) );
  NAND2_X1 U11355 ( .A1(n9637), .A2(n9832), .ZN(n14281) );
  INV_X2 U11356 ( .A(n12721), .ZN(n9575) );
  CLKBUF_X1 U11357 ( .A(n10586), .Z(n13599) );
  INV_X2 U11358 ( .A(n10607), .ZN(n14140) );
  NAND2_X1 U11359 ( .A1(n9591), .A2(n9833), .ZN(n13528) );
  OR2_X1 U11360 ( .A1(n13246), .A2(n13245), .ZN(n13535) );
  OR2_X1 U11361 ( .A1(n13472), .A2(n13471), .ZN(n19019) );
  INV_X2 U11362 ( .A(n14621), .ZN(n9576) );
  INV_X1 U11363 ( .A(n13123), .ZN(n19992) );
  AND4_X2 U11364 ( .A1(n13401), .A2(n13400), .A3(n13399), .A4(n13398), .ZN(
        n14214) );
  AND2_X1 U11365 ( .A1(n13208), .A2(n13205), .ZN(n9832) );
  AND4_X1 U11366 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12307) );
  INV_X2 U11367 ( .A(U212), .ZN(n17366) );
  OR2_X2 U11368 ( .A1(n17369), .A2(n17323), .ZN(n17371) );
  AND4_X1 U11369 ( .A1(n13393), .A2(n13392), .A3(n13391), .A4(n13390), .ZN(
        n13399) );
  CLKBUF_X1 U11370 ( .A(n11702), .Z(n20003) );
  NAND2_X1 U11371 ( .A1(n11646), .A2(n11645), .ZN(n13123) );
  AND2_X1 U11372 ( .A1(n10455), .A2(n10510), .ZN(n10594) );
  AND4_X1 U11373 ( .A1(n13369), .A2(n13368), .A3(n13367), .A4(n13366), .ZN(
        n13380) );
  AND4_X1 U11374 ( .A1(n12305), .A2(n12304), .A3(n12303), .A4(n12302), .ZN(
        n12306) );
  AND4_X1 U11375 ( .A1(n13191), .A2(n13190), .A3(n13189), .A4(n13188), .ZN(
        n13208) );
  AND4_X1 U11376 ( .A1(n13204), .A2(n13203), .A3(n13202), .A4(n13201), .ZN(
        n13205) );
  INV_X2 U11377 ( .A(n18067), .ZN(n18080) );
  INV_X2 U11378 ( .A(n13423), .ZN(n18102) );
  INV_X2 U11379 ( .A(n17112), .ZN(n17897) );
  AND3_X1 U11380 ( .A1(n10489), .A2(n10488), .A3(n10487), .ZN(n10490) );
  AND2_X1 U11381 ( .A1(n10516), .A2(n10515), .ZN(n10519) );
  AND4_X1 U11382 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10509) );
  BUF_X2 U11383 ( .A(n11846), .Z(n12268) );
  INV_X2 U11384 ( .A(n10718), .ZN(n10674) );
  NAND3_X1 U11385 ( .A1(n11609), .A2(n11607), .A3(n11608), .ZN(n9946) );
  NAND2_X1 U11386 ( .A1(n10298), .A2(n11678), .ZN(n9768) );
  OR2_X1 U11387 ( .A1(n19938), .A2(n15837), .ZN(n15814) );
  BUF_X2 U11388 ( .A(n10650), .Z(n10762) );
  INV_X1 U11389 ( .A(n13178), .ZN(n13423) );
  AND4_X1 U11390 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n11609) );
  BUF_X2 U11391 ( .A(n10527), .Z(n11529) );
  AND3_X1 U11392 ( .A1(n11662), .A2(n11661), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11665) );
  INV_X2 U11393 ( .A(n17996), .ZN(n18092) );
  BUF_X4 U11394 ( .A(n18126), .Z(n9580) );
  NAND2_X2 U11395 ( .A1(n20618), .A2(n20507), .ZN(n20562) );
  AND2_X2 U11396 ( .A1(n14597), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9586) );
  INV_X2 U11397 ( .A(n11544), .ZN(n9577) );
  CLKBUF_X1 U11398 ( .A(n11971), .Z(n14592) );
  INV_X2 U11399 ( .A(n17045), .ZN(n18131) );
  INV_X1 U11400 ( .A(n13412), .ZN(n18135) );
  NAND2_X1 U11401 ( .A1(n14389), .A2(n13182), .ZN(n18030) );
  AND2_X2 U11402 ( .A1(n11970), .A2(n11656), .ZN(n11808) );
  NAND2_X1 U11403 ( .A1(n13179), .A2(n13181), .ZN(n17087) );
  NAND2_X1 U11404 ( .A1(n13180), .A2(n13182), .ZN(n10442) );
  AND2_X2 U11405 ( .A1(n10469), .A2(n14409), .ZN(n10650) );
  AND2_X2 U11406 ( .A1(n10050), .A2(n13179), .ZN(n13168) );
  NAND2_X1 U11407 ( .A1(n13177), .A2(n13179), .ZN(n9620) );
  NAND2_X1 U11408 ( .A1(n10050), .A2(n13180), .ZN(n9626) );
  NAND2_X1 U11409 ( .A1(n13177), .A2(n14389), .ZN(n10448) );
  INV_X1 U11410 ( .A(n13200), .ZN(n17996) );
  INV_X2 U11411 ( .A(n17408), .ZN(n17410) );
  AND2_X1 U11412 ( .A1(n13177), .A2(n14215), .ZN(n13178) );
  NAND2_X1 U11413 ( .A1(n14635), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14634) );
  INV_X1 U11414 ( .A(n13172), .ZN(n13182) );
  AND2_X2 U11415 ( .A1(n13925), .A2(n14409), .ZN(n10627) );
  NOR2_X2 U11416 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13181) );
  NOR2_X2 U11417 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14215) );
  AND2_X2 U11418 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13925) );
  INV_X1 U11419 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16797) );
  AND2_X1 U11420 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14635) );
  INV_X2 U11421 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n11005) );
  INV_X1 U11422 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12102) );
  NAND2_X1 U11423 ( .A1(n10050), .A2(n14215), .ZN(n17045) );
  AND2_X1 U11424 ( .A1(n10050), .A2(n14389), .ZN(n18126) );
  OAI21_X2 U11425 ( .B1(n16159), .B2(n16138), .A(n16158), .ZN(n9811) );
  NAND2_X2 U11426 ( .A1(n10801), .A2(n10809), .ZN(n10975) );
  NAND2_X1 U11427 ( .A1(n14484), .A2(n14483), .ZN(n14482) );
  OAI21_X2 U11428 ( .B1(n18697), .B2(n10053), .A(n10052), .ZN(n10051) );
  AND2_X2 U11429 ( .A1(n10097), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9579) );
  INV_X1 U11430 ( .A(n11738), .ZN(n13070) );
  AND3_X1 U11431 ( .A1(n12196), .A2(n12179), .A3(n9575), .ZN(n12215) );
  MUX2_X2 U11432 ( .A(n12581), .B(n12580), .S(n9575), .Z(n12649) );
  NAND2_X2 U11433 ( .A1(n18882), .A2(n18926), .ZN(n18836) );
  NAND2_X1 U11434 ( .A1(n19024), .A2(n19008), .ZN(n14096) );
  OAI21_X1 U11435 ( .B1(n9860), .B2(n16409), .A(n9672), .ZN(n10008) );
  AND2_X1 U11436 ( .A1(n9779), .A2(n13095), .ZN(n11716) );
  OR2_X1 U11437 ( .A1(n12426), .A2(n16665), .ZN(n12427) );
  BUF_X4 U11438 ( .A(n12396), .Z(n12426) );
  NOR2_X1 U11439 ( .A1(n20240), .A2(n12399), .ZN(n9949) );
  AND2_X1 U11440 ( .A1(n19997), .A2(n19992), .ZN(n13127) );
  NAND2_X2 U11441 ( .A1(n12725), .A2(n12724), .ZN(n19633) );
  NOR2_X1 U11442 ( .A1(n16187), .A2(n16186), .ZN(n16185) );
  OAI21_X1 U11443 ( .B1(n10006), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n19918), .ZN(n9931) );
  NAND2_X2 U11444 ( .A1(n15763), .A2(n15938), .ZN(n15932) );
  NOR2_X4 U11445 ( .A1(n15762), .A2(n15764), .ZN(n15763) );
  NOR3_X2 U11446 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17792) );
  AND2_X1 U11447 ( .A1(n13678), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9582) );
  AND2_X4 U11448 ( .A1(n13678), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9583) );
  AND3_X1 U11449 ( .A1(n16656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9584) );
  AND3_X2 U11450 ( .A1(n16656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9585) );
  INV_X4 U11451 ( .A(n12721), .ZN(n12693) );
  INV_X2 U11452 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16837) );
  AND2_X4 U11453 ( .A1(n13678), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12879) );
  INV_X2 U11454 ( .A(n13139), .ZN(n13678) );
  AND2_X1 U11455 ( .A1(n18470), .A2(n13352), .ZN(n13353) );
  AND2_X1 U11456 ( .A1(n10890), .A2(n9634), .ZN(n9859) );
  INV_X1 U11457 ( .A(n12792), .ZN(n10346) );
  NAND2_X1 U11458 ( .A1(n16147), .A2(n16158), .ZN(n12765) );
  INV_X2 U11459 ( .A(n17045), .ZN(n18081) );
  NAND2_X2 U11460 ( .A1(n17119), .A2(n14362), .ZN(n18086) );
  INV_X1 U11461 ( .A(n18379), .ZN(n17422) );
  NAND2_X1 U11462 ( .A1(n10212), .A2(n10146), .ZN(n10145) );
  INV_X1 U11463 ( .A(n15211), .ZN(n10146) );
  INV_X1 U11464 ( .A(n12545), .ZN(n10302) );
  OAI21_X1 U11465 ( .B1(n16315), .B2(n16593), .A(n12544), .ZN(n12545) );
  AOI21_X1 U11466 ( .B1(n10013), .B2(n9590), .A(n13649), .ZN(n10011) );
  NOR2_X1 U11467 ( .A1(n19008), .A2(n19004), .ZN(n14173) );
  NAND2_X1 U11468 ( .A1(n10916), .A2(n10587), .ZN(n10588) );
  NAND2_X1 U11469 ( .A1(n14236), .A2(n10347), .ZN(n10351) );
  NOR2_X1 U11470 ( .A1(n10348), .A2(n19945), .ZN(n10347) );
  NAND2_X1 U11471 ( .A1(n12411), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10348) );
  OAI21_X1 U11472 ( .B1(n10986), .B2(n10092), .A(n9658), .ZN(n10823) );
  INV_X1 U11473 ( .A(n10659), .ZN(n10092) );
  NAND2_X1 U11474 ( .A1(n10659), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U11475 ( .A1(n10609), .A2(n10790), .ZN(n10585) );
  AND2_X2 U11476 ( .A1(n10948), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10469) );
  AND2_X2 U11477 ( .A1(n9923), .A2(n10136), .ZN(n10576) );
  OR2_X1 U11478 ( .A1(n20833), .A2(n10276), .ZN(n10736) );
  AND3_X1 U11479 ( .A1(n14511), .A2(n20833), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10956) );
  INV_X1 U11480 ( .A(n10128), .ZN(n10107) );
  NAND2_X1 U11481 ( .A1(n10163), .A2(n12426), .ZN(n12419) );
  NAND2_X1 U11482 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10355) );
  AND2_X1 U11483 ( .A1(n13749), .A2(n10290), .ZN(n10289) );
  NOR2_X1 U11484 ( .A1(n14746), .A2(n14757), .ZN(n10290) );
  OR2_X1 U11485 ( .A1(n10325), .A2(n10324), .ZN(n10323) );
  INV_X1 U11486 ( .A(n14898), .ZN(n10324) );
  INV_X1 U11487 ( .A(n15285), .ZN(n10081) );
  NOR2_X1 U11488 ( .A1(n9985), .A2(n9984), .ZN(n10892) );
  INV_X1 U11489 ( .A(n15298), .ZN(n9984) );
  NAND2_X1 U11490 ( .A1(n15304), .A2(n10883), .ZN(n15286) );
  NAND2_X1 U11491 ( .A1(n10143), .A2(n9604), .ZN(n10868) );
  NAND2_X1 U11492 ( .A1(n9822), .A2(n10088), .ZN(n11591) );
  INV_X1 U11493 ( .A(n10089), .ZN(n10088) );
  NAND2_X1 U11494 ( .A1(n17240), .A2(n10205), .ZN(n9822) );
  OAI21_X1 U11495 ( .B1(n10864), .B2(n10090), .A(n17231), .ZN(n10089) );
  OR2_X1 U11496 ( .A1(n10657), .A2(n10656), .ZN(n10820) );
  OR2_X1 U11497 ( .A1(n10641), .A2(n10640), .ZN(n10875) );
  INV_X1 U11498 ( .A(n10956), .ZN(n10936) );
  AND2_X1 U11499 ( .A1(n10691), .A2(n10692), .ZN(n10702) );
  INV_X1 U11500 ( .A(n10953), .ZN(n10964) );
  INV_X1 U11501 ( .A(n11723), .ZN(n12779) );
  INV_X1 U11502 ( .A(n13588), .ZN(n12853) );
  INV_X1 U11503 ( .A(n14585), .ZN(n10191) );
  AND2_X1 U11504 ( .A1(n9936), .A2(n9935), .ZN(n12153) );
  INV_X1 U11505 ( .A(n15934), .ZN(n12838) );
  AND2_X1 U11506 ( .A1(n9696), .A2(n10421), .ZN(n10420) );
  INV_X1 U11507 ( .A(n15630), .ZN(n10421) );
  NAND2_X1 U11508 ( .A1(n12758), .A2(n12757), .ZN(n16113) );
  AND2_X1 U11509 ( .A1(n15692), .A2(n12769), .ZN(n12764) );
  NOR2_X1 U11510 ( .A1(n9660), .A2(n10417), .ZN(n10416) );
  INV_X1 U11511 ( .A(n15696), .ZN(n10417) );
  INV_X1 U11512 ( .A(n13978), .ZN(n10375) );
  INV_X1 U11513 ( .A(n13884), .ZN(n12315) );
  AOI21_X1 U11514 ( .B1(n12122), .B2(n12120), .A(n12119), .ZN(n12126) );
  NAND2_X1 U11515 ( .A1(n16853), .A2(n16852), .ZN(n16855) );
  NAND2_X1 U11516 ( .A1(n14188), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10267) );
  NAND2_X1 U11517 ( .A1(n15001), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15004) );
  AND2_X1 U11518 ( .A1(n15001), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13730) );
  NOR2_X1 U11519 ( .A1(n15004), .A2(n13707), .ZN(n13716) );
  XNOR2_X1 U11520 ( .A(n11580), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13731) );
  OR2_X1 U11521 ( .A1(n11579), .A2(n11578), .ZN(n11580) );
  INV_X1 U11522 ( .A(n14771), .ZN(n11460) );
  NAND2_X1 U11523 ( .A1(n10145), .A2(n13623), .ZN(n10144) );
  NOR2_X1 U11524 ( .A1(n9753), .A2(n9752), .ZN(n15389) );
  INV_X1 U11525 ( .A(n13052), .ZN(n9752) );
  NAND2_X1 U11526 ( .A1(n15340), .A2(n10079), .ZN(n10078) );
  AOI21_X1 U11527 ( .B1(n10079), .B2(n9592), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10077) );
  NAND2_X1 U11528 ( .A1(n15555), .A2(n15537), .ZN(n15580) );
  NAND2_X1 U11529 ( .A1(n12919), .A2(n12918), .ZN(n13044) );
  CLKBUF_X1 U11530 ( .A(n12920), .Z(n12921) );
  CLKBUF_X1 U11531 ( .A(n12148), .Z(n12149) );
  NAND2_X1 U11532 ( .A1(n12688), .A2(n9709), .ZN(n12762) );
  OR2_X1 U11533 ( .A1(n10319), .A2(n12693), .ZN(n10318) );
  NAND2_X1 U11534 ( .A1(n16084), .A2(n10374), .ZN(n10372) );
  NAND2_X1 U11535 ( .A1(n12885), .A2(n10339), .ZN(n12886) );
  NAND2_X1 U11536 ( .A1(n10346), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10339) );
  NAND2_X1 U11537 ( .A1(n9588), .A2(n10117), .ZN(n9774) );
  NAND2_X1 U11538 ( .A1(n16576), .A2(n13147), .ZN(n16421) );
  NAND2_X2 U11539 ( .A1(n9758), .A2(n10253), .ZN(n16241) );
  NAND2_X1 U11540 ( .A1(n16262), .A2(n10255), .ZN(n9758) );
  INV_X1 U11541 ( .A(n16250), .ZN(n10254) );
  INV_X1 U11542 ( .A(n13163), .ZN(n13141) );
  INV_X1 U11543 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20392) );
  AND2_X1 U11544 ( .A1(n13520), .A2(n13519), .ZN(n19404) );
  INV_X1 U11545 ( .A(n18264), .ZN(n9965) );
  NAND2_X1 U11546 ( .A1(n13354), .A2(n18659), .ZN(n16960) );
  NAND4_X1 U11547 ( .A1(n13329), .A2(n13328), .A3(n13327), .A4(n13326), .ZN(
        n17130) );
  AND4_X1 U11548 ( .A1(n13312), .A2(n13311), .A3(n13310), .A4(n13309), .ZN(
        n13329) );
  AND4_X1 U11549 ( .A1(n13321), .A2(n13320), .A3(n13319), .A4(n13318), .ZN(
        n13327) );
  NAND2_X1 U11550 ( .A1(n13356), .A2(n13355), .ZN(n18446) );
  NAND2_X1 U11551 ( .A1(n9589), .A2(n16876), .ZN(n13354) );
  NAND2_X1 U11552 ( .A1(n13341), .A2(n10157), .ZN(n10156) );
  NAND2_X1 U11553 ( .A1(n9841), .A2(n10155), .ZN(n9840) );
  AND2_X1 U11554 ( .A1(n16961), .A2(n18302), .ZN(n18878) );
  INV_X1 U11555 ( .A(n19004), .ZN(n14104) );
  NAND2_X1 U11556 ( .A1(n13473), .A2(n14204), .ZN(n9982) );
  INV_X1 U11557 ( .A(n13770), .ZN(n9983) );
  AND2_X1 U11558 ( .A1(n19024), .A2(n14208), .ZN(n13473) );
  INV_X1 U11559 ( .A(n20807), .ZN(n20795) );
  INV_X1 U11560 ( .A(n20488), .ZN(n19771) );
  AND2_X1 U11561 ( .A1(n12526), .A2(n9737), .ZN(n10168) );
  NAND3_X1 U11562 ( .A1(n12521), .A2(n12506), .A3(n12518), .ZN(n10113) );
  NAND2_X1 U11563 ( .A1(n9898), .A2(n9896), .ZN(n12615) );
  NOR2_X1 U11564 ( .A1(n12769), .A2(n9897), .ZN(n9896) );
  INV_X1 U11565 ( .A(n12522), .ZN(n9897) );
  NAND2_X1 U11566 ( .A1(n9628), .A2(n9939), .ZN(n9938) );
  NAND2_X1 U11567 ( .A1(n9951), .A2(n9950), .ZN(n9948) );
  NAND2_X1 U11568 ( .A1(n12402), .A2(n9602), .ZN(n9950) );
  AND2_X2 U11569 ( .A1(n16657), .A2(n16797), .ZN(n11610) );
  NAND2_X1 U11570 ( .A1(n10947), .A2(n10946), .ZN(n10952) );
  XNOR2_X1 U11571 ( .A(n10948), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10951) );
  AND2_X1 U11572 ( .A1(n14428), .A2(n10795), .ZN(n10084) );
  INV_X1 U11573 ( .A(n10801), .ZN(n10085) );
  NAND2_X1 U11574 ( .A1(n15353), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10394) );
  NAND2_X1 U11575 ( .A1(n10995), .A2(n14078), .ZN(n9819) );
  AND2_X1 U11576 ( .A1(n10277), .A2(n10276), .ZN(n10275) );
  NAND2_X1 U11577 ( .A1(n10626), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10515) );
  AOI22_X1 U11578 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10577), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10523) );
  OR2_X1 U11579 ( .A1(n10752), .A2(n10751), .ZN(n10802) );
  NAND2_X1 U11580 ( .A1(n9874), .A2(n9871), .ZN(n9870) );
  NOR2_X1 U11581 ( .A1(n10279), .A2(n9872), .ZN(n9871) );
  INV_X1 U11582 ( .A(n10437), .ZN(n10308) );
  INV_X1 U11583 ( .A(n15883), .ZN(n10018) );
  INV_X1 U11584 ( .A(n10336), .ZN(n10335) );
  OAI21_X1 U11585 ( .B1(n12792), .B2(n20542), .A(n12858), .ZN(n10336) );
  OR2_X1 U11586 ( .A1(n14561), .A2(n10262), .ZN(n10261) );
  INV_X1 U11587 ( .A(n13575), .ZN(n10262) );
  AND2_X1 U11588 ( .A1(n12498), .A2(n9721), .ZN(n10086) );
  NAND2_X1 U11589 ( .A1(n10352), .A2(n10351), .ZN(n12433) );
  NAND2_X1 U11590 ( .A1(n12138), .A2(n16815), .ZN(n11708) );
  NAND2_X1 U11591 ( .A1(n16816), .A2(n9780), .ZN(n9779) );
  AOI21_X1 U11592 ( .B1(n16694), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10020), 
        .ZN(n10019) );
  AND2_X1 U11593 ( .A1(n16830), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10020) );
  INV_X1 U11594 ( .A(n12397), .ZN(n10300) );
  NAND2_X1 U11595 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n9973) );
  INV_X1 U11596 ( .A(n13415), .ZN(n9976) );
  AOI21_X1 U11597 ( .B1(n9573), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(n9975), .ZN(n9974) );
  NOR2_X1 U11598 ( .A1(n18030), .A2(n13410), .ZN(n9975) );
  NOR2_X1 U11599 ( .A1(n14922), .A2(n9927), .ZN(n11599) );
  NAND2_X1 U11600 ( .A1(n9928), .A2(n10424), .ZN(n9927) );
  INV_X1 U11601 ( .A(n14912), .ZN(n9928) );
  NOR2_X1 U11602 ( .A1(n11079), .A2(n21565), .ZN(n11101) );
  NOR2_X1 U11603 ( .A1(n14498), .A2(n14497), .ZN(n10283) );
  NAND2_X1 U11604 ( .A1(n10609), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11196) );
  AND2_X1 U11605 ( .A1(n10601), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11002) );
  OR2_X1 U11606 ( .A1(n10599), .A2(n11005), .ZN(n11537) );
  NAND2_X1 U11607 ( .A1(n15281), .A2(n9596), .ZN(n10037) );
  INV_X1 U11608 ( .A(n14865), .ZN(n10317) );
  NAND2_X1 U11609 ( .A1(n10326), .A2(n12986), .ZN(n10325) );
  INV_X1 U11610 ( .A(n15052), .ZN(n10326) );
  NAND2_X1 U11611 ( .A1(n10868), .A2(n10876), .ZN(n10881) );
  NAND2_X1 U11612 ( .A1(n12968), .A2(n10313), .ZN(n10312) );
  INV_X1 U11613 ( .A(n15073), .ZN(n10313) );
  NAND2_X1 U11614 ( .A1(n14731), .A2(n12941), .ZN(n13020) );
  INV_X1 U11615 ( .A(n14962), .ZN(n12968) );
  INV_X1 U11616 ( .A(n10886), .ZN(n10901) );
  AOI21_X1 U11617 ( .B1(n11028), .B2(n14078), .A(n10872), .ZN(n10873) );
  NAND2_X1 U11618 ( .A1(n10093), .A2(n10861), .ZN(n10863) );
  INV_X1 U11619 ( .A(n14479), .ZN(n12954) );
  INV_X1 U11620 ( .A(n14464), .ZN(n12955) );
  INV_X1 U11621 ( .A(n13020), .ZN(n12995) );
  NOR2_X1 U11622 ( .A1(n20833), .A2(n10587), .ZN(n10600) );
  INV_X1 U11623 ( .A(n10662), .ZN(n10209) );
  INV_X1 U11624 ( .A(n10684), .ZN(n10392) );
  NAND2_X1 U11625 ( .A1(n9875), .A2(n9872), .ZN(n9874) );
  INV_X1 U11626 ( .A(n10277), .ZN(n9875) );
  NAND2_X1 U11627 ( .A1(n10704), .A2(n10278), .ZN(n10277) );
  INV_X1 U11628 ( .A(n10708), .ZN(n10278) );
  AND4_X1 U11629 ( .A1(n10509), .A2(n10508), .A3(n10507), .A4(n10506), .ZN(
        n10510) );
  AND4_X1 U11630 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10456) );
  INV_X1 U11631 ( .A(n14504), .ZN(n21292) );
  OAI21_X1 U11632 ( .B1(n17172), .B2(n17280), .A(n14578), .ZN(n14510) );
  NAND2_X1 U11633 ( .A1(n12600), .A2(n9725), .ZN(n12773) );
  NAND2_X1 U11634 ( .A1(n10039), .A2(n12565), .ZN(n12575) );
  NAND2_X1 U11635 ( .A1(n12563), .A2(n9576), .ZN(n10039) );
  INV_X1 U11636 ( .A(n10334), .ZN(n10333) );
  OAI21_X1 U11637 ( .B1(n12792), .B2(n20533), .A(n12839), .ZN(n10334) );
  CLKBUF_X1 U11638 ( .A(n11977), .Z(n14593) );
  NAND2_X1 U11639 ( .A1(n14369), .A2(n9715), .ZN(n11992) );
  NAND2_X1 U11640 ( .A1(n10346), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U11641 ( .A1(n12838), .A2(n10412), .ZN(n10411) );
  INV_X1 U11642 ( .A(n15928), .ZN(n10412) );
  INV_X1 U11643 ( .A(n15778), .ZN(n10406) );
  NAND2_X1 U11644 ( .A1(n16127), .A2(n16377), .ZN(n16115) );
  NAND2_X1 U11645 ( .A1(n10346), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10344) );
  AND4_X1 U11646 ( .A1(n12287), .A2(n12286), .A3(n12285), .A4(n12284), .ZN(
        n12309) );
  AND4_X1 U11647 ( .A1(n12294), .A2(n12293), .A3(n12292), .A4(n12291), .ZN(
        n12308) );
  NAND2_X1 U11648 ( .A1(n16147), .A2(n16158), .ZN(n10179) );
  NAND2_X1 U11649 ( .A1(n12362), .A2(n10382), .ZN(n10381) );
  INV_X1 U11650 ( .A(n15685), .ZN(n10382) );
  NAND2_X1 U11651 ( .A1(n10134), .A2(n10132), .ZN(n10133) );
  INV_X1 U11652 ( .A(n10135), .ZN(n10134) );
  NOR2_X1 U11653 ( .A1(n10132), .A2(n16136), .ZN(n10131) );
  NAND2_X1 U11654 ( .A1(n10346), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10343) );
  INV_X1 U11655 ( .A(n13668), .ZN(n10418) );
  OR2_X1 U11656 ( .A1(n15717), .A2(n12523), .ZN(n12753) );
  NOR2_X1 U11657 ( .A1(n10264), .A2(n16223), .ZN(n10263) );
  INV_X1 U11658 ( .A(n16231), .ZN(n10264) );
  NAND2_X1 U11659 ( .A1(n10386), .A2(n14224), .ZN(n10385) );
  INV_X1 U11660 ( .A(n16264), .ZN(n9812) );
  NAND2_X1 U11661 ( .A1(n12542), .A2(n12523), .ZN(n16314) );
  NOR2_X1 U11662 ( .A1(n9893), .A2(n9891), .ZN(n9890) );
  INV_X1 U11663 ( .A(n16328), .ZN(n9891) );
  INV_X1 U11664 ( .A(n12527), .ZN(n10066) );
  INV_X1 U11665 ( .A(n12528), .ZN(n10065) );
  NOR2_X1 U11666 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  NOR2_X1 U11667 ( .A1(n12779), .A2(n20513), .ZN(n11741) );
  NAND2_X1 U11668 ( .A1(n14236), .A2(n9652), .ZN(n12499) );
  INV_X1 U11669 ( .A(n12502), .ZN(n20115) );
  INV_X1 U11670 ( .A(n12501), .ZN(n20179) );
  INV_X1 U11671 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16748) );
  NAND2_X1 U11672 ( .A1(n11790), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10181) );
  NAND2_X1 U11673 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10182) );
  NAND2_X1 U11674 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10354) );
  AOI21_X1 U11675 ( .B1(n11790), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n11656), .ZN(n10353) );
  NAND2_X1 U11676 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10356) );
  INV_X1 U11677 ( .A(n11685), .ZN(n11713) );
  NAND2_X1 U11678 ( .A1(n12402), .A2(n12426), .ZN(n16778) );
  AND2_X1 U11679 ( .A1(n12152), .A2(n12572), .ZN(n13786) );
  OR2_X1 U11680 ( .A1(n12569), .A2(n12151), .ZN(n12152) );
  XNOR2_X1 U11681 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12120) );
  NAND2_X1 U11682 ( .A1(n12118), .A2(n12117), .ZN(n12122) );
  NOR2_X1 U11683 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16830) );
  INV_X1 U11684 ( .A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17917) );
  NOR2_X1 U11685 ( .A1(n16848), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10161) );
  NAND2_X1 U11686 ( .A1(n13289), .A2(n18308), .ZN(n13305) );
  NOR2_X1 U11687 ( .A1(n13533), .A2(n18317), .ZN(n13529) );
  NOR2_X1 U11688 ( .A1(n13488), .A2(n13487), .ZN(n13489) );
  OR3_X1 U11689 ( .A1(n13486), .A2(n13485), .A3(n13484), .ZN(n13487) );
  AOI22_X1 U11690 ( .A1(n13178), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13185) );
  NOR2_X1 U11691 ( .A1(n13481), .A2(n18186), .ZN(n13483) );
  NAND2_X1 U11692 ( .A1(n20624), .A2(n10276), .ZN(n11584) );
  INV_X1 U11693 ( .A(n11392), .ZN(n11306) );
  NAND2_X1 U11694 ( .A1(n11306), .A2(n9907), .ZN(n11434) );
  NOR2_X1 U11695 ( .A1(n11371), .A2(n9908), .ZN(n9907) );
  NOR2_X1 U11696 ( .A1(n13040), .A2(n13041), .ZN(n14036) );
  AND2_X1 U11697 ( .A1(n13922), .A2(n13598), .ZN(n13937) );
  INV_X1 U11698 ( .A(n15135), .ZN(n14509) );
  INV_X1 U11699 ( .A(n11537), .ZN(n11575) );
  AND2_X1 U11700 ( .A1(n11489), .A2(n9688), .ZN(n13728) );
  INV_X1 U11701 ( .A(n13729), .ZN(n10288) );
  INV_X1 U11702 ( .A(n11490), .ZN(n11491) );
  NAND2_X1 U11703 ( .A1(n11491), .A2(n9913), .ZN(n11542) );
  NOR2_X1 U11704 ( .A1(n11492), .A2(n14763), .ZN(n9913) );
  AND2_X1 U11705 ( .A1(n11489), .A2(n10290), .ZN(n14745) );
  NAND2_X1 U11706 ( .A1(n11489), .A2(n11488), .ZN(n14755) );
  OR2_X1 U11707 ( .A1(n11436), .A2(n11435), .ZN(n11490) );
  AND2_X1 U11708 ( .A1(n11433), .A2(n9704), .ZN(n10285) );
  NAND2_X1 U11709 ( .A1(n11285), .A2(n9910), .ZN(n11390) );
  NOR2_X1 U11710 ( .A1(n9912), .A2(n9911), .ZN(n9910) );
  OR2_X1 U11711 ( .A1(n11390), .A2(n11389), .ZN(n11392) );
  NAND2_X1 U11712 ( .A1(n11285), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11412) );
  OR2_X1 U11713 ( .A1(n11136), .A2(n11138), .ZN(n11161) );
  OR2_X1 U11714 ( .A1(n15092), .A2(n15091), .ZN(n15094) );
  NAND2_X1 U11715 ( .A1(n14815), .A2(n9714), .ZN(n14758) );
  INV_X1 U11716 ( .A(n14760), .ZN(n10327) );
  OAI21_X1 U11717 ( .B1(n10035), .B2(n13015), .A(n10034), .ZN(n10905) );
  NAND2_X1 U11718 ( .A1(n15281), .A2(n9606), .ZN(n10034) );
  NAND2_X1 U11719 ( .A1(n14815), .A2(n9693), .ZN(n14772) );
  NAND2_X1 U11720 ( .A1(n14815), .A2(n9692), .ZN(n14793) );
  AND2_X1 U11721 ( .A1(n14815), .A2(n14798), .ZN(n14800) );
  AND2_X1 U11722 ( .A1(n13007), .A2(n13006), .ZN(n14816) );
  NOR2_X1 U11723 ( .A1(n10141), .A2(n10139), .ZN(n10902) );
  NAND2_X1 U11724 ( .A1(n10895), .A2(n10140), .ZN(n10139) );
  INV_X1 U11725 ( .A(n10142), .ZN(n10141) );
  INV_X1 U11726 ( .A(n14852), .ZN(n10315) );
  AND2_X1 U11727 ( .A1(n13049), .A2(n15521), .ZN(n15454) );
  INV_X1 U11728 ( .A(n10080), .ZN(n10079) );
  OAI21_X1 U11729 ( .B1(n10082), .B2(n9592), .A(n9671), .ZN(n10080) );
  OR2_X1 U11730 ( .A1(n15340), .A2(n9592), .ZN(n10076) );
  OAI21_X1 U11731 ( .B1(n15341), .B2(n15286), .A(n15285), .ZN(n15296) );
  NAND2_X1 U11732 ( .A1(n10881), .A2(n15531), .ZN(n15316) );
  NAND2_X1 U11733 ( .A1(n10868), .A2(n9712), .ZN(n15302) );
  INV_X1 U11734 ( .A(n10863), .ZN(n17238) );
  NAND2_X1 U11735 ( .A1(n14467), .A2(n10839), .ZN(n17240) );
  OR2_X1 U11736 ( .A1(n11584), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15360) );
  AND2_X1 U11737 ( .A1(n13044), .A2(n17140), .ZN(n14130) );
  AND2_X1 U11738 ( .A1(n13044), .A2(n13036), .ZN(n15428) );
  AND2_X1 U11739 ( .A1(n13044), .A2(n14036), .ZN(n20805) );
  OAI211_X1 U11740 ( .C1(n10936), .C2(n14519), .A(n10661), .B(n10660), .ZN(
        n10984) );
  NAND2_X1 U11741 ( .A1(n10986), .A2(n10276), .ZN(n9925) );
  INV_X1 U11742 ( .A(n10702), .ZN(n9853) );
  INV_X1 U11743 ( .A(n20931), .ZN(n9818) );
  AND2_X1 U11744 ( .A1(n13025), .A2(n10603), .ZN(n12901) );
  INV_X1 U11745 ( .A(n20626), .ZN(n14043) );
  OR2_X1 U11746 ( .A1(n14501), .A2(n14500), .ZN(n20930) );
  INV_X1 U11747 ( .A(n20930), .ZN(n20926) );
  INV_X1 U11748 ( .A(n21064), .ZN(n21059) );
  NOR2_X1 U11749 ( .A1(n14417), .A2(n14502), .ZN(n21215) );
  AND2_X1 U11750 ( .A1(n14417), .A2(n14502), .ZN(n21191) );
  AOI21_X1 U11751 ( .B1(n21264), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20973), 
        .ZN(n21348) );
  NAND2_X1 U11752 ( .A1(n9751), .A2(n10965), .ZN(n9750) );
  INV_X1 U11753 ( .A(n16830), .ZN(n15612) );
  NOR2_X1 U11754 ( .A1(n12598), .A2(n10041), .ZN(n10040) );
  NAND2_X1 U11755 ( .A1(n12624), .A2(n15973), .ZN(n12632) );
  INV_X1 U11756 ( .A(n12644), .ZN(n12583) );
  INV_X1 U11757 ( .A(n15826), .ZN(n15855) );
  NAND2_X1 U11758 ( .A1(n13786), .A2(n13810), .ZN(n13795) );
  NAND2_X1 U11759 ( .A1(n11763), .A2(n11764), .ZN(n11762) );
  AND2_X1 U11760 ( .A1(n12857), .A2(n9707), .ZN(n15741) );
  NAND2_X1 U11761 ( .A1(n12845), .A2(n9646), .ZN(n14569) );
  AND2_X1 U11762 ( .A1(n10031), .A2(n10191), .ZN(n10190) );
  INV_X1 U11763 ( .A(n10192), .ZN(n10188) );
  NAND2_X1 U11764 ( .A1(n15625), .A2(n12374), .ZN(n13113) );
  NAND2_X1 U11765 ( .A1(n10194), .A2(n10196), .ZN(n10025) );
  NAND2_X1 U11766 ( .A1(n14528), .A2(n14527), .ZN(n14526) );
  INV_X1 U11767 ( .A(n15889), .ZN(n11993) );
  NAND2_X1 U11768 ( .A1(n11619), .A2(n11656), .ZN(n11626) );
  NAND2_X1 U11769 ( .A1(n9786), .A2(n15871), .ZN(n19836) );
  NAND2_X1 U11770 ( .A1(n10346), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U11771 ( .A1(n12889), .A2(n9732), .ZN(n13067) );
  AND2_X1 U11772 ( .A1(n14624), .A2(n9705), .ZN(n14660) );
  NAND2_X1 U11773 ( .A1(n14624), .A2(n10247), .ZN(n14659) );
  AND2_X1 U11774 ( .A1(n12837), .A2(n9643), .ZN(n15934) );
  INV_X1 U11775 ( .A(n12766), .ZN(n10213) );
  INV_X1 U11776 ( .A(n13682), .ZN(n10419) );
  INV_X1 U11777 ( .A(n16115), .ZN(n10121) );
  AND2_X1 U11778 ( .A1(n12869), .A2(n12868), .ZN(n15681) );
  OAI211_X1 U11779 ( .C1(n12792), .C2(n20548), .A(n12866), .B(n12865), .ZN(
        n12867) );
  NAND2_X1 U11780 ( .A1(n9922), .A2(n9921), .ZN(n16168) );
  NOR2_X1 U11781 ( .A1(n16186), .A2(n21554), .ZN(n9921) );
  INV_X1 U11782 ( .A(n10263), .ZN(n9994) );
  INV_X1 U11783 ( .A(n14554), .ZN(n13143) );
  AND2_X1 U11784 ( .A1(n10305), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10304) );
  NAND2_X1 U11785 ( .A1(n9761), .A2(n10301), .ZN(n16284) );
  NAND2_X1 U11786 ( .A1(n16241), .A2(n16239), .ZN(n9997) );
  AND2_X1 U11787 ( .A1(n12321), .A2(n12315), .ZN(n10376) );
  AND3_X1 U11788 ( .A1(n12324), .A2(n12323), .A3(n12322), .ZN(n13978) );
  INV_X1 U11789 ( .A(n10370), .ZN(n10369) );
  OAI21_X1 U11790 ( .B1(n9625), .B2(n12310), .A(n13887), .ZN(n10370) );
  NAND2_X1 U11791 ( .A1(n16276), .A2(n16343), .ZN(n9892) );
  NAND2_X1 U11792 ( .A1(n12589), .A2(n12231), .ZN(n10374) );
  AND3_X1 U11793 ( .A1(n12267), .A2(n12266), .A3(n12265), .ZN(n16084) );
  NOR2_X1 U11794 ( .A1(n13099), .A2(n12147), .ZN(n16798) );
  AND2_X1 U11795 ( .A1(n13138), .A2(n13137), .ZN(n16649) );
  NAND2_X1 U11796 ( .A1(n14064), .A2(n14554), .ZN(n16480) );
  NAND2_X1 U11797 ( .A1(n19839), .A2(n20610), .ZN(n12134) );
  INV_X1 U11798 ( .A(n12499), .ZN(n20021) );
  INV_X1 U11799 ( .A(n12515), .ZN(n16717) );
  NAND2_X1 U11800 ( .A1(n16746), .A2(n20601), .ZN(n20247) );
  INV_X1 U11801 ( .A(n16762), .ZN(n16767) );
  INV_X1 U11802 ( .A(n20397), .ZN(n20183) );
  INV_X1 U11803 ( .A(n13786), .ZN(n16800) );
  AND3_X1 U11804 ( .A1(n13787), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13810) );
  AND3_X1 U11805 ( .A1(n13513), .A2(n13519), .A3(n13512), .ZN(n19401) );
  NOR2_X1 U11806 ( .A1(n14398), .A2(n13770), .ZN(n19403) );
  NAND2_X1 U11807 ( .A1(n17469), .A2(n17451), .ZN(n17470) );
  NAND2_X1 U11808 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n9957) );
  INV_X1 U11809 ( .A(n18225), .ZN(n9969) );
  NOR2_X1 U11810 ( .A1(n18428), .A2(n9967), .ZN(n9966) );
  OR2_X1 U11811 ( .A1(n13265), .A2(n13264), .ZN(n13532) );
  NOR2_X1 U11812 ( .A1(n18120), .A2(n14354), .ZN(n14210) );
  AOI21_X1 U11813 ( .B1(n17127), .B2(n10436), .A(n14165), .ZN(n14209) );
  INV_X1 U11814 ( .A(n18183), .ZN(n14279) );
  AND2_X1 U11815 ( .A1(n18431), .A2(n9614), .ZN(n17308) );
  OAI22_X1 U11816 ( .A1(n14293), .A2(n9884), .B1(n13546), .B2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14196) );
  AND2_X1 U11817 ( .A1(n13546), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9884) );
  NOR2_X1 U11818 ( .A1(n13554), .A2(n18458), .ZN(n16978) );
  NAND2_X1 U11819 ( .A1(n13555), .A2(n18741), .ZN(n18458) );
  NAND2_X1 U11820 ( .A1(n13346), .A2(n9885), .ZN(n16891) );
  OAI21_X1 U11821 ( .B1(n16907), .B2(n9841), .A(n9895), .ZN(n18510) );
  AOI21_X1 U11822 ( .B1(n13339), .B2(n18659), .A(n10159), .ZN(n9895) );
  NOR2_X1 U11823 ( .A1(n13340), .A2(n10159), .ZN(n10158) );
  AND2_X1 U11824 ( .A1(n16969), .A2(n16968), .ZN(n18808) );
  NOR2_X1 U11825 ( .A1(n18807), .A2(n18806), .ZN(n18863) );
  NAND2_X1 U11826 ( .A1(n9844), .A2(n13339), .ZN(n18660) );
  NAND2_X1 U11827 ( .A1(n16907), .A2(n18565), .ZN(n9844) );
  NAND2_X1 U11828 ( .A1(n10267), .A2(n10266), .ZN(n18672) );
  AND2_X1 U11829 ( .A1(n13333), .A2(n9678), .ZN(n10266) );
  AND2_X1 U11830 ( .A1(n19404), .A2(n13524), .ZN(n19405) );
  NAND2_X1 U11831 ( .A1(n16932), .A2(n13229), .ZN(n14111) );
  NAND2_X1 U11832 ( .A1(n19574), .A2(n14162), .ZN(n18762) );
  AND4_X1 U11833 ( .A1(n13373), .A2(n13372), .A3(n13371), .A4(n13370), .ZN(
        n13379) );
  AND4_X1 U11834 ( .A1(n13377), .A2(n13376), .A3(n13375), .A4(n13374), .ZN(
        n13378) );
  AND4_X1 U11835 ( .A1(n13365), .A2(n13364), .A3(n13363), .A4(n13362), .ZN(
        n13381) );
  OR2_X1 U11836 ( .A1(n13448), .A2(n13447), .ZN(n19004) );
  INV_X1 U11837 ( .A(n13481), .ZN(n19016) );
  OR2_X1 U11838 ( .A1(n13999), .A2(n13022), .ZN(n14139) );
  NAND2_X1 U11839 ( .A1(n20677), .A2(n9919), .ZN(n20710) );
  NAND2_X1 U11840 ( .A1(n9920), .A2(n13862), .ZN(n9919) );
  INV_X1 U11841 ( .A(n15004), .ZN(n9920) );
  NAND2_X1 U11842 ( .A1(n20710), .A2(n9918), .ZN(n9917) );
  NOR2_X1 U11843 ( .A1(n20693), .A2(n9701), .ZN(n9916) );
  AND2_X1 U11844 ( .A1(n13716), .A2(n13709), .ZN(n20705) );
  INV_X1 U11845 ( .A(n20740), .ZN(n20718) );
  INV_X1 U11846 ( .A(n20784), .ZN(n15274) );
  INV_X1 U11847 ( .A(n20631), .ZN(n20780) );
  NAND2_X1 U11848 ( .A1(n15389), .A2(n13053), .ZN(n15379) );
  OAI21_X1 U11849 ( .B1(n10145), .B2(n9713), .A(n10144), .ZN(n13625) );
  XNOR2_X1 U11850 ( .A(n9862), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15399) );
  NAND2_X1 U11851 ( .A1(n9863), .A2(n10038), .ZN(n9862) );
  OAI21_X1 U11852 ( .B1(n10212), .B2(n9865), .A(n9864), .ZN(n9863) );
  INV_X1 U11853 ( .A(n15220), .ZN(n9865) );
  NAND2_X1 U11854 ( .A1(n13044), .A2(n12926), .ZN(n20807) );
  INV_X1 U11855 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21264) );
  OR2_X1 U11856 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21341) );
  INV_X1 U11857 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21184) );
  INV_X1 U11858 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n21428) );
  NOR2_X1 U11859 ( .A1(n12149), .A2(n13795), .ZN(n19594) );
  OAI211_X1 U11860 ( .C1(n16360), .C2(n19767), .A(n10251), .B(n10250), .ZN(
        n10249) );
  NAND2_X1 U11861 ( .A1(n15616), .A2(n19736), .ZN(n10251) );
  NAND2_X1 U11862 ( .A1(n16369), .A2(n19754), .ZN(n10250) );
  AND2_X1 U11863 ( .A1(n12705), .A2(n12704), .ZN(n19653) );
  NAND2_X1 U11864 ( .A1(n19764), .A2(n19771), .ZN(n19716) );
  AND2_X1 U11865 ( .A1(n19778), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19777) );
  INV_X1 U11866 ( .A(n19767), .ZN(n19785) );
  INV_X1 U11867 ( .A(n13680), .ZN(n10024) );
  NAND2_X1 U11868 ( .A1(n15649), .A2(n9696), .ZN(n15631) );
  AND2_X1 U11869 ( .A1(n13586), .A2(n13589), .ZN(n19621) );
  AND2_X1 U11870 ( .A1(n19832), .A2(n16740), .ZN(n19823) );
  NAND2_X1 U11871 ( .A1(n19832), .A2(n12155), .ZN(n16062) );
  NAND2_X1 U11872 ( .A1(n19905), .A2(n19841), .ZN(n19852) );
  XNOR2_X1 U11873 ( .A(n10005), .B(n16103), .ZN(n16373) );
  OAI21_X1 U11874 ( .B1(n16126), .B2(n10003), .A(n10002), .ZN(n10005) );
  AOI21_X1 U11875 ( .B1(n16097), .B2(n16098), .A(n16099), .ZN(n10002) );
  INV_X1 U11876 ( .A(n9792), .ZN(n9762) );
  NAND2_X1 U11877 ( .A1(n13794), .A2(n12890), .ZN(n19950) );
  NAND2_X1 U11878 ( .A1(n19950), .A2(n13903), .ZN(n19939) );
  NAND2_X1 U11879 ( .A1(n16111), .A2(n16366), .ZN(n9816) );
  INV_X1 U11880 ( .A(n16373), .ZN(n9796) );
  OAI211_X1 U11881 ( .C1(n16159), .C2(n10172), .A(n10173), .B(n10171), .ZN(
        n16408) );
  NAND2_X1 U11882 ( .A1(n10177), .A2(n16139), .ZN(n10172) );
  OAI21_X1 U11883 ( .B1(n16140), .B2(n10177), .A(n10174), .ZN(n10173) );
  NAND2_X1 U11884 ( .A1(n16159), .A2(n9650), .ZN(n10171) );
  INV_X1 U11885 ( .A(n16415), .ZN(n10009) );
  NAND2_X1 U11886 ( .A1(n16416), .A2(n16645), .ZN(n10010) );
  NAND2_X1 U11887 ( .A1(n9861), .A2(n16603), .ZN(n9860) );
  INV_X1 U11888 ( .A(n16141), .ZN(n9861) );
  XNOR2_X1 U11889 ( .A(n9811), .B(n16149), .ZN(n16417) );
  NAND2_X1 U11890 ( .A1(n9792), .A2(n13672), .ZN(n9944) );
  NAND2_X1 U11891 ( .A1(n16196), .A2(n16457), .ZN(n9791) );
  NAND2_X1 U11892 ( .A1(n16205), .A2(n16202), .ZN(n9760) );
  NOR2_X2 U11893 ( .A1(n13163), .A2(n20614), .ZN(n19962) );
  NAND2_X1 U11894 ( .A1(n13141), .A2(n13122), .ZN(n19959) );
  INV_X1 U11895 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20594) );
  AND2_X1 U11896 ( .A1(n16716), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20156) );
  OR2_X1 U11897 ( .A1(n14679), .A2(n14678), .ZN(n20488) );
  NAND2_X1 U11898 ( .A1(n19568), .A2(n19404), .ZN(n18380) );
  INV_X1 U11899 ( .A(n19449), .ZN(n19568) );
  AND2_X1 U11900 ( .A1(n17470), .A2(n14217), .ZN(n17459) );
  NOR2_X1 U11901 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  NOR2_X1 U11902 ( .A1(n17791), .A2(n17457), .ZN(n10237) );
  INV_X1 U11903 ( .A(n17456), .ZN(n10236) );
  INV_X1 U11904 ( .A(n17455), .ZN(n10238) );
  OAI21_X1 U11905 ( .B1(n13767), .B2(n10217), .A(n10216), .ZN(n17562) );
  NAND2_X1 U11906 ( .A1(n18504), .A2(n13764), .ZN(n10217) );
  NAND2_X1 U11907 ( .A1(n17775), .A2(n18504), .ZN(n10216) );
  INV_X1 U11908 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17705) );
  INV_X1 U11909 ( .A(n17816), .ZN(n17796) );
  AND2_X1 U11910 ( .A1(n17885), .A2(n17007), .ZN(n17877) );
  NOR2_X1 U11911 ( .A1(n19024), .A2(n17955), .ZN(n17941) );
  NAND2_X1 U11912 ( .A1(n17972), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17955) );
  NOR2_X1 U11913 ( .A1(n18099), .A2(n17675), .ZN(n18079) );
  NAND2_X1 U11914 ( .A1(n9595), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n18099) );
  NOR2_X1 U11915 ( .A1(n17734), .A2(n9981), .ZN(n9980) );
  INV_X1 U11916 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n9981) );
  INV_X1 U11917 ( .A(n18194), .ZN(n18190) );
  NOR2_X2 U11918 ( .A1(n18186), .A2(n18316), .ZN(n18257) );
  NOR2_X2 U11919 ( .A1(n19016), .A2(n18316), .ZN(n18258) );
  NAND2_X1 U11920 ( .A1(n9965), .A2(n9966), .ZN(n18259) );
  NAND2_X1 U11921 ( .A1(n18184), .A2(n10446), .ZN(n18264) );
  NAND2_X1 U11922 ( .A1(n18444), .A2(n9649), .ZN(n10059) );
  INV_X1 U11923 ( .A(n18442), .ZN(n9880) );
  INV_X1 U11924 ( .A(n18441), .ZN(n9879) );
  OR2_X1 U11925 ( .A1(n18455), .A2(n13355), .ZN(n9883) );
  NOR2_X1 U11926 ( .A1(n18520), .A2(n18438), .ZN(n9882) );
  AND2_X1 U11927 ( .A1(n16923), .A2(n17130), .ZN(n18681) );
  NAND2_X1 U11928 ( .A1(n10273), .A2(n10272), .ZN(n18733) );
  INV_X1 U11929 ( .A(n18450), .ZN(n10272) );
  INV_X1 U11930 ( .A(n18451), .ZN(n10273) );
  NOR2_X1 U11931 ( .A1(n18891), .A2(n18888), .ZN(n18915) );
  INV_X1 U11932 ( .A(n16751), .ZN(n12517) );
  INV_X1 U11933 ( .A(n10594), .ZN(n10203) );
  INV_X1 U11934 ( .A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10756) );
  AND2_X1 U11935 ( .A1(n10919), .A2(n10918), .ZN(n10928) );
  NAND2_X1 U11936 ( .A1(n10610), .A2(n10589), .ZN(n10075) );
  AND2_X1 U11937 ( .A1(n12507), .A2(n12508), .ZN(n9899) );
  AOI22_X1 U11938 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20115), .B1(
        n19976), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12507) );
  NAND2_X1 U11939 ( .A1(n12404), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10124) );
  INV_X1 U11940 ( .A(n11772), .ZN(n11771) );
  INV_X1 U11941 ( .A(n12189), .ZN(n12193) );
  NAND2_X1 U11942 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n9991) );
  AOI21_X1 U11943 ( .B1(n11790), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n11656), .ZN(n9992) );
  NAND2_X1 U11944 ( .A1(n10932), .A2(n10931), .ZN(n10945) );
  INV_X1 U11945 ( .A(n10855), .ZN(n10854) );
  INV_X1 U11946 ( .A(n17232), .ZN(n10090) );
  OR2_X1 U11947 ( .A1(n10853), .A2(n10852), .ZN(n10869) );
  OR2_X1 U11948 ( .A1(n10784), .A2(n10783), .ZN(n10856) );
  INV_X1 U11949 ( .A(n10598), .ZN(n10586) );
  CLKBUF_X1 U11950 ( .A(n10688), .Z(n10707) );
  CLKBUF_X1 U11951 ( .A(n10730), .Z(n10731) );
  NAND2_X1 U11952 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10555) );
  OR2_X1 U11953 ( .A1(n10570), .A2(n10505), .ZN(n10506) );
  NAND2_X1 U11954 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10476) );
  NAND2_X1 U11955 ( .A1(n10956), .A2(n14078), .ZN(n10953) );
  AND2_X1 U11956 ( .A1(n13096), .A2(n12140), .ZN(n9814) );
  INV_X1 U11957 ( .A(n12615), .ZN(n12616) );
  NAND2_X1 U11958 ( .A1(n9898), .A2(n12522), .ZN(n12613) );
  NOR2_X1 U11959 ( .A1(n12415), .A2(n9941), .ZN(n12436) );
  OAI21_X1 U11960 ( .B1(n9940), .B2(n19945), .A(n9938), .ZN(n9941) );
  NAND2_X1 U11961 ( .A1(n9675), .A2(n9947), .ZN(n12407) );
  NOR2_X1 U11962 ( .A1(n16751), .A2(n12455), .ZN(n12458) );
  INV_X1 U11963 ( .A(n12154), .ZN(n13125) );
  NAND2_X1 U11964 ( .A1(n12179), .A2(n19992), .ZN(n13101) );
  AOI21_X1 U11965 ( .B1(n11723), .B2(P2_REIP_REG_1__SCAN_IN), .A(n9717), .ZN(
        n9769) );
  NAND2_X1 U11966 ( .A1(n11699), .A2(n12197), .ZN(n13096) );
  OR2_X1 U11967 ( .A1(n12109), .A2(n12104), .ZN(n12105) );
  NOR2_X1 U11968 ( .A1(n16927), .A2(n10228), .ZN(n10227) );
  NAND2_X1 U11969 ( .A1(n13528), .A2(n14281), .ZN(n13249) );
  NAND2_X1 U11970 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13172) );
  NOR2_X1 U11971 ( .A1(n14863), .A2(n10287), .ZN(n10286) );
  INV_X1 U11972 ( .A(n10423), .ZN(n10287) );
  NAND2_X1 U11973 ( .A1(n10901), .A2(n10893), .ZN(n15311) );
  NAND2_X1 U11974 ( .A1(n10901), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15315) );
  NAND2_X1 U11975 ( .A1(n10840), .A2(n10855), .ZN(n11035) );
  NOR2_X1 U11976 ( .A1(n10996), .A2(n9900), .ZN(n11018) );
  NAND2_X1 U11977 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n9900) );
  AND2_X1 U11978 ( .A1(n15353), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10095) );
  INV_X1 U11979 ( .A(n14774), .ZN(n10328) );
  NOR2_X1 U11980 ( .A1(n15353), .A2(n10036), .ZN(n10035) );
  INV_X1 U11981 ( .A(n10394), .ZN(n10036) );
  NOR2_X1 U11982 ( .A1(n10898), .A2(n10900), .ZN(n10140) );
  NAND2_X1 U11983 ( .A1(n15286), .A2(n10892), .ZN(n9858) );
  OR2_X1 U11984 ( .A1(n15353), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10082) );
  NAND2_X1 U11985 ( .A1(n10800), .A2(n9711), .ZN(n10200) );
  INV_X1 U11986 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10201) );
  NAND2_X1 U11987 ( .A1(n9819), .A2(n9710), .ZN(n9820) );
  NAND2_X1 U11988 ( .A1(n9819), .A2(n10806), .ZN(n14490) );
  XNOR2_X1 U11989 ( .A(n10071), .B(n10727), .ZN(n10808) );
  NAND2_X1 U11990 ( .A1(n9987), .A2(n10606), .ZN(n10692) );
  AND3_X1 U11991 ( .A1(n10621), .A2(n10620), .A3(n10619), .ZN(n10690) );
  INV_X1 U11992 ( .A(n10585), .ZN(n12902) );
  INV_X1 U11993 ( .A(n10279), .ZN(n9869) );
  NAND2_X1 U11994 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n9757) );
  NOR2_X1 U11995 ( .A1(n9659), .A2(n10087), .ZN(n10532) );
  AND2_X1 U11996 ( .A1(n10635), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10087) );
  AOI22_X1 U11997 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10650), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10522) );
  NAND2_X1 U11998 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10541) );
  INV_X1 U11999 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21216) );
  OAI211_X1 U12000 ( .C1(n9873), .C2(n9627), .A(n10276), .B(n9870), .ZN(n9876)
         );
  NAND2_X1 U12001 ( .A1(n9874), .A2(n10279), .ZN(n9873) );
  INV_X1 U12002 ( .A(n21265), .ZN(n21339) );
  OAI21_X1 U12003 ( .B1(n10961), .B2(n10960), .A(n9667), .ZN(n9751) );
  INV_X1 U12004 ( .A(n11698), .ZN(n9998) );
  AND2_X1 U12005 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11669) );
  INV_X1 U12006 ( .A(n11705), .ZN(n11710) );
  INV_X1 U12007 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U12008 ( .A1(n10307), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U12009 ( .A1(n12594), .A2(n10308), .ZN(n10307) );
  OR2_X1 U12010 ( .A1(n19764), .A2(n20488), .ZN(n15826) );
  INV_X1 U12011 ( .A(n10338), .ZN(n10337) );
  OAI21_X1 U12012 ( .B1(n12792), .B2(n20540), .A(n12855), .ZN(n10338) );
  NAND2_X1 U12013 ( .A1(n10346), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10341) );
  CLKBUF_X1 U12014 ( .A(n12037), .Z(n14598) );
  CLKBUF_X1 U12015 ( .A(n12089), .Z(n14599) );
  NOR2_X1 U12016 ( .A1(n15865), .A2(n10193), .ZN(n10192) );
  INV_X1 U12017 ( .A(n10184), .ZN(n10183) );
  NAND2_X1 U12018 ( .A1(n15889), .A2(n10018), .ZN(n10017) );
  AND2_X1 U12019 ( .A1(n14566), .A2(n16067), .ZN(n10377) );
  INV_X1 U12020 ( .A(n15917), .ZN(n10197) );
  NOR2_X1 U12021 ( .A1(n9601), .A2(n9651), .ZN(n10298) );
  NAND2_X1 U12022 ( .A1(n11790), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U12023 ( .A1(n10346), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10345) );
  AND2_X1 U12024 ( .A1(n12860), .A2(n9645), .ZN(n13668) );
  AND2_X1 U12025 ( .A1(n9705), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10247) );
  INV_X1 U12026 ( .A(n10332), .ZN(n10331) );
  OAI21_X1 U12027 ( .B1(n12792), .B2(n20531), .A(n12835), .ZN(n10332) );
  NOR2_X1 U12028 ( .A1(n10405), .A2(n10403), .ZN(n10400) );
  INV_X1 U12029 ( .A(n15962), .ZN(n10403) );
  NOR2_X1 U12030 ( .A1(n9594), .A2(n10243), .ZN(n10242) );
  INV_X1 U12031 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10243) );
  INV_X1 U12032 ( .A(n10330), .ZN(n10329) );
  OAI21_X1 U12033 ( .B1(n12792), .B2(n20520), .A(n12795), .ZN(n10330) );
  NOR2_X1 U12034 ( .A1(n19748), .A2(n10245), .ZN(n10244) );
  INV_X1 U12035 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10245) );
  NAND2_X1 U12036 ( .A1(n12530), .A2(n9706), .ZN(n12533) );
  NOR2_X1 U12037 ( .A1(n12211), .A2(n12212), .ZN(n12563) );
  OAI21_X1 U12038 ( .B1(n16248), .B2(n10438), .A(n10116), .ZN(n10001) );
  INV_X1 U12039 ( .A(n10117), .ZN(n10116) );
  AOI21_X1 U12040 ( .B1(n16097), .B2(n16098), .A(n16099), .ZN(n10047) );
  NOR2_X1 U12041 ( .A1(n10381), .A2(n10379), .ZN(n10378) );
  INV_X1 U12042 ( .A(n15676), .ZN(n10379) );
  INV_X1 U12043 ( .A(n15698), .ZN(n10380) );
  INV_X1 U12044 ( .A(n16238), .ZN(n10015) );
  NAND2_X1 U12045 ( .A1(n10257), .A2(n16232), .ZN(n10256) );
  INV_X1 U12046 ( .A(n10261), .ZN(n10257) );
  INV_X1 U12047 ( .A(n10014), .ZN(n10013) );
  OAI21_X1 U12048 ( .B1(n9590), .B2(n16239), .A(n10259), .ZN(n10014) );
  INV_X1 U12049 ( .A(n10260), .ZN(n10259) );
  OAI21_X1 U12050 ( .B1(n10263), .B2(n10261), .A(n13578), .ZN(n10260) );
  NOR2_X1 U12051 ( .A1(n10385), .A2(n10387), .ZN(n10384) );
  INV_X1 U12052 ( .A(n10450), .ZN(n10387) );
  AND2_X1 U12053 ( .A1(n16249), .A2(n16263), .ZN(n10255) );
  AND3_X1 U12054 ( .A1(n12336), .A2(n12335), .A3(n12334), .ZN(n14185) );
  NOR2_X1 U12055 ( .A1(n12310), .A2(n10367), .ZN(n10366) );
  INV_X1 U12056 ( .A(n10374), .ZN(n10367) );
  NAND2_X1 U12057 ( .A1(n12543), .A2(n12547), .ZN(n16313) );
  INV_X1 U12058 ( .A(n12547), .ZN(n12548) );
  NOR2_X1 U12059 ( .A1(n12264), .A2(n12263), .ZN(n12586) );
  OR2_X1 U12060 ( .A1(n12248), .A2(n12247), .ZN(n12585) );
  NAND2_X1 U12061 ( .A1(n11707), .A2(n11706), .ZN(n9809) );
  INV_X1 U12062 ( .A(n11708), .ZN(n9810) );
  INV_X1 U12063 ( .A(n11716), .ZN(n13119) );
  AND2_X1 U12064 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11759) );
  OR2_X1 U12065 ( .A1(n12230), .A2(n12229), .ZN(n12579) );
  NAND2_X1 U12066 ( .A1(n12148), .A2(n9804), .ZN(n11724) );
  NAND2_X1 U12067 ( .A1(n12153), .A2(n9662), .ZN(n9804) );
  AND2_X1 U12068 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U12069 ( .A1(n10110), .A2(n10108), .ZN(n11702) );
  NOR2_X1 U12070 ( .A1(n20183), .A2(n20589), .ZN(n16715) );
  NOR2_X1 U12071 ( .A1(n13511), .A2(n13521), .ZN(n13518) );
  AND2_X1 U12072 ( .A1(n13509), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13515) );
  AOI21_X1 U12073 ( .B1(n13507), .B2(n13506), .A(n13505), .ZN(n13519) );
  AND4_X1 U12074 ( .A1(n13255), .A2(n13254), .A3(n13253), .A4(n13252), .ZN(
        n13259) );
  AND2_X1 U12075 ( .A1(n13177), .A2(n13180), .ZN(n13256) );
  NAND2_X1 U12076 ( .A1(n18431), .A2(n9612), .ZN(n17439) );
  NAND2_X1 U12077 ( .A1(n18431), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n18433) );
  AND2_X1 U12078 ( .A1(n16896), .A2(n16881), .ZN(n18431) );
  NAND2_X1 U12079 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n10222), .ZN(
        n10221) );
  AND4_X1 U12080 ( .A1(n13316), .A2(n13315), .A3(n13314), .A4(n13313), .ZN(
        n13328) );
  AND2_X1 U12081 ( .A1(n13343), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9846) );
  NOR2_X1 U12082 ( .A1(n9845), .A2(n18659), .ZN(n9843) );
  AND2_X1 U12083 ( .A1(n18565), .A2(n18818), .ZN(n18530) );
  AND2_X1 U12084 ( .A1(n18670), .A2(n10057), .ZN(n10056) );
  NAND2_X1 U12085 ( .A1(n13479), .A2(n17413), .ZN(n14160) );
  NOR2_X1 U12086 ( .A1(n19016), .A2(n18186), .ZN(n14098) );
  AOI21_X1 U12087 ( .B1(n13287), .B2(n18942), .A(n10153), .ZN(n10052) );
  INV_X1 U12088 ( .A(n14301), .ZN(n10153) );
  AND2_X1 U12089 ( .A1(n14173), .A2(n14098), .ZN(n14204) );
  NOR2_X1 U12090 ( .A1(n13172), .A2(n14393), .ZN(n17119) );
  AND3_X1 U12091 ( .A1(n13437), .A2(n13436), .A3(n13435), .ZN(n13441) );
  AND2_X1 U12092 ( .A1(n9971), .A2(n9656), .ZN(n13474) );
  NOR2_X1 U12093 ( .A1(n13414), .A2(n9972), .ZN(n9971) );
  NOR2_X1 U12094 ( .A1(n13434), .A2(n13433), .ZN(n13481) );
  AOI221_X1 U12095 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n21628), .C1(n19451), 
        .C2(P3_STATE2_REG_2__SCAN_IN), .A(n19444), .ZN(n18991) );
  CLKBUF_X1 U12096 ( .A(n10616), .Z(n13862) );
  OR3_X1 U12097 ( .A1(n21505), .A2(n13706), .A3(n13705), .ZN(n15001) );
  OR2_X1 U12098 ( .A1(n10312), .A2(n10310), .ZN(n10309) );
  INV_X1 U12099 ( .A(n14947), .ZN(n10310) );
  NAND2_X1 U12100 ( .A1(n10274), .A2(n14039), .ZN(n13914) );
  OR2_X1 U12101 ( .A1(n11542), .A2(n9914), .ZN(n11579) );
  OR2_X1 U12102 ( .A1(n11434), .A2(n9909), .ZN(n11436) );
  OR2_X1 U12103 ( .A1(n15214), .A2(n11573), .ZN(n11459) );
  AND2_X1 U12104 ( .A1(n11284), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11285) );
  AND2_X1 U12105 ( .A1(n11305), .A2(n11304), .ZN(n14849) );
  OR2_X1 U12106 ( .A1(n15262), .A2(n11573), .ZN(n11305) );
  NAND2_X1 U12107 ( .A1(n11239), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11283) );
  NOR2_X1 U12108 ( .A1(n11238), .A2(n14901), .ZN(n11239) );
  OR2_X1 U12109 ( .A1(n11199), .A2(n17191), .ZN(n11200) );
  OR2_X1 U12110 ( .A1(n11200), .A2(n14914), .ZN(n11238) );
  NAND2_X1 U12111 ( .A1(n9903), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11199) );
  INV_X1 U12112 ( .A(n11193), .ZN(n9903) );
  INV_X1 U12113 ( .A(n10424), .ZN(n9926) );
  NAND2_X1 U12114 ( .A1(n11102), .A2(n9901), .ZN(n11193) );
  NOR2_X1 U12115 ( .A1(n14932), .A2(n9902), .ZN(n9901) );
  AND3_X1 U12116 ( .A1(n14927), .A2(n14926), .A3(n14943), .ZN(n15054) );
  NAND2_X1 U12117 ( .A1(n11029), .A2(n9904), .ZN(n11079) );
  NOR2_X1 U12118 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  INV_X1 U12119 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9905) );
  INV_X1 U12120 ( .A(n11036), .ZN(n11029) );
  NAND2_X1 U12121 ( .A1(n11029), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11074) );
  NAND2_X1 U12122 ( .A1(n11037), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11036) );
  AND2_X1 U12123 ( .A1(n11018), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11037) );
  NAND3_X1 U12124 ( .A1(n14450), .A2(n14449), .A3(n11016), .ZN(n14498) );
  INV_X1 U12125 ( .A(n14459), .ZN(n11016) );
  INV_X1 U12126 ( .A(n11017), .ZN(n11027) );
  INV_X1 U12127 ( .A(n10283), .ZN(n10284) );
  OAI21_X1 U12128 ( .B1(n10975), .B2(n10825), .A(n10813), .ZN(n14484) );
  OAI21_X1 U12129 ( .B1(n10975), .B2(n11196), .A(n10974), .ZN(n10280) );
  NAND2_X1 U12130 ( .A1(n15203), .A2(n13735), .ZN(n12898) );
  NOR2_X1 U12131 ( .A1(n15204), .A2(n13062), .ZN(n13739) );
  NAND2_X1 U12132 ( .A1(n9989), .A2(n9742), .ZN(n10102) );
  NAND2_X1 U12133 ( .A1(n15333), .A2(n15219), .ZN(n9864) );
  INV_X1 U12134 ( .A(n10903), .ZN(n9988) );
  AND2_X1 U12135 ( .A1(n14814), .A2(n13008), .ZN(n14815) );
  AND2_X1 U12136 ( .A1(n12998), .A2(n12997), .ZN(n14852) );
  NAND2_X1 U12137 ( .A1(n10142), .A2(n10137), .ZN(n15252) );
  NOR2_X1 U12138 ( .A1(n10138), .A2(n10898), .ZN(n10137) );
  INV_X1 U12139 ( .A(n10895), .ZN(n10138) );
  AND2_X1 U12140 ( .A1(n12994), .A2(n12993), .ZN(n14865) );
  OR2_X1 U12141 ( .A1(n10323), .A2(n14891), .ZN(n10322) );
  NOR2_X1 U12142 ( .A1(n15061), .A2(n10325), .ZN(n10434) );
  XNOR2_X1 U12143 ( .A(n10885), .B(n15493), .ZN(n15289) );
  INV_X1 U12144 ( .A(n10892), .ZN(n15287) );
  NAND2_X1 U12145 ( .A1(n14929), .A2(n14930), .ZN(n15063) );
  OR2_X1 U12146 ( .A1(n15063), .A2(n15064), .ZN(n15061) );
  NAND2_X1 U12147 ( .A1(n15341), .A2(n15285), .ZN(n15305) );
  AND2_X1 U12148 ( .A1(n12973), .A2(n12972), .ZN(n15073) );
  NAND2_X1 U12149 ( .A1(n10311), .A2(n12968), .ZN(n15074) );
  INV_X1 U12150 ( .A(n15086), .ZN(n10311) );
  AND2_X1 U12151 ( .A1(n12955), .A2(n9687), .ZN(n15084) );
  INV_X1 U12152 ( .A(n15580), .ZN(n17255) );
  AOI21_X1 U12153 ( .B1(n14073), .B2(n12959), .A(n12939), .ZN(n14256) );
  INV_X1 U12154 ( .A(n20889), .ZN(n14502) );
  OAI21_X1 U12155 ( .B1(n10819), .B2(n10209), .A(n10207), .ZN(n9924) );
  INV_X1 U12156 ( .A(n10208), .ZN(n10207) );
  OAI21_X1 U12157 ( .B1(n10984), .B2(n10209), .A(n10684), .ZN(n10208) );
  INV_X1 U12158 ( .A(n14576), .ZN(n15595) );
  NAND2_X1 U12160 ( .A1(n13925), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13928) );
  NAND2_X1 U12161 ( .A1(n9867), .A2(n9866), .ZN(n21088) );
  NAND2_X1 U12162 ( .A1(n9627), .A2(n10279), .ZN(n9866) );
  AND2_X1 U12163 ( .A1(n9868), .A2(n9874), .ZN(n9867) );
  NAND2_X1 U12164 ( .A1(n9869), .A2(n9872), .ZN(n9868) );
  OR3_X1 U12165 ( .A1(n13944), .A2(n13943), .A3(n13942), .ZN(n17143) );
  AND3_X1 U12166 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n10276), .A3(n14510), 
        .ZN(n20854) );
  NOR2_X1 U12167 ( .A1(n14417), .A2(n20889), .ZN(n21263) );
  AND2_X1 U12168 ( .A1(n14417), .A2(n20889), .ZN(n21295) );
  INV_X1 U12169 ( .A(n21341), .ZN(n21349) );
  OR2_X1 U12170 ( .A1(n14037), .A2(n12922), .ZN(n17155) );
  NAND2_X2 U12171 ( .A1(n11689), .A2(n14621), .ZN(n10293) );
  OR2_X1 U12172 ( .A1(n12445), .A2(n15607), .ZN(n11689) );
  NAND2_X1 U12173 ( .A1(n15607), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15606) );
  NOR2_X1 U12174 ( .A1(n15733), .A2(n10240), .ZN(n10239) );
  INV_X1 U12175 ( .A(n16199), .ZN(n10240) );
  NAND2_X1 U12176 ( .A1(n12718), .A2(n12596), .ZN(n12719) );
  NAND2_X1 U12177 ( .A1(n12693), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U12178 ( .A1(n12575), .A2(n12721), .ZN(n12577) );
  INV_X1 U12179 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15842) );
  AND2_X1 U12180 ( .A1(n12884), .A2(n12883), .ZN(n15630) );
  OAI211_X1 U12181 ( .C1(n12779), .C2(n16117), .A(n12881), .B(n12880), .ZN(
        n12882) );
  AND2_X1 U12182 ( .A1(n12874), .A2(n12873), .ZN(n15663) );
  OAI211_X1 U12183 ( .C1(n12779), .C2(n20550), .A(n12871), .B(n12870), .ZN(
        n12872) );
  CLKBUF_X1 U12184 ( .A(n13585), .Z(n13586) );
  AND2_X1 U12185 ( .A1(n12841), .A2(n9644), .ZN(n15928) );
  INV_X1 U12186 ( .A(n13113), .ZN(n13116) );
  AND2_X1 U12187 ( .A1(n15894), .A2(n15910), .ZN(n15912) );
  AND2_X1 U12188 ( .A1(n12347), .A2(n12346), .ZN(n16497) );
  AND3_X1 U12189 ( .A1(n12330), .A2(n12329), .A3(n12328), .ZN(n14119) );
  INV_X2 U12190 ( .A(n16714), .ZN(n16713) );
  INV_X1 U12191 ( .A(n15606), .ZN(n19839) );
  NOR2_X1 U12192 ( .A1(n10004), .A2(n16097), .ZN(n10003) );
  INV_X1 U12193 ( .A(n16100), .ZN(n10004) );
  NAND2_X1 U12194 ( .A1(n14667), .A2(n9613), .ZN(n14670) );
  NAND2_X1 U12195 ( .A1(n9801), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9800) );
  INV_X1 U12196 ( .A(n16315), .ZN(n9801) );
  AND2_X1 U12197 ( .A1(n14667), .A2(n9728), .ZN(n14669) );
  AND2_X1 U12198 ( .A1(n14624), .A2(n10246), .ZN(n14663) );
  AND2_X1 U12199 ( .A1(n10247), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10246) );
  NOR2_X1 U12200 ( .A1(n15740), .A2(n13668), .ZN(n15714) );
  NAND2_X1 U12201 ( .A1(n12847), .A2(n9647), .ZN(n15915) );
  NAND2_X1 U12202 ( .A1(n10409), .A2(n14569), .ZN(n10408) );
  INV_X1 U12203 ( .A(n10411), .ZN(n10409) );
  NAND2_X1 U12204 ( .A1(n14643), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14646) );
  INV_X1 U12205 ( .A(n15932), .ZN(n10410) );
  AND2_X1 U12206 ( .A1(n12831), .A2(n12830), .ZN(n15764) );
  INV_X1 U12207 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12891) );
  NAND2_X1 U12208 ( .A1(n14625), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14644) );
  AND2_X1 U12209 ( .A1(n12824), .A2(n12823), .ZN(n15950) );
  CLKBUF_X1 U12210 ( .A(n14628), .Z(n14640) );
  INV_X1 U12211 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16296) );
  INV_X1 U12212 ( .A(n15792), .ZN(n10404) );
  OR2_X1 U12213 ( .A1(n14375), .A2(n10405), .ZN(n10402) );
  NOR2_X1 U12214 ( .A1(n14636), .A2(n9594), .ZN(n14641) );
  NAND2_X1 U12215 ( .A1(n10241), .A2(n10244), .ZN(n14638) );
  NOR2_X1 U12216 ( .A1(n14636), .A2(n19748), .ZN(n14639) );
  NAND2_X1 U12217 ( .A1(n16837), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12894) );
  INV_X1 U12218 ( .A(n13079), .ZN(n13081) );
  NAND2_X1 U12219 ( .A1(n14531), .A2(n10388), .ZN(n10391) );
  AND2_X1 U12220 ( .A1(n10389), .A2(n15623), .ZN(n10388) );
  NOR2_X1 U12221 ( .A1(n13114), .A2(n10390), .ZN(n10389) );
  INV_X1 U12222 ( .A(n12374), .ZN(n10390) );
  NAND2_X1 U12223 ( .A1(n12878), .A2(n9708), .ZN(n14540) );
  NAND2_X1 U12224 ( .A1(n9607), .A2(n12590), .ZN(n16127) );
  AND2_X1 U12225 ( .A1(n12367), .A2(n12366), .ZN(n15660) );
  CLKBUF_X1 U12226 ( .A(n14529), .Z(n14530) );
  CLKBUF_X1 U12227 ( .A(n15658), .Z(n15678) );
  INV_X1 U12228 ( .A(n10179), .ZN(n10176) );
  NAND2_X1 U12229 ( .A1(n10175), .A2(n10177), .ZN(n10174) );
  NAND2_X1 U12230 ( .A1(n16139), .A2(n10179), .ZN(n10175) );
  INV_X1 U12231 ( .A(n10178), .ZN(n10177) );
  OAI21_X1 U12232 ( .B1(n10179), .B2(n16157), .A(n16148), .ZN(n10178) );
  OR2_X1 U12233 ( .A1(n16421), .A2(n13148), .ZN(n16412) );
  NAND2_X1 U12234 ( .A1(n10415), .A2(n9615), .ZN(n15683) );
  INV_X1 U12235 ( .A(n15681), .ZN(n10414) );
  AND2_X1 U12236 ( .A1(n12364), .A2(n12363), .ZN(n15685) );
  NOR2_X1 U12237 ( .A1(n15698), .A2(n10381), .ZN(n15675) );
  NAND2_X1 U12238 ( .A1(n9771), .A2(n10129), .ZN(n16174) );
  INV_X1 U12239 ( .A(n16179), .ZN(n10130) );
  NAND2_X1 U12240 ( .A1(n12864), .A2(n9648), .ZN(n15696) );
  INV_X1 U12241 ( .A(n10416), .ZN(n10413) );
  AND2_X1 U12242 ( .A1(n12358), .A2(n12357), .ZN(n13666) );
  NAND2_X1 U12243 ( .A1(n9813), .A2(n9772), .ZN(n16262) );
  CLKBUF_X1 U12244 ( .A(n14021), .Z(n14022) );
  NAND2_X1 U12245 ( .A1(n9888), .A2(n9887), .ZN(n16305) );
  NAND2_X1 U12246 ( .A1(n9889), .A2(n16279), .ZN(n9888) );
  NAND2_X1 U12247 ( .A1(n9890), .A2(n16319), .ZN(n9889) );
  AND3_X1 U12248 ( .A1(n12314), .A2(n12313), .A3(n12312), .ZN(n13884) );
  XNOR2_X1 U12249 ( .A(n9849), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16334) );
  NAND2_X1 U12250 ( .A1(n12641), .A2(n12786), .ZN(n16634) );
  INV_X1 U12251 ( .A(n16347), .ZN(n10068) );
  XNOR2_X1 U12252 ( .A(n11743), .B(n12806), .ZN(n11744) );
  INV_X1 U12253 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13142) );
  NOR2_X1 U12254 ( .A1(n12341), .A2(n12173), .ZN(n12176) );
  XNOR2_X1 U12255 ( .A(n16654), .B(n11777), .ZN(n14012) );
  CLKBUF_X1 U12256 ( .A(n14048), .Z(n14049) );
  OAI21_X1 U12257 ( .B1(n16735), .B2(n9587), .A(n20581), .ZN(n11773) );
  CLKBUF_X1 U12258 ( .A(n16660), .Z(n16661) );
  CLKBUF_X1 U12259 ( .A(n12556), .Z(n16693) );
  INV_X1 U12260 ( .A(n12516), .ZN(n16728) );
  INV_X1 U12261 ( .A(n20576), .ZN(n20182) );
  AND2_X1 U12262 ( .A1(n20386), .A2(n20385), .ZN(n20390) );
  INV_X1 U12263 ( .A(n20390), .ZN(n20396) );
  AND3_X1 U12264 ( .A1(n10182), .A2(n10181), .A3(n11656), .ZN(n11614) );
  AND2_X1 U12265 ( .A1(n20302), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11752) );
  OR2_X1 U12266 ( .A1(n20247), .A2(n20574), .ZN(n19972) );
  NAND2_X2 U12267 ( .A1(n16715), .A2(n16714), .ZN(n20005) );
  NAND2_X2 U12268 ( .A1(n16713), .A2(n16715), .ZN(n20007) );
  NOR2_X1 U12269 ( .A1(n20582), .A2(n19970), .ZN(n20306) );
  AND2_X1 U12270 ( .A1(n12104), .A2(n12103), .ZN(n12566) );
  NAND2_X1 U12271 ( .A1(n12124), .A2(n12123), .ZN(n12569) );
  NOR2_X1 U12272 ( .A1(n20392), .A2(n13787), .ZN(n14151) );
  AND4_X1 U12273 ( .A1(n13389), .A2(n13388), .A3(n13387), .A4(n13386), .ZN(
        n13400) );
  AND4_X1 U12274 ( .A1(n13385), .A2(n13384), .A3(n13383), .A4(n13382), .ZN(
        n13401) );
  AND4_X1 U12275 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13398) );
  NAND2_X1 U12276 ( .A1(n10215), .A2(n14217), .ZN(n17469) );
  OR2_X1 U12277 ( .A1(n17486), .A2(n17487), .ZN(n10215) );
  NOR2_X1 U12278 ( .A1(n18452), .A2(n17495), .ZN(n17494) );
  INV_X1 U12279 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17540) );
  AND2_X1 U12280 ( .A1(n17551), .A2(n14217), .ZN(n17539) );
  OR2_X1 U12281 ( .A1(n17553), .A2(n18496), .ZN(n17551) );
  NOR2_X1 U12282 ( .A1(n17823), .A2(n17824), .ZN(n9961) );
  NAND2_X1 U12283 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18079), .ZN(n17117) );
  NOR2_X1 U12284 ( .A1(n18327), .A2(n18329), .ZN(n9970) );
  NOR2_X1 U12285 ( .A1(n19001), .A2(n18992), .ZN(n14208) );
  AOI21_X1 U12286 ( .B1(n14160), .B2(n19442), .A(n19569), .ZN(n18322) );
  INV_X1 U12287 ( .A(n18380), .ZN(n18378) );
  NOR2_X1 U12288 ( .A1(n10441), .A2(n17540), .ZN(n16896) );
  NAND2_X1 U12289 ( .A1(n17574), .A2(n9699), .ZN(n18497) );
  NOR2_X1 U12290 ( .A1(n18538), .A2(n10231), .ZN(n10230) );
  NAND2_X1 U12291 ( .A1(n17574), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18537) );
  NOR2_X1 U12292 ( .A1(n18904), .A2(n10159), .ZN(n13555) );
  NAND3_X1 U12293 ( .A1(n13558), .A2(n10218), .A3(n10220), .ZN(n18571) );
  INV_X1 U12294 ( .A(n10221), .ZN(n10220) );
  NOR2_X1 U12295 ( .A1(n16911), .A2(n17634), .ZN(n10218) );
  AND2_X1 U12296 ( .A1(n13558), .A2(n10219), .ZN(n18596) );
  NOR2_X1 U12297 ( .A1(n16911), .A2(n10221), .ZN(n10219) );
  NAND2_X1 U12298 ( .A1(n16901), .A2(n13558), .ZN(n18638) );
  NOR2_X1 U12299 ( .A1(n16911), .A2(n18685), .ZN(n16901) );
  NAND2_X1 U12300 ( .A1(n18701), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16911) );
  NAND2_X1 U12301 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10214) );
  INV_X1 U12302 ( .A(n16878), .ZN(n10055) );
  NAND2_X1 U12303 ( .A1(n16891), .A2(n18565), .ZN(n18469) );
  NAND2_X1 U12304 ( .A1(n13351), .A2(n18659), .ZN(n18470) );
  AND2_X1 U12305 ( .A1(n18548), .A2(n13343), .ZN(n18476) );
  INV_X1 U12306 ( .A(n18861), .ZN(n18858) );
  OR2_X1 U12307 ( .A1(n13338), .A2(n18659), .ZN(n13556) );
  NOR2_X1 U12308 ( .A1(n14260), .A2(n13334), .ZN(n14259) );
  NAND2_X1 U12309 ( .A1(n18694), .A2(n13545), .ZN(n14293) );
  NAND2_X1 U12310 ( .A1(n16924), .A2(n13544), .ZN(n18695) );
  NAND2_X1 U12311 ( .A1(n18695), .A2(n18696), .ZN(n18694) );
  NAND2_X1 U12312 ( .A1(n14087), .A2(n13542), .ZN(n18704) );
  NAND2_X1 U12313 ( .A1(n18704), .A2(n18705), .ZN(n18706) );
  XNOR2_X1 U12314 ( .A(n13541), .B(n9877), .ZN(n14088) );
  NAND2_X1 U12315 ( .A1(n14089), .A2(n14088), .ZN(n14087) );
  NAND2_X1 U12316 ( .A1(n13187), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9829) );
  NOR2_X2 U12317 ( .A1(n14102), .A2(n18836), .ZN(n16961) );
  INV_X1 U12318 ( .A(n18762), .ZN(n19400) );
  NAND2_X1 U12319 ( .A1(n13769), .A2(n14388), .ZN(n17127) );
  NOR3_X1 U12320 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n19571), .ZN(n19271) );
  NOR2_X1 U12321 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18991), .ZN(n19323) );
  INV_X1 U12322 ( .A(n19323), .ZN(n19179) );
  INV_X1 U12323 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19452) );
  NAND2_X1 U12324 ( .A1(n14139), .A2(n13802), .ZN(n21505) );
  NAND2_X1 U12325 ( .A1(n11306), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11372) );
  NOR2_X1 U12326 ( .A1(n20687), .A2(n14869), .ZN(n20652) );
  NAND2_X1 U12327 ( .A1(n13731), .A2(n13730), .ZN(n20677) );
  INV_X1 U12328 ( .A(n20710), .ZN(n20692) );
  INV_X1 U12329 ( .A(n15099), .ZN(n15107) );
  NAND2_X1 U12330 ( .A1(n14044), .A2(n14043), .ZN(n15096) );
  NAND2_X1 U12331 ( .A1(n14042), .A2(n14041), .ZN(n14044) );
  INV_X1 U12332 ( .A(n15105), .ZN(n15097) );
  OR2_X1 U12333 ( .A1(n15096), .A2(n10599), .ZN(n15105) );
  INV_X1 U12334 ( .A(n15107), .ZN(n15079) );
  CLKBUF_X1 U12335 ( .A(n11600), .Z(n11601) );
  AND2_X1 U12336 ( .A1(n15177), .A2(n14031), .ZN(n17225) );
  OR2_X1 U12337 ( .A1(n13999), .A2(n13998), .ZN(n20740) );
  AND2_X1 U12338 ( .A1(n14137), .A2(n21501), .ZN(n14138) );
  XNOR2_X1 U12339 ( .A(n13728), .B(n11576), .ZN(n14729) );
  NAND2_X1 U12340 ( .A1(n13727), .A2(n13750), .ZN(n14710) );
  NAND2_X1 U12341 ( .A1(n11491), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11493) );
  INV_X1 U12342 ( .A(n11489), .ZN(n14754) );
  NAND2_X1 U12343 ( .A1(n11102), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11142) );
  OAI21_X1 U12344 ( .B1(n14975), .B2(n14974), .A(n14973), .ZN(n15365) );
  AND2_X1 U12345 ( .A1(n15094), .A2(n15093), .ZN(n20668) );
  XNOR2_X1 U12346 ( .A(n14736), .B(n14735), .ZN(n15376) );
  AOI21_X1 U12347 ( .B1(n15368), .B2(n13062), .A(n15379), .ZN(n13742) );
  OAI21_X1 U12348 ( .B1(n15203), .B2(n15333), .A(n10397), .ZN(n10396) );
  OR2_X1 U12349 ( .A1(n15419), .A2(n15218), .ZN(n15400) );
  INV_X1 U12350 ( .A(n9753), .ZN(n15408) );
  INV_X1 U12351 ( .A(n10393), .ZN(n15243) );
  OAI21_X1 U12352 ( .B1(n15251), .B2(n10897), .A(n15333), .ZN(n10393) );
  NAND2_X1 U12353 ( .A1(n9631), .A2(n15454), .ZN(n15446) );
  XNOR2_X1 U12354 ( .A(n11598), .B(n11597), .ZN(n15491) );
  NAND2_X1 U12355 ( .A1(n10078), .A2(n10077), .ZN(n11595) );
  XNOR2_X1 U12356 ( .A(n9823), .B(n9703), .ZN(n15503) );
  NOR2_X1 U12357 ( .A1(n15296), .A2(n9985), .ZN(n9823) );
  NAND2_X1 U12358 ( .A1(n20811), .A2(n15464), .ZN(n9755) );
  NAND2_X1 U12359 ( .A1(n15302), .A2(n10880), .ZN(n15318) );
  NAND2_X1 U12360 ( .A1(n10083), .A2(n11593), .ZN(n9824) );
  NAND2_X1 U12361 ( .A1(n10206), .A2(n10864), .ZN(n17234) );
  INV_X1 U12362 ( .A(n15360), .ZN(n20786) );
  OR2_X1 U12363 ( .A1(n15428), .A2(n14130), .ZN(n20811) );
  OR2_X1 U12364 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14130), .ZN(
        n20810) );
  XNOR2_X1 U12365 ( .A(n10819), .B(n10984), .ZN(n20889) );
  INV_X1 U12366 ( .A(n11574), .ZN(n14429) );
  INV_X1 U12367 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20818) );
  OAI21_X1 U12368 ( .B1(n14416), .B2(n17285), .A(n20973), .ZN(n20817) );
  CLKBUF_X1 U12369 ( .A(n10933), .Z(n10934) );
  NOR2_X1 U12370 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20624) );
  INV_X1 U12371 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14519) );
  INV_X1 U12372 ( .A(n20851), .ZN(n20859) );
  OAI22_X1 U12373 ( .A1(n14516), .A2(n14515), .B1(n21154), .B2(n20970), .ZN(
        n20858) );
  INV_X1 U12374 ( .A(n20920), .ZN(n20891) );
  OAI21_X1 U12375 ( .B1(n20898), .B2(n20896), .A(n20895), .ZN(n20923) );
  OAI21_X1 U12376 ( .B1(n20939), .B2(n20937), .A(n20936), .ZN(n20965) );
  OAI21_X1 U12377 ( .B1(n20992), .B2(n20975), .A(n21301), .ZN(n20994) );
  INV_X1 U12378 ( .A(n21016), .ZN(n21019) );
  INV_X1 U12379 ( .A(n21087), .ZN(n21077) );
  INV_X1 U12380 ( .A(n21135), .ZN(n21138) );
  OAI21_X1 U12381 ( .B1(n21156), .B2(n21153), .A(n21152), .ZN(n21180) );
  NAND2_X1 U12382 ( .A1(n20854), .A2(n10587), .ZN(n21250) );
  OAI211_X1 U12383 ( .C1(n21223), .C2(n21222), .A(n21301), .B(n21221), .ZN(
        n21259) );
  INV_X1 U12384 ( .A(n21285), .ZN(n21288) );
  INV_X1 U12385 ( .A(n21217), .ZN(n21343) );
  INV_X1 U12386 ( .A(n21230), .ZN(n21356) );
  INV_X1 U12387 ( .A(n21234), .ZN(n21362) );
  INV_X1 U12388 ( .A(n21238), .ZN(n21368) );
  INV_X1 U12389 ( .A(n21242), .ZN(n21374) );
  INV_X1 U12390 ( .A(n21246), .ZN(n21380) );
  INV_X1 U12391 ( .A(n21250), .ZN(n21386) );
  INV_X1 U12392 ( .A(n21391), .ZN(n21397) );
  INV_X1 U12393 ( .A(n21256), .ZN(n21396) );
  INV_X1 U12394 ( .A(n21503), .ZN(n17172) );
  AND2_X1 U12395 ( .A1(n21403), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n17170) );
  NOR2_X1 U12396 ( .A1(n11005), .A2(n21403), .ZN(n17280) );
  INV_X1 U12397 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21222) );
  OAI211_X1 U12398 ( .C1(n16802), .C2(n9786), .A(n9785), .B(n9784), .ZN(n20607) );
  NAND2_X1 U12399 ( .A1(n16799), .A2(n16800), .ZN(n9784) );
  NAND2_X1 U12400 ( .A1(n9786), .A2(n16801), .ZN(n9785) );
  NAND2_X1 U12401 ( .A1(n12574), .A2(n13810), .ZN(n13794) );
  NAND2_X1 U12402 ( .A1(n12763), .A2(n10314), .ZN(n15671) );
  AOI21_X1 U12403 ( .B1(n12762), .B2(n12761), .A(n12760), .ZN(n10314) );
  NAND2_X1 U12404 ( .A1(n12688), .A2(n10040), .ZN(n12751) );
  NAND2_X1 U12405 ( .A1(n15743), .A2(n16199), .ZN(n15725) );
  OR2_X1 U12406 ( .A1(n12631), .A2(n12630), .ZN(n15803) );
  BUF_X1 U12407 ( .A(n14700), .Z(n19764) );
  OR3_X1 U12408 ( .A1(n19594), .A2(n19771), .A3(n14681), .ZN(n19778) );
  NAND2_X1 U12409 ( .A1(n19594), .A2(n14618), .ZN(n19767) );
  AND2_X1 U12410 ( .A1(n19594), .A2(n14615), .ZN(n19754) );
  OR2_X1 U12411 ( .A1(n11878), .A2(n11877), .ZN(n15940) );
  OR2_X1 U12412 ( .A1(n15990), .A2(n15924), .ZN(n15955) );
  OR2_X1 U12413 ( .A1(n11831), .A2(n11830), .ZN(n15960) );
  OR2_X1 U12414 ( .A1(n11841), .A2(n11840), .ZN(n15968) );
  OR2_X1 U12415 ( .A1(n11807), .A2(n11806), .ZN(n15972) );
  NOR2_X1 U12416 ( .A1(n15977), .A2(n15951), .ZN(n15978) );
  OR2_X1 U12417 ( .A1(n11819), .A2(n11818), .ZN(n15980) );
  NOR2_X1 U12418 ( .A1(n15990), .A2(n14451), .ZN(n15991) );
  INV_X1 U12419 ( .A(n15975), .ZN(n15992) );
  XNOR2_X1 U12420 ( .A(n10195), .B(n14606), .ZN(n14614) );
  NOR2_X1 U12421 ( .A1(n15884), .A2(n15883), .ZN(n15882) );
  AND2_X1 U12422 ( .A1(n11993), .A2(n11994), .ZN(n15884) );
  INV_X1 U12423 ( .A(n19799), .ZN(n16077) );
  NOR2_X1 U12424 ( .A1(n13879), .A2(n16713), .ZN(n19799) );
  AND2_X1 U12425 ( .A1(n19832), .A2(n9731), .ZN(n19798) );
  INV_X1 U12426 ( .A(n10368), .ZN(n13888) );
  AOI21_X1 U12427 ( .B1(n10373), .B2(n9625), .A(n12310), .ZN(n10368) );
  NAND2_X1 U12428 ( .A1(n16083), .A2(n10374), .ZN(n10373) );
  AOI21_X2 U12429 ( .B1(n13808), .B2(n13129), .A(n20481), .ZN(n19832) );
  OR2_X1 U12430 ( .A1(n16654), .A2(n13907), .ZN(n16745) );
  INV_X1 U12431 ( .A(n19832), .ZN(n19813) );
  INV_X1 U12432 ( .A(n19821), .ZN(n19824) );
  OAI21_X1 U12433 ( .B1(n19836), .B2(n19835), .A(n19834), .ZN(n19837) );
  INV_X2 U12434 ( .A(n19852), .ZN(n19903) );
  NAND2_X1 U12435 ( .A1(n13068), .A2(n10340), .ZN(n13069) );
  NOR2_X1 U12436 ( .A1(n19941), .A2(n10361), .ZN(n10360) );
  INV_X1 U12437 ( .A(n10364), .ZN(n10361) );
  INV_X1 U12438 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16169) );
  AND2_X1 U12439 ( .A1(n10301), .A2(n10303), .ZN(n9933) );
  AND2_X1 U12440 ( .A1(n10304), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10303) );
  INV_X1 U12441 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16257) );
  INV_X1 U12442 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19748) );
  INV_X1 U12443 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19934) );
  INV_X1 U12444 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19949) );
  INV_X1 U12445 ( .A(n19939), .ZN(n19917) );
  XNOR2_X1 U12446 ( .A(n9847), .B(n13066), .ZN(n13648) );
  NAND2_X1 U12447 ( .A1(n10363), .A2(n9744), .ZN(n10362) );
  NAND2_X1 U12448 ( .A1(n16366), .A2(n13635), .ZN(n10364) );
  XNOR2_X1 U12449 ( .A(n12777), .B(n12776), .ZN(n13164) );
  OAI21_X1 U12450 ( .B1(n9778), .B2(n16375), .A(n9776), .ZN(n9775) );
  INV_X1 U12451 ( .A(n16379), .ZN(n9778) );
  XNOR2_X1 U12452 ( .A(n10119), .B(n9639), .ZN(n16382) );
  OAI21_X1 U12453 ( .B1(n16126), .B2(n10121), .A(n10120), .ZN(n10119) );
  NAND2_X1 U12454 ( .A1(n16114), .A2(n9607), .ZN(n10120) );
  NAND2_X1 U12455 ( .A1(n16248), .A2(n10135), .ZN(n10115) );
  NAND2_X1 U12456 ( .A1(n10258), .A2(n13575), .ZN(n14562) );
  OAI21_X1 U12457 ( .B1(n16241), .B2(n9996), .A(n9993), .ZN(n10258) );
  AOI21_X1 U12458 ( .B1(n9995), .B2(n13574), .A(n9994), .ZN(n9993) );
  XNOR2_X1 U12459 ( .A(n10049), .B(n10048), .ZN(n16502) );
  INV_X1 U12460 ( .A(n16223), .ZN(n10048) );
  NAND2_X1 U12461 ( .A1(n10265), .A2(n16231), .ZN(n10049) );
  NAND2_X1 U12462 ( .A1(n9997), .A2(n9995), .ZN(n10265) );
  INV_X1 U12463 ( .A(n16284), .ZN(n13581) );
  NAND2_X1 U12464 ( .A1(n9997), .A2(n16238), .ZN(n16230) );
  NAND2_X1 U12465 ( .A1(n16578), .A2(n13670), .ZN(n16543) );
  NAND2_X1 U12466 ( .A1(n12316), .A2(n10376), .ZN(n13979) );
  NAND2_X1 U12467 ( .A1(n9783), .A2(n16549), .ZN(n16576) );
  INV_X1 U12468 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16593) );
  AND2_X1 U12469 ( .A1(n9892), .A2(n9894), .ZN(n16327) );
  OR2_X1 U12470 ( .A1(n16083), .A2(n16084), .ZN(n10371) );
  NAND2_X1 U12471 ( .A1(n13141), .A2(n13140), .ZN(n14554) );
  INV_X1 U12472 ( .A(n16480), .ZN(n14559) );
  INV_X1 U12473 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20604) );
  INV_X1 U12474 ( .A(n14151), .ZN(n20597) );
  INV_X1 U12475 ( .A(n16744), .ZN(n19968) );
  OAI21_X1 U12476 ( .B1(n20023), .B2(n20575), .A(n20022), .ZN(n20043) );
  OAI21_X1 U12477 ( .B1(n20084), .B2(n20057), .A(n20056), .ZN(n20077) );
  OAI21_X1 U12478 ( .B1(n20136), .B2(n20581), .A(n20121), .ZN(n20138) );
  AOI21_X1 U12479 ( .B1(n20392), .B2(n20116), .A(n20118), .ZN(n20137) );
  OAI21_X1 U12480 ( .B1(n16719), .B2(n20114), .A(n16718), .ZN(n20158) );
  AND2_X1 U12481 ( .A1(n20181), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20213) );
  NOR2_X1 U12482 ( .A1(n20184), .A2(n20180), .ZN(n20201) );
  NOR2_X1 U12483 ( .A1(n20295), .A2(n20382), .ZN(n10125) );
  OAI21_X1 U12484 ( .B1(n20307), .B2(n20575), .A(n20304), .ZN(n20334) );
  AOI21_X1 U12485 ( .B1(n20392), .B2(n16757), .A(n16756), .ZN(n20357) );
  OAI21_X1 U12486 ( .B1(n16769), .B2(n20575), .A(n16768), .ZN(n20377) );
  INV_X1 U12487 ( .A(n20401), .ZN(n20434) );
  INV_X1 U12488 ( .A(n20404), .ZN(n20441) );
  INV_X1 U12489 ( .A(n20407), .ZN(n20448) );
  INV_X1 U12490 ( .A(n20410), .ZN(n20455) );
  INV_X1 U12491 ( .A(n20413), .ZN(n20462) );
  INV_X1 U12492 ( .A(n20419), .ZN(n20373) );
  INV_X1 U12493 ( .A(n20425), .ZN(n20376) );
  INV_X1 U12494 ( .A(n20384), .ZN(n20473) );
  INV_X1 U12495 ( .A(n19972), .ZN(n20475) );
  NOR2_X1 U12496 ( .A1(n16783), .A2(n16782), .ZN(n20471) );
  NAND2_X2 U12497 ( .A1(n20618), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20558) );
  NAND2_X1 U12498 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20496), .ZN(n20619) );
  NAND2_X1 U12499 ( .A1(n10225), .A2(n17441), .ZN(n10223) );
  OAI21_X1 U12500 ( .B1(n17528), .B2(n17517), .A(n10224), .ZN(n10226) );
  NOR2_X1 U12501 ( .A1(n17516), .A2(n17517), .ZN(n17515) );
  AND2_X1 U12502 ( .A1(n17528), .A2(n14217), .ZN(n17516) );
  NOR2_X1 U12503 ( .A1(n17562), .A2(n17775), .ZN(n17553) );
  NOR2_X1 U12504 ( .A1(n17775), .A2(n13766), .ZN(n13767) );
  NOR2_X1 U12505 ( .A1(n13767), .A2(n18519), .ZN(n17446) );
  NOR2_X1 U12506 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17626), .ZN(n17609) );
  INV_X1 U12507 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17754) );
  NOR2_X1 U12508 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17785), .ZN(n17759) );
  INV_X1 U12509 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17787) );
  OR2_X1 U12510 ( .A1(n13777), .A2(n13776), .ZN(n17812) );
  INV_X1 U12511 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n16927) );
  OR2_X1 U12512 ( .A1(n19586), .A2(n13772), .ZN(n17816) );
  NAND2_X1 U12513 ( .A1(n9962), .A2(n9961), .ZN(n9960) );
  NOR2_X1 U12514 ( .A1(n17822), .A2(n17825), .ZN(n9962) );
  INV_X1 U12515 ( .A(n9961), .ZN(n9959) );
  NOR2_X1 U12516 ( .A1(n17927), .A2(n17823), .ZN(n17890) );
  NOR2_X1 U12517 ( .A1(n18026), .A2(n9958), .ZN(n17972) );
  NAND2_X1 U12518 ( .A1(n9740), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U12519 ( .A1(n9570), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n18026) );
  NOR2_X1 U12520 ( .A1(n9978), .A2(n17705), .ZN(n9977) );
  INV_X1 U12521 ( .A(n9980), .ZN(n9978) );
  AND3_X1 U12522 ( .A1(n9957), .A2(n9956), .A3(n9955), .ZN(n9953) );
  NAND2_X1 U12523 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n9956) );
  NOR2_X1 U12524 ( .A1(n18152), .A2(n17734), .ZN(n18121) );
  NAND2_X1 U12525 ( .A1(n18180), .A2(n19024), .ZN(n18163) );
  INV_X1 U12526 ( .A(n18177), .ZN(n18171) );
  NAND2_X1 U12527 ( .A1(n18206), .A2(n9618), .ZN(n18194) );
  NAND2_X1 U12528 ( .A1(n18206), .A2(P3_EAX_REG_27__SCAN_IN), .ZN(n18202) );
  NOR2_X1 U12529 ( .A1(n18331), .A2(n18211), .ZN(n18206) );
  INV_X1 U12530 ( .A(n18216), .ZN(n18212) );
  NAND2_X1 U12531 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n18212), .ZN(n18211) );
  NOR2_X1 U12532 ( .A1(n19024), .A2(n18221), .ZN(n18217) );
  NOR2_X1 U12533 ( .A1(n9968), .A2(n9964), .ZN(n9963) );
  INV_X1 U12534 ( .A(n9966), .ZN(n9964) );
  NAND2_X1 U12535 ( .A1(n9969), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12536 ( .A1(n9638), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n18221) );
  NOR2_X1 U12537 ( .A1(n18183), .A2(n18301), .ZN(n18296) );
  INV_X1 U12538 ( .A(n13306), .ZN(n18305) );
  OR2_X1 U12539 ( .A1(n13284), .A2(n13283), .ZN(n18308) );
  AND2_X1 U12540 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n14287), .ZN(n18315) );
  NOR3_X1 U12541 ( .A1(n14278), .A2(n18372), .A3(n18300), .ZN(n14287) );
  AOI22_X1 U12542 ( .A1(n19568), .A2(n14209), .B1(n14208), .B2(n17005), .ZN(
        n18183) );
  INV_X1 U12543 ( .A(n18318), .ZN(n18309) );
  NAND2_X1 U12546 ( .A1(n17574), .A2(n10229), .ZN(n10441) );
  AND2_X1 U12547 ( .A1(n9699), .A2(n10232), .ZN(n10229) );
  INV_X1 U12548 ( .A(n18498), .ZN(n10232) );
  NOR2_X2 U12549 ( .A1(n18571), .A2(n18572), .ZN(n17574) );
  INV_X1 U12550 ( .A(n13555), .ZN(n18843) );
  INV_X1 U12551 ( .A(n18529), .ZN(n18622) );
  INV_X1 U12552 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17721) );
  NOR2_X1 U12553 ( .A1(n17713), .A2(n17721), .ZN(n18637) );
  INV_X2 U12554 ( .A(n19351), .ZN(n19180) );
  INV_X1 U12555 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17713) );
  NOR2_X1 U12556 ( .A1(n10214), .A2(n17761), .ZN(n18701) );
  INV_X1 U12557 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19451) );
  NOR4_X1 U12558 ( .A1(n16982), .A2(n18736), .A3(n16981), .A4(n16980), .ZN(
        n18728) );
  NAND2_X1 U12559 ( .A1(n13346), .A2(n13347), .ZN(n16893) );
  INV_X1 U12560 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21628) );
  NAND2_X1 U12561 ( .A1(n18660), .A2(n10158), .ZN(n10160) );
  INV_X1 U12562 ( .A(n18808), .ZN(n18809) );
  NAND2_X1 U12563 ( .A1(n13335), .A2(n18670), .ZN(n18632) );
  NAND2_X1 U12564 ( .A1(n14110), .A2(n19568), .ZN(n18888) );
  OR2_X1 U12565 ( .A1(n14161), .A2(n14109), .ZN(n14110) );
  NAND2_X1 U12566 ( .A1(n10154), .A2(n13287), .ZN(n14302) );
  NAND2_X1 U12567 ( .A1(n18697), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10154) );
  INV_X1 U12568 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19430) );
  INV_X1 U12569 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14362) );
  INV_X1 U12570 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19412) );
  NOR2_X1 U12571 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19584) );
  NOR2_X1 U12572 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19552), .ZN(
        n19444) );
  NOR2_X1 U12573 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19452), .ZN(n19456) );
  NAND2_X1 U12574 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n19572) );
  INV_X1 U12575 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19479) );
  INV_X2 U12576 ( .A(n19581), .ZN(n19583) );
  NOR2_X1 U12577 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13763), .ZN(n17393)
         );
  CLKBUF_X1 U12578 ( .A(n17393), .Z(n17405) );
  INV_X1 U12579 ( .A(n9915), .ZN(n20694) );
  OAI211_X1 U12580 ( .C1(n20691), .C2(n20783), .A(n9917), .B(n9916), .ZN(n9915) );
  INV_X1 U12581 ( .A(n9855), .ZN(n9854) );
  AND2_X1 U12582 ( .A1(n13631), .A2(n13630), .ZN(n13632) );
  AND2_X1 U12583 ( .A1(n15404), .A2(n9718), .ZN(n9856) );
  NAND2_X1 U12584 ( .A1(n9754), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15470) );
  NAND2_X1 U12585 ( .A1(n10252), .A2(n10248), .ZN(P2_U2826) );
  INV_X1 U12586 ( .A(n15620), .ZN(n10252) );
  AOI21_X1 U12587 ( .B1(n15621), .B2(n15622), .A(n10249), .ZN(n10248) );
  NAND2_X1 U12588 ( .A1(n10022), .A2(n13686), .ZN(P2_U2858) );
  NAND2_X1 U12589 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U12590 ( .B1(n16360), .B2(n16081), .A(n12392), .ZN(n12393) );
  INV_X1 U12591 ( .A(n9794), .ZN(n9793) );
  OAI21_X1 U12592 ( .B1(n16373), .B2(n17292), .A(n16109), .ZN(n9794) );
  INV_X1 U12593 ( .A(n10170), .ZN(n10169) );
  OAI21_X1 U12594 ( .B1(n16397), .B2(n19941), .A(n10180), .ZN(n10170) );
  AOI21_X1 U12595 ( .B1(n16146), .B2(n19946), .A(n16145), .ZN(n10180) );
  AOI21_X1 U12596 ( .B1(n16427), .B2(n16335), .A(n16166), .ZN(n16167) );
  INV_X1 U12597 ( .A(n13692), .ZN(n9943) );
  NAND2_X1 U12598 ( .A1(n9569), .A2(n19936), .ZN(n9817) );
  NAND2_X1 U12599 ( .A1(n10064), .A2(n19936), .ZN(n10063) );
  AOI211_X1 U12600 ( .C1(n16369), .C2(n19952), .A(n16368), .B(n16367), .ZN(
        n16372) );
  NAND2_X1 U12601 ( .A1(n9796), .A2(n19962), .ZN(n9795) );
  OAI21_X1 U12602 ( .B1(n16408), .B2(n16648), .A(n10150), .ZN(P2_U3020) );
  INV_X1 U12603 ( .A(n9827), .ZN(n10150) );
  OAI21_X1 U12604 ( .B1(n16397), .B2(n19967), .A(n10151), .ZN(n9827) );
  AOI21_X1 U12605 ( .B1(n16407), .B2(n16645), .A(n16406), .ZN(n10151) );
  OAI21_X1 U12606 ( .B1(n16417), .B2(n16648), .A(n10007), .ZN(P2_U3021) );
  INV_X1 U12607 ( .A(n10008), .ZN(n10007) );
  OAI211_X1 U12608 ( .C1(n13693), .C2(n19967), .A(n13677), .B(n10016), .ZN(
        P2_U3025) );
  NAND2_X1 U12609 ( .A1(n13687), .A2(n19962), .ZN(n10016) );
  NOR2_X1 U12610 ( .A1(n16465), .A2(n16464), .ZN(n9788) );
  NAND2_X1 U12611 ( .A1(n16466), .A2(n16603), .ZN(n9790) );
  NAND2_X1 U12612 ( .A1(n9569), .A2(n19962), .ZN(n9789) );
  INV_X1 U12613 ( .A(n10064), .ZN(n16479) );
  OAI21_X1 U12614 ( .B1(n17459), .B2(n9729), .A(n10233), .ZN(P3_U2640) );
  AOI21_X1 U12615 ( .B1(n17466), .B2(n17830), .A(n10234), .ZN(n10233) );
  NAND2_X1 U12616 ( .A1(n10238), .A2(n10235), .ZN(n10234) );
  NOR2_X1 U12617 ( .A1(n18264), .A2(n18428), .ZN(n18260) );
  NAND2_X1 U12618 ( .A1(n13527), .A2(n18681), .ZN(n13573) );
  NAND2_X1 U12619 ( .A1(n9883), .A2(n9882), .ZN(n9881) );
  NAND2_X1 U12620 ( .A1(n9880), .A2(n9879), .ZN(n9878) );
  AOI21_X1 U12621 ( .B1(n18456), .B2(n18443), .A(n10059), .ZN(n10058) );
  OAI21_X1 U12622 ( .B1(n18733), .B2(n18653), .A(n10268), .ZN(P3_U2803) );
  AOI21_X1 U12623 ( .B1(n18455), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10270), .ZN(n10269) );
  NAND2_X1 U12624 ( .A1(n18456), .A2(n13355), .ZN(n10271) );
  INV_X2 U12625 ( .A(n13921), .ZN(n11323) );
  AND2_X2 U12626 ( .A1(n10474), .A2(n15593), .ZN(n10622) );
  AND2_X2 U12627 ( .A1(n16740), .A2(n20581), .ZN(n12327) );
  AND3_X1 U12628 ( .A1(n16157), .A2(n16137), .A3(n16179), .ZN(n9588) );
  AND2_X1 U12629 ( .A1(n14369), .A2(n9700), .ZN(n15894) );
  INV_X1 U12630 ( .A(n13168), .ZN(n18138) );
  INV_X1 U12631 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10276) );
  OR2_X1 U12632 ( .A1(n10256), .A2(n10015), .ZN(n9590) );
  NAND2_X1 U12633 ( .A1(n14563), .A2(n10377), .ZN(n16058) );
  OR2_X1 U12634 ( .A1(n15287), .A2(n10081), .ZN(n9592) );
  NAND2_X1 U12635 ( .A1(n12688), .A2(n12746), .ZN(n12744) );
  NAND2_X1 U12636 ( .A1(n14369), .A2(n9689), .ZN(n15916) );
  OR2_X1 U12637 ( .A1(n14118), .A2(n10385), .ZN(n14223) );
  NAND2_X1 U12638 ( .A1(n10244), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9594) );
  AND2_X1 U12639 ( .A1(n9979), .A2(n9977), .ZN(n9595) );
  AND2_X1 U12640 ( .A1(n15280), .A2(n9738), .ZN(n9596) );
  AND3_X1 U12641 ( .A1(n9842), .A2(n18565), .A3(n9840), .ZN(n9597) );
  NAND2_X1 U12642 ( .A1(n11262), .A2(n10423), .ZN(n14862) );
  NAND2_X1 U12643 ( .A1(n10410), .A2(n12838), .ZN(n15927) );
  OR2_X1 U12644 ( .A1(n9661), .A2(n9787), .ZN(n9598) );
  NOR2_X1 U12645 ( .A1(n15740), .A2(n9660), .ZN(n15695) );
  INV_X1 U12646 ( .A(n13339), .ZN(n9841) );
  INV_X1 U12647 ( .A(n15244), .ZN(n9989) );
  OR2_X1 U12648 ( .A1(n12609), .A2(n10320), .ZN(n12608) );
  AND2_X1 U12649 ( .A1(n16187), .A2(n16335), .ZN(n9599) );
  XNOR2_X1 U12650 ( .A(n10391), .B(n13641), .ZN(n14695) );
  OR2_X1 U12651 ( .A1(n9619), .A2(n10316), .ZN(n9600) );
  NOR2_X1 U12652 ( .A1(n12278), .A2(n12277), .ZN(n12588) );
  AND2_X1 U12653 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n9601) );
  AND2_X1 U12654 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n9602) );
  AND2_X1 U12655 ( .A1(n12426), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n9603) );
  INV_X1 U12656 ( .A(n12426), .ZN(n14063) );
  INV_X1 U12657 ( .A(n12418), .ZN(n12425) );
  AND2_X1 U12658 ( .A1(n16652), .A2(n12401), .ZN(n12418) );
  AND2_X1 U12659 ( .A1(n9676), .A2(n10795), .ZN(n9604) );
  NAND2_X1 U12660 ( .A1(n9576), .A2(n13127), .ZN(n9605) );
  INV_X1 U12661 ( .A(n13332), .ZN(n9838) );
  AND2_X1 U12662 ( .A1(n9596), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9606) );
  AND2_X1 U12663 ( .A1(n12601), .A2(n12605), .ZN(n9607) );
  AND2_X1 U12664 ( .A1(n9813), .A2(n10132), .ZN(n9608) );
  NAND2_X1 U12665 ( .A1(n12718), .A2(n9698), .ZN(n9609) );
  AND2_X1 U12666 ( .A1(n12958), .A2(n12954), .ZN(n9610) );
  AND2_X1 U12667 ( .A1(n10376), .A2(n10375), .ZN(n9611) );
  INV_X1 U12668 ( .A(n15822), .ZN(n14236) );
  INV_X1 U12669 ( .A(n9808), .ZN(n16740) );
  NAND2_X2 U12670 ( .A1(n11625), .A2(n11626), .ZN(n9808) );
  INV_X1 U12671 ( .A(n10742), .ZN(n11528) );
  INV_X1 U12672 ( .A(n10634), .ZN(n10742) );
  INV_X1 U12673 ( .A(n16639), .ZN(n19952) );
  NAND2_X1 U12674 ( .A1(n12316), .A2(n12315), .ZN(n13882) );
  AND2_X1 U12675 ( .A1(n10227), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9612) );
  AND2_X1 U12676 ( .A1(n9728), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9613) );
  AND2_X1 U12677 ( .A1(n9612), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9614) );
  AND2_X1 U12678 ( .A1(n10416), .A2(n10414), .ZN(n9615) );
  INV_X1 U12679 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20509) );
  INV_X1 U12680 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18685) );
  INV_X1 U12681 ( .A(n10321), .ZN(n14890) );
  INV_X1 U12682 ( .A(n12156), .ZN(n10193) );
  AND2_X1 U12683 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9616) );
  AND2_X1 U12684 ( .A1(n9616), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9617) );
  AND2_X1 U12685 ( .A1(n9970), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n9618) );
  BUF_X2 U12686 ( .A(n12779), .Z(n12792) );
  OR2_X1 U12687 ( .A1(n15061), .A2(n10322), .ZN(n9619) );
  AND2_X2 U12688 ( .A1(n12037), .A2(n11656), .ZN(n11851) );
  NAND2_X1 U12689 ( .A1(n10709), .A2(n20862), .ZN(n14504) );
  NOR2_X1 U12690 ( .A1(n14646), .A2(n19671), .ZN(n14624) );
  NAND2_X1 U12691 ( .A1(n12700), .A2(n12592), .ZN(n12624) );
  INV_X1 U12692 ( .A(n10293), .ZN(n13799) );
  XNOR2_X1 U12693 ( .A(n10186), .B(n10185), .ZN(n15868) );
  INV_X1 U12694 ( .A(n20778), .ZN(n9918) );
  NAND2_X1 U12695 ( .A1(n10380), .A2(n12362), .ZN(n15684) );
  OR2_X1 U12696 ( .A1(n14922), .A2(n9926), .ZN(n14910) );
  AND2_X1 U12697 ( .A1(n14563), .A2(n14566), .ZN(n14564) );
  NAND2_X1 U12698 ( .A1(n10292), .A2(n10293), .ZN(n13118) );
  NOR2_X1 U12699 ( .A1(n14629), .A2(n12891), .ZN(n14625) );
  AND2_X2 U12700 ( .A1(n10469), .A2(n15593), .ZN(n10577) );
  NAND2_X1 U12701 ( .A1(n16174), .A2(n16173), .ZN(n16175) );
  OR2_X1 U12702 ( .A1(n15740), .A2(n10413), .ZN(n9621) );
  AND2_X1 U12703 ( .A1(n13181), .A2(n13180), .ZN(n13297) );
  NAND2_X1 U12704 ( .A1(n9593), .A2(n9761), .ZN(n9622) );
  AND2_X1 U12705 ( .A1(n18206), .A2(n9970), .ZN(n9623) );
  NAND2_X1 U12706 ( .A1(n17574), .A2(n10230), .ZN(n9624) );
  AND2_X1 U12707 ( .A1(n10372), .A2(n13878), .ZN(n9625) );
  AND2_X1 U12708 ( .A1(n11262), .A2(n10286), .ZN(n14848) );
  NOR2_X1 U12709 ( .A1(n15932), .A2(n10408), .ZN(n14567) );
  AND2_X1 U12710 ( .A1(n10277), .A2(n20968), .ZN(n9627) );
  AND2_X1 U12711 ( .A1(n14063), .A2(n9942), .ZN(n9628) );
  NAND2_X1 U12712 ( .A1(n11783), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n9629) );
  AND2_X1 U12713 ( .A1(n16313), .A2(n10302), .ZN(n9630) );
  NAND2_X1 U12714 ( .A1(n15580), .A2(n15433), .ZN(n9631) );
  INV_X1 U12715 ( .A(n9932), .ZN(n16206) );
  OR2_X1 U12716 ( .A1(n17927), .A2(n9960), .ZN(n9632) );
  AND2_X1 U12717 ( .A1(n10800), .A2(n10799), .ZN(n9633) );
  AND2_X1 U12718 ( .A1(n15297), .A2(n15289), .ZN(n9634) );
  AND2_X1 U12719 ( .A1(n10968), .A2(n10073), .ZN(n9635) );
  INV_X1 U12720 ( .A(n17996), .ZN(n18124) );
  AND2_X1 U12721 ( .A1(n9772), .A2(n9812), .ZN(n9636) );
  AND2_X1 U12722 ( .A1(n13207), .A2(n13206), .ZN(n9637) );
  AND2_X1 U12723 ( .A1(n9965), .A2(n9963), .ZN(n9638) );
  XOR2_X1 U12724 ( .A(n16116), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(
        n9639) );
  NOR2_X1 U12725 ( .A1(n14758), .A2(n13626), .ZN(n13697) );
  NAND2_X1 U12726 ( .A1(n13581), .A2(n10304), .ZN(n16224) );
  AND2_X1 U12727 ( .A1(n11750), .A2(n14370), .ZN(n14233) );
  AND4_X1 U12728 ( .A1(n13123), .A2(n11702), .A3(n9808), .A4(n19997), .ZN(
        n9640) );
  XOR2_X1 U12729 ( .A(n15353), .B(n15565), .Z(n9641) );
  NAND2_X1 U12730 ( .A1(n14637), .A2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14636) );
  NAND2_X1 U12731 ( .A1(n12619), .A2(n12684), .ZN(n12683) );
  AND2_X1 U12732 ( .A1(n10279), .A2(n10277), .ZN(n9642) );
  INV_X1 U12733 ( .A(n16380), .ZN(n9777) );
  AND2_X1 U12734 ( .A1(n12836), .A2(n10331), .ZN(n9643) );
  AND2_X1 U12735 ( .A1(n12840), .A2(n10333), .ZN(n9644) );
  AND2_X1 U12736 ( .A1(n12859), .A2(n10335), .ZN(n9645) );
  AND2_X1 U12737 ( .A1(n12844), .A2(n10341), .ZN(n9646) );
  AND2_X1 U12738 ( .A1(n12846), .A2(n10342), .ZN(n9647) );
  AND2_X1 U12739 ( .A1(n12863), .A2(n10343), .ZN(n9648) );
  OR2_X1 U12740 ( .A1(n18622), .A2(n18445), .ZN(n9649) );
  AND2_X1 U12741 ( .A1(n16140), .A2(n10176), .ZN(n9650) );
  AND2_X1 U12742 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n9651)
         );
  AND2_X1 U12743 ( .A1(n14063), .A2(n12411), .ZN(n9652) );
  INV_X1 U12744 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14393) );
  NAND2_X1 U12745 ( .A1(n10585), .A2(n10811), .ZN(n10617) );
  OR2_X1 U12746 ( .A1(n13585), .A2(n15741), .ZN(n15740) );
  INV_X1 U12747 ( .A(n15740), .ZN(n10415) );
  AND2_X1 U12748 ( .A1(n12180), .A2(n9807), .ZN(n9653) );
  AND3_X1 U12749 ( .A1(n11651), .A2(n9992), .A3(n9991), .ZN(n9654) );
  AND2_X1 U12750 ( .A1(n14977), .A2(n15095), .ZN(n9655) );
  INV_X1 U12751 ( .A(n13574), .ZN(n16239) );
  AND2_X1 U12752 ( .A1(n12738), .A2(n12832), .ZN(n13574) );
  NAND2_X1 U12753 ( .A1(n10037), .A2(n10035), .ZN(n10038) );
  AND4_X1 U12754 ( .A1(n13419), .A2(n13418), .A3(n13417), .A4(n13416), .ZN(
        n9656) );
  AND2_X1 U12755 ( .A1(n10594), .A2(n10811), .ZN(n10969) );
  AND2_X1 U12756 ( .A1(n10392), .A2(n10662), .ZN(n9657) );
  AND2_X1 U12757 ( .A1(n10091), .A2(n10984), .ZN(n9658) );
  AND2_X1 U12758 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n9659) );
  INV_X1 U12759 ( .A(n14388), .ZN(n14392) );
  NAND2_X1 U12760 ( .A1(n10418), .A2(n15713), .ZN(n9660) );
  AND2_X1 U12761 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n9661) );
  AND2_X1 U12762 ( .A1(n11693), .A2(n9808), .ZN(n9662) );
  AND2_X1 U12763 ( .A1(n13269), .A2(n13285), .ZN(n9663) );
  AND2_X1 U12764 ( .A1(n11648), .A2(n11647), .ZN(n9664) );
  AND2_X1 U12765 ( .A1(n13032), .A2(n10074), .ZN(n9665) );
  INV_X1 U12766 ( .A(n12412), .ZN(n10198) );
  OR2_X1 U12767 ( .A1(n13111), .A2(n19928), .ZN(n9666) );
  AND2_X1 U12768 ( .A1(n10958), .A2(n10959), .ZN(n9667) );
  AND3_X1 U12769 ( .A1(n13463), .A2(n13462), .A3(n13461), .ZN(n9668) );
  INV_X1 U12770 ( .A(n10155), .ZN(n9845) );
  AND2_X1 U12771 ( .A1(n10158), .A2(n13341), .ZN(n10155) );
  INV_X1 U12772 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19721) );
  AND2_X1 U12773 ( .A1(n13031), .A2(n9665), .ZN(n9669) );
  INV_X1 U12774 ( .A(n14530), .ZN(n15659) );
  OR2_X1 U12775 ( .A1(n18035), .A2(n18014), .ZN(n9670) );
  INV_X1 U12776 ( .A(n12426), .ZN(n10164) );
  AND2_X1 U12777 ( .A1(n9858), .A2(n9634), .ZN(n9671) );
  AND2_X1 U12778 ( .A1(n10010), .A2(n10009), .ZN(n9672) );
  OAI21_X1 U12779 ( .B1(n15671), .B2(n12523), .A(n16401), .ZN(n16147) );
  INV_X1 U12780 ( .A(n9996), .ZN(n9995) );
  NAND2_X1 U12781 ( .A1(n16232), .A2(n16238), .ZN(n9996) );
  XNOR2_X1 U12782 ( .A(n12773), .B(n12771), .ZN(n15616) );
  NAND2_X1 U12783 ( .A1(n13692), .A2(n13672), .ZN(n9673) );
  NAND2_X1 U12784 ( .A1(n16141), .A2(n9616), .ZN(n16110) );
  AND2_X1 U12785 ( .A1(n19945), .A2(n16665), .ZN(n9674) );
  OR2_X1 U12786 ( .A1(n20305), .A2(n12403), .ZN(n9675) );
  AND2_X1 U12787 ( .A1(n10854), .A2(n10785), .ZN(n9676) );
  OR2_X1 U12788 ( .A1(n12753), .A2(n16186), .ZN(n16179) );
  NOR2_X1 U12789 ( .A1(n15891), .A2(n15890), .ZN(n15889) );
  OR2_X1 U12790 ( .A1(n10810), .A2(n10736), .ZN(n9677) );
  NAND2_X2 U12791 ( .A1(n9764), .A2(n9763), .ZN(n15607) );
  INV_X2 U12792 ( .A(n15607), .ZN(n16815) );
  OR2_X1 U12793 ( .A1(n10539), .A2(n10538), .ZN(n10811) );
  INV_X1 U12794 ( .A(n10811), .ZN(n10202) );
  NAND2_X1 U12795 ( .A1(n10770), .A2(n10769), .ZN(n10795) );
  AND2_X1 U12796 ( .A1(n18565), .A2(n13334), .ZN(n9678) );
  AND2_X2 U12797 ( .A1(n11977), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12288) );
  AND3_X1 U12798 ( .A1(n10708), .A2(n10440), .A3(n10422), .ZN(n9679) );
  AND2_X2 U12799 ( .A1(n11977), .A2(n11656), .ZN(n12282) );
  NAND2_X1 U12800 ( .A1(n12747), .A2(n13087), .ZN(n12688) );
  AND2_X1 U12801 ( .A1(n13791), .A2(n13793), .ZN(n9680) );
  AND2_X1 U12802 ( .A1(n10115), .A2(n10132), .ZN(n9681) );
  AND2_X1 U12803 ( .A1(n12614), .A2(n12523), .ZN(n9682) );
  OR2_X1 U12804 ( .A1(n18457), .A2(n10228), .ZN(n9683) );
  AND2_X1 U12805 ( .A1(n12796), .A2(n10329), .ZN(n9684) );
  AND2_X1 U12806 ( .A1(n9588), .A2(n10047), .ZN(n9685) );
  AND2_X1 U12807 ( .A1(n11699), .A2(n9808), .ZN(n9686) );
  AND2_X1 U12808 ( .A1(n9610), .A2(n9655), .ZN(n9687) );
  AND2_X1 U12809 ( .A1(n10288), .A2(n10289), .ZN(n9688) );
  INV_X1 U12810 ( .A(n10438), .ZN(n10132) );
  INV_X1 U12811 ( .A(n9894), .ZN(n9893) );
  INV_X1 U12812 ( .A(n10576), .ZN(n11468) );
  INV_X1 U12813 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9830) );
  NAND2_X1 U12814 ( .A1(n12955), .A2(n9610), .ZN(n14976) );
  INV_X1 U12815 ( .A(n10577), .ZN(n13921) );
  NOR2_X1 U12816 ( .A1(n14375), .A2(n14376), .ZN(n14452) );
  NOR2_X1 U12817 ( .A1(n9619), .A2(n14865), .ZN(n14851) );
  NAND2_X1 U12818 ( .A1(n14369), .A2(n11891), .ZN(n15919) );
  AND2_X1 U12819 ( .A1(n14667), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14665) );
  AND2_X1 U12820 ( .A1(n11891), .A2(n11902), .ZN(n9689) );
  NAND2_X1 U12821 ( .A1(n13141), .A2(n20609), .ZN(n19967) );
  INV_X1 U12822 ( .A(n19967), .ZN(n16603) );
  INV_X1 U12823 ( .A(n20968), .ZN(n9872) );
  NAND2_X1 U12824 ( .A1(n13335), .A2(n10056), .ZN(n9690) );
  NAND2_X1 U12825 ( .A1(n14624), .A2(n10429), .ZN(n9691) );
  AND2_X1 U12826 ( .A1(n14798), .A2(n14794), .ZN(n9692) );
  AND2_X1 U12827 ( .A1(n9692), .A2(n10328), .ZN(n9693) );
  NOR2_X1 U12828 ( .A1(n15086), .A2(n10312), .ZN(n14946) );
  NOR3_X1 U12829 ( .A1(n9619), .A2(n14865), .A3(n10315), .ZN(n14843) );
  NOR2_X1 U12830 ( .A1(n15932), .A2(n10411), .ZN(n14568) );
  NOR2_X1 U12831 ( .A1(n15086), .A2(n10309), .ZN(n14929) );
  AND2_X1 U12832 ( .A1(n13596), .A2(n13595), .ZN(n9694) );
  NOR2_X1 U12833 ( .A1(n10404), .A2(n10402), .ZN(n15779) );
  OR2_X1 U12834 ( .A1(n15061), .A2(n15052), .ZN(n9695) );
  AND2_X1 U12835 ( .A1(n15648), .A2(n14540), .ZN(n9696) );
  OR3_X1 U12836 ( .A1(n12013), .A2(n12012), .A3(n15886), .ZN(n9697) );
  AND2_X1 U12837 ( .A1(n12596), .A2(n10306), .ZN(n9698) );
  AND2_X1 U12838 ( .A1(n10230), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9699) );
  OAI21_X1 U12839 ( .B1(n18568), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10160), .ZN(n18555) );
  NAND2_X1 U12840 ( .A1(n10371), .A2(n10374), .ZN(n13877) );
  AND2_X1 U12841 ( .A1(n9689), .A2(n10197), .ZN(n9700) );
  AND2_X1 U12842 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9701) );
  XNOR2_X1 U12843 ( .A(n13579), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9702) );
  AND2_X1 U12844 ( .A1(n15298), .A2(n15297), .ZN(n9703) );
  INV_X1 U12845 ( .A(n12684), .ZN(n10044) );
  INV_X1 U12846 ( .A(n14404), .ZN(n17129) );
  AOI21_X1 U12847 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19452), .A(n14166), 
        .ZN(n14404) );
  NOR2_X1 U12848 ( .A1(n14259), .A2(n13553), .ZN(n18904) );
  AND2_X1 U12849 ( .A1(n14849), .A2(n10286), .ZN(n9704) );
  AND2_X1 U12850 ( .A1(n10429), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9705) );
  AND2_X2 U12851 ( .A1(n10811), .A2(n10607), .ZN(n12932) );
  AND2_X1 U12852 ( .A1(n13890), .A2(n19985), .ZN(n9706) );
  AND2_X1 U12853 ( .A1(n12856), .A2(n10337), .ZN(n9707) );
  AND2_X1 U12854 ( .A1(n12877), .A2(n10344), .ZN(n9708) );
  AND2_X1 U12855 ( .A1(n10040), .A2(n10042), .ZN(n9709) );
  AND2_X1 U12856 ( .A1(n10806), .A2(n12946), .ZN(n9710) );
  AND2_X1 U12857 ( .A1(n10799), .A2(n10201), .ZN(n9711) );
  OR2_X1 U12858 ( .A1(n12172), .A2(n12171), .ZN(n13890) );
  AND2_X1 U12859 ( .A1(n10876), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9712) );
  NOR2_X1 U12860 ( .A1(n15061), .A2(n10323), .ZN(n10321) );
  NOR3_X1 U12861 ( .A1(n9619), .A2(n14828), .A3(n10316), .ZN(n14814) );
  AND3_X1 U12862 ( .A1(n15333), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9713) );
  AND2_X1 U12863 ( .A1(n9693), .A2(n10327), .ZN(n9714) );
  AND2_X1 U12864 ( .A1(n9700), .A2(n11959), .ZN(n9715) );
  INV_X1 U12865 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n17474) );
  AND2_X1 U12866 ( .A1(n18847), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18810) );
  INV_X1 U12867 ( .A(n18810), .ZN(n10159) );
  NAND2_X1 U12868 ( .A1(n14498), .A2(n14497), .ZN(n9716) );
  AND2_X1 U12869 ( .A1(n20819), .A2(n20838), .ZN(n14078) );
  NAND2_X1 U12870 ( .A1(n15302), .A2(n10884), .ZN(n9985) );
  AND2_X1 U12871 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n9717) );
  INV_X1 U12872 ( .A(n10225), .ZN(n10224) );
  OAI21_X1 U12873 ( .B1(n14217), .B2(n17517), .A(n14217), .ZN(n10225) );
  OR2_X1 U12874 ( .A1(n15406), .A2(n15571), .ZN(n9718) );
  OR2_X1 U12875 ( .A1(n17517), .A2(n17506), .ZN(n9719) );
  AND2_X1 U12876 ( .A1(n13096), .A2(n9808), .ZN(n9720) );
  AND2_X1 U12877 ( .A1(n12585), .A2(n12497), .ZN(n9721) );
  AND2_X1 U12878 ( .A1(n10420), .A2(n10419), .ZN(n9722) );
  AND2_X1 U12879 ( .A1(n10377), .A2(n12352), .ZN(n9723) );
  AND2_X1 U12880 ( .A1(n9698), .A2(n12597), .ZN(n9724) );
  INV_X1 U12881 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15728) );
  INV_X1 U12882 ( .A(n12069), .ZN(n10032) );
  INV_X1 U12883 ( .A(n19941), .ZN(n16335) );
  OR2_X1 U12884 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n11573) );
  NAND2_X1 U12885 ( .A1(n9575), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n9725) );
  INV_X1 U12886 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9877) );
  INV_X1 U12887 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9902) );
  AND2_X1 U12888 ( .A1(n14256), .A2(n14255), .ZN(n14254) );
  NAND2_X1 U12889 ( .A1(n14254), .A2(n12950), .ZN(n14464) );
  INV_X1 U12890 ( .A(n10622), .ZN(n10718) );
  AND2_X1 U12891 ( .A1(n18431), .A2(n10227), .ZN(n9726) );
  OR2_X1 U12892 ( .A1(n10996), .A2(n10997), .ZN(n9727) );
  INV_X1 U12893 ( .A(n12047), .ZN(n10185) );
  AND2_X1 U12894 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9728) );
  INV_X1 U12895 ( .A(n12746), .ZN(n10041) );
  AND2_X1 U12896 ( .A1(n12778), .A2(n15871), .ZN(n19936) );
  NAND2_X1 U12897 ( .A1(n12955), .A2(n12954), .ZN(n14477) );
  XNOR2_X1 U12898 ( .A(n13074), .B(n13073), .ZN(n14623) );
  OR2_X1 U12899 ( .A1(n17738), .A2(n17460), .ZN(n9729) );
  NOR2_X1 U12900 ( .A1(n17446), .A2(n17775), .ZN(n9730) );
  AND2_X1 U12901 ( .A1(n12693), .A2(n9808), .ZN(n9731) );
  AND2_X1 U12902 ( .A1(n12888), .A2(n10345), .ZN(n9732) );
  NAND2_X1 U12903 ( .A1(n18158), .A2(P3_EBX_REG_6__SCAN_IN), .ZN(n18152) );
  INV_X1 U12904 ( .A(n18152), .ZN(n9979) );
  AND2_X1 U12905 ( .A1(n10056), .A2(n13336), .ZN(n9733) );
  NOR2_X1 U12906 ( .A1(n12893), .A2(n15643), .ZN(n9734) );
  AND2_X1 U12907 ( .A1(n9979), .A2(n9980), .ZN(n9735) );
  AND2_X1 U12908 ( .A1(n9734), .A2(n9613), .ZN(n9736) );
  INV_X1 U12909 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10228) );
  INV_X1 U12910 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10231) );
  INV_X1 U12911 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10057) );
  INV_X1 U12912 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9908) );
  INV_X1 U12913 ( .A(n20382), .ZN(n20575) );
  NOR2_X2 U12914 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20382) );
  AND2_X1 U12915 ( .A1(n12552), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9737) );
  INV_X1 U12916 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9911) );
  INV_X1 U12917 ( .A(n15865), .ZN(n10196) );
  AND2_X1 U12918 ( .A1(n10395), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9738) );
  AND2_X1 U12919 ( .A1(n9737), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9739) );
  NOR2_X1 U12920 ( .A1(n14553), .A2(n16551), .ZN(n10305) );
  AND2_X1 U12921 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .ZN(n9740) );
  AND2_X1 U12922 ( .A1(n12526), .A2(n9739), .ZN(n9741) );
  INV_X1 U12923 ( .A(n20480), .ZN(n10291) );
  INV_X1 U12924 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10157) );
  INV_X1 U12925 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10054) );
  AND2_X1 U12926 ( .A1(n15221), .A2(n13621), .ZN(n9742) );
  NAND2_X1 U12927 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18611) );
  INV_X1 U12928 ( .A(n18611), .ZN(n10222) );
  AND2_X1 U12929 ( .A1(n9617), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9743) );
  INV_X1 U12930 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n9967) );
  INV_X1 U12931 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9886) );
  AND2_X1 U12932 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9744) );
  INV_X1 U12933 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9914) );
  INV_X1 U12934 ( .A(n10897), .ZN(n10395) );
  AND2_X1 U12935 ( .A1(n9743), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9745) );
  OAI21_X1 U12936 ( .B1(n15226), .B2(n17244), .A(n15224), .ZN(n9855) );
  NOR2_X2 U12937 ( .A1(n17244), .A2(n14509), .ZN(n9746) );
  NOR2_X1 U12938 ( .A1(n17244), .A2(n14509), .ZN(n20852) );
  NAND2_X1 U12939 ( .A1(n21349), .A2(n11577), .ZN(n17244) );
  INV_X1 U12940 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19552) );
  INV_X1 U12941 ( .A(n21336), .ZN(n9747) );
  INV_X1 U12942 ( .A(n9747), .ZN(n9748) );
  AOI22_X2 U12943 ( .A1(DATAI_16_), .A2(n9567), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9746), .ZN(n21354) );
  AOI22_X2 U12944 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9746), .B1(DATAI_23_), 
        .B2(n9567), .ZN(n21402) );
  NOR3_X2 U12945 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19318), .A3(
        n19158), .ZN(n19173) );
  AND2_X2 U12946 ( .A1(n14684), .A2(n19985), .ZN(n13850) );
  NOR2_X1 U12947 ( .A1(n13788), .A2(n13795), .ZN(n14684) );
  NOR2_X1 U12948 ( .A1(n20004), .A2(n19997), .ZN(n9749) );
  NAND2_X1 U12949 ( .A1(n20397), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20004) );
  OR2_X2 U12950 ( .A1(n14037), .A2(n20626), .ZN(n13999) );
  NAND2_X2 U12951 ( .A1(n9750), .A2(n10967), .ZN(n14037) );
  NAND2_X1 U12952 ( .A1(n15417), .A2(n13051), .ZN(n9753) );
  INV_X1 U12953 ( .A(n15454), .ZN(n9754) );
  NAND2_X1 U12954 ( .A1(n13043), .A2(n9755), .ZN(n13047) );
  NOR2_X1 U12955 ( .A1(n10607), .A2(n14511), .ZN(n10616) );
  NAND2_X1 U12956 ( .A1(n10202), .A2(n14511), .ZN(n12945) );
  NAND2_X1 U12957 ( .A1(n14140), .A2(n14511), .ZN(n14137) );
  OR2_X4 U12958 ( .A1(n10583), .A2(n10582), .ZN(n14511) );
  AND2_X2 U12959 ( .A1(n10933), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10474) );
  AND2_X2 U12960 ( .A1(n9825), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9923) );
  OAI211_X1 U12961 ( .C1(n10570), .C2(n10569), .A(n9757), .B(n9756), .ZN(
        n10571) );
  NAND2_X1 U12962 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n9756) );
  NAND2_X1 U12963 ( .A1(n9761), .A2(n10166), .ZN(n16123) );
  NAND2_X1 U12964 ( .A1(n9761), .A2(n13664), .ZN(n16187) );
  AND2_X4 U12966 ( .A1(n9761), .A2(n10167), .ZN(n16141) );
  AND2_X2 U12967 ( .A1(n9761), .A2(n13583), .ZN(n9799) );
  AND2_X1 U12968 ( .A1(n9761), .A2(n9826), .ZN(n16161) );
  NAND2_X1 U12969 ( .A1(n9933), .A2(n9761), .ZN(n9932) );
  NAND2_X2 U12970 ( .A1(n9934), .A2(n9761), .ZN(n16268) );
  NAND2_X4 U12971 ( .A1(n9850), .A2(n9630), .ZN(n9761) );
  NAND2_X2 U12972 ( .A1(n11688), .A2(n15607), .ZN(n14621) );
  NAND2_X1 U12973 ( .A1(n9766), .A2(n11656), .ZN(n9763) );
  NAND2_X1 U12974 ( .A1(n9765), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9764) );
  NAND4_X1 U12975 ( .A1(n11670), .A2(n11672), .A3(n11671), .A4(n11673), .ZN(
        n9765) );
  NAND4_X1 U12976 ( .A1(n11674), .A2(n11675), .A3(n11676), .A4(n11677), .ZN(
        n9766) );
  NAND2_X2 U12977 ( .A1(n9767), .A2(n11684), .ZN(n11688) );
  OAI21_X2 U12978 ( .B1(n9598), .B2(n9768), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U12979 ( .A1(n9583), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n9770) );
  NAND3_X1 U12980 ( .A1(n16248), .A2(n16178), .A3(n10133), .ZN(n9771) );
  NAND3_X1 U12981 ( .A1(n9773), .A2(n12766), .A3(n9774), .ZN(n16126) );
  NAND3_X1 U12982 ( .A1(n9608), .A2(n9588), .A3(n9636), .ZN(n9773) );
  AOI21_X1 U12983 ( .B1(n9777), .B2(n19952), .A(n16378), .ZN(n9776) );
  AND2_X1 U12984 ( .A1(n12445), .A2(n19992), .ZN(n9780) );
  NAND3_X1 U12985 ( .A1(n11710), .A2(n9999), .A3(n12140), .ZN(n16816) );
  INV_X1 U12986 ( .A(n16278), .ZN(n16277) );
  NAND2_X1 U12987 ( .A1(n12616), .A2(n12617), .ZN(n9781) );
  NAND2_X1 U12988 ( .A1(n12613), .A2(n9682), .ZN(n9782) );
  NAND2_X1 U12989 ( .A1(n16591), .A2(n16590), .ZN(n9783) );
  NOR2_X1 U12990 ( .A1(n9786), .A2(n16676), .ZN(n13806) );
  NAND2_X1 U12991 ( .A1(n9786), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16836) );
  AOI21_X1 U12992 ( .B1(n9786), .B2(n16798), .A(n9680), .ZN(n13808) );
  NAND3_X1 U12993 ( .A1(n10299), .A2(n10296), .A3(n10297), .ZN(n9787) );
  NOR2_X4 U12994 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16657) );
  NAND3_X1 U12995 ( .A1(n9790), .A2(n9789), .A3(n9788), .ZN(P2_U3026) );
  INV_X1 U12996 ( .A(n16111), .ZN(n10363) );
  NAND2_X1 U12997 ( .A1(n16111), .A2(n13635), .ZN(n10359) );
  NAND2_X1 U12998 ( .A1(n16108), .A2(n9793), .ZN(P2_U2985) );
  NAND3_X1 U12999 ( .A1(n16371), .A2(n16372), .A3(n9795), .ZN(P2_U3017) );
  XNOR2_X2 U13000 ( .A(n12617), .B(n9797), .ZN(n12641) );
  INV_X1 U13001 ( .A(n12614), .ZN(n9797) );
  NAND2_X1 U13002 ( .A1(n13095), .A2(n15607), .ZN(n9803) );
  NAND2_X1 U13003 ( .A1(n9803), .A2(n11708), .ZN(n12148) );
  NAND2_X1 U13004 ( .A1(n11724), .A2(n19985), .ZN(n10000) );
  NAND2_X1 U13005 ( .A1(n10063), .A2(n9805), .ZN(P2_U2995) );
  INV_X1 U13006 ( .A(n9806), .ZN(n9805) );
  OAI21_X1 U13007 ( .B1(n16467), .B2(n19941), .A(n9694), .ZN(n9806) );
  NAND2_X1 U13008 ( .A1(n9808), .A2(n20581), .ZN(n12177) );
  NOR2_X1 U13009 ( .A1(n9808), .A2(n11699), .ZN(n11692) );
  AND2_X2 U13010 ( .A1(n13135), .A2(n9808), .ZN(n12140) );
  NAND2_X1 U13011 ( .A1(n12135), .A2(n9808), .ZN(n12136) );
  AOI21_X1 U13012 ( .B1(n16740), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U13013 ( .A1(n16002), .A2(n9808), .ZN(n15975) );
  NAND2_X2 U13014 ( .A1(n16175), .A2(n16137), .ZN(n16159) );
  NAND2_X1 U13015 ( .A1(n9814), .A2(n12137), .ZN(n10204) );
  NAND2_X1 U13016 ( .A1(n12137), .A2(n9720), .ZN(n13133) );
  NAND2_X1 U13017 ( .A1(n16141), .A2(n9743), .ZN(n9815) );
  NAND2_X1 U13018 ( .A1(n16141), .A2(n9745), .ZN(n9847) );
  NAND2_X1 U13019 ( .A1(n16201), .A2(n9817), .ZN(P2_U2994) );
  XNOR2_X2 U13020 ( .A(n10689), .B(n10707), .ZN(n20931) );
  NAND3_X1 U13021 ( .A1(n20775), .A2(n9820), .A3(n10200), .ZN(n10199) );
  XNOR2_X1 U13022 ( .A(n10833), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14483) );
  NAND2_X1 U13023 ( .A1(n13040), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10605) );
  NAND3_X1 U13024 ( .A1(n9821), .A2(n10597), .A3(n10596), .ZN(n13040) );
  NOR2_X1 U13025 ( .A1(n13026), .A2(n10615), .ZN(n9821) );
  OAI211_X1 U13026 ( .C1(n14137), .C2(n13599), .A(n10592), .B(n13913), .ZN(
        n10615) );
  NAND3_X2 U13027 ( .A1(n10083), .A2(n11594), .A3(n11593), .ZN(n15340) );
  XNOR2_X1 U13028 ( .A(n9824), .B(n9641), .ZN(n15570) );
  INV_X1 U13029 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9825) );
  INV_X2 U13030 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10933) );
  NOR2_X1 U13031 ( .A1(n16161), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16409) );
  NAND2_X1 U13032 ( .A1(n16933), .A2(n16936), .ZN(n16932) );
  NAND3_X1 U13033 ( .A1(n9833), .A2(n9591), .A3(n9830), .ZN(n9828) );
  NAND2_X1 U13034 ( .A1(n13249), .A2(n9831), .ZN(n13230) );
  NAND4_X1 U13035 ( .A1(n9591), .A2(n9833), .A3(n9637), .A4(n9832), .ZN(n9831)
         );
  INV_X1 U13036 ( .A(n13187), .ZN(n9833) );
  NAND2_X1 U13037 ( .A1(n14112), .A2(n14111), .ZN(n13233) );
  XNOR2_X1 U13038 ( .A(n13230), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14112) );
  NAND2_X1 U13039 ( .A1(n10051), .A2(n13308), .ZN(n18567) );
  OAI211_X1 U13040 ( .C1(n10051), .C2(n9838), .A(n9835), .B(n9834), .ZN(n14188) );
  NAND2_X1 U13041 ( .A1(n13332), .A2(n9837), .ZN(n9834) );
  NAND2_X1 U13042 ( .A1(n10051), .A2(n9836), .ZN(n9835) );
  NOR2_X1 U13043 ( .A1(n13332), .A2(n9837), .ZN(n9836) );
  INV_X1 U13044 ( .A(n13308), .ZN(n9837) );
  NAND2_X1 U13045 ( .A1(n18710), .A2(n18709), .ZN(n9839) );
  OAI21_X2 U13046 ( .B1(n18568), .B2(n10156), .A(n9597), .ZN(n13347) );
  NAND2_X1 U13047 ( .A1(n16907), .A2(n9843), .ZN(n9842) );
  NAND3_X1 U13048 ( .A1(n16891), .A2(n18548), .A3(n9846), .ZN(n13351) );
  NAND3_X1 U13049 ( .A1(n9589), .A2(n16876), .A3(n16851), .ZN(n16852) );
  INV_X1 U13050 ( .A(n13354), .ZN(n18447) );
  NOR2_X1 U13051 ( .A1(n16332), .A2(n9848), .ZN(n16317) );
  AND2_X1 U13052 ( .A1(n9849), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9848) );
  NAND2_X1 U13053 ( .A1(n9850), .A2(n16313), .ZN(n9849) );
  OAI21_X1 U13054 ( .B1(n16340), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n9850), .ZN(n16626) );
  NAND2_X2 U13055 ( .A1(n16340), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9850) );
  NAND4_X2 U13056 ( .A1(n10617), .A2(n9929), .A3(n9852), .A4(n9851), .ZN(
        n10618) );
  NAND2_X1 U13057 ( .A1(n10590), .A2(n13028), .ZN(n9851) );
  NAND2_X1 U13058 ( .A1(n10203), .A2(n10602), .ZN(n9852) );
  OR2_X2 U13059 ( .A1(n10554), .A2(n10553), .ZN(n10599) );
  NAND2_X1 U13060 ( .A1(n15225), .A2(n9854), .ZN(P1_U2974) );
  NAND2_X1 U13061 ( .A1(n15405), .A2(n9856), .ZN(P1_U3006) );
  AND2_X2 U13062 ( .A1(n14583), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10468) );
  OAI21_X2 U13064 ( .B1(n11591), .B2(n10891), .A(n9857), .ZN(n10142) );
  NAND3_X1 U13065 ( .A1(n10058), .A2(n9881), .A3(n9878), .ZN(P3_U2802) );
  INV_X1 U13066 ( .A(n13287), .ZN(n10053) );
  NAND3_X1 U13067 ( .A1(n16343), .A2(n16276), .A3(n16279), .ZN(n9887) );
  INV_X1 U13068 ( .A(n16331), .ZN(n16320) );
  NAND2_X1 U13069 ( .A1(n16278), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9894) );
  XNOR2_X2 U13070 ( .A(n13338), .B(n13334), .ZN(n16907) );
  NAND2_X1 U13071 ( .A1(n10112), .A2(n9899), .ZN(n9898) );
  INV_X1 U13072 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n9906) );
  INV_X1 U13073 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n9909) );
  INV_X1 U13074 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n9912) );
  INV_X1 U13075 ( .A(n16187), .ZN(n9922) );
  NAND3_X1 U13076 ( .A1(n10474), .A2(n9923), .A3(
        P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10529) );
  NAND3_X1 U13077 ( .A1(n10474), .A2(n9923), .A3(
        P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10512) );
  AND2_X2 U13078 ( .A1(n10469), .A2(n9923), .ZN(n10633) );
  NAND2_X1 U13079 ( .A1(n10695), .A2(n9924), .ZN(n10977) );
  NAND2_X1 U13080 ( .A1(n11599), .A2(n11602), .ZN(n11600) );
  NAND3_X1 U13081 ( .A1(n10594), .A2(n10790), .A3(n10587), .ZN(n9929) );
  NAND2_X1 U13082 ( .A1(n14450), .A2(n14449), .ZN(n14448) );
  INV_X1 U13083 ( .A(n16632), .ZN(n12549) );
  NAND2_X2 U13084 ( .A1(n16633), .A2(n16634), .ZN(n16632) );
  NAND2_X1 U13085 ( .A1(n9931), .A2(n9930), .ZN(n16633) );
  NAND2_X1 U13086 ( .A1(n10006), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9930) );
  AND2_X4 U13087 ( .A1(n10147), .A2(n12532), .ZN(n12527) );
  NAND2_X1 U13088 ( .A1(n10067), .A2(n12538), .ZN(n19918) );
  NAND2_X1 U13089 ( .A1(n10066), .A2(n10065), .ZN(n10069) );
  BUF_X4 U13090 ( .A(n12426), .Z(n19945) );
  OAI22_X1 U13091 ( .A1(n10123), .A2(n10124), .B1(n20446), .B2(n16778), .ZN(
        n12442) );
  NOR3_X1 U13092 ( .A1(n16858), .A2(n18659), .A3(n16940), .ZN(n16859) );
  NOR2_X1 U13093 ( .A1(n16298), .A2(n15783), .ZN(n19712) );
  OR2_X1 U13094 ( .A1(n19719), .A2(n19717), .ZN(n15796) );
  INV_X1 U13095 ( .A(n15796), .ZN(n15795) );
  INV_X1 U13096 ( .A(n15814), .ZN(n15813) );
  NOR2_X1 U13097 ( .A1(n19916), .A2(n19789), .ZN(n19763) );
  OAI21_X2 U13098 ( .B1(n15617), .B2(n15622), .A(n19790), .ZN(n14702) );
  NOR2_X1 U13099 ( .A1(n14642), .A2(n19687), .ZN(n15768) );
  NOR2_X2 U13100 ( .A1(n14649), .A2(n19645), .ZN(n15755) );
  OR2_X2 U13101 ( .A1(n20240), .A2(n12444), .ZN(n12446) );
  NOR2_X1 U13102 ( .A1(n12448), .A2(n10149), .ZN(n10148) );
  NAND3_X2 U13103 ( .A1(n12528), .A2(n12527), .A3(n12585), .ZN(n12617) );
  NAND2_X1 U13104 ( .A1(n10046), .A2(n10045), .ZN(n13084) );
  NAND3_X2 U13105 ( .A1(n9998), .A2(n9999), .A3(n12140), .ZN(n13095) );
  NOR2_X1 U13106 ( .A1(n13135), .A2(n15607), .ZN(n9935) );
  INV_X1 U13107 ( .A(n13101), .ZN(n9936) );
  NOR2_X1 U13108 ( .A1(n15822), .A2(n12408), .ZN(n9939) );
  NAND3_X1 U13109 ( .A1(n14236), .A2(n10198), .A3(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9940) );
  INV_X1 U13110 ( .A(n12417), .ZN(n9942) );
  NAND2_X1 U13111 ( .A1(n9944), .A2(n16187), .ZN(n13693) );
  INV_X2 U13112 ( .A(n19997), .ZN(n13135) );
  NAND4_X1 U13113 ( .A1(n11614), .A2(n11613), .A3(n11611), .A4(n11612), .ZN(
        n9945) );
  NOR2_X1 U13114 ( .A1(n9949), .A2(n9948), .ZN(n9947) );
  NAND2_X1 U13115 ( .A1(n10300), .A2(n9603), .ZN(n9951) );
  NOR2_X1 U13116 ( .A1(n13408), .A2(n9952), .ZN(n9954) );
  NAND3_X1 U13117 ( .A1(n9670), .A2(n13402), .A3(n13403), .ZN(n9952) );
  NAND2_X1 U13118 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n9955) );
  NOR2_X2 U13119 ( .A1(n17927), .A2(n9959), .ZN(n17885) );
  NAND4_X1 U13120 ( .A1(n9976), .A2(n13409), .A3(n9974), .A4(n9973), .ZN(n9972) );
  AND2_X2 U13121 ( .A1(n9983), .A2(n9982), .ZN(n14388) );
  NAND3_X1 U13122 ( .A1(n14045), .A2(n10587), .A3(n13599), .ZN(n14038) );
  INV_X1 U13123 ( .A(n10794), .ZN(n10143) );
  NAND3_X1 U13124 ( .A1(n10729), .A2(n10728), .A3(n14428), .ZN(n10794) );
  NAND2_X2 U13125 ( .A1(n10729), .A2(n10728), .ZN(n10801) );
  AND4_X2 U13126 ( .A1(n15285), .A2(n10894), .A3(n11594), .A4(n10892), .ZN(
        n10895) );
  OR2_X2 U13127 ( .A1(n10977), .A2(n10978), .ZN(n10976) );
  NAND3_X1 U13128 ( .A1(n10709), .A2(n20862), .A3(n10276), .ZN(n9986) );
  NAND2_X1 U13129 ( .A1(n10730), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9987) );
  NOR2_X2 U13130 ( .A1(n9990), .A2(n10439), .ZN(n11714) );
  NAND2_X1 U13131 ( .A1(n9990), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10021) );
  NAND2_X1 U13132 ( .A1(n9990), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11731) );
  AOI21_X1 U13133 ( .B1(n9990), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11737), .ZN(n11743) );
  NAND2_X2 U13134 ( .A1(n10060), .A2(n11711), .ZN(n9990) );
  AND2_X4 U13135 ( .A1(n16660), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11972) );
  AND2_X4 U13136 ( .A1(n16660), .A2(n16797), .ZN(n11790) );
  AND2_X2 U13137 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16660) );
  OR2_X2 U13138 ( .A1(n11686), .A2(n11685), .ZN(n11698) );
  NOR2_X2 U13139 ( .A1(n11699), .A2(n13123), .ZN(n9999) );
  NAND2_X2 U13140 ( .A1(n13112), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11738) );
  NAND2_X2 U13141 ( .A1(n10000), .A2(n16673), .ZN(n13112) );
  NAND2_X1 U13142 ( .A1(n10001), .A2(n9685), .ZN(n10045) );
  XNOR2_X2 U13143 ( .A(n10127), .B(n12585), .ZN(n10006) );
  XNOR2_X1 U13144 ( .A(n19919), .B(n10006), .ZN(n19966) );
  NAND2_X1 U13145 ( .A1(n16241), .A2(n10013), .ZN(n10012) );
  NOR2_X1 U13146 ( .A1(n14586), .A2(n15975), .ZN(n10023) );
  INV_X1 U13147 ( .A(n14373), .ZN(n10026) );
  NAND2_X1 U13148 ( .A1(n10030), .A2(n10027), .ZN(n14528) );
  NAND3_X1 U13149 ( .A1(n10029), .A2(n10028), .A3(n10032), .ZN(n10027) );
  INV_X1 U13150 ( .A(n12054), .ZN(n10028) );
  INV_X1 U13151 ( .A(n12055), .ZN(n10029) );
  OAI21_X1 U13152 ( .B1(n12055), .B2(n12054), .A(n12069), .ZN(n10030) );
  OAI21_X1 U13153 ( .B1(n12055), .B2(n12054), .A(n10032), .ZN(n10031) );
  NAND3_X1 U13154 ( .A1(n10275), .A2(n10033), .A3(n10279), .ZN(n10072) );
  NAND2_X1 U13155 ( .A1(n9642), .A2(n10033), .ZN(n13984) );
  NAND2_X1 U13156 ( .A1(n10709), .A2(n9679), .ZN(n10033) );
  XNOR2_X1 U13157 ( .A(n10868), .B(n10867), .ZN(n11028) );
  NAND2_X1 U13158 ( .A1(n15281), .A2(n15280), .ZN(n15251) );
  INV_X1 U13159 ( .A(n10038), .ZN(n15210) );
  INV_X1 U13160 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10042) );
  AND2_X2 U13161 ( .A1(n12619), .A2(n10043), .ZN(n12698) );
  AND2_X2 U13162 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12556) );
  AND2_X4 U13163 ( .A1(n12556), .A2(n12102), .ZN(n14597) );
  NOR2_X2 U13164 ( .A1(n14167), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10050) );
  NAND2_X1 U13165 ( .A1(n11718), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10060) );
  NAND2_X1 U13166 ( .A1(n10062), .A2(n10061), .ZN(n11718) );
  NAND2_X1 U13167 ( .A1(n11701), .A2(n13124), .ZN(n10062) );
  NAND2_X2 U13168 ( .A1(n12527), .A2(n12528), .ZN(n10127) );
  XNOR2_X1 U13169 ( .A(n12527), .B(n12528), .ZN(n16348) );
  NAND2_X2 U13170 ( .A1(n10070), .A2(n12439), .ZN(n12528) );
  NAND3_X1 U13171 ( .A1(n10127), .A2(n10069), .A3(n10068), .ZN(n10067) );
  NAND2_X1 U13172 ( .A1(n12438), .A2(n12445), .ZN(n10070) );
  NAND2_X1 U13173 ( .A1(n10072), .A2(n9677), .ZN(n10071) );
  NOR2_X1 U13174 ( .A1(n10075), .A2(n10595), .ZN(n10073) );
  NAND2_X1 U13175 ( .A1(n10075), .A2(n12951), .ZN(n10074) );
  NAND2_X1 U13176 ( .A1(n10076), .A2(n10079), .ZN(n11596) );
  NAND2_X1 U13177 ( .A1(n15340), .A2(n10082), .ZN(n15341) );
  INV_X1 U13178 ( .A(n10788), .ZN(n10786) );
  NAND2_X1 U13179 ( .A1(n11710), .A2(n9640), .ZN(n12138) );
  AND2_X2 U13180 ( .A1(n10136), .A2(n15593), .ZN(n10635) );
  AND2_X2 U13181 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15593) );
  XNOR2_X2 U13182 ( .A(n10692), .B(n10690), .ZN(n10986) );
  NAND3_X1 U13183 ( .A1(n11035), .A2(n10868), .A3(n14078), .ZN(n10093) );
  NAND3_X1 U13184 ( .A1(n10128), .A2(n11763), .A3(n11764), .ZN(n10104) );
  AND2_X4 U13185 ( .A1(n10097), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11970) );
  NAND2_X1 U13186 ( .A1(n10098), .A2(n16335), .ZN(n16261) );
  NAND2_X1 U13187 ( .A1(n10098), .A2(n16603), .ZN(n16536) );
  AND2_X2 U13188 ( .A1(n10100), .A2(n10099), .ZN(n10098) );
  INV_X1 U13189 ( .A(n16253), .ZN(n10099) );
  NAND2_X1 U13190 ( .A1(n16539), .A2(n16254), .ZN(n10100) );
  AND2_X2 U13191 ( .A1(n12410), .A2(n12418), .ZN(n12402) );
  NOR2_X4 U13192 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14409) );
  NAND2_X1 U13193 ( .A1(n10104), .A2(n11771), .ZN(n10106) );
  NAND2_X1 U13194 ( .A1(n10106), .A2(n10105), .ZN(n11751) );
  NAND2_X1 U13195 ( .A1(n11762), .A2(n10107), .ZN(n10105) );
  NAND4_X1 U13196 ( .A1(n10109), .A2(n11629), .A3(n11628), .A4(n11630), .ZN(
        n10108) );
  AND2_X1 U13197 ( .A1(n11627), .A2(n11656), .ZN(n10109) );
  NAND4_X1 U13198 ( .A1(n10111), .A2(n11634), .A3(n11632), .A4(n11633), .ZN(
        n10110) );
  AND2_X1 U13199 ( .A1(n11631), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10111) );
  NOR2_X1 U13200 ( .A1(n10114), .A2(n10113), .ZN(n10112) );
  NAND3_X1 U13201 ( .A1(n12519), .A2(n12520), .A3(n12509), .ZN(n10114) );
  NAND3_X1 U13202 ( .A1(n12404), .A2(n19945), .A3(n15847), .ZN(n16751) );
  NAND2_X1 U13203 ( .A1(n12549), .A2(n12548), .ZN(n10122) );
  INV_X1 U13204 ( .A(n12429), .ZN(n10123) );
  NAND2_X1 U13205 ( .A1(n12429), .A2(n12404), .ZN(n10126) );
  OAI22_X1 U13206 ( .A1(n10126), .A2(n12430), .B1(n20216), .B2(n12431), .ZN(
        n12432) );
  OAI22_X1 U13207 ( .A1(n10126), .A2(n12503), .B1(n20216), .B2(n12504), .ZN(
        n12505) );
  OAI22_X1 U13208 ( .A1(n10126), .A2(n12480), .B1(n20216), .B2(n12479), .ZN(
        n12481) );
  OAI21_X1 U13209 ( .B1(n10126), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10125), 
        .ZN(n20278) );
  AOI21_X1 U13210 ( .B1(n10126), .B2(n20277), .A(n20392), .ZN(n20275) );
  NAND3_X1 U13211 ( .A1(n9576), .A2(n13127), .A3(n12154), .ZN(n13139) );
  OR2_X2 U13212 ( .A1(n12743), .A2(n13655), .ZN(n10135) );
  NOR2_X1 U13213 ( .A1(n20388), .A2(n12488), .ZN(n12492) );
  MUX2_X1 U13214 ( .A(n10136), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15593), .Z(n13924) );
  INV_X1 U13215 ( .A(n10885), .ZN(n15342) );
  NAND2_X2 U13216 ( .A1(n10142), .A2(n10895), .ZN(n15281) );
  NAND4_X1 U13217 ( .A1(n10148), .A2(n12465), .A3(n12466), .A4(n12467), .ZN(
        n10147) );
  OAI21_X1 U13218 ( .B1(n16959), .B2(n18653), .A(n10152), .ZN(P3_U2799) );
  AND2_X1 U13219 ( .A1(n16875), .A2(n16874), .ZN(n10152) );
  AND2_X2 U13220 ( .A1(n14393), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13180) );
  NAND2_X1 U13221 ( .A1(n13356), .A2(n10161), .ZN(n16850) );
  NAND2_X1 U13222 ( .A1(n16850), .A2(n18565), .ZN(n16853) );
  NAND2_X1 U13223 ( .A1(n11751), .A2(n10162), .ZN(n11736) );
  XNOR2_X1 U13224 ( .A(n11751), .B(n10162), .ZN(n12396) );
  INV_X1 U13225 ( .A(n11738), .ZN(n12783) );
  NAND2_X1 U13226 ( .A1(n12783), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10398) );
  AND3_X4 U13227 ( .A1(n16656), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11784) );
  INV_X1 U13228 ( .A(n12410), .ZN(n10163) );
  INV_X1 U13229 ( .A(n11688), .ZN(n12179) );
  NOR2_X1 U13230 ( .A1(n11688), .A2(n16815), .ZN(n14617) );
  NAND2_X1 U13231 ( .A1(n11699), .A2(n19985), .ZN(n12145) );
  NAND2_X1 U13232 ( .A1(n12159), .A2(n12179), .ZN(n12341) );
  NAND2_X1 U13233 ( .A1(n12588), .A2(n19985), .ZN(n12522) );
  NOR2_X1 U13234 ( .A1(n12012), .A2(n19985), .ZN(n11990) );
  NAND2_X1 U13235 ( .A1(n12029), .A2(n19985), .ZN(n15879) );
  AND2_X1 U13236 ( .A1(n12070), .A2(n19985), .ZN(n14527) );
  NAND2_X1 U13237 ( .A1(n12008), .A2(n19985), .ZN(n15890) );
  NAND2_X1 U13238 ( .A1(n12011), .A2(n19985), .ZN(n15886) );
  NAND2_X1 U13239 ( .A1(n16829), .A2(n19985), .ZN(n16832) );
  NAND2_X2 U13240 ( .A1(n14684), .A2(n10165), .ZN(n13961) );
  NAND2_X1 U13241 ( .A1(n11688), .A2(n10291), .ZN(n10165) );
  AND2_X1 U13242 ( .A1(n13580), .A2(n9741), .ZN(n10166) );
  AND2_X1 U13243 ( .A1(n13580), .A2(n10168), .ZN(n10167) );
  OAI21_X1 U13244 ( .B1(n16408), .B2(n17292), .A(n10169), .ZN(P2_U2988) );
  NAND2_X1 U13245 ( .A1(n14526), .A2(n10031), .ZN(n10194) );
  NAND2_X1 U13246 ( .A1(n10189), .A2(n10187), .ZN(n10195) );
  NAND2_X1 U13247 ( .A1(n10188), .A2(n10191), .ZN(n10187) );
  NAND2_X1 U13248 ( .A1(n14526), .A2(n10190), .ZN(n10189) );
  AOI22_X1 U13249 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9568), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10494) );
  AND3_X2 U13250 ( .A1(n10600), .A2(n14030), .A3(n10969), .ZN(n13936) );
  NAND4_X1 U13251 ( .A1(n10600), .A2(n14030), .A3(n14511), .A4(n10969), .ZN(
        n13022) );
  NAND2_X1 U13252 ( .A1(n13936), .A2(n12941), .ZN(n12925) );
  NAND2_X1 U13253 ( .A1(n10204), .A2(n13125), .ZN(n11700) );
  NAND2_X1 U13254 ( .A1(n17240), .A2(n10862), .ZN(n10206) );
  NOR2_X2 U13255 ( .A1(n10902), .A2(n15333), .ZN(n15244) );
  OR2_X1 U13256 ( .A1(n10903), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10210) );
  NAND2_X1 U13257 ( .A1(n15416), .A2(n9742), .ZN(n10211) );
  XNOR2_X1 U13258 ( .A(n10794), .B(n10795), .ZN(n11015) );
  NOR2_X1 U13259 ( .A1(n10214), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17767) );
  NOR2_X1 U13260 ( .A1(n16927), .A2(n10214), .ZN(n17774) );
  AOI21_X1 U13261 ( .B1(n18606), .B2(n10214), .A(n18722), .ZN(n18712) );
  INV_X1 U13262 ( .A(n10215), .ZN(n17485) );
  NOR2_X1 U13263 ( .A1(n17494), .A2(n17775), .ZN(n17486) );
  OAI21_X1 U13264 ( .B1(n17528), .B2(n9719), .A(n10223), .ZN(n17504) );
  INV_X1 U13265 ( .A(n10226), .ZN(n17505) );
  NAND2_X1 U13266 ( .A1(n15743), .A2(n10239), .ZN(n14662) );
  NAND2_X2 U13267 ( .A1(n19790), .A2(n14658), .ZN(n15743) );
  INV_X1 U13268 ( .A(n14636), .ZN(n10241) );
  NAND2_X1 U13269 ( .A1(n10241), .A2(n10242), .ZN(n14628) );
  AOI21_X1 U13270 ( .B1(n10255), .B2(n16264), .A(n10254), .ZN(n10253) );
  NAND2_X1 U13271 ( .A1(n16876), .A2(n13353), .ZN(n13356) );
  NAND3_X1 U13272 ( .A1(n18454), .A2(n18453), .A3(n9683), .ZN(n10270) );
  NAND3_X1 U13273 ( .A1(n11589), .A2(n11590), .A3(n11588), .ZN(P1_U2968) );
  NAND2_X1 U13274 ( .A1(n10280), .A2(n10994), .ZN(n14251) );
  INV_X1 U13275 ( .A(n14498), .ZN(n10282) );
  INV_X1 U13276 ( .A(n14497), .ZN(n10281) );
  NAND4_X1 U13277 ( .A1(n10282), .A2(n14957), .A3(n11100), .A4(n10281), .ZN(
        n14922) );
  NAND2_X1 U13278 ( .A1(n10283), .A2(n15100), .ZN(n15092) );
  NAND2_X1 U13279 ( .A1(n9716), .A2(n10284), .ZN(n17245) );
  XNOR2_X1 U13280 ( .A(n10284), .B(n15100), .ZN(n17241) );
  NAND2_X1 U13281 ( .A1(n11262), .A2(n10285), .ZN(n14770) );
  AND2_X2 U13282 ( .A1(n11262), .A2(n9704), .ZN(n14783) );
  NAND2_X1 U13283 ( .A1(n11489), .A2(n10289), .ZN(n13727) );
  NOR2_X1 U13284 ( .A1(n13799), .A2(n10291), .ZN(n13791) );
  NAND2_X1 U13285 ( .A1(n13126), .A2(n10293), .ZN(n13128) );
  NAND2_X1 U13286 ( .A1(n16492), .A2(n10294), .ZN(P2_U3028) );
  NAND2_X1 U13287 ( .A1(n10295), .A2(n19962), .ZN(n10294) );
  INV_X1 U13288 ( .A(n16493), .ZN(n10295) );
  NAND2_X1 U13289 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10296) );
  NAND2_X1 U13290 ( .A1(n11977), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U13291 ( .A1(n12718), .A2(n9724), .ZN(n12747) );
  NOR2_X2 U13292 ( .A1(n12683), .A2(n10437), .ZN(n12707) );
  NAND3_X1 U13293 ( .A1(n14731), .A2(n12941), .A3(n12933), .ZN(n12936) );
  NAND3_X1 U13294 ( .A1(n10317), .A2(n14852), .A3(n14844), .ZN(n10316) );
  NOR2_X2 U13295 ( .A1(n12609), .A2(n10319), .ZN(n12625) );
  OR2_X2 U13296 ( .A1(n12609), .A2(n10318), .ZN(n12700) );
  INV_X1 U13297 ( .A(n12610), .ZN(n10320) );
  AND3_X2 U13298 ( .A1(n13925), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U13299 ( .A1(n14063), .A2(n12418), .ZN(n10349) );
  OR2_X1 U13300 ( .A1(n15822), .A2(n10350), .ZN(n10352) );
  NAND3_X1 U13301 ( .A1(n14063), .A2(n12418), .A3(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10350) );
  NAND2_X1 U13302 ( .A1(n13164), .A2(n19936), .ZN(n10358) );
  NAND3_X1 U13303 ( .A1(n10358), .A2(n10426), .A3(n10357), .ZN(P2_U2984) );
  NAND3_X1 U13304 ( .A1(n10362), .A2(n10360), .A3(n10359), .ZN(n10357) );
  NAND3_X1 U13305 ( .A1(n10362), .A2(n10364), .A3(n10359), .ZN(n13167) );
  NAND2_X1 U13306 ( .A1(n16083), .A2(n10366), .ZN(n10365) );
  NAND2_X1 U13307 ( .A1(n10365), .A2(n10369), .ZN(n13883) );
  NAND2_X1 U13308 ( .A1(n14563), .A2(n9723), .ZN(n15737) );
  NAND2_X1 U13309 ( .A1(n10380), .A2(n10378), .ZN(n15658) );
  INV_X1 U13310 ( .A(n14118), .ZN(n10383) );
  NAND2_X1 U13311 ( .A1(n10383), .A2(n10384), .ZN(n14323) );
  NOR2_X1 U13312 ( .A1(n14118), .A2(n14185), .ZN(n14184) );
  INV_X1 U13313 ( .A(n14185), .ZN(n10386) );
  INV_X1 U13314 ( .A(n10391), .ZN(n13642) );
  AND2_X2 U13315 ( .A1(n14531), .A2(n15623), .ZN(n15625) );
  OAI21_X1 U13316 ( .B1(n15388), .B2(n20807), .A(n15387), .ZN(P1_U3004) );
  XNOR2_X1 U13317 ( .A(n10396), .B(n15383), .ZN(n15388) );
  NAND2_X1 U13318 ( .A1(n15204), .A2(n15333), .ZN(n10397) );
  NAND2_X1 U13319 ( .A1(n10905), .A2(n13622), .ZN(n15204) );
  NAND2_X1 U13320 ( .A1(n10786), .A2(n10785), .ZN(n10840) );
  INV_X1 U13321 ( .A(n11762), .ZN(n11770) );
  INV_X1 U13322 ( .A(n14375), .ZN(n10401) );
  NAND3_X1 U13323 ( .A1(n10401), .A2(n15792), .A3(n10400), .ZN(n15948) );
  NAND4_X1 U13324 ( .A1(n10401), .A2(n15792), .A3(n10407), .A4(n12804), .ZN(
        n15777) );
  NAND3_X1 U13325 ( .A1(n10407), .A2(n12804), .A3(n10406), .ZN(n10405) );
  INV_X1 U13326 ( .A(n14376), .ZN(n10407) );
  NAND2_X1 U13327 ( .A1(n15649), .A2(n10420), .ZN(n15633) );
  AND2_X1 U13328 ( .A1(n15649), .A2(n15648), .ZN(n14539) );
  NAND2_X1 U13329 ( .A1(n16113), .A2(n12759), .ZN(n16139) );
  INV_X1 U13330 ( .A(n12620), .ZN(n12621) );
  INV_X1 U13331 ( .A(n13685), .ZN(n13686) );
  AOI21_X1 U13333 ( .B1(n13747), .B2(n20801), .A(n13746), .ZN(n13748) );
  NOR2_X1 U13334 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  XNOR2_X1 U13335 ( .A(n13625), .B(n13624), .ZN(n15202) );
  XNOR2_X1 U13336 ( .A(n10801), .B(n14428), .ZN(n10995) );
  XNOR2_X1 U13337 ( .A(n12900), .B(n10430), .ZN(n13758) );
  CLKBUF_X1 U13338 ( .A(n14323), .Z(n16496) );
  INV_X1 U13339 ( .A(n13078), .ZN(n13093) );
  NOR2_X1 U13340 ( .A1(n16751), .A2(n12405), .ZN(n12406) );
  NAND2_X1 U13341 ( .A1(n14369), .A2(n14371), .ZN(n15990) );
  AOI21_X1 U13342 ( .B1(n12898), .B2(n15353), .A(n13739), .ZN(n12900) );
  CLKBUF_X1 U13343 ( .A(n13139), .Z(n16672) );
  CLKBUF_X1 U13344 ( .A(n11599), .Z(n14911) );
  XNOR2_X1 U13345 ( .A(n11992), .B(n12013), .ZN(n15891) );
  OAI211_X1 U13346 ( .C1(n16191), .C2(n13662), .A(n13661), .B(n13660), .ZN(
        n13687) );
  NAND2_X1 U13347 ( .A1(n16191), .A2(n13653), .ZN(n13661) );
  XNOR2_X1 U13348 ( .A(n13681), .B(n13067), .ZN(n13111) );
  OR2_X1 U13349 ( .A1(n16206), .A2(n14550), .ZN(n14558) );
  OR2_X1 U13350 ( .A1(n10975), .A2(n14428), .ZN(n21064) );
  OR2_X1 U13351 ( .A1(n10975), .A2(n14427), .ZN(n21345) );
  OAI21_X1 U13352 ( .B1(n15202), .B2(n20807), .A(n13632), .ZN(P1_U3003) );
  NAND2_X1 U13353 ( .A1(n13645), .A2(n19936), .ZN(n13092) );
  INV_X1 U13354 ( .A(n13111), .ZN(n14612) );
  AOI22_X1 U13355 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13356 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10524) );
  OR2_X1 U13357 ( .A1(n11738), .A2(n13142), .ZN(n11729) );
  NAND2_X1 U13358 ( .A1(n14729), .A2(n13604), .ZN(n13620) );
  NAND2_X1 U13359 ( .A1(n14729), .A2(n20779), .ZN(n11589) );
  INV_X1 U13360 ( .A(n13587), .ZN(n12854) );
  NOR2_X1 U13361 ( .A1(n20004), .A2(n19997), .ZN(n20454) );
  NAND2_X1 U13362 ( .A1(n11790), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11662) );
  AOI22_X1 U13363 ( .A1(n9571), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U13364 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11627) );
  INV_X1 U13365 ( .A(n18163), .ZN(n18177) );
  AND2_X1 U13366 ( .A1(n13603), .A2(n13602), .ZN(n15123) );
  INV_X2 U13367 ( .A(n15123), .ZN(n17230) );
  INV_X1 U13368 ( .A(n12628), .ZN(n12591) );
  AND2_X1 U13369 ( .A1(n14686), .A2(n14685), .ZN(n19651) );
  OR2_X2 U13370 ( .A1(n14139), .A2(n14138), .ZN(n20765) );
  AND2_X2 U13371 ( .A1(n20631), .A2(n11581), .ZN(n20773) );
  AND2_X1 U13372 ( .A1(n10701), .A2(n10700), .ZN(n10422) );
  AND2_X1 U13373 ( .A1(n11261), .A2(n11260), .ZN(n10423) );
  AND2_X1 U13374 ( .A1(n11198), .A2(n15055), .ZN(n10424) );
  AND2_X1 U13375 ( .A1(n9574), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10425) );
  AND2_X1 U13376 ( .A1(n9666), .A2(n12897), .ZN(n10426) );
  OR2_X1 U13377 ( .A1(n15879), .A2(n15870), .ZN(n10427) );
  OR2_X1 U13378 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n17454), .ZN(n10428) );
  INV_X1 U13379 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14555) );
  AND2_X1 U13380 ( .A1(n12892), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10429) );
  AND2_X1 U13381 ( .A1(n12899), .A2(n13737), .ZN(n10430) );
  INV_X1 U13382 ( .A(n11587), .ZN(n11588) );
  INV_X1 U13383 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10899) );
  OR4_X1 U13384 ( .A1(n15333), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n10431) );
  NAND3_X1 U13385 ( .A1(n14103), .A2(n19404), .A3(n17420), .ZN(n10432) );
  NOR2_X1 U13386 ( .A1(n14254), .A2(n14257), .ZN(n10433) );
  AND3_X1 U13387 ( .A1(n18834), .A2(n18868), .A3(n18890), .ZN(n10435) );
  OR2_X1 U13388 ( .A1(n17422), .A2(n19570), .ZN(n10436) );
  AND2_X1 U13389 ( .A1(n12693), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10437) );
  INV_X1 U13390 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17605) );
  INV_X1 U13391 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11597) );
  INV_X1 U13392 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16551) );
  INV_X1 U13393 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13066) );
  OR2_X1 U13394 ( .A1(n12728), .A2(n13649), .ZN(n10438) );
  AND2_X1 U13395 ( .A1(n11723), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10439) );
  INV_X1 U13396 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12127) );
  OR2_X1 U13397 ( .A1(n20765), .A2(n20819), .ZN(n14326) );
  INV_X2 U13398 ( .A(n14326), .ZN(n20770) );
  INV_X1 U13399 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18931) );
  OR2_X1 U13400 ( .A1(n17170), .A2(n21143), .ZN(n10440) );
  AND2_X1 U13401 ( .A1(n11657), .A2(n11656), .ZN(n10444) );
  AND2_X1 U13402 ( .A1(n11650), .A2(n11649), .ZN(n10445) );
  INV_X1 U13403 ( .A(n18316), .ZN(n18312) );
  AND3_X1 U13404 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .A3(P3_EAX_REG_14__SCAN_IN), .ZN(n10446) );
  AND4_X1 U13405 ( .A1(n12188), .A2(n12187), .A3(n12186), .A4(n12185), .ZN(
        n10447) );
  INV_X1 U13406 ( .A(n12613), .ZN(n12546) );
  INV_X1 U13407 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13787) );
  INV_X1 U13408 ( .A(n20685), .ZN(n17214) );
  INV_X1 U13409 ( .A(n13850), .ZN(n19834) );
  AND2_X1 U13410 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10449) );
  NAND3_X1 U13411 ( .A1(n12344), .A2(n12343), .A3(n12342), .ZN(n10450) );
  AND2_X1 U13412 ( .A1(n15807), .A2(n13964), .ZN(n10451) );
  AND2_X1 U13413 ( .A1(n19950), .A2(n14146), .ZN(n19946) );
  INV_X1 U13414 ( .A(n19946), .ZN(n19928) );
  NOR2_X2 U13415 ( .A1(n20178), .A2(n16765), .ZN(n10453) );
  OR2_X1 U13416 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20597), .ZN(n19841) );
  NAND2_X1 U13417 ( .A1(n12410), .A2(n13909), .ZN(n12428) );
  AND3_X1 U13418 ( .A1(n10530), .A2(n10529), .A3(n10528), .ZN(n10454) );
  AND4_X1 U13419 ( .A1(n10500), .A2(n10499), .A3(n10498), .A4(n10497), .ZN(
        n10455) );
  NAND2_X1 U13420 ( .A1(n10693), .A2(n10875), .ZN(n10662) );
  INV_X1 U13421 ( .A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10485) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n16717), .B1(
        n16728), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12520) );
  INV_X1 U13423 ( .A(n10633), .ZN(n10717) );
  INV_X1 U13424 ( .A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10477) );
  INV_X1 U13425 ( .A(n10736), .ZN(n10693) );
  AOI22_X1 U13426 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11649) );
  INV_X1 U13427 ( .A(n11739), .ZN(n11740) );
  NAND2_X1 U13428 ( .A1(n12191), .A2(n12190), .ZN(n12192) );
  NOR2_X1 U13429 ( .A1(n11656), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12119) );
  INV_X1 U13430 ( .A(n10952), .ZN(n10949) );
  NAND2_X1 U13431 ( .A1(n21143), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10946) );
  INV_X1 U13432 ( .A(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10569) );
  NOR2_X1 U13433 ( .A1(n10725), .A2(n10724), .ZN(n10810) );
  NAND2_X1 U13434 ( .A1(n10598), .A2(n10599), .ZN(n10590) );
  NAND2_X1 U13435 ( .A1(n16100), .A2(n16116), .ZN(n12606) );
  NOR2_X1 U13436 ( .A1(n12193), .A2(n12192), .ZN(n12194) );
  INV_X1 U13437 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16656) );
  INV_X1 U13438 ( .A(n14097), .ZN(n13482) );
  NOR2_X1 U13439 ( .A1(n10949), .A2(n10951), .ZN(n10950) );
  OR2_X1 U13440 ( .A1(n10922), .A2(n10921), .ZN(n10932) );
  OR2_X1 U13441 ( .A1(n10768), .A2(n10767), .ZN(n10796) );
  AND4_X1 U13442 ( .A1(n15100), .A2(n14959), .A3(n14974), .A4(n15081), .ZN(
        n11100) );
  OR2_X1 U13443 ( .A1(n10680), .A2(n10679), .ZN(n10815) );
  OR2_X1 U13444 ( .A1(n10707), .A2(n10706), .ZN(n10708) );
  AND4_X1 U13445 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        n10480) );
  INV_X1 U13446 ( .A(n15950), .ZN(n12825) );
  OR2_X1 U13447 ( .A1(n11734), .A2(n11733), .ZN(n11735) );
  INV_X1 U13448 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n13509) );
  INV_X1 U13449 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13334) );
  AOI21_X1 U13450 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21184), .A(
        n10950), .ZN(n10963) );
  AOI22_X1 U13451 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10549) );
  INV_X1 U13452 ( .A(n11283), .ZN(n11284) );
  NAND2_X1 U13453 ( .A1(n15595), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11570) );
  INV_X1 U13454 ( .A(n11161), .ZN(n11102) );
  NAND2_X1 U13455 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10904) );
  NAND2_X1 U13456 ( .A1(n10896), .A2(n10899), .ZN(n10900) );
  INV_X1 U13457 ( .A(n14913), .ZN(n12986) );
  INV_X1 U13458 ( .A(n15101), .ZN(n12958) );
  INV_X1 U13459 ( .A(n13028), .ZN(n10601) );
  NAND2_X1 U13460 ( .A1(n10735), .A2(n10734), .ZN(n20968) );
  OR2_X1 U13461 ( .A1(n12129), .A2(n12128), .ZN(n12131) );
  INV_X1 U13462 ( .A(n14119), .ZN(n12331) );
  NAND2_X1 U13463 ( .A1(n11683), .A2(n11656), .ZN(n11684) );
  INV_X1 U13464 ( .A(n16101), .ZN(n13080) );
  NOR2_X1 U13465 ( .A1(n12523), .A2(n16399), .ZN(n12757) );
  AND2_X1 U13466 ( .A1(n16190), .A2(n16193), .ZN(n13651) );
  INV_X1 U13467 ( .A(n12523), .ZN(n12769) );
  NOR2_X1 U13468 ( .A1(n19945), .A2(n15847), .ZN(n12429) );
  INV_X1 U13469 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13491) );
  NOR2_X1 U13470 ( .A1(n13476), .A2(n13475), .ZN(n13488) );
  INV_X1 U13471 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n21549) );
  AOI221_X1 U13472 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10963), 
        .C1(n17275), .C2(n10963), .A(n10962), .ZN(n12910) );
  INV_X1 U13473 ( .A(n11196), .ZN(n11026) );
  INV_X1 U13474 ( .A(n14757), .ZN(n11488) );
  INV_X1 U13475 ( .A(n11570), .ZN(n11539) );
  INV_X1 U13476 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17191) );
  NAND2_X1 U13477 ( .A1(n12910), .A2(n10966), .ZN(n10967) );
  NOR2_X1 U13478 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13735) );
  AND2_X1 U13479 ( .A1(n11005), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11574) );
  NAND2_X1 U13480 ( .A1(n12131), .A2(n12130), .ZN(n12572) );
  AND2_X1 U13481 ( .A1(n12852), .A2(n12851), .ZN(n13588) );
  INV_X1 U13482 ( .A(n14595), .ZN(n14587) );
  INV_X1 U13483 ( .A(n16059), .ZN(n12352) );
  INV_X1 U13484 ( .A(n13911), .ZN(n12321) );
  AND2_X1 U13485 ( .A1(n13652), .A2(n13651), .ZN(n13653) );
  AND2_X1 U13486 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16552) );
  NOR2_X1 U13487 ( .A1(n16589), .A2(n13153), .ZN(n16578) );
  INV_X1 U13488 ( .A(n12894), .ZN(n11776) );
  AND2_X1 U13489 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19433), .ZN(
        n13505) );
  INV_X1 U13490 ( .A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17081) );
  NOR2_X1 U13491 ( .A1(n19570), .A2(n18992), .ZN(n13479) );
  INV_X1 U13492 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21565) );
  INV_X1 U13493 ( .A(n21419), .ZN(n21501) );
  INV_X1 U13494 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n14914) );
  INV_X1 U13495 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14932) );
  INV_X1 U13496 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U13497 ( .A1(n13716), .A2(n13715), .ZN(n20687) );
  AND2_X1 U13498 ( .A1(n12976), .A2(n12975), .ZN(n14947) );
  AOI21_X1 U13499 ( .B1(n11027), .B2(n11026), .A(n11025), .ZN(n14497) );
  OR2_X1 U13500 ( .A1(n13999), .A2(n13937), .ZN(n13603) );
  INV_X1 U13501 ( .A(n11573), .ZN(n11431) );
  INV_X1 U13502 ( .A(n15054), .ZN(n15059) );
  INV_X1 U13503 ( .A(n14250), .ZN(n10992) );
  INV_X1 U13504 ( .A(n20773), .ZN(n15271) );
  AND2_X1 U13505 ( .A1(n15333), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13738) );
  INV_X1 U13506 ( .A(n20811), .ZN(n15555) );
  OR3_X1 U13507 ( .A1(n13999), .A2(n12917), .A3(n20824), .ZN(n12918) );
  INV_X1 U13508 ( .A(n17173), .ZN(n14578) );
  AND2_X1 U13509 ( .A1(n20934), .A2(n20961), .ZN(n20940) );
  NOR2_X1 U13510 ( .A1(n20973), .A2(n14505), .ZN(n21149) );
  NOR2_X1 U13511 ( .A1(n20974), .A2(n20973), .ZN(n21301) );
  NOR2_X1 U13512 ( .A1(n14037), .A2(n21222), .ZN(n17173) );
  INV_X1 U13513 ( .A(n12572), .ZN(n20610) );
  NOR2_X1 U13514 ( .A1(n14688), .A2(n10449), .ZN(n14689) );
  NAND2_X1 U13515 ( .A1(n19594), .A2(n14622), .ZN(n19782) );
  NOR2_X1 U13516 ( .A1(n13116), .A2(n13115), .ZN(n13117) );
  AND2_X1 U13517 ( .A1(n12354), .A2(n12353), .ZN(n15736) );
  INV_X1 U13518 ( .A(n13594), .ZN(n13595) );
  AND2_X1 U13519 ( .A1(n12361), .A2(n12360), .ZN(n15700) );
  OR3_X1 U13520 ( .A1(n16562), .A2(n16551), .A3(n16563), .ZN(n14552) );
  AND2_X1 U13521 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20302) );
  OR2_X1 U13522 ( .A1(n20590), .A2(n16744), .ZN(n16765) );
  OR2_X1 U13523 ( .A1(n20247), .A2(n16765), .ZN(n20383) );
  OR2_X1 U13524 ( .A1(n20269), .A2(n20574), .ZN(n20384) );
  INV_X1 U13525 ( .A(n17127), .ZN(n14398) );
  NOR2_X1 U13526 ( .A1(n18480), .A2(n17539), .ZN(n17538) );
  NAND2_X1 U13527 ( .A1(n19586), .A2(n18992), .ZN(n13778) );
  AND4_X1 U13528 ( .A1(n13325), .A2(n13324), .A3(n13323), .A4(n13322), .ZN(
        n13326) );
  AND4_X1 U13529 ( .A1(n13195), .A2(n13194), .A3(n13193), .A4(n13192), .ZN(
        n13207) );
  NAND2_X1 U13530 ( .A1(n16883), .A2(n18708), .ZN(n18495) );
  NOR2_X1 U13531 ( .A1(n18889), .A2(n18890), .ZN(n18617) );
  AND2_X1 U13532 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18858), .ZN(
        n18847) );
  OR2_X1 U13533 ( .A1(n18890), .A2(n18634), .ZN(n18615) );
  NOR2_X1 U13534 ( .A1(n18863), .A2(n18809), .ZN(n18891) );
  INV_X1 U13535 ( .A(n18978), .ZN(n18927) );
  INV_X1 U13536 ( .A(n19270), .ZN(n19246) );
  OAI211_X1 U13537 ( .C1(n14165), .C2(n14164), .A(n14163), .B(n14207), .ZN(
        n19418) );
  NOR2_X1 U13538 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21403), .ZN(n21508) );
  INV_X1 U13539 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14901) );
  INV_X1 U13540 ( .A(n20687), .ZN(n20672) );
  NOR2_X1 U13541 ( .A1(n15181), .A2(n17324), .ZN(n13617) );
  INV_X1 U13542 ( .A(n15181), .ZN(n15171) );
  NAND2_X1 U13543 ( .A1(n17230), .A2(n10601), .ZN(n14031) );
  NAND2_X1 U13544 ( .A1(n17170), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n20626) );
  NOR2_X1 U13545 ( .A1(n15094), .A2(n14958), .ZN(n15082) );
  INV_X1 U13546 ( .A(n17244), .ZN(n20779) );
  INV_X1 U13547 ( .A(n17278), .ZN(n11577) );
  NOR2_X1 U13548 ( .A1(n20799), .A2(n15529), .ZN(n17266) );
  AND2_X1 U13549 ( .A1(n20811), .A2(n20810), .ZN(n15539) );
  NAND2_X1 U13550 ( .A1(n10276), .A2(n14510), .ZN(n20973) );
  OR2_X1 U13551 ( .A1(n20933), .A2(n21292), .ZN(n14515) );
  OAI22_X1 U13552 ( .A1(n20898), .A2(n20897), .B1(n21154), .B2(n21029), .ZN(
        n20922) );
  OAI22_X1 U13553 ( .A1(n20940), .A2(n20939), .B1(n11005), .B2(n20938), .ZN(
        n20964) );
  OAI21_X1 U13554 ( .B1(n21293), .B2(n20970), .A(n20969), .ZN(n20991) );
  OAI22_X1 U13555 ( .A1(n21031), .A2(n21030), .B1(n21029), .B2(n21293), .ZN(
        n21054) );
  OAI211_X1 U13556 ( .C1(n21027), .C2(n21222), .A(n21301), .B(n21026), .ZN(
        n21055) );
  OAI211_X1 U13557 ( .C1(n21111), .C2(n21222), .A(n21149), .B(n21095), .ZN(
        n21112) );
  INV_X1 U13558 ( .A(n21183), .ZN(n21145) );
  OAI22_X1 U13559 ( .A1(n21156), .A2(n21155), .B1(n21154), .B2(n21294), .ZN(
        n21179) );
  INV_X1 U13560 ( .A(n21262), .ZN(n21210) );
  OAI22_X1 U13561 ( .A1(n21227), .A2(n21226), .B1(n21225), .B2(n21293), .ZN(
        n21258) );
  NAND2_X1 U13562 ( .A1(n14501), .A2(n10975), .ZN(n21193) );
  OAI211_X1 U13563 ( .C1(n21330), .C2(n21302), .A(n21301), .B(n21300), .ZN(
        n21332) );
  INV_X1 U13564 ( .A(n21345), .ZN(n21296) );
  NOR2_X1 U13565 ( .A1(n12906), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n17186) );
  INV_X1 U13566 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n21415) );
  INV_X1 U13567 ( .A(n19782), .ZN(n19736) );
  INV_X1 U13568 ( .A(n12333), .ZN(n15944) );
  INV_X1 U13569 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n15973) );
  OAI21_X1 U13570 ( .B1(n13678), .B2(n13806), .A(n13810), .ZN(n13679) );
  XNOR2_X1 U13571 ( .A(n14012), .B(n14011), .ZN(n16744) );
  AND2_X1 U13572 ( .A1(n12351), .A2(n12350), .ZN(n16059) );
  AND3_X1 U13573 ( .A1(n12320), .A2(n12319), .A3(n12318), .ZN(n13911) );
  INV_X1 U13574 ( .A(n16062), .ZN(n19828) );
  INV_X1 U13575 ( .A(n13876), .ZN(n19909) );
  AND2_X1 U13576 ( .A1(n16830), .A2(n20382), .ZN(n16341) );
  INV_X1 U13577 ( .A(n19950), .ZN(n17289) );
  INV_X1 U13578 ( .A(n16485), .ZN(n16512) );
  AND2_X1 U13579 ( .A1(n14552), .A2(n14551), .ZN(n16545) );
  INV_X1 U13580 ( .A(n19959), .ZN(n16645) );
  NOR2_X1 U13581 ( .A1(n16816), .A2(n12562), .ZN(n20609) );
  INV_X1 U13582 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14633) );
  INV_X1 U13583 ( .A(n16745), .ZN(n20601) );
  NOR2_X2 U13584 ( .A1(n20246), .A2(n20178), .ZN(n20078) );
  AND2_X1 U13585 ( .A1(n20090), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20109) );
  OAI21_X1 U13586 ( .B1(n16730), .B2(n20575), .A(n16729), .ZN(n20174) );
  OAI21_X1 U13587 ( .B1(n20213), .B2(n20581), .A(n20186), .ZN(n20203) );
  NOR2_X2 U13588 ( .A1(n20247), .A2(n20246), .ZN(n20296) );
  NOR2_X2 U13589 ( .A1(n20269), .A2(n20308), .ZN(n20335) );
  NOR2_X1 U13590 ( .A1(n20247), .A2(n20308), .ZN(n20358) );
  AND2_X1 U13591 ( .A1(n16766), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20387) );
  INV_X1 U13592 ( .A(n19822), .ZN(n19995) );
  INV_X1 U13593 ( .A(n20383), .ZN(n20427) );
  INV_X1 U13594 ( .A(n20431), .ZN(n20470) );
  NAND2_X1 U13595 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20480) );
  AND3_X1 U13596 ( .A1(n20496), .A2(n20558), .A3(n20501), .ZN(n20495) );
  INV_X1 U13597 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20507) );
  INV_X1 U13598 ( .A(n18983), .ZN(n19567) );
  OAI211_X1 U13599 ( .C1(n17464), .C2(n19459), .A(n10428), .B(n17463), .ZN(
        n17465) );
  NOR2_X1 U13600 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17519), .ZN(n17503) );
  NOR2_X1 U13601 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17543), .ZN(n17527) );
  INV_X1 U13602 ( .A(n17786), .ZN(n17811) );
  NOR2_X1 U13603 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17650), .ZN(n17632) );
  OR3_X1 U13604 ( .A1(n19504), .A2(n19501), .A3(n17631), .ZN(n17608) );
  NOR2_X1 U13605 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17753), .ZN(n17735) );
  INV_X1 U13606 ( .A(n17812), .ZN(n17764) );
  INV_X1 U13607 ( .A(n17822), .ZN(n17007) );
  INV_X1 U13608 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n18006) );
  INV_X1 U13609 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17675) );
  NOR2_X1 U13610 ( .A1(n19570), .A2(n14214), .ZN(n17006) );
  OR4_X1 U13611 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17874) );
  NOR3_X1 U13612 ( .A1(n19024), .A2(n18259), .A3(n18383), .ZN(n18251) );
  OR2_X1 U13613 ( .A1(n13303), .A2(n13302), .ZN(n13306) );
  INV_X1 U13614 ( .A(n18321), .ZN(n18310) );
  INV_X1 U13615 ( .A(n18376), .ZN(n18323) );
  OAI211_X1 U13616 ( .C1(n19572), .C2(n19570), .A(n18379), .B(n18378), .ZN(
        n18417) );
  OR2_X1 U13617 ( .A1(n13568), .A2(n13567), .ZN(n13569) );
  NOR2_X2 U13618 ( .A1(n18674), .A2(n19451), .ZN(n18529) );
  AND2_X1 U13619 ( .A1(n19323), .A2(n19271), .ZN(n19351) );
  NAND2_X1 U13620 ( .A1(n18708), .A2(n16928), .ZN(n18674) );
  INV_X1 U13621 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18800) );
  OR2_X1 U13622 ( .A1(n18661), .A2(n10057), .ZN(n18634) );
  INV_X1 U13623 ( .A(n18913), .ZN(n18936) );
  AND2_X1 U13624 ( .A1(n19399), .A2(n18958), .ZN(n18870) );
  INV_X1 U13625 ( .A(n18888), .ZN(n18958) );
  INV_X1 U13626 ( .A(n19344), .ZN(n19324) );
  INV_X1 U13627 ( .A(n19050), .ZN(n19104) );
  INV_X1 U13628 ( .A(n21669), .ZN(n19127) );
  INV_X1 U13629 ( .A(n19109), .ZN(n19150) );
  INV_X1 U13630 ( .A(n19132), .ZN(n19198) );
  INV_X1 U13631 ( .A(n19154), .ZN(n19220) );
  INV_X1 U13632 ( .A(n19178), .ZN(n19241) );
  INV_X1 U13633 ( .A(n19272), .ZN(n19340) );
  INV_X1 U13634 ( .A(n19318), .ZN(n19454) );
  INV_X1 U13635 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19480) );
  NAND2_X1 U13636 ( .A1(n12386), .A2(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n16714)
         );
  INV_X1 U13637 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21497) );
  AOI21_X1 U13638 ( .B1(n15376), .B2(n20705), .A(n14742), .ZN(n14743) );
  INV_X1 U13639 ( .A(n20705), .ZN(n20650) );
  OR2_X1 U13640 ( .A1(n15096), .A2(n14045), .ZN(n15099) );
  INV_X1 U13641 ( .A(n15096), .ZN(n15104) );
  OR2_X1 U13642 ( .A1(n14031), .A2(n14509), .ZN(n15181) );
  AND2_X1 U13643 ( .A1(n14312), .A2(n14311), .ZN(n20857) );
  NAND2_X2 U13644 ( .A1(n17230), .A2(n14029), .ZN(n15195) );
  NAND2_X1 U13645 ( .A1(n20718), .A2(n14511), .ZN(n14248) );
  INV_X1 U13646 ( .A(n20765), .ZN(n14327) );
  NOR2_X1 U13647 ( .A1(n13756), .A2(n13755), .ZN(n13757) );
  OR2_X1 U13648 ( .A1(n14783), .A2(n14850), .ZN(n15266) );
  OR2_X1 U13649 ( .A1(n17155), .A2(n20626), .ZN(n20631) );
  INV_X1 U13650 ( .A(n20801), .ZN(n15571) );
  AOI22_X1 U13651 ( .A1(n15539), .A2(n14471), .B1(n20805), .B2(n14470), .ZN(
        n20799) );
  INV_X1 U13652 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21143) );
  INV_X1 U13653 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n17275) );
  AOI211_X1 U13654 ( .C1(n14508), .C2(n14515), .A(n20894), .B(n14507), .ZN(
        n20851) );
  NAND2_X1 U13655 ( .A1(n20926), .A2(n21215), .ZN(n20888) );
  NAND2_X1 U13656 ( .A1(n20926), .A2(n21263), .ZN(n20920) );
  NAND2_X1 U13657 ( .A1(n20926), .A2(n21295), .ZN(n20962) );
  NAND2_X1 U13658 ( .A1(n20926), .A2(n21191), .ZN(n20990) );
  NAND2_X1 U13659 ( .A1(n21059), .A2(n21215), .ZN(n21016) );
  NAND2_X1 U13660 ( .A1(n21059), .A2(n21263), .ZN(n21058) );
  NAND2_X1 U13661 ( .A1(n21059), .A2(n21295), .ZN(n21087) );
  NAND2_X1 U13662 ( .A1(n21059), .A2(n21191), .ZN(n21115) );
  OR2_X1 U13663 ( .A1(n21193), .A2(n21091), .ZN(n21135) );
  OR2_X1 U13664 ( .A1(n21193), .A2(n21116), .ZN(n21183) );
  OR2_X1 U13665 ( .A1(n21193), .A2(n21142), .ZN(n21214) );
  OR2_X1 U13666 ( .A1(n21193), .A2(n21192), .ZN(n21262) );
  NAND2_X1 U13667 ( .A1(n21296), .A2(n21215), .ZN(n21285) );
  INV_X1 U13668 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21403) );
  OAI21_X1 U13669 ( .B1(n21415), .B2(n21418), .A(n21495), .ZN(n21407) );
  INV_X1 U13670 ( .A(n21407), .ZN(n21486) );
  NAND2_X1 U13671 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n21419) );
  INV_X1 U13672 ( .A(n21474), .ZN(n21468) );
  NAND2_X1 U13673 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21511), .ZN(n21472) );
  INV_X1 U13674 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20496) );
  INV_X1 U13675 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19970) );
  INV_X1 U13676 ( .A(n19754), .ZN(n19786) );
  INV_X1 U13677 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19671) );
  INV_X1 U13678 ( .A(n19777), .ZN(n19775) );
  INV_X1 U13679 ( .A(n13679), .ZN(n16002) );
  AND2_X1 U13680 ( .A1(n16081), .A2(n16062), .ZN(n16096) );
  AND2_X1 U13681 ( .A1(n13880), .A2(n13879), .ZN(n19821) );
  INV_X1 U13682 ( .A(n19823), .ZN(n16081) );
  NAND2_X1 U13683 ( .A1(n19840), .A2(n19839), .ZN(n19871) );
  NAND2_X1 U13684 ( .A1(n19837), .A2(n20495), .ZN(n19905) );
  INV_X1 U13685 ( .A(n13961), .ZN(n13874) );
  INV_X1 U13686 ( .A(n19936), .ZN(n17292) );
  NAND2_X1 U13687 ( .A1(n12778), .A2(n19985), .ZN(n19941) );
  INV_X1 U13688 ( .A(n19962), .ZN(n16648) );
  INV_X1 U13689 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17306) );
  INV_X1 U13690 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20586) );
  OAI22_X1 U13691 ( .A1(n19975), .A2(n20014), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19979), .ZN(n20018) );
  AOI211_X2 U13692 ( .C1(n20020), .C2(n20023), .A(n20019), .B(n20183), .ZN(
        n20048) );
  AOI21_X1 U13693 ( .B1(n20054), .B2(n20382), .A(n20053), .ZN(n20082) );
  AOI21_X1 U13694 ( .B1(n20092), .B2(n20090), .A(n20087), .ZN(n20113) );
  AOI211_X2 U13695 ( .C1(n16711), .C2(n16710), .A(n20183), .B(n16709), .ZN(
        n20162) );
  AOI211_X2 U13696 ( .C1(n16727), .C2(n16730), .A(n16726), .B(n20183), .ZN(
        n20177) );
  INV_X1 U13697 ( .A(n10443), .ZN(n20206) );
  OAI22_X1 U13698 ( .A1(n20211), .A2(n20210), .B1(n20209), .B2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n20236) );
  AOI21_X1 U13699 ( .B1(n20243), .B2(n20241), .A(n20238), .ZN(n20267) );
  AOI21_X1 U13700 ( .B1(n20276), .B2(n20279), .A(n20275), .ZN(n20300) );
  INV_X1 U13701 ( .A(n20358), .ZN(n20339) );
  AOI21_X1 U13702 ( .B1(n16754), .B2(n16753), .A(n16752), .ZN(n20362) );
  OAI22_X1 U13703 ( .A1(n20391), .A2(n20426), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n20396), .ZN(n20432) );
  NOR2_X1 U13704 ( .A1(n16780), .A2(n16779), .ZN(n20479) );
  INV_X1 U13705 ( .A(n13810), .ZN(n20481) );
  OAI21_X1 U13706 ( .B1(n20496), .B2(n20500), .A(n20497), .ZN(n20573) );
  INV_X1 U13707 ( .A(n20573), .ZN(n20570) );
  NOR2_X1 U13708 ( .A1(n19403), .A2(n18380), .ZN(n19586) );
  OR2_X2 U13709 ( .A1(n19409), .A2(n19449), .ZN(n17423) );
  INV_X1 U13710 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17734) );
  NAND2_X1 U13711 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n17816), .ZN(n17791) );
  NOR2_X1 U13712 ( .A1(n17830), .A2(n17829), .ZN(n17860) );
  INV_X1 U13713 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17653) );
  AND2_X1 U13714 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n18284), .ZN(n18281) );
  INV_X1 U13715 ( .A(n17130), .ZN(n18302) );
  INV_X1 U13716 ( .A(n13532), .ZN(n18317) );
  NAND2_X1 U13717 ( .A1(n14354), .A2(n14279), .ZN(n18318) );
  NAND2_X1 U13718 ( .A1(n18323), .A2(n18992), .ZN(n18348) );
  NAND2_X1 U13719 ( .A1(n18378), .A2(n18322), .ZN(n18376) );
  INV_X1 U13720 ( .A(n18425), .ZN(n18419) );
  AOI21_X1 U13721 ( .B1(n13571), .B2(n13570), .A(n13569), .ZN(n13572) );
  NOR2_X1 U13722 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18670) );
  INV_X1 U13723 ( .A(n18681), .ZN(n18653) );
  INV_X1 U13724 ( .A(n18714), .ZN(n18720) );
  OR2_X1 U13725 ( .A1(n18971), .A2(n18302), .ZN(n18913) );
  INV_X1 U13726 ( .A(n18870), .ZN(n18973) );
  NAND2_X1 U13727 ( .A1(n16961), .A2(n18958), .ZN(n18971) );
  INV_X1 U13728 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19433) );
  INV_X1 U13729 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n19410) );
  INV_X1 U13730 ( .A(n19175), .ZN(n19108) );
  INV_X1 U13731 ( .A(n19395), .ZN(n19317) );
  NAND2_X1 U13732 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19456), .ZN(n19449) );
  INV_X1 U13733 ( .A(n17784), .ZN(n19459) );
  INV_X1 U13734 ( .A(n19550), .ZN(n19547) );
  INV_X1 U13735 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19501) );
  INV_X1 U13736 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n21548) );
  NAND2_X1 U13737 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19479), .ZN(n19581) );
  INV_X1 U13738 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n19020) );
  INV_X1 U13739 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20512) );
  OAI21_X1 U13740 ( .B1(n15491), .B2(n20631), .A(n11605), .ZN(P1_U2982) );
  OAI21_X1 U13741 ( .B1(n13758), .B2(n20807), .A(n13065), .ZN(P1_U3002) );
  OR4_X1 U13742 ( .A1(n13784), .A2(n13783), .A3(n13782), .A4(n13781), .ZN(
        P3_U2651) );
  NAND2_X1 U13743 ( .A1(n13573), .A2(n13572), .ZN(P3_U2801) );
  AND2_X4 U13744 ( .A1(n10469), .A2(n10468), .ZN(n10634) );
  NAND2_X1 U13745 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13746 ( .A1(n10626), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10459) );
  NAND2_X1 U13747 ( .A1(n10635), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10458) );
  INV_X2 U13748 ( .A(n11465), .ZN(n10527) );
  NAND2_X1 U13749 ( .A1(n10527), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10457) );
  NAND4_X1 U13750 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10463) );
  INV_X1 U13751 ( .A(n10544), .ZN(n10461) );
  NOR2_X1 U13752 ( .A1(n10461), .A2(n10756), .ZN(n10462) );
  NOR2_X1 U13753 ( .A1(n10463), .A2(n10462), .ZN(n10482) );
  NAND2_X1 U13754 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13755 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13756 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10465) );
  NAND2_X1 U13757 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13758 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10473) );
  AND2_X2 U13759 ( .A1(n10474), .A2(n14409), .ZN(n10632) );
  NAND2_X1 U13760 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U13761 ( .A1(n10650), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10471) );
  NAND2_X1 U13762 ( .A1(n10627), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13763 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10475) );
  OAI211_X1 U13764 ( .C1(n10570), .C2(n10477), .A(n10476), .B(n10475), .ZN(
        n10478) );
  INV_X1 U13765 ( .A(n10478), .ZN(n10479) );
  NAND2_X1 U13766 ( .A1(n10650), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10484) );
  NAND2_X1 U13767 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10483) );
  OAI211_X1 U13768 ( .C1(n10570), .C2(n10485), .A(n10484), .B(n10483), .ZN(
        n10486) );
  INV_X1 U13769 ( .A(n10486), .ZN(n10491) );
  AOI22_X1 U13770 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10626), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10489) );
  AOI22_X1 U13771 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10488) );
  NAND2_X1 U13772 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10487) );
  AOI22_X1 U13773 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10527), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U13774 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10632), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10493) );
  AOI22_X1 U13775 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10492) );
  AOI22_X1 U13776 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10663), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U13777 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10622), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U13778 ( .A1(n10626), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10527), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10498) );
  AOI22_X1 U13779 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10497) );
  NAND2_X1 U13780 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13781 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13782 ( .A1(n10576), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13783 ( .A1(n10635), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10501) );
  AOI22_X1 U13784 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10650), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U13785 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n10507) );
  INV_X1 U13786 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10505) );
  INV_X1 U13787 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10513) );
  NAND2_X1 U13788 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10511) );
  OAI211_X1 U13789 ( .C1(n10570), .C2(n10513), .A(n10512), .B(n10511), .ZN(
        n10514) );
  INV_X1 U13790 ( .A(n10514), .ZN(n10520) );
  NAND2_X1 U13791 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10516) );
  AOI22_X1 U13792 ( .A1(n10527), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U13793 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n10517) );
  NAND4_X1 U13794 ( .A1(n10520), .A2(n10519), .A3(n10518), .A4(n10517), .ZN(
        n10526) );
  AOI22_X1 U13795 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10521) );
  NAND4_X1 U13796 ( .A1(n10524), .A2(n10523), .A3(n10522), .A4(n10521), .ZN(
        n10525) );
  OR2_X2 U13797 ( .A1(n10526), .A2(n10525), .ZN(n10587) );
  AOI22_X1 U13798 ( .A1(n10626), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10527), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13799 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10530) );
  NAND2_X1 U13800 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10528) );
  INV_X2 U13801 ( .A(n10570), .ZN(n11472) );
  NAND2_X1 U13802 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10531) );
  NAND4_X1 U13803 ( .A1(n10533), .A2(n10454), .A3(n10532), .A4(n10531), .ZN(
        n10539) );
  AOI22_X1 U13804 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10650), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13805 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10634), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13806 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10663), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13807 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13808 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10538) );
  INV_X1 U13809 ( .A(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10542) );
  NAND2_X1 U13810 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10540) );
  OAI211_X1 U13811 ( .C1(n10570), .C2(n10542), .A(n10541), .B(n10540), .ZN(
        n10543) );
  INV_X1 U13812 ( .A(n10543), .ZN(n10548) );
  AOI22_X1 U13813 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10626), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13814 ( .A1(n10527), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10546) );
  NAND2_X1 U13815 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10545) );
  NAND4_X1 U13816 ( .A1(n10548), .A2(n10547), .A3(n10546), .A4(n10545), .ZN(
        n10554) );
  AOI22_X1 U13817 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10552) );
  AOI22_X1 U13818 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10577), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13819 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10650), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10550) );
  NAND4_X1 U13820 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10553) );
  INV_X1 U13821 ( .A(n14039), .ZN(n13986) );
  INV_X1 U13822 ( .A(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10557) );
  NAND2_X1 U13823 ( .A1(n10663), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10556) );
  OAI211_X1 U13824 ( .C1(n10570), .C2(n10557), .A(n10556), .B(n10555), .ZN(
        n10558) );
  INV_X1 U13825 ( .A(n10558), .ZN(n10562) );
  AOI22_X1 U13826 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10626), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13827 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10527), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10560) );
  NAND2_X1 U13828 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10559) );
  NAND4_X1 U13829 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n10568) );
  AOI22_X1 U13830 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10632), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13831 ( .A1(n10650), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10564) );
  AOI22_X1 U13832 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10563) );
  NAND4_X1 U13833 ( .A1(n10566), .A2(n10565), .A3(n10564), .A4(n10563), .ZN(
        n10567) );
  NAND2_X1 U13834 ( .A1(n13986), .A2(n14140), .ZN(n10584) );
  AOI22_X1 U13835 ( .A1(n10527), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U13836 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10626), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10574) );
  INV_X1 U13837 ( .A(n10571), .ZN(n10573) );
  NAND2_X1 U13838 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10572) );
  NAND4_X1 U13839 ( .A1(n10575), .A2(n10574), .A3(n10573), .A4(n10572), .ZN(
        n10583) );
  AOI22_X1 U13840 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10576), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10581) );
  AOI22_X1 U13841 ( .A1(n10633), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10577), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10580) );
  AOI22_X1 U13842 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10650), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13843 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10578) );
  NAND4_X1 U13844 ( .A1(n10581), .A2(n10580), .A3(n10579), .A4(n10578), .ZN(
        n10582) );
  NAND2_X1 U13845 ( .A1(n12902), .A2(n13599), .ZN(n10589) );
  INV_X2 U13846 ( .A(n10790), .ZN(n10916) );
  INV_X1 U13847 ( .A(n10590), .ZN(n10591) );
  NAND2_X1 U13848 ( .A1(n12904), .A2(n14576), .ZN(n10596) );
  INV_X1 U13849 ( .A(n10602), .ZN(n10970) );
  INV_X1 U13850 ( .A(n10594), .ZN(n20824) );
  NAND2_X1 U13851 ( .A1(n20824), .A2(n14511), .ZN(n10592) );
  INV_X1 U13852 ( .A(n12932), .ZN(n10593) );
  NAND2_X1 U13853 ( .A1(n12945), .A2(n10593), .ZN(n12927) );
  INV_X1 U13854 ( .A(n10969), .ZN(n10595) );
  AND2_X2 U13855 ( .A1(n10916), .A2(n10599), .ZN(n14030) );
  XNOR2_X1 U13856 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12906) );
  OAI211_X1 U13857 ( .C1(n13022), .C2(n12906), .A(n12925), .B(n13023), .ZN(
        n10604) );
  NOR2_X1 U13858 ( .A1(n10602), .A2(n14511), .ZN(n10603) );
  OAI21_X1 U13859 ( .B1(n10604), .B2(n12920), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n10688) );
  NAND2_X1 U13860 ( .A1(n10605), .A2(n10688), .ZN(n10730) );
  MUX2_X1 U13861 ( .A(n11584), .B(n17170), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n10606) );
  AND2_X1 U13862 ( .A1(n14576), .A2(n20819), .ZN(n10608) );
  NAND2_X1 U13863 ( .A1(n12904), .A2(n10608), .ZN(n10621) );
  NAND2_X1 U13864 ( .A1(n14039), .A2(n10609), .ZN(n13034) );
  INV_X1 U13865 ( .A(n10610), .ZN(n10611) );
  NAND2_X1 U13866 ( .A1(n10611), .A2(n21499), .ZN(n10613) );
  AND2_X1 U13867 ( .A1(n20624), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13868 ( .A1(n13707), .A2(n20819), .ZN(n15003) );
  NAND4_X1 U13869 ( .A1(n13034), .A2(n10613), .A3(n10612), .A4(n15003), .ZN(
        n10614) );
  NOR2_X1 U13870 ( .A1(n10615), .A2(n10614), .ZN(n10620) );
  OAI21_X1 U13871 ( .B1(n13862), .B2(n10617), .A(n10618), .ZN(n10619) );
  INV_X1 U13872 ( .A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11324) );
  NAND2_X1 U13873 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13874 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10623) );
  OAI211_X1 U13875 ( .C1(n11555), .C2(n11324), .A(n10624), .B(n10623), .ZN(
        n10625) );
  INV_X1 U13876 ( .A(n10625), .ZN(n10631) );
  INV_X1 U13877 ( .A(n10626), .ZN(n11544) );
  AOI22_X1 U13878 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10630) );
  INV_X2 U13879 ( .A(n11468), .ZN(n11316) );
  INV_X1 U13880 ( .A(n10627), .ZN(n11325) );
  AOI22_X1 U13881 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10629) );
  NAND2_X1 U13882 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10628) );
  NAND4_X1 U13883 ( .A1(n10631), .A2(n10630), .A3(n10629), .A4(n10628), .ZN(
        n10641) );
  AOI22_X1 U13884 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10639) );
  INV_X1 U13885 ( .A(n10632), .ZN(n10719) );
  INV_X1 U13886 ( .A(n10719), .ZN(n10664) );
  AOI22_X1 U13887 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10664), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10638) );
  INV_X2 U13888 ( .A(n10717), .ZN(n10669) );
  AOI22_X1 U13889 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10637) );
  INV_X1 U13890 ( .A(n10635), .ZN(n11352) );
  AOI22_X1 U13891 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10636) );
  NAND4_X1 U13892 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10640) );
  INV_X1 U13893 ( .A(n10875), .ZN(n10877) );
  INV_X1 U13894 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10644) );
  NAND2_X1 U13895 ( .A1(n9568), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10643) );
  NAND2_X1 U13896 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10642) );
  OAI211_X1 U13897 ( .C1(n11555), .C2(n10644), .A(n10643), .B(n10642), .ZN(
        n10645) );
  INV_X1 U13898 ( .A(n10645), .ZN(n10649) );
  AOI22_X1 U13899 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10648) );
  AOI22_X1 U13900 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13901 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10646) );
  NAND4_X1 U13902 ( .A1(n10649), .A2(n10648), .A3(n10647), .A4(n10646), .ZN(
        n10657) );
  AOI22_X1 U13903 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n11400), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10655) );
  AOI22_X1 U13904 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10654) );
  AOI22_X1 U13905 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10653) );
  AOI22_X1 U13906 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10652) );
  NAND4_X1 U13907 ( .A1(n10655), .A2(n10654), .A3(n10653), .A4(n10652), .ZN(
        n10656) );
  XNOR2_X1 U13908 ( .A(n10877), .B(n10820), .ZN(n10658) );
  NAND2_X1 U13909 ( .A1(n10658), .A2(n10693), .ZN(n10659) );
  AOI21_X1 U13910 ( .B1(n13599), .B2(n10875), .A(n10276), .ZN(n10661) );
  NAND2_X1 U13911 ( .A1(n13707), .A2(n10820), .ZN(n10660) );
  NAND2_X1 U13912 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10683) );
  INV_X1 U13913 ( .A(n10737), .ZN(n10681) );
  INV_X1 U13914 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10667) );
  NAND2_X1 U13915 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10666) );
  NAND2_X1 U13916 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10665) );
  OAI211_X1 U13917 ( .C1(n11555), .C2(n10667), .A(n10666), .B(n10665), .ZN(
        n10668) );
  INV_X1 U13918 ( .A(n10668), .ZN(n10673) );
  AOI22_X1 U13919 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10672) );
  AOI22_X1 U13920 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10671) );
  NAND2_X1 U13921 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10670) );
  NAND4_X1 U13922 ( .A1(n10673), .A2(n10672), .A3(n10671), .A4(n10670), .ZN(
        n10680) );
  AOI22_X1 U13923 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11400), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13924 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13925 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10676) );
  AOI22_X1 U13926 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10635), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10675) );
  NAND4_X1 U13927 ( .A1(n10678), .A2(n10677), .A3(n10676), .A4(n10675), .ZN(
        n10679) );
  NAND2_X1 U13928 ( .A1(n10681), .A2(n10815), .ZN(n10682) );
  OAI211_X1 U13929 ( .C1(n10736), .C2(n10875), .A(n10683), .B(n10682), .ZN(
        n10684) );
  NAND2_X1 U13930 ( .A1(n10730), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10687) );
  NAND2_X1 U13931 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10697) );
  OAI21_X1 U13932 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10697), .ZN(n21148) );
  OR2_X1 U13933 ( .A1(n17170), .A2(n21216), .ZN(n10705) );
  OAI21_X1 U13934 ( .B1(n11584), .B2(n21148), .A(n10705), .ZN(n10685) );
  INV_X1 U13935 ( .A(n10685), .ZN(n10686) );
  NAND2_X1 U13936 ( .A1(n10687), .A2(n10686), .ZN(n10689) );
  INV_X1 U13937 ( .A(n10690), .ZN(n10691) );
  NAND2_X1 U13938 ( .A1(n10693), .A2(n10815), .ZN(n10694) );
  NAND2_X1 U13939 ( .A1(n10976), .A2(n10695), .ZN(n10807) );
  INV_X1 U13940 ( .A(n10807), .ZN(n10729) );
  NAND2_X1 U13941 ( .A1(n10730), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10701) );
  INV_X1 U13942 ( .A(n11584), .ZN(n10699) );
  INV_X1 U13943 ( .A(n10697), .ZN(n10696) );
  NAND2_X1 U13944 ( .A1(n10696), .A2(n21143), .ZN(n21185) );
  NAND2_X1 U13945 ( .A1(n10697), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10698) );
  NAND2_X1 U13946 ( .A1(n21185), .A2(n10698), .ZN(n14514) );
  NAND2_X1 U13947 ( .A1(n10699), .A2(n14514), .ZN(n10700) );
  NAND2_X1 U13948 ( .A1(n10422), .A2(n10440), .ZN(n10704) );
  AND2_X1 U13949 ( .A1(n10702), .A2(n10704), .ZN(n10703) );
  INV_X1 U13950 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15596) );
  AND2_X1 U13951 ( .A1(n10705), .A2(n15596), .ZN(n10706) );
  INV_X1 U13952 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U13953 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10711) );
  NAND2_X1 U13954 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n10710) );
  OAI211_X1 U13955 ( .C1(n11555), .C2(n11355), .A(n10711), .B(n10710), .ZN(
        n10712) );
  INV_X1 U13956 ( .A(n10712), .ZN(n10716) );
  AOI22_X1 U13957 ( .A1(n10634), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13958 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10714) );
  NAND2_X1 U13959 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10713) );
  NAND4_X1 U13960 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        n10725) );
  AOI22_X1 U13961 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10723) );
  AOI22_X1 U13962 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10722) );
  INV_X1 U13963 ( .A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21612) );
  AOI22_X1 U13964 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10721) );
  AOI22_X1 U13965 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10627), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10720) );
  NAND4_X1 U13966 ( .A1(n10723), .A2(n10722), .A3(n10721), .A4(n10720), .ZN(
        n10724) );
  INV_X1 U13967 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10726) );
  OAI22_X1 U13968 ( .A1(n10737), .A2(n10810), .B1(n10936), .B2(n10726), .ZN(
        n10727) );
  INV_X1 U13969 ( .A(n10808), .ZN(n10728) );
  NAND2_X1 U13970 ( .A1(n10731), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10735) );
  NOR3_X1 U13971 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21143), .A3(
        n21216), .ZN(n21066) );
  NAND2_X1 U13972 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21066), .ZN(
        n21060) );
  NAND2_X1 U13973 ( .A1(n21184), .A2(n21060), .ZN(n10732) );
  NAND3_X1 U13974 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21340) );
  INV_X1 U13975 ( .A(n21340), .ZN(n21350) );
  NAND2_X1 U13976 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21350), .ZN(
        n21337) );
  NAND2_X1 U13977 ( .A1(n10732), .A2(n21337), .ZN(n21089) );
  OAI22_X1 U13978 ( .A1(n11584), .A2(n21089), .B1(n17170), .B2(n21184), .ZN(
        n10733) );
  INV_X1 U13979 ( .A(n10733), .ZN(n10734) );
  INV_X1 U13980 ( .A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13981 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13982 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10738) );
  OAI211_X1 U13983 ( .C1(n11555), .C2(n10740), .A(n10739), .B(n10738), .ZN(
        n10741) );
  INV_X1 U13984 ( .A(n10741), .ZN(n10746) );
  AOI22_X1 U13985 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13986 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10744) );
  NAND2_X1 U13987 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10743) );
  NAND4_X1 U13988 ( .A1(n10746), .A2(n10745), .A3(n10744), .A4(n10743), .ZN(
        n10752) );
  AOI22_X1 U13989 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10750) );
  AOI22_X1 U13990 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13991 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13992 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10747) );
  NAND4_X1 U13993 ( .A1(n10750), .A2(n10749), .A3(n10748), .A4(n10747), .ZN(
        n10751) );
  AOI22_X1 U13994 ( .A1(n10966), .A2(n10802), .B1(n10956), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10753) );
  NAND2_X1 U13995 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10755) );
  NAND2_X1 U13996 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10754) );
  OAI211_X1 U13997 ( .C1(n11555), .C2(n10756), .A(n10755), .B(n10754), .ZN(
        n10757) );
  INV_X1 U13998 ( .A(n10757), .ZN(n10761) );
  AOI22_X1 U13999 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U14000 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U14001 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10758) );
  NAND4_X1 U14002 ( .A1(n10761), .A2(n10760), .A3(n10759), .A4(n10758), .ZN(
        n10768) );
  AOI22_X1 U14003 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10766) );
  AOI22_X1 U14004 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10765) );
  AOI22_X1 U14005 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U14006 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10763) );
  NAND4_X1 U14007 ( .A1(n10766), .A2(n10765), .A3(n10764), .A4(n10763), .ZN(
        n10767) );
  NAND2_X1 U14008 ( .A1(n10966), .A2(n10796), .ZN(n10770) );
  NAND2_X1 U14009 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10769) );
  INV_X1 U14010 ( .A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U14011 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10772) );
  NAND2_X1 U14012 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10771) );
  OAI211_X1 U14013 ( .C1(n11555), .C2(n10773), .A(n10772), .B(n10771), .ZN(
        n10774) );
  INV_X1 U14014 ( .A(n10774), .ZN(n10778) );
  AOI22_X1 U14015 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10777) );
  INV_X1 U14016 ( .A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n21536) );
  AOI22_X1 U14017 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10776) );
  NAND2_X1 U14018 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10775) );
  NAND4_X1 U14019 ( .A1(n10778), .A2(n10777), .A3(n10776), .A4(n10775), .ZN(
        n10784) );
  AOI22_X1 U14020 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10782) );
  AOI22_X1 U14021 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10781) );
  AOI22_X1 U14022 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10780) );
  AOI22_X1 U14023 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10779) );
  NAND4_X1 U14024 ( .A1(n10782), .A2(n10781), .A3(n10780), .A4(n10779), .ZN(
        n10783) );
  AOI22_X1 U14025 ( .A1(n10966), .A2(n10856), .B1(n10956), .B2(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10787) );
  INV_X1 U14026 ( .A(n10787), .ZN(n10785) );
  NAND2_X1 U14027 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  NAND2_X1 U14028 ( .A1(n10840), .A2(n10789), .ZN(n11017) );
  INV_X1 U14029 ( .A(n14078), .ZN(n10825) );
  NAND2_X1 U14030 ( .A1(n10820), .A2(n10815), .ZN(n10814) );
  NAND2_X1 U14031 ( .A1(n10814), .A2(n10810), .ZN(n10804) );
  AND2_X1 U14032 ( .A1(n10802), .A2(n10796), .ZN(n10791) );
  NAND2_X1 U14033 ( .A1(n10804), .A2(n10791), .ZN(n10858) );
  XNOR2_X1 U14034 ( .A(n10858), .B(n10856), .ZN(n10792) );
  NAND2_X1 U14035 ( .A1(n10792), .A2(n21499), .ZN(n10793) );
  OAI21_X2 U14036 ( .B1(n11017), .B2(n10825), .A(n10793), .ZN(n10838) );
  INV_X1 U14037 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13037) );
  XNOR2_X1 U14038 ( .A(n10838), .B(n13037), .ZN(n14469) );
  NAND2_X1 U14039 ( .A1(n11015), .A2(n14078), .ZN(n10800) );
  NAND2_X1 U14040 ( .A1(n10804), .A2(n10802), .ZN(n10797) );
  XNOR2_X1 U14041 ( .A(n10797), .B(n10796), .ZN(n10798) );
  NAND2_X1 U14042 ( .A1(n10798), .A2(n21499), .ZN(n10799) );
  INV_X1 U14043 ( .A(n10802), .ZN(n10803) );
  XNOR2_X1 U14044 ( .A(n10804), .B(n10803), .ZN(n10805) );
  NAND2_X1 U14045 ( .A1(n10805), .A2(n21499), .ZN(n10806) );
  NAND2_X1 U14046 ( .A1(n10807), .A2(n10808), .ZN(n10809) );
  XNOR2_X1 U14047 ( .A(n10814), .B(n10810), .ZN(n10812) );
  AND2_X1 U14048 ( .A1(n13707), .A2(n10811), .ZN(n10822) );
  AOI21_X1 U14049 ( .B1(n10812), .B2(n21499), .A(n10822), .ZN(n10813) );
  OAI21_X1 U14050 ( .B1(n10820), .B2(n10815), .A(n10814), .ZN(n10818) );
  OR2_X1 U14051 ( .A1(n10978), .A2(n14140), .ZN(n10817) );
  AND2_X1 U14052 ( .A1(n10969), .A2(n20838), .ZN(n10816) );
  OAI211_X1 U14053 ( .C1(n10818), .C2(n14137), .A(n10817), .B(n10816), .ZN(
        n14437) );
  INV_X1 U14054 ( .A(n10820), .ZN(n10821) );
  NAND2_X1 U14055 ( .A1(n21499), .A2(n10821), .ZN(n14076) );
  INV_X1 U14056 ( .A(n10822), .ZN(n14075) );
  NAND2_X1 U14057 ( .A1(n14076), .A2(n14075), .ZN(n10824) );
  OR2_X1 U14058 ( .A1(n10824), .A2(n10984), .ZN(n10829) );
  OR2_X1 U14059 ( .A1(n10823), .A2(n10824), .ZN(n10828) );
  INV_X1 U14060 ( .A(n10824), .ZN(n10826) );
  AOI21_X1 U14061 ( .B1(n10826), .B2(n10825), .A(n15426), .ZN(n10827) );
  OAI211_X1 U14062 ( .C1(n10819), .C2(n10829), .A(n10828), .B(n10827), .ZN(
        n14079) );
  INV_X1 U14063 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14473) );
  NOR2_X1 U14064 ( .A1(n14079), .A2(n14473), .ZN(n10830) );
  NAND2_X1 U14065 ( .A1(n14079), .A2(n14473), .ZN(n10831) );
  NAND2_X1 U14066 ( .A1(n10832), .A2(n10831), .ZN(n10833) );
  INV_X1 U14067 ( .A(n10833), .ZN(n10834) );
  NAND2_X1 U14068 ( .A1(n10834), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10835) );
  AOI21_X1 U14069 ( .B1(n14490), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10837) );
  NAND3_X1 U14070 ( .A1(n14490), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U14071 ( .A1(n10838), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10839) );
  INV_X1 U14072 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11522) );
  NAND2_X1 U14073 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U14074 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10841) );
  OAI211_X1 U14075 ( .C1(n11555), .C2(n11522), .A(n10842), .B(n10841), .ZN(
        n10843) );
  INV_X1 U14076 ( .A(n10843), .ZN(n10847) );
  AOI22_X1 U14077 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U14078 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10845) );
  NAND2_X1 U14079 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10844) );
  NAND4_X1 U14080 ( .A1(n10847), .A2(n10846), .A3(n10845), .A4(n10844), .ZN(
        n10853) );
  AOI22_X1 U14081 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10851) );
  AOI22_X1 U14082 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U14083 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10849) );
  AOI22_X1 U14084 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10848) );
  NAND4_X1 U14085 ( .A1(n10851), .A2(n10850), .A3(n10849), .A4(n10848), .ZN(
        n10852) );
  AOI22_X1 U14086 ( .A1(n10966), .A2(n10869), .B1(n10956), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10855) );
  INV_X1 U14087 ( .A(n10856), .ZN(n10857) );
  NOR2_X1 U14088 ( .A1(n10858), .A2(n10857), .ZN(n10870) );
  INV_X1 U14089 ( .A(n10870), .ZN(n10859) );
  XNOR2_X1 U14090 ( .A(n10859), .B(n10869), .ZN(n10860) );
  NAND2_X1 U14091 ( .A1(n10860), .A2(n21499), .ZN(n10861) );
  INV_X1 U14092 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17237) );
  NAND2_X1 U14093 ( .A1(n17238), .A2(n17237), .ZN(n10862) );
  NAND2_X1 U14094 ( .A1(n10863), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10864) );
  NAND2_X1 U14095 ( .A1(n10966), .A2(n10875), .ZN(n10866) );
  NAND2_X1 U14096 ( .A1(n10956), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10865) );
  NAND2_X1 U14097 ( .A1(n10866), .A2(n10865), .ZN(n10867) );
  NAND2_X1 U14098 ( .A1(n10870), .A2(n10869), .ZN(n10878) );
  XNOR2_X1 U14099 ( .A(n10878), .B(n10875), .ZN(n10871) );
  AND2_X1 U14100 ( .A1(n10871), .A2(n21499), .ZN(n10872) );
  INV_X1 U14101 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17251) );
  NAND2_X1 U14102 ( .A1(n10873), .A2(n17251), .ZN(n17232) );
  INV_X1 U14103 ( .A(n10873), .ZN(n10874) );
  NAND2_X1 U14104 ( .A1(n10874), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17231) );
  AND2_X1 U14105 ( .A1(n14078), .A2(n10875), .ZN(n10876) );
  OR3_X1 U14106 ( .A1(n10878), .A2(n10877), .A3(n14137), .ZN(n10887) );
  NAND2_X1 U14107 ( .A1(n10886), .A2(n10887), .ZN(n15357) );
  AND2_X1 U14108 ( .A1(n15357), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10891) );
  INV_X1 U14109 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10879) );
  NAND2_X1 U14110 ( .A1(n10881), .A2(n10879), .ZN(n10880) );
  INV_X1 U14111 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15531) );
  NAND2_X1 U14112 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U14113 ( .A1(n15342), .A2(n10882), .ZN(n15313) );
  INV_X1 U14114 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15475) );
  NAND2_X1 U14115 ( .A1(n10886), .A2(n15475), .ZN(n10883) );
  NAND2_X1 U14116 ( .A1(n10885), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10884) );
  NAND2_X1 U14117 ( .A1(n10885), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15298) );
  INV_X1 U14118 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15492) );
  NAND2_X1 U14119 ( .A1(n10886), .A2(n15492), .ZN(n15297) );
  INV_X1 U14120 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11592) );
  NAND2_X1 U14121 ( .A1(n10887), .A2(n11592), .ZN(n10888) );
  NAND3_X1 U14122 ( .A1(n10888), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10889) );
  NAND2_X1 U14123 ( .A1(n10886), .A2(n10889), .ZN(n10890) );
  INV_X1 U14124 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15564) );
  INV_X1 U14125 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15548) );
  NAND2_X1 U14126 ( .A1(n15564), .A2(n15548), .ZN(n10893) );
  OAI21_X1 U14127 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n10901), .ZN(n10894) );
  NAND2_X1 U14128 ( .A1(n10901), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11594) );
  XNOR2_X1 U14129 ( .A(n15342), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15280) );
  NAND2_X1 U14130 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15433) );
  INV_X1 U14131 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10896) );
  OR2_X1 U14132 ( .A1(n15433), .A2(n10896), .ZN(n10897) );
  INV_X1 U14133 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13015) );
  OR2_X1 U14134 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10898) );
  INV_X1 U14135 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15416) );
  INV_X1 U14136 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15221) );
  INV_X1 U14137 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13621) );
  OAI21_X1 U14138 ( .B1(n12898), .B2(n10431), .A(n10904), .ZN(n10907) );
  NAND2_X1 U14139 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15218) );
  NOR2_X1 U14140 ( .A1(n15218), .A2(n15221), .ZN(n13622) );
  NAND2_X1 U14141 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13062) );
  INV_X1 U14142 ( .A(n13739), .ZN(n10906) );
  NAND2_X1 U14143 ( .A1(n10907), .A2(n10906), .ZN(n10912) );
  INV_X1 U14144 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13054) );
  NAND2_X1 U14145 ( .A1(n15353), .A2(n13054), .ZN(n13737) );
  NAND2_X1 U14146 ( .A1(n13738), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10908) );
  OAI211_X1 U14147 ( .C1(n12898), .C2(n13737), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n10908), .ZN(n10911) );
  INV_X1 U14148 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10909) );
  NOR2_X1 U14149 ( .A1(n10909), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15367) );
  NAND3_X1 U14150 ( .A1(n13739), .A2(n13738), .A3(n15367), .ZN(n10910) );
  NAND3_X1 U14151 ( .A1(n10912), .A2(n10911), .A3(n10910), .ZN(n15366) );
  NAND2_X1 U14152 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21264), .ZN(
        n10921) );
  OAI21_X1 U14153 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21264), .A(
        n10921), .ZN(n10915) );
  INV_X1 U14154 ( .A(n10915), .ZN(n10913) );
  NAND2_X1 U14155 ( .A1(n10966), .A2(n10913), .ZN(n10914) );
  NAND2_X1 U14156 ( .A1(n10914), .A2(n10953), .ZN(n10919) );
  NAND2_X1 U14157 ( .A1(n10916), .A2(n14511), .ZN(n10917) );
  NAND2_X1 U14158 ( .A1(n10917), .A2(n14140), .ZN(n10938) );
  OAI211_X1 U14159 ( .C1(n10602), .C2(n13707), .A(n10913), .B(n10938), .ZN(
        n10918) );
  NAND2_X1 U14160 ( .A1(n21216), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10931) );
  NAND2_X1 U14161 ( .A1(n15596), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10920) );
  NAND2_X1 U14162 ( .A1(n10931), .A2(n10920), .ZN(n10922) );
  NAND2_X1 U14163 ( .A1(n10922), .A2(n10921), .ZN(n10923) );
  AND2_X1 U14164 ( .A1(n10932), .A2(n10923), .ZN(n12908) );
  NAND2_X1 U14165 ( .A1(n10966), .A2(n20819), .ZN(n10924) );
  NAND2_X1 U14166 ( .A1(n10916), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10925) );
  OAI211_X1 U14167 ( .C1(n12908), .C2(n10936), .A(n10924), .B(n10925), .ZN(
        n10927) );
  NAND2_X1 U14168 ( .A1(n10925), .A2(n20819), .ZN(n10926) );
  NOR2_X1 U14169 ( .A1(n10966), .A2(n10926), .ZN(n10957) );
  OAI22_X1 U14170 ( .A1(n10928), .A2(n10927), .B1(n10957), .B2(n12908), .ZN(
        n10930) );
  NAND2_X1 U14171 ( .A1(n10928), .A2(n10927), .ZN(n10929) );
  NAND2_X1 U14172 ( .A1(n10930), .A2(n10929), .ZN(n10942) );
  NAND2_X1 U14173 ( .A1(n10934), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10935) );
  NAND2_X1 U14174 ( .A1(n10946), .A2(n10935), .ZN(n10943) );
  XNOR2_X1 U14175 ( .A(n10945), .B(n10943), .ZN(n12909) );
  NAND2_X1 U14176 ( .A1(n10966), .A2(n12909), .ZN(n10937) );
  OAI211_X1 U14177 ( .C1(n12909), .C2(n10936), .A(n10937), .B(n10938), .ZN(
        n10941) );
  INV_X1 U14178 ( .A(n10937), .ZN(n10940) );
  INV_X1 U14179 ( .A(n10938), .ZN(n10939) );
  AOI22_X1 U14180 ( .A1(n10942), .A2(n10941), .B1(n10940), .B2(n10939), .ZN(
        n10961) );
  INV_X1 U14181 ( .A(n10943), .ZN(n10944) );
  NAND2_X1 U14182 ( .A1(n10945), .A2(n10944), .ZN(n10947) );
  NAND3_X1 U14183 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10963), .A3(
        n17275), .ZN(n12911) );
  XNOR2_X1 U14184 ( .A(n10952), .B(n10951), .ZN(n12907) );
  AOI21_X1 U14185 ( .B1(n12911), .B2(n12907), .A(n10956), .ZN(n10960) );
  INV_X1 U14186 ( .A(n12907), .ZN(n10954) );
  AOI22_X1 U14187 ( .A1(n10964), .A2(n10954), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10276), .ZN(n10959) );
  INV_X1 U14188 ( .A(n12911), .ZN(n10955) );
  NAND3_X1 U14189 ( .A1(n10957), .A2(n10956), .A3(n10955), .ZN(n10958) );
  NOR2_X1 U14190 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20818), .ZN(
        n10962) );
  NAND2_X1 U14191 ( .A1(n12910), .A2(n10964), .ZN(n10965) );
  NAND2_X1 U14192 ( .A1(n14576), .A2(n13707), .ZN(n10968) );
  NAND2_X1 U14193 ( .A1(n9635), .A2(n10970), .ZN(n12922) );
  NAND2_X1 U14194 ( .A1(n15366), .A2(n20780), .ZN(n11590) );
  INV_X1 U14195 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n10972) );
  XNOR2_X1 U14196 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15009) );
  AOI21_X1 U14197 ( .B1(n11431), .B2(n15009), .A(n11574), .ZN(n10971) );
  OAI21_X1 U14198 ( .B1(n11537), .B2(n10972), .A(n10971), .ZN(n10973) );
  AOI21_X1 U14199 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n11002), .A(
        n10973), .ZN(n10974) );
  NAND2_X1 U14200 ( .A1(n11574), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10994) );
  INV_X1 U14201 ( .A(n14251), .ZN(n10993) );
  NAND2_X1 U14202 ( .A1(n10977), .A2(n10978), .ZN(n10979) );
  NAND2_X1 U14203 ( .A1(n14417), .A2(n11026), .ZN(n10983) );
  INV_X1 U14204 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n10980) );
  INV_X1 U14205 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15020) );
  OAI22_X1 U14206 ( .A1(n11537), .A2(n10980), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15020), .ZN(n10981) );
  AOI21_X1 U14207 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11002), .A(
        n10981), .ZN(n10982) );
  NAND2_X1 U14208 ( .A1(n10983), .A2(n10982), .ZN(n14072) );
  NAND2_X1 U14209 ( .A1(n20889), .A2(n10609), .ZN(n10985) );
  NAND2_X1 U14210 ( .A1(n10985), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14025) );
  INV_X1 U14211 ( .A(n11002), .ZN(n11008) );
  NAND2_X1 U14212 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10988) );
  NAND2_X1 U14213 ( .A1(n11575), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n10987) );
  OAI211_X1 U14214 ( .C1(n11008), .C2(n14583), .A(n10988), .B(n10987), .ZN(
        n10989) );
  AOI21_X1 U14215 ( .B1(n10986), .B2(n11026), .A(n10989), .ZN(n10990) );
  OR2_X1 U14216 ( .A1(n14025), .A2(n10990), .ZN(n14026) );
  INV_X1 U14217 ( .A(n10990), .ZN(n14027) );
  OR2_X1 U14218 ( .A1(n14027), .A2(n11573), .ZN(n10991) );
  NAND2_X1 U14219 ( .A1(n14026), .A2(n10991), .ZN(n14071) );
  NAND2_X1 U14220 ( .A1(n14072), .A2(n14071), .ZN(n14250) );
  NAND2_X1 U14221 ( .A1(n10993), .A2(n10992), .ZN(n14253) );
  NAND2_X1 U14222 ( .A1(n14501), .A2(n11026), .ZN(n11004) );
  INV_X1 U14223 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11000) );
  NAND2_X1 U14224 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10996) );
  INV_X1 U14225 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U14226 ( .A1(n10997), .A2(n10996), .ZN(n10998) );
  NAND2_X1 U14227 ( .A1(n9727), .A2(n10998), .ZN(n20707) );
  AOI22_X1 U14228 ( .A1(n20707), .A2(n11431), .B1(n11574), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10999) );
  OAI21_X1 U14229 ( .B1(n11537), .B2(n11000), .A(n10999), .ZN(n11001) );
  AOI21_X1 U14230 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11002), .A(
        n11001), .ZN(n11003) );
  NAND2_X1 U14231 ( .A1(n11004), .A2(n11003), .ZN(n14449) );
  NAND2_X1 U14232 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U14233 ( .A1(n11575), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11006) );
  OAI211_X1 U14234 ( .C1(n11008), .C2(n17275), .A(n11007), .B(n11006), .ZN(
        n11009) );
  NAND2_X1 U14235 ( .A1(n11009), .A2(n11573), .ZN(n11013) );
  INV_X1 U14236 ( .A(n11018), .ZN(n11020) );
  INV_X1 U14237 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11010) );
  NAND2_X1 U14238 ( .A1(n9727), .A2(n11010), .ZN(n11011) );
  NAND2_X1 U14239 ( .A1(n11020), .A2(n11011), .ZN(n20783) );
  NAND2_X1 U14240 ( .A1(n20783), .A2(n11431), .ZN(n11012) );
  NAND2_X1 U14241 ( .A1(n11013), .A2(n11012), .ZN(n11014) );
  AOI21_X1 U14242 ( .B1(n11015), .B2(n11026), .A(n11014), .ZN(n14459) );
  INV_X1 U14243 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n11024) );
  INV_X1 U14244 ( .A(n11037), .ZN(n11022) );
  INV_X1 U14245 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11019) );
  NAND2_X1 U14246 ( .A1(n11020), .A2(n11019), .ZN(n11021) );
  NAND2_X1 U14247 ( .A1(n11022), .A2(n11021), .ZN(n17250) );
  AOI22_X1 U14248 ( .A1(n17250), .A2(n11431), .B1(n11574), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11023) );
  OAI21_X1 U14249 ( .B1(n11537), .B2(n11024), .A(n11023), .ZN(n11025) );
  NAND2_X1 U14250 ( .A1(n11028), .A2(n11026), .ZN(n11034) );
  INV_X1 U14251 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11031) );
  OAI21_X1 U14252 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11029), .A(
        n11074), .ZN(n20666) );
  AOI22_X1 U14253 ( .A1(n11431), .A2(n20666), .B1(n11574), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11030) );
  OAI21_X1 U14254 ( .B1(n11537), .B2(n11031), .A(n11030), .ZN(n11032) );
  INV_X1 U14255 ( .A(n11032), .ZN(n11033) );
  NAND2_X1 U14256 ( .A1(n11034), .A2(n11033), .ZN(n14957) );
  NAND2_X1 U14257 ( .A1(n11035), .A2(n11026), .ZN(n11042) );
  INV_X1 U14258 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11039) );
  OAI21_X1 U14259 ( .B1(n11037), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n11036), .ZN(n20683) );
  AOI22_X1 U14260 ( .A1(n20683), .A2(n11431), .B1(n11574), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11038) );
  OAI21_X1 U14261 ( .B1(n11537), .B2(n11039), .A(n11038), .ZN(n11040) );
  INV_X1 U14262 ( .A(n11040), .ZN(n11041) );
  INV_X1 U14263 ( .A(n11101), .ZN(n11081) );
  INV_X1 U14264 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14966) );
  XNOR2_X1 U14265 ( .A(n11081), .B(n14966), .ZN(n15349) );
  NAND2_X1 U14266 ( .A1(n15349), .A2(n11431), .ZN(n11060) );
  INV_X1 U14267 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n15190) );
  OAI22_X1 U14268 ( .A1(n11537), .A2(n15190), .B1(n14966), .B2(n14429), .ZN(
        n11058) );
  CLKBUF_X1 U14269 ( .A(n10544), .Z(n11550) );
  NAND2_X1 U14270 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14271 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14272 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11043) );
  AND3_X1 U14273 ( .A1(n11045), .A2(n11044), .A3(n11043), .ZN(n11049) );
  AOI22_X1 U14274 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U14275 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11047) );
  NAND2_X1 U14276 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11046) );
  NAND4_X1 U14277 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n11055) );
  AOI22_X1 U14278 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10664), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U14279 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11052) );
  AOI22_X1 U14280 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11051) );
  AOI22_X1 U14281 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11050) );
  NAND4_X1 U14282 ( .A1(n11053), .A2(n11052), .A3(n11051), .A4(n11050), .ZN(
        n11054) );
  NOR2_X1 U14283 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NOR2_X1 U14284 ( .A1(n11196), .A2(n11056), .ZN(n11057) );
  NOR2_X1 U14285 ( .A1(n11058), .A2(n11057), .ZN(n11059) );
  NAND2_X1 U14286 ( .A1(n11060), .A2(n11059), .ZN(n14959) );
  AOI22_X1 U14287 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11064) );
  AOI22_X1 U14288 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n10664), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11063) );
  AOI22_X1 U14289 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n11528), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U14290 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11061) );
  NAND4_X1 U14291 ( .A1(n11064), .A2(n11063), .A3(n11062), .A4(n11061), .ZN(
        n11073) );
  NAND2_X1 U14292 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11066) );
  NAND2_X1 U14293 ( .A1(n11551), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11065) );
  OAI211_X1 U14294 ( .C1(n11555), .C2(n14519), .A(n11066), .B(n11065), .ZN(
        n11067) );
  INV_X1 U14295 ( .A(n11067), .ZN(n11071) );
  AOI22_X1 U14296 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U14297 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U14298 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11068) );
  NAND4_X1 U14299 ( .A1(n11071), .A2(n11070), .A3(n11069), .A4(n11068), .ZN(
        n11072) );
  NOR2_X1 U14300 ( .A1(n11073), .A2(n11072), .ZN(n11078) );
  NAND2_X1 U14301 ( .A1(n11575), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11077) );
  INV_X1 U14302 ( .A(n11074), .ZN(n11075) );
  XNOR2_X1 U14303 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11075), .ZN(
        n15361) );
  AOI22_X1 U14304 ( .A1(n11431), .A2(n15361), .B1(n11574), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11076) );
  OAI211_X1 U14305 ( .C1(n11078), .C2(n11196), .A(n11077), .B(n11076), .ZN(
        n14974) );
  NAND2_X1 U14306 ( .A1(n11079), .A2(n21565), .ZN(n11080) );
  NAND2_X1 U14307 ( .A1(n11081), .A2(n11080), .ZN(n20655) );
  NAND2_X1 U14308 ( .A1(n20655), .A2(n11431), .ZN(n11099) );
  NAND2_X1 U14309 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11084) );
  NAND2_X1 U14310 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11083) );
  NAND2_X1 U14311 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11082) );
  AND3_X1 U14312 ( .A1(n11084), .A2(n11083), .A3(n11082), .ZN(n11088) );
  AOI22_X1 U14313 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14314 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11086) );
  NAND2_X1 U14315 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11085) );
  NAND4_X1 U14316 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11094) );
  AOI22_X1 U14317 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14318 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10664), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14319 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14320 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11089) );
  NAND4_X1 U14321 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n11093) );
  NOR2_X1 U14322 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  OAI22_X1 U14323 ( .A1(n11196), .A2(n11095), .B1(n21565), .B2(n14429), .ZN(
        n11097) );
  INV_X1 U14324 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n15192) );
  NOR2_X1 U14325 ( .A1(n11537), .A2(n15192), .ZN(n11096) );
  NOR2_X1 U14326 ( .A1(n11097), .A2(n11096), .ZN(n11098) );
  NAND2_X1 U14327 ( .A1(n11099), .A2(n11098), .ZN(n15081) );
  NAND2_X1 U14328 ( .A1(n11101), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11136) );
  INV_X1 U14329 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11103) );
  XNOR2_X1 U14330 ( .A(n11193), .B(n11103), .ZN(n17207) );
  AOI22_X1 U14331 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U14332 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14333 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14334 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11104) );
  NAND4_X1 U14335 ( .A1(n11107), .A2(n11106), .A3(n11105), .A4(n11104), .ZN(
        n11116) );
  INV_X1 U14336 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20850) );
  NAND2_X1 U14337 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14338 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11108) );
  OAI211_X1 U14339 ( .C1(n11555), .C2(n20850), .A(n11109), .B(n11108), .ZN(
        n11110) );
  INV_X1 U14340 ( .A(n11110), .ZN(n11114) );
  AOI22_X1 U14341 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14342 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11112) );
  NAND2_X1 U14343 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11111) );
  NAND4_X1 U14344 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n11115) );
  OAI21_X1 U14345 ( .B1(n11116), .B2(n11115), .A(n11026), .ZN(n11119) );
  NAND2_X1 U14346 ( .A1(n11575), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11118) );
  NAND2_X1 U14347 ( .A1(n11574), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11117) );
  NAND3_X1 U14348 ( .A1(n11119), .A2(n11118), .A3(n11117), .ZN(n11120) );
  AOI21_X1 U14349 ( .B1(n17207), .B2(n11431), .A(n11120), .ZN(n15060) );
  AOI22_X1 U14350 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11124) );
  AOI22_X1 U14351 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14352 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14353 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11121) );
  NAND4_X1 U14354 ( .A1(n11124), .A2(n11123), .A3(n11122), .A4(n11121), .ZN(
        n11134) );
  INV_X1 U14355 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14356 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11126) );
  NAND2_X1 U14357 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11125) );
  OAI211_X1 U14358 ( .C1(n11555), .C2(n11127), .A(n11126), .B(n11125), .ZN(
        n11128) );
  INV_X1 U14359 ( .A(n11128), .ZN(n11132) );
  AOI22_X1 U14360 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14361 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11130) );
  NAND2_X1 U14362 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11129) );
  NAND4_X1 U14363 ( .A1(n11132), .A2(n11131), .A3(n11130), .A4(n11129), .ZN(
        n11133) );
  NOR2_X1 U14364 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  NOR2_X1 U14365 ( .A1(n11196), .A2(n11135), .ZN(n15071) );
  NAND2_X1 U14366 ( .A1(n11136), .A2(n11138), .ZN(n11137) );
  NAND2_X1 U14367 ( .A1(n11161), .A2(n11137), .ZN(n17223) );
  NAND2_X1 U14368 ( .A1(n17223), .A2(n11431), .ZN(n11141) );
  INV_X1 U14369 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n15187) );
  OAI22_X1 U14370 ( .A1(n11537), .A2(n15187), .B1(n11138), .B2(n14429), .ZN(
        n11139) );
  INV_X1 U14371 ( .A(n11139), .ZN(n11140) );
  NAND2_X1 U14372 ( .A1(n11141), .A2(n11140), .ZN(n14923) );
  XNOR2_X1 U14373 ( .A(n11142), .B(n14932), .ZN(n15320) );
  NAND2_X1 U14374 ( .A1(n15320), .A2(n11431), .ZN(n11160) );
  INV_X1 U14375 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n15184) );
  OAI22_X1 U14376 ( .A1(n11537), .A2(n15184), .B1(n14429), .B2(n14932), .ZN(
        n11158) );
  NAND2_X1 U14377 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U14378 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14379 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11143) );
  AND3_X1 U14380 ( .A1(n11145), .A2(n11144), .A3(n11143), .ZN(n11149) );
  AOI22_X1 U14381 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11148) );
  AOI22_X1 U14382 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14383 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11146) );
  NAND4_X1 U14384 ( .A1(n11149), .A2(n11148), .A3(n11147), .A4(n11146), .ZN(
        n11155) );
  AOI22_X1 U14385 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11153) );
  AOI22_X1 U14386 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10664), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14387 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U14388 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11150) );
  NAND4_X1 U14389 ( .A1(n11153), .A2(n11152), .A3(n11151), .A4(n11150), .ZN(
        n11154) );
  NOR2_X1 U14390 ( .A1(n11155), .A2(n11154), .ZN(n11156) );
  NOR2_X1 U14391 ( .A1(n11196), .A2(n11156), .ZN(n11157) );
  NOR2_X1 U14392 ( .A1(n11158), .A2(n11157), .ZN(n11159) );
  NAND2_X1 U14393 ( .A1(n11160), .A2(n11159), .ZN(n14926) );
  XNOR2_X1 U14394 ( .A(n11161), .B(n9902), .ZN(n15328) );
  NAND2_X1 U14395 ( .A1(n15328), .A2(n11431), .ZN(n11179) );
  INV_X1 U14396 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n15186) );
  OAI22_X1 U14397 ( .A1(n11537), .A2(n15186), .B1(n9902), .B2(n14429), .ZN(
        n11177) );
  NAND2_X1 U14398 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11164) );
  NAND2_X1 U14399 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11163) );
  NAND2_X1 U14400 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11162) );
  AND3_X1 U14401 ( .A1(n11164), .A2(n11163), .A3(n11162), .ZN(n11168) );
  AOI22_X1 U14402 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U14403 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U14404 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11165) );
  NAND4_X1 U14405 ( .A1(n11168), .A2(n11167), .A3(n11166), .A4(n11165), .ZN(
        n11174) );
  AOI22_X1 U14406 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11172) );
  AOI22_X1 U14407 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14408 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14409 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11169) );
  NAND4_X1 U14410 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11173) );
  NOR2_X1 U14411 ( .A1(n11174), .A2(n11173), .ZN(n11175) );
  NOR2_X1 U14412 ( .A1(n11196), .A2(n11175), .ZN(n11176) );
  NOR2_X1 U14413 ( .A1(n11177), .A2(n11176), .ZN(n11178) );
  NAND2_X1 U14414 ( .A1(n11179), .A2(n11178), .ZN(n14943) );
  OAI211_X1 U14415 ( .C1(n15071), .C2(n14923), .A(n14926), .B(n14943), .ZN(
        n11180) );
  NOR2_X1 U14416 ( .A1(n15060), .A2(n11180), .ZN(n11198) );
  AOI22_X1 U14417 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11182) );
  NAND2_X1 U14418 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11181) );
  AND2_X1 U14419 ( .A1(n11182), .A2(n11181), .ZN(n11186) );
  AOI22_X1 U14420 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U14421 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11184) );
  NAND2_X1 U14422 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11183) );
  NAND4_X1 U14423 ( .A1(n11186), .A2(n11185), .A3(n11184), .A4(n11183), .ZN(
        n11192) );
  AOI22_X1 U14424 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11190) );
  AOI22_X1 U14425 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U14426 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U14427 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11187) );
  NAND4_X1 U14428 ( .A1(n11190), .A2(n11189), .A3(n11188), .A4(n11187), .ZN(
        n11191) );
  NOR2_X1 U14429 ( .A1(n11192), .A2(n11191), .ZN(n11197) );
  XNOR2_X1 U14430 ( .A(n11199), .B(n17191), .ZN(n17197) );
  NAND2_X1 U14431 ( .A1(n17197), .A2(n11431), .ZN(n11195) );
  AOI22_X1 U14432 ( .A1(n11575), .A2(P1_EAX_REG_15__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n11574), .ZN(n11194) );
  OAI211_X1 U14433 ( .C1(n11197), .C2(n11196), .A(n11195), .B(n11194), .ZN(
        n15055) );
  NAND2_X1 U14434 ( .A1(n11200), .A2(n14914), .ZN(n11201) );
  NAND2_X1 U14435 ( .A1(n11238), .A2(n11201), .ZN(n15292) );
  AOI22_X1 U14436 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14437 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n10632), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U14438 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n11528), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14439 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11202) );
  NAND4_X1 U14440 ( .A1(n11205), .A2(n11204), .A3(n11203), .A4(n11202), .ZN(
        n11215) );
  INV_X1 U14441 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14442 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14443 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11206) );
  OAI211_X1 U14444 ( .C1(n11555), .C2(n11208), .A(n11207), .B(n11206), .ZN(
        n11209) );
  INV_X1 U14445 ( .A(n11209), .ZN(n11213) );
  AOI22_X1 U14446 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n9577), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14447 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11211) );
  NAND2_X1 U14448 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11210) );
  NAND4_X1 U14449 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11214) );
  NOR2_X1 U14450 ( .A1(n11215), .A2(n11214), .ZN(n11216) );
  NOR2_X1 U14451 ( .A1(n11570), .A2(n11216), .ZN(n11219) );
  INV_X1 U14452 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n15175) );
  NAND2_X1 U14453 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11217) );
  OAI211_X1 U14454 ( .C1(n11537), .C2(n15175), .A(n11573), .B(n11217), .ZN(
        n11218) );
  OAI22_X1 U14455 ( .A1(n15292), .A2(n11573), .B1(n11219), .B2(n11218), .ZN(
        n14912) );
  XNOR2_X1 U14456 ( .A(n11238), .B(n14901), .ZN(n14909) );
  NAND2_X1 U14457 ( .A1(n14909), .A2(n11431), .ZN(n11237) );
  INV_X1 U14458 ( .A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U14459 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11221) );
  NAND2_X1 U14460 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11220) );
  OAI211_X1 U14461 ( .C1(n11555), .C2(n11222), .A(n11221), .B(n11220), .ZN(
        n11223) );
  INV_X1 U14462 ( .A(n11223), .ZN(n11227) );
  AOI22_X1 U14463 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14464 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11225) );
  NAND2_X1 U14465 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11224) );
  NAND4_X1 U14466 ( .A1(n11227), .A2(n11226), .A3(n11225), .A4(n11224), .ZN(
        n11233) );
  AOI22_X1 U14467 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14468 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14469 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14470 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14471 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11232) );
  OR2_X1 U14472 ( .A1(n11233), .A2(n11232), .ZN(n11235) );
  INV_X1 U14473 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15169) );
  OAI22_X1 U14474 ( .A1(n11537), .A2(n15169), .B1(n14901), .B2(n14429), .ZN(
        n11234) );
  AOI21_X1 U14475 ( .B1(n11539), .B2(n11235), .A(n11234), .ZN(n11236) );
  NAND2_X1 U14476 ( .A1(n11237), .A2(n11236), .ZN(n11602) );
  INV_X1 U14477 ( .A(n11600), .ZN(n11262) );
  INV_X1 U14478 ( .A(n11239), .ZN(n11241) );
  INV_X1 U14479 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U14480 ( .A1(n11241), .A2(n11240), .ZN(n11242) );
  NAND2_X1 U14481 ( .A1(n11283), .A2(n11242), .ZN(n15278) );
  OR2_X1 U14482 ( .A1(n15278), .A2(n11573), .ZN(n11261) );
  AOI22_X1 U14483 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14484 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14485 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14486 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11243) );
  NAND4_X1 U14487 ( .A1(n11246), .A2(n11245), .A3(n11244), .A4(n11243), .ZN(
        n11256) );
  INV_X1 U14488 ( .A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11249) );
  NAND2_X1 U14489 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n11248) );
  NAND2_X1 U14490 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11247) );
  OAI211_X1 U14491 ( .C1(n11555), .C2(n11249), .A(n11248), .B(n11247), .ZN(
        n11250) );
  INV_X1 U14492 ( .A(n11250), .ZN(n11254) );
  AOI22_X1 U14493 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10527), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14494 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11252) );
  NAND2_X1 U14495 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11251) );
  NAND4_X1 U14496 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11255) );
  NOR2_X1 U14497 ( .A1(n11256), .A2(n11255), .ZN(n11259) );
  OAI21_X1 U14498 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21497), .A(
        n11005), .ZN(n11258) );
  NAND2_X1 U14499 ( .A1(n11575), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n11257) );
  OAI211_X1 U14500 ( .C1(n11570), .C2(n11259), .A(n11258), .B(n11257), .ZN(
        n11260) );
  XNOR2_X1 U14501 ( .A(n11283), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15273) );
  NAND2_X1 U14502 ( .A1(n15273), .A2(n11431), .ZN(n11282) );
  AOI22_X1 U14503 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14504 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14505 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14506 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14507 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11276) );
  INV_X1 U14508 ( .A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14509 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14510 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11267) );
  OAI211_X1 U14511 ( .C1(n11555), .C2(n11269), .A(n11268), .B(n11267), .ZN(
        n11270) );
  INV_X1 U14512 ( .A(n11270), .ZN(n11274) );
  AOI22_X1 U14513 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11273) );
  AOI22_X1 U14514 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11272) );
  NAND2_X1 U14515 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11271) );
  NAND4_X1 U14516 ( .A1(n11274), .A2(n11273), .A3(n11272), .A4(n11271), .ZN(
        n11275) );
  NOR2_X1 U14517 ( .A1(n11276), .A2(n11275), .ZN(n11280) );
  NAND2_X1 U14518 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14519 ( .A1(n11573), .A2(n11277), .ZN(n11278) );
  AOI21_X1 U14520 ( .B1(n11575), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11278), .ZN(
        n11279) );
  OAI21_X1 U14521 ( .B1(n11570), .B2(n11280), .A(n11279), .ZN(n11281) );
  NAND2_X1 U14522 ( .A1(n11282), .A2(n11281), .ZN(n14863) );
  INV_X1 U14523 ( .A(n11285), .ZN(n11286) );
  NAND2_X1 U14524 ( .A1(n11286), .A2(n9911), .ZN(n11287) );
  NAND2_X1 U14525 ( .A1(n11412), .A2(n11287), .ZN(n15262) );
  AOI22_X1 U14526 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U14527 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11288) );
  AND2_X1 U14528 ( .A1(n11289), .A2(n11288), .ZN(n11293) );
  AOI22_X1 U14529 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14530 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14531 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11290) );
  NAND4_X1 U14532 ( .A1(n11293), .A2(n11292), .A3(n11291), .A4(n11290), .ZN(
        n11299) );
  AOI22_X1 U14533 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11297) );
  AOI22_X1 U14534 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14535 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11528), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14536 ( .A1(n10577), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11294) );
  NAND4_X1 U14537 ( .A1(n11297), .A2(n11296), .A3(n11295), .A4(n11294), .ZN(
        n11298) );
  NOR2_X1 U14538 ( .A1(n11299), .A2(n11298), .ZN(n11303) );
  NAND2_X1 U14539 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11300) );
  NAND2_X1 U14540 ( .A1(n11573), .A2(n11300), .ZN(n11301) );
  AOI21_X1 U14541 ( .B1(n11575), .B2(P1_EAX_REG_20__SCAN_IN), .A(n11301), .ZN(
        n11302) );
  OAI21_X1 U14542 ( .B1(n11570), .B2(n11303), .A(n11302), .ZN(n11304) );
  INV_X1 U14543 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11389) );
  INV_X1 U14544 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n11371) );
  XNOR2_X1 U14545 ( .A(n11434), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15223) );
  INV_X1 U14546 ( .A(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11315) );
  INV_X1 U14547 ( .A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11308) );
  INV_X1 U14548 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11307) );
  OAI22_X1 U14549 ( .A1(n11308), .A2(n11465), .B1(n11352), .B2(n11307), .ZN(
        n11312) );
  INV_X1 U14550 ( .A(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11310) );
  INV_X1 U14551 ( .A(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11309) );
  OAI22_X1 U14552 ( .A1(n11310), .A2(n10742), .B1(n11544), .B2(n11309), .ZN(
        n11311) );
  AOI211_X1 U14553 ( .C1(n11550), .C2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n11312), .B(n11311), .ZN(n11314) );
  AOI22_X1 U14554 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11313) );
  OAI211_X1 U14555 ( .C1(n11555), .C2(n11315), .A(n11314), .B(n11313), .ZN(
        n11322) );
  AOI22_X1 U14556 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n11316), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14557 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n10664), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14558 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n11497), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11318) );
  AOI22_X1 U14559 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11317) );
  NAND4_X1 U14560 ( .A1(n11320), .A2(n11319), .A3(n11318), .A4(n11317), .ZN(
        n11321) );
  NOR2_X1 U14561 ( .A1(n11322), .A2(n11321), .ZN(n11382) );
  INV_X1 U14562 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11554) );
  INV_X1 U14563 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11545) );
  OAI22_X1 U14564 ( .A1(n13921), .A2(n11545), .B1(n11325), .B2(n11324), .ZN(
        n11328) );
  INV_X1 U14565 ( .A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11547) );
  INV_X1 U14566 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11326) );
  OAI22_X1 U14567 ( .A1(n10742), .A2(n11547), .B1(n11465), .B2(n11326), .ZN(
        n11327) );
  AOI211_X1 U14568 ( .C1(n11472), .C2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11328), .B(n11327), .ZN(n11330) );
  AOI22_X1 U14569 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11329) );
  OAI211_X1 U14570 ( .C1(n10461), .C2(n11554), .A(n11330), .B(n11329), .ZN(
        n11336) );
  AOI22_X1 U14571 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14572 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14573 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10664), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14574 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14575 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11335) );
  NOR2_X1 U14576 ( .A1(n11336), .A2(n11335), .ZN(n11381) );
  NOR2_X1 U14577 ( .A1(n11382), .A2(n11381), .ZN(n11376) );
  INV_X1 U14578 ( .A(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11339) );
  NAND2_X1 U14579 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14580 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11337) );
  OAI211_X1 U14581 ( .C1(n11555), .C2(n11339), .A(n11338), .B(n11337), .ZN(
        n11340) );
  INV_X1 U14582 ( .A(n11340), .ZN(n11344) );
  AOI22_X1 U14583 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14584 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14585 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11341) );
  NAND4_X1 U14586 ( .A1(n11344), .A2(n11343), .A3(n11342), .A4(n11341), .ZN(
        n11350) );
  AOI22_X1 U14587 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11348) );
  AOI22_X1 U14588 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14589 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14590 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11345) );
  NAND4_X1 U14591 ( .A1(n11348), .A2(n11347), .A3(n11346), .A4(n11345), .ZN(
        n11349) );
  OR2_X1 U14592 ( .A1(n11350), .A2(n11349), .ZN(n11374) );
  NAND2_X1 U14593 ( .A1(n11376), .A2(n11374), .ZN(n11438) );
  INV_X1 U14594 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11360) );
  INV_X1 U14595 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11353) );
  INV_X1 U14596 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11351) );
  OAI22_X1 U14597 ( .A1(n13921), .A2(n11353), .B1(n11352), .B2(n11351), .ZN(
        n11357) );
  INV_X1 U14598 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11354) );
  OAI22_X1 U14599 ( .A1(n10718), .A2(n11355), .B1(n11468), .B2(n11354), .ZN(
        n11356) );
  AOI211_X1 U14600 ( .C1(n11550), .C2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n11357), .B(n11356), .ZN(n11359) );
  AOI22_X1 U14601 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11358) );
  OAI211_X1 U14602 ( .C1(n11555), .C2(n11360), .A(n11359), .B(n11358), .ZN(
        n11366) );
  AOI22_X1 U14603 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14604 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14605 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11362) );
  AOI22_X1 U14606 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11361) );
  NAND4_X1 U14607 ( .A1(n11364), .A2(n11363), .A3(n11362), .A4(n11361), .ZN(
        n11365) );
  NOR2_X1 U14608 ( .A1(n11366), .A2(n11365), .ZN(n11439) );
  XOR2_X1 U14609 ( .A(n11438), .B(n11439), .Z(n11369) );
  INV_X1 U14610 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n15138) );
  NAND2_X1 U14611 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11367) );
  OAI211_X1 U14612 ( .C1(n11537), .C2(n15138), .A(n11573), .B(n11367), .ZN(
        n11368) );
  AOI21_X1 U14613 ( .B1(n11369), .B2(n11539), .A(n11368), .ZN(n11370) );
  AOI21_X1 U14614 ( .B1(n15223), .B2(n11431), .A(n11370), .ZN(n14786) );
  NAND2_X1 U14615 ( .A1(n11372), .A2(n11371), .ZN(n11373) );
  AND2_X1 U14616 ( .A1(n11434), .A2(n11373), .ZN(n15230) );
  INV_X1 U14617 ( .A(n11374), .ZN(n11375) );
  XNOR2_X1 U14618 ( .A(n11376), .B(n11375), .ZN(n11379) );
  INV_X1 U14619 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n15142) );
  NAND2_X1 U14620 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11377) );
  OAI211_X1 U14621 ( .C1(n11537), .C2(n15142), .A(n11573), .B(n11377), .ZN(
        n11378) );
  AOI21_X1 U14622 ( .B1(n11379), .B2(n11539), .A(n11378), .ZN(n11380) );
  AOI21_X1 U14623 ( .B1(n15230), .B2(n11431), .A(n11380), .ZN(n14804) );
  INV_X1 U14624 ( .A(n14804), .ZN(n11411) );
  XNOR2_X1 U14625 ( .A(n11392), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15238) );
  NAND2_X1 U14626 ( .A1(n15238), .A2(n11431), .ZN(n11388) );
  XOR2_X1 U14627 ( .A(n11382), .B(n11381), .Z(n11383) );
  NAND2_X1 U14628 ( .A1(n11383), .A2(n11539), .ZN(n11386) );
  AOI21_X1 U14629 ( .B1(n9908), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11384) );
  AOI21_X1 U14630 ( .B1(n11575), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11384), .ZN(
        n11385) );
  NAND2_X1 U14631 ( .A1(n11386), .A2(n11385), .ZN(n11387) );
  NAND2_X1 U14632 ( .A1(n11388), .A2(n11387), .ZN(n14813) );
  NAND2_X1 U14633 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  NAND2_X1 U14634 ( .A1(n11392), .A2(n11391), .ZN(n15247) );
  NAND2_X1 U14635 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14636 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11394) );
  NAND2_X1 U14637 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11393) );
  AND3_X1 U14638 ( .A1(n11395), .A2(n11394), .A3(n11393), .ZN(n11399) );
  AOI22_X1 U14639 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11398) );
  AOI22_X1 U14640 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11397) );
  NAND2_X1 U14641 ( .A1(n11472), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11396) );
  NAND4_X1 U14642 ( .A1(n11399), .A2(n11398), .A3(n11397), .A4(n11396), .ZN(
        n11406) );
  AOI22_X1 U14643 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11404) );
  AOI22_X1 U14644 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14645 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14646 ( .A1(n11323), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11401) );
  NAND4_X1 U14647 ( .A1(n11404), .A2(n11403), .A3(n11402), .A4(n11401), .ZN(
        n11405) );
  NOR2_X1 U14648 ( .A1(n11406), .A2(n11405), .ZN(n11407) );
  NOR2_X1 U14649 ( .A1(n11570), .A2(n11407), .ZN(n11410) );
  INV_X1 U14650 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n15150) );
  NAND2_X1 U14651 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11408) );
  OAI211_X1 U14652 ( .C1(n11537), .C2(n15150), .A(n11573), .B(n11408), .ZN(
        n11409) );
  OAI22_X1 U14653 ( .A1(n15247), .A2(n11573), .B1(n11410), .B2(n11409), .ZN(
        n14826) );
  OR2_X1 U14654 ( .A1(n14813), .A2(n14826), .ZN(n14801) );
  NOR2_X1 U14655 ( .A1(n11411), .A2(n14801), .ZN(n14784) );
  AND2_X1 U14656 ( .A1(n14786), .A2(n14784), .ZN(n11432) );
  XNOR2_X1 U14657 ( .A(n11412), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15255) );
  INV_X1 U14658 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11415) );
  NAND2_X1 U14659 ( .A1(n10762), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11414) );
  NAND2_X1 U14660 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11413) );
  OAI211_X1 U14661 ( .C1(n11555), .C2(n11415), .A(n11414), .B(n11413), .ZN(
        n11416) );
  INV_X1 U14662 ( .A(n11416), .ZN(n11420) );
  AOI22_X1 U14663 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14664 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11529), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14665 ( .A1(n11550), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11417) );
  NAND4_X1 U14666 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(
        n11426) );
  AOI22_X1 U14667 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14668 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14669 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14670 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14671 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11425) );
  OR2_X1 U14672 ( .A1(n11426), .A2(n11425), .ZN(n11429) );
  INV_X1 U14673 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n15155) );
  NAND2_X1 U14674 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11427) );
  OAI211_X1 U14675 ( .C1(n11537), .C2(n15155), .A(n11573), .B(n11427), .ZN(
        n11428) );
  AOI21_X1 U14676 ( .B1(n11539), .B2(n11429), .A(n11428), .ZN(n11430) );
  AOI21_X1 U14677 ( .B1(n15255), .B2(n11431), .A(n11430), .ZN(n14838) );
  AND2_X1 U14678 ( .A1(n11432), .A2(n14838), .ZN(n11433) );
  INV_X1 U14679 ( .A(n14770), .ZN(n11461) );
  INV_X1 U14680 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U14681 ( .A1(n11436), .A2(n11435), .ZN(n11437) );
  NAND2_X1 U14682 ( .A1(n11490), .A2(n11437), .ZN(n15214) );
  NOR2_X1 U14683 ( .A1(n11439), .A2(n11438), .ZN(n11463) );
  INV_X1 U14684 ( .A(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11442) );
  NAND2_X1 U14685 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11441) );
  NAND2_X1 U14686 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11440) );
  OAI211_X1 U14687 ( .C1(n11555), .C2(n11442), .A(n11441), .B(n11440), .ZN(
        n11443) );
  INV_X1 U14688 ( .A(n11443), .ZN(n11447) );
  AOI22_X1 U14689 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14690 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11445) );
  NAND2_X1 U14691 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11444) );
  NAND4_X1 U14692 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11453) );
  AOI22_X1 U14693 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11323), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14694 ( .A1(n10622), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14695 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14696 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14697 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11452) );
  OR2_X1 U14698 ( .A1(n11453), .A2(n11452), .ZN(n11462) );
  XNOR2_X1 U14699 ( .A(n11463), .B(n11462), .ZN(n11457) );
  NAND2_X1 U14700 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11454) );
  NAND2_X1 U14701 ( .A1(n11573), .A2(n11454), .ZN(n11455) );
  AOI21_X1 U14702 ( .B1(n11575), .B2(P1_EAX_REG_26__SCAN_IN), .A(n11455), .ZN(
        n11456) );
  OAI21_X1 U14703 ( .B1(n11457), .B2(n11570), .A(n11456), .ZN(n11458) );
  NAND2_X1 U14704 ( .A1(n11459), .A2(n11458), .ZN(n14771) );
  XNOR2_X1 U14705 ( .A(n11490), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14761) );
  NAND2_X1 U14706 ( .A1(n14761), .A2(n11431), .ZN(n11487) );
  NAND2_X1 U14707 ( .A1(n11463), .A2(n11462), .ZN(n11495) );
  INV_X1 U14708 ( .A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11475) );
  INV_X1 U14709 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11466) );
  INV_X1 U14710 ( .A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11464) );
  OAI22_X1 U14711 ( .A1(n10742), .A2(n11466), .B1(n11465), .B2(n11464), .ZN(
        n11471) );
  INV_X1 U14712 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11469) );
  INV_X1 U14713 ( .A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11467) );
  OAI22_X1 U14714 ( .A1(n13921), .A2(n11469), .B1(n11468), .B2(n11467), .ZN(
        n11470) );
  AOI211_X1 U14715 ( .C1(n11472), .C2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11471), .B(n11470), .ZN(n11474) );
  AOI22_X1 U14716 ( .A1(n11400), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11473) );
  OAI211_X1 U14717 ( .C1(n10461), .C2(n11475), .A(n11474), .B(n11473), .ZN(
        n11481) );
  AOI22_X1 U14718 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10622), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11479) );
  AOI22_X1 U14719 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14720 ( .A1(n9577), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11477) );
  AOI22_X1 U14721 ( .A1(n10664), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11476) );
  NAND4_X1 U14722 ( .A1(n11479), .A2(n11478), .A3(n11477), .A4(n11476), .ZN(
        n11480) );
  NOR2_X1 U14723 ( .A1(n11481), .A2(n11480), .ZN(n11496) );
  XOR2_X1 U14724 ( .A(n11495), .B(n11496), .Z(n11482) );
  NAND2_X1 U14725 ( .A1(n11482), .A2(n11539), .ZN(n11485) );
  INV_X1 U14726 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14763) );
  AOI21_X1 U14727 ( .B1(n14763), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11483) );
  AOI21_X1 U14728 ( .B1(n11575), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11483), .ZN(
        n11484) );
  NAND2_X1 U14729 ( .A1(n11485), .A2(n11484), .ZN(n11486) );
  NAND2_X1 U14730 ( .A1(n11487), .A2(n11486), .ZN(n14757) );
  INV_X1 U14731 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U14732 ( .A1(n11493), .A2(n11492), .ZN(n11494) );
  NAND2_X1 U14733 ( .A1(n11542), .A2(n11494), .ZN(n15198) );
  NOR2_X1 U14734 ( .A1(n11496), .A2(n11495), .ZN(n11518) );
  INV_X1 U14735 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U14736 ( .A1(n10651), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14737 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11498) );
  OAI211_X1 U14738 ( .C1(n11555), .C2(n11500), .A(n11499), .B(n11498), .ZN(
        n11501) );
  INV_X1 U14739 ( .A(n11501), .ZN(n11505) );
  AOI22_X1 U14740 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14741 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14742 ( .A1(n10544), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11502) );
  NAND4_X1 U14743 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11511) );
  AOI22_X1 U14744 ( .A1(n10669), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10577), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14745 ( .A1(n10674), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11316), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11508) );
  AOI22_X1 U14746 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14747 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14748 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11510) );
  OR2_X1 U14749 ( .A1(n11511), .A2(n11510), .ZN(n11517) );
  XNOR2_X1 U14750 ( .A(n11518), .B(n11517), .ZN(n11515) );
  NAND2_X1 U14751 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11512) );
  NAND2_X1 U14752 ( .A1(n11573), .A2(n11512), .ZN(n11513) );
  AOI21_X1 U14753 ( .B1(n11575), .B2(P1_EAX_REG_28__SCAN_IN), .A(n11513), .ZN(
        n11514) );
  OAI21_X1 U14754 ( .B1(n11515), .B2(n11570), .A(n11514), .ZN(n11516) );
  OAI21_X1 U14755 ( .B1(n15198), .B2(n11573), .A(n11516), .ZN(n14746) );
  XNOR2_X1 U14756 ( .A(n11542), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14723) );
  NAND2_X1 U14757 ( .A1(n11518), .A2(n11517), .ZN(n11564) );
  INV_X1 U14758 ( .A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11527) );
  INV_X1 U14759 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11520) );
  INV_X1 U14760 ( .A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11519) );
  OAI22_X1 U14761 ( .A1(n10717), .A2(n11520), .B1(n13921), .B2(n11519), .ZN(
        n11524) );
  INV_X1 U14762 ( .A(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11521) );
  OAI22_X1 U14763 ( .A1(n10718), .A2(n11522), .B1(n10719), .B2(n11521), .ZN(
        n11523) );
  AOI211_X1 U14764 ( .C1(n10544), .C2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n11524), .B(n11523), .ZN(n11526) );
  AOI22_X1 U14765 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11525) );
  OAI211_X1 U14766 ( .C1(n11555), .C2(n11527), .A(n11526), .B(n11525), .ZN(
        n11535) );
  AOI22_X1 U14767 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14768 ( .A1(n11528), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9577), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14769 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14770 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14771 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  NOR2_X1 U14772 ( .A1(n11535), .A2(n11534), .ZN(n11565) );
  XOR2_X1 U14773 ( .A(n11564), .B(n11565), .Z(n11540) );
  INV_X1 U14774 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n14714) );
  NAND2_X1 U14775 ( .A1(n11005), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11536) );
  OAI211_X1 U14776 ( .C1(n11537), .C2(n14714), .A(n11573), .B(n11536), .ZN(
        n11538) );
  AOI21_X1 U14777 ( .B1(n11540), .B2(n11539), .A(n11538), .ZN(n11541) );
  AOI21_X1 U14778 ( .B1(n14723), .B2(n11431), .A(n11541), .ZN(n13749) );
  INV_X1 U14779 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11578) );
  XNOR2_X1 U14780 ( .A(n11579), .B(n11578), .ZN(n14522) );
  INV_X1 U14781 ( .A(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11543) );
  OAI22_X1 U14782 ( .A1(n10742), .A2(n11545), .B1(n11544), .B2(n11543), .ZN(
        n11549) );
  INV_X1 U14783 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11546) );
  OAI22_X1 U14784 ( .A1(n10717), .A2(n11547), .B1(n13921), .B2(n11546), .ZN(
        n11548) );
  AOI211_X1 U14785 ( .C1(n11550), .C2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n11549), .B(n11548), .ZN(n11553) );
  AOI22_X1 U14786 ( .A1(n11316), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11551), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11552) );
  OAI211_X1 U14787 ( .C1(n11555), .C2(n11554), .A(n11553), .B(n11552), .ZN(
        n11563) );
  AOI22_X1 U14788 ( .A1(n11556), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10674), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14789 ( .A1(n10632), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10762), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11560) );
  AOI22_X1 U14790 ( .A1(n11497), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10651), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11559) );
  AOI22_X1 U14791 ( .A1(n11529), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11557), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11558) );
  NAND4_X1 U14792 ( .A1(n11561), .A2(n11560), .A3(n11559), .A4(n11558), .ZN(
        n11562) );
  NOR2_X1 U14793 ( .A1(n11563), .A2(n11562), .ZN(n11567) );
  NOR2_X1 U14794 ( .A1(n11565), .A2(n11564), .ZN(n11566) );
  XOR2_X1 U14795 ( .A(n11567), .B(n11566), .Z(n11571) );
  AOI21_X1 U14796 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n11005), .A(
        n11431), .ZN(n11569) );
  NAND2_X1 U14797 ( .A1(n11575), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11568) );
  OAI211_X1 U14798 ( .C1(n11571), .C2(n11570), .A(n11569), .B(n11568), .ZN(
        n11572) );
  OAI21_X1 U14799 ( .B1(n14522), .B2(n11573), .A(n11572), .ZN(n13729) );
  AOI22_X1 U14800 ( .A1(n11575), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11574), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11576) );
  NAND2_X1 U14801 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n21508), .ZN(n17278) );
  INV_X1 U14802 ( .A(n13731), .ZN(n11586) );
  NAND2_X1 U14803 ( .A1(n21341), .A2(n11584), .ZN(n21506) );
  NAND2_X1 U14804 ( .A1(n21506), .A2(n10276), .ZN(n11581) );
  NAND2_X1 U14805 ( .A1(n10276), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11583) );
  NAND2_X1 U14806 ( .A1(n21497), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11582) );
  AND2_X1 U14807 ( .A1(n11583), .A2(n11582), .ZN(n14082) );
  OR2_X2 U14808 ( .A1(n20773), .A2(n14082), .ZN(n20784) );
  INV_X1 U14809 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14740) );
  NOR2_X1 U14810 ( .A1(n15360), .A2(n14740), .ZN(n15370) );
  AOI21_X1 U14811 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n15370), .ZN(n11585) );
  OAI21_X1 U14812 ( .B1(n11586), .B2(n20784), .A(n11585), .ZN(n11587) );
  NAND2_X1 U14813 ( .A1(n15359), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11593) );
  INV_X1 U14814 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15493) );
  MUX2_X1 U14815 ( .A(n11596), .B(n11595), .S(n15353), .Z(n11598) );
  OAI21_X1 U14816 ( .B1(n14911), .B2(n11602), .A(n11601), .ZN(n15174) );
  INV_X1 U14817 ( .A(n15174), .ZN(n14897) );
  INV_X1 U14818 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14904) );
  NOR2_X1 U14819 ( .A1(n15360), .A2(n14904), .ZN(n15488) );
  AOI21_X1 U14820 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15488), .ZN(n11603) );
  OAI21_X1 U14821 ( .B1(n20784), .B2(n14909), .A(n11603), .ZN(n11604) );
  AOI21_X1 U14822 ( .B1(n14897), .B2(n20779), .A(n11604), .ZN(n11605) );
  BUF_X4 U14823 ( .A(n11610), .Z(n11971) );
  AND2_X4 U14824 ( .A1(n11606), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11977) );
  AOI22_X1 U14825 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11608) );
  AND2_X4 U14826 ( .A1(n16657), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12037) );
  AOI22_X1 U14827 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11607) );
  BUF_X4 U14828 ( .A(n11610), .Z(n11785) );
  AOI22_X1 U14829 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14830 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U14831 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U14832 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11972), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14833 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14834 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11616) );
  AOI22_X1 U14835 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11615) );
  NAND4_X1 U14836 ( .A1(n11618), .A2(n11617), .A3(n11616), .A4(n11615), .ZN(
        n11619) );
  AOI22_X1 U14837 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11971), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14838 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14839 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9571), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14840 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11620) );
  NAND4_X1 U14841 ( .A1(n11623), .A2(n11622), .A3(n11621), .A4(n11620), .ZN(
        n11624) );
  NAND2_X1 U14842 ( .A1(n11624), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11625) );
  AOI22_X1 U14843 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11628) );
  AOI22_X1 U14844 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14845 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14846 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U14847 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U14848 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14849 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9571), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14850 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14851 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14852 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U14853 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11635) );
  NAND4_X1 U14854 ( .A1(n11638), .A2(n11637), .A3(n11636), .A4(n11635), .ZN(
        n11639) );
  NAND2_X1 U14855 ( .A1(n11639), .A2(n11656), .ZN(n11646) );
  AOI22_X1 U14856 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14857 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11642) );
  AOI22_X1 U14858 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14859 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11640) );
  NAND4_X1 U14860 ( .A1(n11643), .A2(n11642), .A3(n11641), .A4(n11640), .ZN(
        n11644) );
  NAND2_X1 U14861 ( .A1(n11644), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11645) );
  AOI22_X1 U14862 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U14863 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14864 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11650) );
  NAND3_X1 U14865 ( .A1(n9664), .A2(n11656), .A3(n10445), .ZN(n11655) );
  AOI22_X1 U14866 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14867 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14868 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11652) );
  NAND3_X1 U14869 ( .A1(n9654), .A2(n11653), .A3(n11652), .ZN(n11654) );
  AND2_X2 U14870 ( .A1(n11655), .A2(n11654), .ZN(n11686) );
  AOI22_X1 U14871 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11972), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14872 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11659) );
  AOI22_X1 U14873 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11658) );
  NAND4_X1 U14874 ( .A1(n10444), .A2(n11660), .A3(n11659), .A4(n11658), .ZN(
        n11668) );
  AOI22_X1 U14875 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11666) );
  NAND2_X1 U14876 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11661) );
  AOI22_X1 U14877 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11664) );
  AOI22_X1 U14878 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9571), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11663) );
  NAND4_X1 U14879 ( .A1(n11666), .A2(n11665), .A3(n11664), .A4(n11663), .ZN(
        n11667) );
  AND2_X2 U14880 ( .A1(n11668), .A2(n11667), .ZN(n11685) );
  AOI22_X1 U14881 ( .A1(n9585), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12037), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14882 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14883 ( .A1(n11785), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11671) );
  BUF_X2 U14884 ( .A(n11790), .Z(n12089) );
  AOI21_X1 U14885 ( .B1(n12089), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n11669), .ZN(n11670) );
  AOI22_X1 U14886 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11971), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14887 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11972), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11677) );
  AOI22_X1 U14888 ( .A1(n9572), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14889 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14890 ( .A1(n11685), .A2(n11686), .ZN(n11705) );
  AOI22_X1 U14891 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9572), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11678) );
  AOI22_X1 U14892 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9571), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14893 ( .A1(n11971), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11977), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14894 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14895 ( .A1(n11972), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11790), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11679) );
  NAND4_X1 U14896 ( .A1(n11682), .A2(n11681), .A3(n11680), .A4(n11679), .ZN(
        n11683) );
  CLKBUF_X3 U14897 ( .A(n12179), .Z(n19985) );
  NAND2_X2 U14898 ( .A1(n11686), .A2(n11713), .ZN(n12197) );
  NAND2_X1 U14899 ( .A1(n12197), .A2(n13135), .ZN(n11687) );
  NAND2_X1 U14900 ( .A1(n11687), .A2(n9686), .ZN(n11704) );
  INV_X1 U14901 ( .A(n11704), .ZN(n11691) );
  OAI21_X1 U14902 ( .B1(n11698), .B2(n15607), .A(n19997), .ZN(n11690) );
  BUF_X4 U14903 ( .A(n11688), .Z(n12445) );
  INV_X1 U14904 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14632) );
  NAND2_X1 U14905 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11694) );
  NAND2_X1 U14906 ( .A1(n15612), .A2(n11694), .ZN(n11695) );
  AOI21_X1 U14907 ( .B1(n9582), .B2(P2_EBX_REG_0__SCAN_IN), .A(n11695), .ZN(
        n11696) );
  OAI21_X1 U14908 ( .B1(n11738), .B2(n14632), .A(n11696), .ZN(n11697) );
  INV_X1 U14909 ( .A(n11697), .ZN(n11715) );
  NAND2_X1 U14910 ( .A1(n11698), .A2(n11705), .ZN(n12135) );
  OR2_X2 U14911 ( .A1(n12135), .A2(n11699), .ZN(n12137) );
  NAND2_X1 U14912 ( .A1(n11700), .A2(n15607), .ZN(n11701) );
  NAND2_X1 U14913 ( .A1(n12197), .A2(n19985), .ZN(n13124) );
  NAND3_X1 U14914 ( .A1(n20003), .A2(n19997), .A3(n11685), .ZN(n11703) );
  NAND2_X1 U14915 ( .A1(n11704), .A2(n11703), .ZN(n11707) );
  AND2_X1 U14916 ( .A1(n11705), .A2(n19992), .ZN(n11706) );
  OAI21_X1 U14917 ( .B1(n16815), .B2(n13135), .A(n12154), .ZN(n11709) );
  NAND2_X1 U14918 ( .A1(n11716), .A2(n19839), .ZN(n11711) );
  INV_X1 U14919 ( .A(n13095), .ZN(n11712) );
  NAND2_X1 U14920 ( .A1(n11712), .A2(n15607), .ZN(n13788) );
  OAI21_X1 U14921 ( .B1(n13119), .B2(n16815), .A(n9605), .ZN(n11719) );
  AND2_X1 U14922 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n11717) );
  OAI22_X1 U14923 ( .A1(n11719), .A2(n11718), .B1(n9583), .B2(n11717), .ZN(
        n11722) );
  OAI22_X1 U14924 ( .A1(n16673), .A2(n16837), .B1(n20604), .B2(n15612), .ZN(
        n11720) );
  INV_X1 U14925 ( .A(n11720), .ZN(n11721) );
  NAND2_X1 U14926 ( .A1(n11722), .A2(n11721), .ZN(n11764) );
  INV_X1 U14927 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20511) );
  NAND2_X1 U14928 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14929 ( .A1(n12879), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11725) );
  OAI211_X1 U14930 ( .C1(n12779), .C2(n20511), .A(n11726), .B(n11725), .ZN(
        n11727) );
  INV_X1 U14931 ( .A(n11727), .ZN(n11728) );
  AOI21_X1 U14932 ( .B1(n16837), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11730) );
  INV_X1 U14933 ( .A(n11732), .ZN(n11733) );
  NOR2_X1 U14934 ( .A1(n15612), .A2(n20586), .ZN(n11737) );
  AOI22_X1 U14935 ( .A1(n12879), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11739) );
  OAI21_X1 U14936 ( .B1(n12887), .B2(n17306), .A(n11742), .ZN(n12806) );
  XNOR2_X2 U14937 ( .A(n12805), .B(n11744), .ZN(n12410) );
  NAND2_X1 U14938 ( .A1(n12410), .A2(n11776), .ZN(n11748) );
  NAND2_X1 U14939 ( .A1(n11752), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19978) );
  OAI211_X1 U14940 ( .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n11752), .A(
        n19978), .B(n20382), .ZN(n11745) );
  INV_X1 U14941 ( .A(n11745), .ZN(n11746) );
  AOI21_X1 U14942 ( .B1(n11773), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n11746), .ZN(n11747) );
  NAND2_X1 U14943 ( .A1(n11748), .A2(n11747), .ZN(n11783) );
  OR2_X1 U14944 ( .A1(n11783), .A2(n11749), .ZN(n11750) );
  NAND2_X1 U14945 ( .A1(n11783), .A2(n11749), .ZN(n14370) );
  NAND2_X1 U14946 ( .A1(n12396), .A2(n11776), .ZN(n11758) );
  INV_X1 U14947 ( .A(n11752), .ZN(n11755) );
  INV_X1 U14948 ( .A(n20302), .ZN(n11753) );
  NAND2_X1 U14949 ( .A1(n11753), .A2(n20594), .ZN(n11754) );
  NAND2_X1 U14950 ( .A1(n11755), .A2(n11754), .ZN(n16747) );
  NOR2_X1 U14951 ( .A1(n16747), .A2(n20575), .ZN(n11756) );
  AOI21_X1 U14952 ( .B1(n11773), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11756), .ZN(n11757) );
  NAND2_X1 U14953 ( .A1(n11758), .A2(n11757), .ZN(n11760) );
  OR2_X1 U14954 ( .A1(n11760), .A2(n11759), .ZN(n11761) );
  NAND2_X1 U14955 ( .A1(n11760), .A2(n11759), .ZN(n11780) );
  INV_X1 U14956 ( .A(n11763), .ZN(n11766) );
  INV_X1 U14957 ( .A(n11764), .ZN(n11765) );
  NAND2_X1 U14958 ( .A1(n11766), .A2(n11765), .ZN(n11767) );
  NAND2_X1 U14959 ( .A1(n16652), .A2(n11776), .ZN(n11769) );
  AOI22_X1 U14960 ( .A1(n11773), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20382), .B2(n20604), .ZN(n11768) );
  NAND2_X1 U14961 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U14962 ( .A1(n11773), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14963 ( .A1(n16748), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20237) );
  NAND2_X1 U14964 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20604), .ZN(
        n20274) );
  NAND2_X1 U14965 ( .A1(n20237), .A2(n20274), .ZN(n20272) );
  NAND2_X1 U14966 ( .A1(n20272), .A2(n20382), .ZN(n20057) );
  NAND2_X1 U14967 ( .A1(n11774), .A2(n20057), .ZN(n11775) );
  INV_X1 U14968 ( .A(n11777), .ZN(n11778) );
  NOR2_X1 U14969 ( .A1(n16654), .A2(n11778), .ZN(n11779) );
  NAND2_X1 U14970 ( .A1(n14229), .A2(n14228), .ZN(n11781) );
  NAND2_X1 U14971 ( .A1(n11781), .A2(n11780), .ZN(n14234) );
  NAND2_X1 U14972 ( .A1(n14233), .A2(n14234), .ZN(n14232) );
  NAND2_X1 U14973 ( .A1(n11685), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11782) );
  NAND2_X1 U14974 ( .A1(n14232), .A2(n11782), .ZN(n14373) );
  AOI22_X1 U14975 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11789) );
  NAND2_X1 U14976 ( .A1(n9585), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12557) );
  INV_X4 U14977 ( .A(n12557), .ZN(n12281) );
  AOI22_X1 U14978 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11788) );
  AND2_X2 U14979 ( .A1(n11785), .A2(n11656), .ZN(n11846) );
  AND2_X2 U14980 ( .A1(n11971), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11821) );
  AOI22_X1 U14981 ( .A1(n11846), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14982 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U14983 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11796) );
  AND2_X2 U14984 ( .A1(n12037), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11951) );
  AOI22_X1 U14985 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14986 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11793) );
  AND2_X2 U14987 ( .A1(n11972), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12166) );
  AOI22_X1 U14988 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11792) );
  AND2_X2 U14989 ( .A1(n12089), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11917) );
  AOI22_X1 U14990 ( .A1(n12295), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14991 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11795) );
  NOR2_X1 U14992 ( .A1(n11796), .A2(n11795), .ZN(n15953) );
  INV_X1 U14993 ( .A(n15953), .ZN(n11845) );
  AOI22_X1 U14994 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12160), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11801) );
  AOI22_X1 U14995 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n12282), .ZN(n11800) );
  AOI22_X1 U14996 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12268), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14997 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n12288), .ZN(n11798) );
  NAND4_X1 U14998 ( .A1(n11801), .A2(n11800), .A3(n11799), .A4(n11798), .ZN(
        n11807) );
  AOI22_X1 U14999 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11851), .B1(
        n11951), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11805) );
  AOI22_X1 U15000 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9586), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11804) );
  AOI22_X1 U15001 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12166), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11803) );
  AOI22_X1 U15002 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11813), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11802) );
  NAND4_X1 U15003 ( .A1(n11805), .A2(n11804), .A3(n11803), .A4(n11802), .ZN(
        n11806) );
  AOI22_X1 U15004 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11808), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15005 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U15006 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U15007 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11809) );
  NAND4_X1 U15008 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n11819) );
  AOI22_X1 U15009 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11817) );
  AOI22_X1 U15010 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U15011 ( .A1(n12166), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15012 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11814) );
  NAND4_X1 U15013 ( .A1(n11817), .A2(n11816), .A3(n11815), .A4(n11814), .ZN(
        n11818) );
  AND2_X1 U15014 ( .A1(n15972), .A2(n15980), .ZN(n11844) );
  NAND2_X1 U15015 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14451) );
  INV_X1 U15016 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11820) );
  NOR2_X1 U15017 ( .A1(n14451), .A2(n11820), .ZN(n11843) );
  AOI22_X1 U15018 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U15019 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U15020 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U15021 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11822) );
  NAND4_X1 U15022 ( .A1(n11825), .A2(n11824), .A3(n11823), .A4(n11822), .ZN(
        n11831) );
  AOI22_X1 U15023 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U15024 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U15025 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U15026 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U15027 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11830) );
  AOI22_X1 U15028 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11835) );
  AOI22_X1 U15029 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U15030 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n11951), .B1(
        n11846), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15031 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11832) );
  NAND4_X1 U15032 ( .A1(n11835), .A2(n11834), .A3(n11833), .A4(n11832), .ZN(
        n11841) );
  AOI22_X1 U15033 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11851), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U15034 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n11872), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U15035 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12166), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15036 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11917), .B1(
        n11813), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11836) );
  NAND4_X1 U15037 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11840) );
  AND2_X1 U15038 ( .A1(n15960), .A2(n15968), .ZN(n11842) );
  NAND4_X1 U15039 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n15924) );
  INV_X1 U15040 ( .A(n14368), .ZN(n12050) );
  AOI22_X1 U15041 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15042 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U15043 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U15044 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11847) );
  NAND4_X1 U15045 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11857) );
  AOI22_X1 U15046 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U15047 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U15048 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U15049 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11852) );
  NAND4_X1 U15050 ( .A1(n11855), .A2(n11854), .A3(n11853), .A4(n11852), .ZN(
        n11856) );
  OR2_X1 U15051 ( .A1(n11857), .A2(n11856), .ZN(n15925) );
  AND2_X1 U15052 ( .A1(n15925), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11889) );
  AOI22_X1 U15053 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U15054 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U15055 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U15056 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U15057 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11867) );
  AOI22_X1 U15058 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U15059 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11864) );
  AOI22_X1 U15060 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11863) );
  AOI22_X1 U15061 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11862) );
  NAND4_X1 U15062 ( .A1(n11865), .A2(n11864), .A3(n11863), .A4(n11862), .ZN(
        n11866) );
  OR2_X1 U15063 ( .A1(n11867), .A2(n11866), .ZN(n12340) );
  AOI22_X1 U15064 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U15065 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U15066 ( .A1(n11846), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U15067 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U15068 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11878) );
  AOI22_X1 U15069 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U15070 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U15071 ( .A1(n12295), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U15072 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11873) );
  NAND4_X1 U15073 ( .A1(n11876), .A2(n11875), .A3(n11874), .A4(n11873), .ZN(
        n11877) );
  AOI22_X1 U15074 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U15075 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11881) );
  AOI22_X1 U15076 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U15077 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11879) );
  NAND4_X1 U15078 ( .A1(n11882), .A2(n11881), .A3(n11880), .A4(n11879), .ZN(
        n11888) );
  AOI22_X1 U15079 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U15080 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U15081 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U15082 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U15083 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11887) );
  OR2_X1 U15084 ( .A1(n11888), .A2(n11887), .ZN(n12333) );
  NAND4_X1 U15085 ( .A1(n11889), .A2(n12340), .A3(n15940), .A4(n12333), .ZN(
        n11890) );
  NOR3_X1 U15086 ( .A1(n15924), .A2(n12050), .A3(n11890), .ZN(n11891) );
  AOI22_X1 U15087 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12160), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U15088 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n12282), .ZN(n11894) );
  AOI22_X1 U15089 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12268), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U15090 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n12288), .ZN(n11892) );
  NAND4_X1 U15091 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11901) );
  AOI22_X1 U15092 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11851), .B1(
        n11951), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U15093 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9586), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U15094 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12166), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11897) );
  AOI22_X1 U15095 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11813), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11896) );
  NAND4_X1 U15096 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11900) );
  NOR2_X1 U15097 ( .A1(n11901), .A2(n11900), .ZN(n15921) );
  INV_X1 U15098 ( .A(n15921), .ZN(n11902) );
  AOI22_X1 U15099 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U15100 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U15101 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11846), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U15102 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11903) );
  NAND4_X1 U15103 ( .A1(n11906), .A2(n11905), .A3(n11904), .A4(n11903), .ZN(
        n11912) );
  AOI22_X1 U15104 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U15105 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n9586), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U15106 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11872), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U15107 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11813), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11907) );
  NAND4_X1 U15108 ( .A1(n11910), .A2(n11909), .A3(n11908), .A4(n11907), .ZN(
        n11911) );
  NOR2_X1 U15109 ( .A1(n11912), .A2(n11911), .ZN(n15917) );
  AOI22_X1 U15110 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15111 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15112 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15113 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U15114 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11923) );
  AOI22_X1 U15115 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U15116 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15117 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15118 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11918) );
  NAND4_X1 U15119 ( .A1(n11921), .A2(n11920), .A3(n11919), .A4(n11918), .ZN(
        n11922) );
  OR2_X1 U15120 ( .A1(n11923), .A2(n11922), .ZN(n15900) );
  AOI22_X1 U15121 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11927) );
  AOI22_X1 U15122 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11926) );
  AOI22_X1 U15123 ( .A1(n11846), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15124 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11924) );
  NAND4_X1 U15125 ( .A1(n11927), .A2(n11926), .A3(n11925), .A4(n11924), .ZN(
        n11933) );
  AOI22_X1 U15126 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15127 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15128 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15129 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U15130 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11932) );
  OR2_X1 U15131 ( .A1(n11933), .A2(n11932), .ZN(n15904) );
  AND2_X1 U15132 ( .A1(n15900), .A2(n15904), .ZN(n15895) );
  AOI22_X1 U15133 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15134 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15135 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15136 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11934) );
  NAND4_X1 U15137 ( .A1(n11937), .A2(n11936), .A3(n11935), .A4(n11934), .ZN(
        n11943) );
  AOI22_X1 U15138 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11941) );
  AOI22_X1 U15139 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11940) );
  AOI22_X1 U15140 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15141 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11938) );
  NAND4_X1 U15142 ( .A1(n11941), .A2(n11940), .A3(n11939), .A4(n11938), .ZN(
        n11942) );
  NOR2_X1 U15143 ( .A1(n11943), .A2(n11942), .ZN(n15897) );
  INV_X1 U15144 ( .A(n15897), .ZN(n11944) );
  AND2_X1 U15145 ( .A1(n15895), .A2(n11944), .ZN(n11958) );
  AOI22_X1 U15146 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11950) );
  NAND2_X1 U15147 ( .A1(n12282), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11945) );
  OAI21_X1 U15148 ( .B1(n12557), .B2(n12409), .A(n11945), .ZN(n11946) );
  INV_X1 U15149 ( .A(n11946), .ZN(n11949) );
  AOI22_X1 U15150 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15151 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15152 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11957) );
  AOI22_X1 U15153 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U15154 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15155 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15156 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U15157 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11956) );
  OR2_X1 U15158 ( .A1(n11957), .A2(n11956), .ZN(n15910) );
  AND2_X1 U15159 ( .A1(n11958), .A2(n15910), .ZN(n11959) );
  INV_X1 U15160 ( .A(n11992), .ZN(n15896) );
  AOI22_X1 U15161 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11963) );
  AOI22_X1 U15162 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15163 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15164 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U15165 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11969) );
  AOI22_X1 U15166 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U15167 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15168 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15169 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11964) );
  NAND4_X1 U15170 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11968) );
  NOR2_X1 U15171 ( .A1(n11969), .A2(n11968), .ZN(n12007) );
  AOI22_X1 U15172 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11980) );
  XNOR2_X1 U15173 ( .A(n11656), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14595) );
  NAND2_X1 U15174 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11976) );
  NAND2_X1 U15175 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11975) );
  INV_X1 U15176 ( .A(n11972), .ZN(n16674) );
  INV_X1 U15177 ( .A(n16674), .ZN(n16692) );
  NAND2_X1 U15178 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11974) );
  NAND2_X1 U15179 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11973) );
  AND4_X1 U15180 ( .A1(n11976), .A2(n11975), .A3(n11974), .A4(n11973), .ZN(
        n11979) );
  AOI22_X1 U15181 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U15182 ( .A1(n11980), .A2(n14595), .A3(n11979), .A4(n11978), .ZN(
        n11989) );
  AOI22_X1 U15183 ( .A1(n11784), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14592), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11987) );
  NAND2_X1 U15184 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11984) );
  NAND2_X1 U15185 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U15186 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11982) );
  NAND2_X1 U15187 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11981) );
  AND4_X1 U15188 ( .A1(n11984), .A2(n11983), .A3(n11982), .A4(n11981), .ZN(
        n11986) );
  AOI22_X1 U15189 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11985) );
  NAND4_X1 U15190 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n14587), .ZN(
        n11988) );
  NAND2_X1 U15191 ( .A1(n11989), .A2(n11988), .ZN(n12012) );
  XOR2_X1 U15192 ( .A(n12007), .B(n11990), .Z(n12013) );
  INV_X1 U15193 ( .A(n12013), .ZN(n11991) );
  NAND2_X1 U15194 ( .A1(n15896), .A2(n11991), .ZN(n11994) );
  INV_X1 U15195 ( .A(n12012), .ZN(n12008) );
  AOI22_X1 U15196 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15197 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11995) );
  AND2_X1 U15198 ( .A1(n11996), .A2(n11995), .ZN(n11999) );
  AOI22_X1 U15199 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9585), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15200 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11997) );
  NAND4_X1 U15201 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n14587), .ZN(
        n12006) );
  AOI22_X1 U15202 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15203 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12000) );
  AND2_X1 U15204 ( .A1(n12001), .A2(n12000), .ZN(n12004) );
  AOI22_X1 U15205 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15206 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U15207 ( .A1(n12004), .A2(n14595), .A3(n12003), .A4(n12002), .ZN(
        n12005) );
  NAND2_X1 U15208 ( .A1(n12006), .A2(n12005), .ZN(n12014) );
  INV_X1 U15209 ( .A(n12007), .ZN(n12009) );
  NAND2_X1 U15210 ( .A1(n12009), .A2(n12008), .ZN(n12015) );
  XOR2_X1 U15211 ( .A(n12014), .B(n12015), .Z(n12010) );
  NAND2_X1 U15212 ( .A1(n12010), .A2(n14368), .ZN(n15883) );
  INV_X1 U15213 ( .A(n12014), .ZN(n12011) );
  NOR2_X1 U15214 ( .A1(n12015), .A2(n12014), .ZN(n12028) );
  AOI22_X1 U15215 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16692), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15216 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12089), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12016) );
  AND2_X1 U15217 ( .A1(n12017), .A2(n12016), .ZN(n12020) );
  AOI22_X1 U15218 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9585), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15219 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15220 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n14587), .ZN(
        n12027) );
  AOI22_X1 U15221 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12022) );
  INV_X1 U15222 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20453) );
  AOI22_X1 U15223 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12021) );
  AND2_X1 U15224 ( .A1(n12022), .A2(n12021), .ZN(n12025) );
  AOI22_X1 U15225 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12024) );
  INV_X1 U15226 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n21641) );
  AOI22_X1 U15227 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12023) );
  NAND4_X1 U15228 ( .A1(n12025), .A2(n14595), .A3(n12024), .A4(n12023), .ZN(
        n12026) );
  AND2_X1 U15229 ( .A1(n12027), .A2(n12026), .ZN(n12029) );
  NAND2_X1 U15230 ( .A1(n12028), .A2(n12029), .ZN(n12051) );
  OAI211_X1 U15231 ( .C1(n12028), .C2(n12029), .A(n12051), .B(n14368), .ZN(
        n12047) );
  AOI22_X1 U15232 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9585), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U15233 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12033) );
  NAND2_X1 U15234 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n12032) );
  NAND2_X1 U15235 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12031) );
  NAND2_X1 U15236 ( .A1(n12089), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12030) );
  AND4_X1 U15237 ( .A1(n12033), .A2(n12032), .A3(n12031), .A4(n12030), .ZN(
        n12035) );
  AOI22_X1 U15238 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U15239 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n14587), .ZN(
        n12046) );
  AOI22_X1 U15240 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U15241 ( .A1(n12037), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12041) );
  NAND2_X1 U15242 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12040) );
  NAND2_X1 U15243 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n12039) );
  NAND2_X1 U15244 ( .A1(n14599), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12038) );
  AND4_X1 U15245 ( .A1(n12041), .A2(n12040), .A3(n12039), .A4(n12038), .ZN(
        n12043) );
  AOI22_X1 U15246 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12042) );
  NAND4_X1 U15247 ( .A1(n12044), .A2(n14595), .A3(n12043), .A4(n12042), .ZN(
        n12045) );
  NAND2_X1 U15248 ( .A1(n12046), .A2(n12045), .ZN(n15870) );
  NOR2_X1 U15249 ( .A1(n15868), .A2(n10427), .ZN(n12055) );
  INV_X1 U15250 ( .A(n15869), .ZN(n12053) );
  INV_X1 U15251 ( .A(n12051), .ZN(n12049) );
  INV_X1 U15252 ( .A(n15870), .ZN(n12048) );
  AND2_X1 U15253 ( .A1(n12049), .A2(n12048), .ZN(n12068) );
  AOI211_X1 U15254 ( .C1(n15870), .C2(n12051), .A(n12050), .B(n12068), .ZN(
        n15873) );
  INV_X1 U15255 ( .A(n15873), .ZN(n12052) );
  NOR2_X2 U15256 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  AOI22_X1 U15257 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16692), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12057) );
  AOI22_X1 U15258 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12056) );
  AND2_X1 U15259 ( .A1(n12057), .A2(n12056), .ZN(n12060) );
  AOI22_X1 U15260 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15261 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12058) );
  NAND4_X1 U15262 ( .A1(n12060), .A2(n12059), .A3(n12058), .A4(n14587), .ZN(
        n12067) );
  INV_X1 U15263 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n21647) );
  AOI22_X1 U15264 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n16692), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U15265 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12061) );
  AND2_X1 U15266 ( .A1(n12062), .A2(n12061), .ZN(n12065) );
  AOI22_X1 U15267 ( .A1(n9584), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12064) );
  INV_X1 U15268 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n20372) );
  AOI22_X1 U15269 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14592), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15270 ( .A1(n12065), .A2(n14595), .A3(n12064), .A4(n12063), .ZN(
        n12066) );
  AND2_X1 U15271 ( .A1(n12067), .A2(n12066), .ZN(n12070) );
  NAND2_X1 U15272 ( .A1(n12068), .A2(n12070), .ZN(n15863) );
  OAI211_X1 U15273 ( .C1(n12068), .C2(n12070), .A(n14368), .B(n15863), .ZN(
        n12069) );
  AOI22_X1 U15274 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15275 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12071) );
  AND2_X1 U15276 ( .A1(n12072), .A2(n12071), .ZN(n12075) );
  AOI22_X1 U15277 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15278 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12073) );
  NAND4_X1 U15279 ( .A1(n12075), .A2(n12074), .A3(n12073), .A4(n14587), .ZN(
        n12083) );
  AOI22_X1 U15280 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15281 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12077) );
  AND2_X1 U15282 ( .A1(n12078), .A2(n12077), .ZN(n12081) );
  AOI22_X1 U15283 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9585), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15284 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12079) );
  NAND4_X1 U15285 ( .A1(n12081), .A2(n14595), .A3(n12080), .A4(n12079), .ZN(
        n12082) );
  NAND2_X1 U15286 ( .A1(n12083), .A2(n12082), .ZN(n15865) );
  AOI22_X1 U15287 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15288 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12084) );
  AND2_X1 U15289 ( .A1(n12085), .A2(n12084), .ZN(n12088) );
  AOI22_X1 U15290 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12087) );
  INV_X1 U15291 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n21585) );
  AOI22_X1 U15292 ( .A1(n9585), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14592), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12086) );
  NAND4_X1 U15293 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n14587), .ZN(
        n12096) );
  AOI22_X1 U15294 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16692), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U15295 ( .A1(n14597), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12089), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12090) );
  AND2_X1 U15296 ( .A1(n12091), .A2(n12090), .ZN(n12094) );
  AOI22_X1 U15297 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9584), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15298 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12092) );
  NAND4_X1 U15299 ( .A1(n12094), .A2(n14595), .A3(n12093), .A4(n12092), .ZN(
        n12095) );
  NAND2_X1 U15300 ( .A1(n12096), .A2(n12095), .ZN(n12098) );
  OR3_X1 U15301 ( .A1(n15863), .A2(n19985), .A3(n15865), .ZN(n12097) );
  NOR2_X1 U15302 ( .A1(n12097), .A2(n12098), .ZN(n14585) );
  AOI21_X1 U15303 ( .B1(n12098), .B2(n12097), .A(n14585), .ZN(n12156) );
  NAND2_X1 U15304 ( .A1(n16748), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12100) );
  NAND2_X1 U15305 ( .A1(n16656), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12099) );
  NAND2_X1 U15306 ( .A1(n12100), .A2(n12099), .ZN(n12109) );
  NAND2_X1 U15307 ( .A1(n20604), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12104) );
  NAND2_X1 U15308 ( .A1(n12105), .A2(n12100), .ZN(n12116) );
  XNOR2_X1 U15309 ( .A(n20594), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12101) );
  XNOR2_X1 U15310 ( .A(n12116), .B(n12101), .ZN(n12553) );
  INV_X1 U15311 ( .A(n12553), .ZN(n12564) );
  NAND2_X1 U15312 ( .A1(n12102), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12103) );
  NAND2_X1 U15313 ( .A1(n12109), .A2(n12104), .ZN(n12567) );
  AND2_X1 U15314 ( .A1(n12105), .A2(n12567), .ZN(n12150) );
  OAI21_X1 U15315 ( .B1(n12445), .B2(n12566), .A(n12150), .ZN(n12106) );
  OAI21_X1 U15316 ( .B1(n12564), .B2(n15871), .A(n12106), .ZN(n12107) );
  NAND2_X1 U15317 ( .A1(n12107), .A2(n16815), .ZN(n12111) );
  INV_X1 U15318 ( .A(n12566), .ZN(n12108) );
  OAI21_X1 U15319 ( .B1(n12109), .B2(n12108), .A(n9576), .ZN(n12110) );
  NAND2_X1 U15320 ( .A1(n12111), .A2(n12110), .ZN(n12114) );
  NAND2_X1 U15321 ( .A1(n15606), .A2(n12445), .ZN(n12112) );
  MUX2_X1 U15322 ( .A(n12112), .B(n14621), .S(n12553), .Z(n12113) );
  NAND2_X1 U15323 ( .A1(n12114), .A2(n12113), .ZN(n12125) );
  NAND2_X1 U15324 ( .A1(n16797), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12115) );
  NAND2_X1 U15325 ( .A1(n12116), .A2(n12115), .ZN(n12118) );
  NAND2_X1 U15326 ( .A1(n20594), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12117) );
  NAND3_X1 U15327 ( .A1(n12126), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n12127), .ZN(n12124) );
  INV_X1 U15328 ( .A(n12120), .ZN(n12121) );
  XNOR2_X1 U15329 ( .A(n12122), .B(n12121), .ZN(n12123) );
  MUX2_X1 U15330 ( .A(n12125), .B(n14621), .S(n12569), .Z(n12132) );
  INV_X1 U15331 ( .A(n12126), .ZN(n12129) );
  NOR2_X1 U15332 ( .A1(n12127), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12128) );
  NAND2_X1 U15333 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12127), .ZN(
        n12130) );
  NAND2_X1 U15334 ( .A1(n12132), .A2(n12572), .ZN(n12133) );
  MUX2_X1 U15335 ( .A(n12133), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n9587), .Z(n13094) );
  NAND2_X1 U15336 ( .A1(n12136), .A2(n14617), .ZN(n13134) );
  AND2_X1 U15337 ( .A1(n13134), .A2(n12137), .ZN(n12144) );
  INV_X1 U15338 ( .A(n12138), .ZN(n12139) );
  NAND2_X1 U15339 ( .A1(n12139), .A2(n16815), .ZN(n19833) );
  NAND2_X1 U15340 ( .A1(n12145), .A2(n16815), .ZN(n12141) );
  NAND3_X1 U15341 ( .A1(n12141), .A2(n19992), .A3(n12140), .ZN(n12142) );
  NAND2_X1 U15342 ( .A1(n19833), .A2(n12142), .ZN(n12143) );
  NAND2_X1 U15343 ( .A1(n12144), .A2(n12143), .ZN(n13099) );
  INV_X1 U15344 ( .A(n12197), .ZN(n12155) );
  INV_X1 U15345 ( .A(n12145), .ZN(n12146) );
  NAND2_X1 U15346 ( .A1(n12155), .A2(n12146), .ZN(n12147) );
  NAND2_X1 U15347 ( .A1(n12553), .A2(n12150), .ZN(n12151) );
  NOR2_X1 U15348 ( .A1(n12149), .A2(n16800), .ZN(n13793) );
  NAND2_X1 U15349 ( .A1(n12154), .A2(n12153), .ZN(n13129) );
  NOR2_X1 U15350 ( .A1(n13680), .A2(n16062), .ZN(n12158) );
  INV_X1 U15351 ( .A(n14586), .ZN(n12157) );
  NAND2_X1 U15352 ( .A1(n12158), .A2(n12157), .ZN(n12395) );
  NOR2_X1 U15353 ( .A1(n12178), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15354 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15355 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15356 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15357 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12161) );
  NAND4_X1 U15358 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12172) );
  AOI22_X1 U15359 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15360 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15361 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15362 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12167) );
  NAND4_X1 U15363 ( .A1(n12170), .A2(n12169), .A3(n12168), .A4(n12167), .ZN(
        n12171) );
  INV_X1 U15364 ( .A(n13890), .ZN(n12173) );
  NAND2_X1 U15365 ( .A1(n12445), .A2(n20581), .ZN(n12183) );
  OR2_X1 U15366 ( .A1(n12197), .A2(n12183), .ZN(n12213) );
  NAND2_X1 U15367 ( .A1(n20604), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20596) );
  NAND2_X1 U15368 ( .A1(n12177), .A2(n20596), .ZN(n12174) );
  NAND2_X1 U15369 ( .A1(n12213), .A2(n12174), .ZN(n12175) );
  INV_X1 U15370 ( .A(n12177), .ZN(n12196) );
  NAND2_X1 U15371 ( .A1(n12215), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12182) );
  INV_X1 U15372 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12181) );
  NAND2_X1 U15373 ( .A1(n12445), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12180) );
  NAND2_X1 U15374 ( .A1(n12182), .A2(n9653), .ZN(n13892) );
  NAND2_X1 U15375 ( .A1(n13893), .A2(n13892), .ZN(n12201) );
  INV_X2 U15376 ( .A(n12215), .ZN(n12373) );
  AOI22_X1 U15377 ( .A1(n12327), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12184) );
  XNOR2_X1 U15378 ( .A(n12201), .B(n12200), .ZN(n13965) );
  AOI22_X1 U15379 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12160), .B1(
        n11797), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15380 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n12282), .ZN(n12187) );
  AOI22_X1 U15381 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11846), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15382 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n12288), .ZN(n12185) );
  AOI22_X1 U15383 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n11813), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15384 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n12165), .B1(
        n9586), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15385 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n11851), .B1(
        n11951), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15386 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12166), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12190) );
  NAND3_X1 U15387 ( .A1(n10447), .A2(n12195), .A3(n12194), .ZN(n12468) );
  INV_X1 U15388 ( .A(n12468), .ZN(n12581) );
  OR2_X1 U15389 ( .A1(n12341), .A2(n12581), .ZN(n12199) );
  AOI22_X1 U15390 ( .A1(n12197), .A2(n12196), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12198) );
  AND2_X1 U15391 ( .A1(n12199), .A2(n12198), .ZN(n13964) );
  NAND2_X1 U15392 ( .A1(n13965), .A2(n13964), .ZN(n13967) );
  INV_X1 U15393 ( .A(n12200), .ZN(n12202) );
  NAND2_X1 U15394 ( .A1(n12202), .A2(n12201), .ZN(n12220) );
  NAND2_X1 U15395 ( .A1(n13967), .A2(n12220), .ZN(n15808) );
  AOI22_X1 U15396 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12160), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15397 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n12282), .ZN(n12205) );
  AOI22_X1 U15398 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n11846), .B1(
        n11951), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15399 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n12288), .ZN(n12203) );
  NAND4_X1 U15400 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n12212) );
  AOI22_X1 U15401 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n11821), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15402 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n9586), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15403 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n11813), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15404 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12166), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15405 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12211) );
  OR2_X1 U15406 ( .A1(n12341), .A2(n12563), .ZN(n12214) );
  OAI211_X1 U15407 ( .C1(n20581), .C2(n20594), .A(n12214), .B(n12213), .ZN(
        n12219) );
  XNOR2_X1 U15408 ( .A(n15808), .B(n12219), .ZN(n14051) );
  NAND2_X1 U15409 ( .A1(n13640), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12218) );
  AOI22_X1 U15410 ( .A1(n12327), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12217) );
  AND2_X1 U15411 ( .A1(n12218), .A2(n12217), .ZN(n14050) );
  INV_X1 U15412 ( .A(n12219), .ZN(n15807) );
  AND2_X1 U15413 ( .A1(n13965), .A2(n10451), .ZN(n12238) );
  OR2_X1 U15414 ( .A1(n12219), .A2(n12220), .ZN(n12236) );
  INV_X1 U15415 ( .A(n12341), .ZN(n12231) );
  AOI22_X1 U15416 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15417 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15418 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15419 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12221) );
  NAND4_X1 U15420 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12230) );
  AOI22_X1 U15421 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15422 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15423 ( .A1(n12166), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15424 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12165), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15425 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  AOI22_X1 U15426 ( .A1(n12231), .A2(n12579), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n12327), .ZN(n12234) );
  OAI22_X1 U15427 ( .A1(n12183), .A2(n17306), .B1(n20586), .B2(n20581), .ZN(
        n12232) );
  AOI21_X1 U15428 ( .B1(n13640), .B2(P2_REIP_REG_3__SCAN_IN), .A(n12232), .ZN(
        n12233) );
  AND2_X1 U15429 ( .A1(n12234), .A2(n12233), .ZN(n15810) );
  INV_X1 U15430 ( .A(n15810), .ZN(n12235) );
  NAND2_X1 U15431 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  NAND2_X1 U15432 ( .A1(n13640), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15433 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15434 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11808), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15435 ( .A1(n12282), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15436 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12239) );
  NAND4_X1 U15437 ( .A1(n12242), .A2(n12241), .A3(n12240), .A4(n12239), .ZN(
        n12248) );
  AOI22_X1 U15438 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15439 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15440 ( .A1(n12165), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15441 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U15442 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12247) );
  INV_X1 U15443 ( .A(n12585), .ZN(n12249) );
  OR2_X1 U15444 ( .A1(n12341), .A2(n12249), .ZN(n12251) );
  AOI22_X1 U15445 ( .A1(n12327), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12250) );
  AND3_X1 U15446 ( .A1(n12252), .A2(n12251), .A3(n12250), .ZN(n16089) );
  INV_X1 U15447 ( .A(n16089), .ZN(n12253) );
  AND2_X1 U15448 ( .A1(n15806), .A2(n12253), .ZN(n12254) );
  NAND2_X1 U15449 ( .A1(n13640), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15450 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11808), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15451 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15452 ( .A1(n11846), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15453 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12255) );
  NAND4_X1 U15454 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12264) );
  AOI22_X1 U15455 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15456 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11872), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15457 ( .A1(n12295), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15458 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12259) );
  NAND4_X1 U15459 ( .A1(n12262), .A2(n12261), .A3(n12260), .A4(n12259), .ZN(
        n12263) );
  OR2_X1 U15460 ( .A1(n12341), .A2(n12586), .ZN(n12266) );
  AOI22_X1 U15461 ( .A1(n12327), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15462 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9581), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15463 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12282), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15464 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11821), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15465 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12288), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12269) );
  NAND4_X1 U15466 ( .A1(n12272), .A2(n12271), .A3(n12270), .A4(n12269), .ZN(
        n12278) );
  AOI22_X1 U15467 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11851), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15468 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12295), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15469 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12166), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15470 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11917), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12273) );
  NAND4_X1 U15471 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12277) );
  INV_X1 U15472 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20516) );
  AOI22_X1 U15473 ( .A1(n12327), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12279) );
  OAI21_X1 U15474 ( .B1(n12373), .B2(n20516), .A(n12279), .ZN(n13878) );
  NAND2_X1 U15475 ( .A1(n9581), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12287) );
  NAND2_X1 U15476 ( .A1(n12160), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15477 ( .A1(n12281), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12285) );
  INV_X1 U15478 ( .A(n12282), .ZN(n12283) );
  INV_X1 U15479 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n21630) );
  OR2_X1 U15480 ( .A1(n12283), .A2(n21630), .ZN(n12284) );
  NAND2_X1 U15481 ( .A1(n11808), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n12294) );
  INV_X1 U15482 ( .A(n12288), .ZN(n12290) );
  INV_X1 U15483 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12289) );
  OR2_X1 U15484 ( .A1(n12290), .A2(n12289), .ZN(n12293) );
  NAND2_X1 U15485 ( .A1(n11821), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12292) );
  NAND2_X1 U15486 ( .A1(n12268), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12291) );
  NAND2_X1 U15487 ( .A1(n11951), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n12299) );
  NAND2_X1 U15488 ( .A1(n11851), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12298) );
  NAND2_X1 U15489 ( .A1(n12295), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12297) );
  NAND2_X1 U15490 ( .A1(n9586), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12296) );
  NAND2_X1 U15491 ( .A1(n11872), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n12305) );
  NAND2_X1 U15492 ( .A1(n12166), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12304) );
  NAND2_X1 U15493 ( .A1(n11917), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n12303) );
  NAND2_X1 U15494 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12302) );
  INV_X1 U15495 ( .A(n12590), .ZN(n12523) );
  INV_X1 U15496 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20518) );
  AOI22_X1 U15497 ( .A1(n12327), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12311) );
  OAI21_X1 U15498 ( .B1(n12373), .B2(n20518), .A(n12311), .ZN(n13887) );
  INV_X1 U15499 ( .A(n13883), .ZN(n12316) );
  NAND2_X1 U15500 ( .A1(n13640), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n12314) );
  INV_X1 U15501 ( .A(n15980), .ZN(n15951) );
  OR2_X1 U15502 ( .A1(n12341), .A2(n15951), .ZN(n12313) );
  AOI22_X1 U15503 ( .A1(n12327), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U15504 ( .A1(n13640), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12320) );
  INV_X1 U15505 ( .A(n15972), .ZN(n12317) );
  OR2_X1 U15506 ( .A1(n12341), .A2(n12317), .ZN(n12319) );
  AOI22_X1 U15507 ( .A1(n12327), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12216), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12318) );
  NAND2_X1 U15508 ( .A1(n13640), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12324) );
  INV_X1 U15509 ( .A(n15968), .ZN(n15952) );
  OR2_X1 U15510 ( .A1(n12341), .A2(n15952), .ZN(n12323) );
  AOI22_X1 U15511 ( .A1(n12327), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12322) );
  INV_X1 U15512 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19703) );
  INV_X1 U15513 ( .A(n15960), .ZN(n15954) );
  OR2_X1 U15514 ( .A1(n12341), .A2(n15954), .ZN(n12326) );
  AOI22_X1 U15515 ( .A1(n12327), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12325) );
  OAI211_X1 U15516 ( .C1(n12373), .C2(n19703), .A(n12326), .B(n12325), .ZN(
        n14023) );
  NAND2_X1 U15517 ( .A1(n13977), .A2(n14023), .ZN(n14021) );
  INV_X1 U15518 ( .A(n14021), .ZN(n12332) );
  NAND2_X1 U15519 ( .A1(n13640), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n12330) );
  OR2_X1 U15520 ( .A1(n12341), .A2(n15953), .ZN(n12329) );
  AOI22_X1 U15521 ( .A1(n12327), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U15522 ( .A1(n12332), .A2(n12331), .ZN(n14118) );
  NAND2_X1 U15523 ( .A1(n13640), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12336) );
  OR2_X1 U15524 ( .A1(n12341), .A2(n15944), .ZN(n12335) );
  AOI22_X1 U15525 ( .A1(n12327), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12334) );
  INV_X1 U15526 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n20529) );
  INV_X1 U15527 ( .A(n15940), .ZN(n12337) );
  OR2_X1 U15528 ( .A1(n12341), .A2(n12337), .ZN(n12339) );
  AOI22_X1 U15529 ( .A1(n12327), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12338) );
  OAI211_X1 U15530 ( .C1(n12373), .C2(n20529), .A(n12339), .B(n12338), .ZN(
        n14224) );
  NAND2_X1 U15531 ( .A1(n13640), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12344) );
  INV_X1 U15532 ( .A(n12340), .ZN(n15931) );
  OR2_X1 U15533 ( .A1(n12341), .A2(n15931), .ZN(n12343) );
  AOI22_X1 U15534 ( .A1(n12327), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12342) );
  NAND2_X1 U15535 ( .A1(n13640), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15536 ( .A1(n12327), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12346) );
  NOR2_X2 U15537 ( .A1(n14323), .A2(n16497), .ZN(n14563) );
  INV_X1 U15538 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20535) );
  AOI22_X1 U15539 ( .A1(n12327), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12348) );
  OAI21_X1 U15540 ( .B1(n12373), .B2(n20535), .A(n12348), .ZN(n14566) );
  INV_X1 U15541 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19630) );
  AOI22_X1 U15542 ( .A1(n12327), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12349) );
  OAI21_X1 U15543 ( .B1(n12373), .B2(n19630), .A(n12349), .ZN(n16067) );
  NAND2_X1 U15544 ( .A1(n13640), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15545 ( .A1(n12327), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12350) );
  INV_X1 U15546 ( .A(n15737), .ZN(n12356) );
  NAND2_X1 U15547 ( .A1(n13640), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15548 ( .A1(n12327), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12353) );
  INV_X1 U15549 ( .A(n15736), .ZN(n12355) );
  NAND2_X1 U15550 ( .A1(n12356), .A2(n12355), .ZN(n15739) );
  NAND2_X1 U15551 ( .A1(n13640), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15552 ( .A1(n12327), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12357) );
  NOR2_X2 U15553 ( .A1(n15739), .A2(n13666), .ZN(n13665) );
  INV_X1 U15554 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20544) );
  AOI22_X1 U15555 ( .A1(n12327), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12359) );
  OAI21_X1 U15556 ( .B1(n12373), .B2(n20544), .A(n12359), .ZN(n15711) );
  NAND2_X1 U15557 ( .A1(n13665), .A2(n15711), .ZN(n15698) );
  NAND2_X1 U15558 ( .A1(n13640), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15559 ( .A1(n12327), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12360) );
  INV_X1 U15560 ( .A(n15700), .ZN(n12362) );
  NAND2_X1 U15561 ( .A1(n13640), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15562 ( .A1(n12327), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12363) );
  INV_X1 U15563 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20550) );
  AOI22_X1 U15564 ( .A1(n12327), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12365) );
  OAI21_X1 U15565 ( .B1(n12373), .B2(n20550), .A(n12365), .ZN(n15676) );
  NAND2_X1 U15566 ( .A1(n13640), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15567 ( .A1(n12327), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12366) );
  NOR2_X2 U15568 ( .A1(n15658), .A2(n15660), .ZN(n14529) );
  NAND2_X1 U15569 ( .A1(n13640), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12369) );
  AOI22_X1 U15570 ( .A1(n12327), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12368) );
  AND2_X1 U15571 ( .A1(n12369), .A2(n12368), .ZN(n14532) );
  INV_X1 U15572 ( .A(n14532), .ZN(n12370) );
  AND2_X2 U15573 ( .A1(n14529), .A2(n12370), .ZN(n14531) );
  INV_X1 U15574 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U15575 ( .A1(n12327), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12371) );
  OAI21_X1 U15576 ( .B1(n12373), .B2(n16117), .A(n12371), .ZN(n15623) );
  INV_X1 U15577 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20556) );
  AOI22_X1 U15578 ( .A1(n12327), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12216), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12372) );
  OAI21_X1 U15579 ( .B1(n12373), .B2(n20556), .A(n12372), .ZN(n12374) );
  NOR2_X1 U15580 ( .A1(n16740), .A2(n16735), .ZN(n12376) );
  NAND2_X1 U15581 ( .A1(n19832), .A2(n12376), .ZN(n13879) );
  NOR4_X1 U15582 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12380) );
  NOR4_X1 U15583 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12379) );
  NOR4_X1 U15584 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12378) );
  NOR4_X1 U15585 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12377) );
  AND4_X1 U15586 ( .A1(n12380), .A2(n12379), .A3(n12378), .A4(n12377), .ZN(
        n12385) );
  NOR4_X1 U15587 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12383) );
  NOR4_X1 U15588 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12382) );
  NOR4_X1 U15589 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12381) );
  AND4_X1 U15590 ( .A1(n12383), .A2(n12382), .A3(n12381), .A4(n20512), .ZN(
        n12384) );
  NAND2_X1 U15591 ( .A1(n12385), .A2(n12384), .ZN(n12386) );
  NOR2_X2 U15592 ( .A1(n13879), .A2(n16714), .ZN(n19800) );
  INV_X1 U15593 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n12390) );
  INV_X1 U15594 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n12388) );
  NAND2_X1 U15595 ( .A1(n16713), .A2(BUF1_REG_13__SCAN_IN), .ZN(n12387) );
  OAI21_X1 U15596 ( .B1(n16713), .B2(n12388), .A(n12387), .ZN(n14186) );
  AOI22_X1 U15597 ( .A1(n19798), .A2(n14186), .B1(n19813), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n12389) );
  OAI21_X1 U15598 ( .B1(n16077), .B2(n12390), .A(n12389), .ZN(n12391) );
  AOI21_X1 U15599 ( .B1(n19800), .B2(BUF1_REG_29__SCAN_IN), .A(n12391), .ZN(
        n12392) );
  INV_X1 U15600 ( .A(n12393), .ZN(n12394) );
  NAND2_X1 U15601 ( .A1(n12395), .A2(n12394), .ZN(P2_U2890) );
  INV_X1 U15602 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16611) );
  INV_X1 U15603 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12399) );
  AND2_X1 U15604 ( .A1(n16652), .A2(n12400), .ZN(n12411) );
  NAND2_X1 U15605 ( .A1(n12410), .A2(n12411), .ZN(n12397) );
  OR2_X2 U15606 ( .A1(n12397), .A2(n12426), .ZN(n20240) );
  INV_X1 U15607 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12398) );
  INV_X1 U15608 ( .A(n12400), .ZN(n12401) );
  INV_X1 U15609 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12403) );
  INV_X1 U15610 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12405) );
  NOR2_X1 U15611 ( .A1(n12407), .A2(n12406), .ZN(n12437) );
  INV_X1 U15612 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12409) );
  NAND2_X1 U15613 ( .A1(n15847), .A2(n13909), .ZN(n12412) );
  NAND2_X1 U15614 ( .A1(n16665), .A2(n13909), .ZN(n12417) );
  INV_X1 U15615 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12408) );
  INV_X1 U15616 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12414) );
  INV_X1 U15617 ( .A(n12411), .ZN(n12424) );
  INV_X1 U15618 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12413) );
  INV_X1 U15619 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12416) );
  NOR2_X1 U15620 ( .A1(n20388), .A2(n12416), .ZN(n12423) );
  INV_X1 U15621 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12421) );
  INV_X1 U15622 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12420) );
  NOR2_X1 U15623 ( .A1(n12423), .A2(n12422), .ZN(n12435) );
  INV_X1 U15624 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20034) );
  INV_X1 U15625 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12431) );
  INV_X1 U15626 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12430) );
  NOR2_X1 U15627 ( .A1(n12433), .A2(n12432), .ZN(n12434) );
  NAND4_X1 U15628 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12438) );
  NAND2_X1 U15629 ( .A1(n12579), .A2(n19985), .ZN(n12439) );
  INV_X1 U15630 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12441) );
  INV_X1 U15631 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12440) );
  OAI22_X1 U15632 ( .A1(n12441), .A2(n16762), .B1(n20305), .B2(n12440), .ZN(
        n12443) );
  INV_X1 U15633 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n20446) );
  INV_X1 U15634 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12447) );
  INV_X1 U15635 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12444) );
  OAI211_X1 U15636 ( .C1(n12501), .C2(n12447), .A(n12446), .B(n12445), .ZN(
        n12448) );
  INV_X1 U15637 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12450) );
  INV_X1 U15638 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12449) );
  OAI22_X1 U15639 ( .A1(n12450), .A2(n12515), .B1(n19973), .B2(n12449), .ZN(
        n12454) );
  INV_X1 U15640 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12452) );
  INV_X1 U15641 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12451) );
  OAI22_X1 U15642 ( .A1(n12452), .A2(n12516), .B1(n12502), .B2(n12451), .ZN(
        n12453) );
  NOR2_X1 U15643 ( .A1(n12454), .A2(n12453), .ZN(n12467) );
  INV_X1 U15644 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12455) );
  INV_X1 U15645 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12456) );
  INV_X1 U15646 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12460) );
  INV_X1 U15647 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12459) );
  OAI22_X1 U15648 ( .A1(n12460), .A2(n20051), .B1(n20089), .B2(n12459), .ZN(
        n12464) );
  INV_X1 U15649 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12462) );
  INV_X1 U15650 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12461) );
  OAI22_X1 U15651 ( .A1(n12462), .A2(n12499), .B1(n20216), .B2(n12461), .ZN(
        n12463) );
  NOR2_X1 U15652 ( .A1(n12464), .A2(n12463), .ZN(n12465) );
  NAND2_X1 U15653 ( .A1(n12533), .A2(n12563), .ZN(n12532) );
  INV_X1 U15654 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12470) );
  INV_X1 U15655 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12469) );
  OAI22_X1 U15656 ( .A1(n12470), .A2(n16762), .B1(n20240), .B2(n12469), .ZN(
        n12473) );
  INV_X1 U15657 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12471) );
  INV_X1 U15658 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16789) );
  OAI22_X1 U15659 ( .A1(n12471), .A2(n20305), .B1(n16778), .B2(n16789), .ZN(
        n12472) );
  OR2_X1 U15660 ( .A1(n12473), .A2(n12472), .ZN(n12476) );
  INV_X1 U15661 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12474) );
  NOR2_X1 U15662 ( .A1(n16751), .A2(n12474), .ZN(n12475) );
  NOR2_X1 U15663 ( .A1(n12476), .A2(n12475), .ZN(n12496) );
  INV_X1 U15664 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12478) );
  INV_X1 U15665 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12477) );
  OAI22_X1 U15666 ( .A1(n12478), .A2(n12499), .B1(n20089), .B2(n12477), .ZN(
        n12482) );
  INV_X1 U15667 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12480) );
  INV_X1 U15668 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12479) );
  NOR2_X1 U15669 ( .A1(n12482), .A2(n12481), .ZN(n12495) );
  INV_X1 U15670 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12483) );
  INV_X1 U15671 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15989) );
  OAI22_X1 U15672 ( .A1(n12483), .A2(n20051), .B1(n19973), .B2(n15989), .ZN(
        n12487) );
  INV_X1 U15673 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12485) );
  INV_X1 U15674 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12484) );
  OAI22_X1 U15675 ( .A1(n12485), .A2(n12515), .B1(n12502), .B2(n12484), .ZN(
        n12486) );
  NOR2_X1 U15676 ( .A1(n12487), .A2(n12486), .ZN(n12494) );
  INV_X1 U15677 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12488) );
  INV_X1 U15678 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12490) );
  INV_X1 U15679 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12489) );
  OAI22_X1 U15680 ( .A1(n12490), .A2(n12516), .B1(n12501), .B2(n12489), .ZN(
        n12491) );
  NOR2_X1 U15681 ( .A1(n12492), .A2(n12491), .ZN(n12493) );
  NAND4_X1 U15682 ( .A1(n12496), .A2(n12495), .A3(n12494), .A4(n12493), .ZN(
        n12498) );
  NAND2_X1 U15683 ( .A1(n12586), .A2(n19985), .ZN(n12497) );
  INV_X1 U15684 ( .A(n20089), .ZN(n12500) );
  AOI22_X1 U15685 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20021), .B1(
        n12500), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12509) );
  INV_X1 U15686 ( .A(n20051), .ZN(n20055) );
  AOI22_X1 U15687 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20055), .B1(
        n20179), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12508) );
  INV_X1 U15688 ( .A(n19973), .ZN(n19976) );
  INV_X1 U15689 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12504) );
  INV_X1 U15690 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12503) );
  INV_X1 U15691 ( .A(n12505), .ZN(n12506) );
  INV_X1 U15692 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12510) );
  INV_X1 U15693 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16794) );
  OAI22_X1 U15694 ( .A1(n12510), .A2(n16762), .B1(n16778), .B2(n16794), .ZN(
        n12514) );
  INV_X1 U15695 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12512) );
  INV_X1 U15696 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12511) );
  OAI22_X1 U15697 ( .A1(n12512), .A2(n20240), .B1(n20305), .B2(n12511), .ZN(
        n12513) );
  NOR2_X1 U15698 ( .A1(n12514), .A2(n12513), .ZN(n12521) );
  NAND2_X1 U15699 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12519) );
  INV_X1 U15700 ( .A(n20388), .ZN(n20393) );
  NAND2_X1 U15701 ( .A1(n20393), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12518) );
  OAI21_X1 U15702 ( .B1(n16314), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12524) );
  AND2_X1 U15703 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14548) );
  NAND2_X1 U15704 ( .A1(n14548), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16484) );
  INV_X1 U15705 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16481) );
  NOR2_X1 U15706 ( .A1(n16484), .A2(n16481), .ZN(n13583) );
  AND2_X1 U15707 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16527) );
  AND2_X1 U15708 ( .A1(n16527), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13582) );
  NAND2_X1 U15709 ( .A1(n13583), .A2(n13582), .ZN(n16458) );
  NAND2_X1 U15710 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12525) );
  OR2_X1 U15711 ( .A1(n16458), .A2(n12525), .ZN(n13671) );
  NAND2_X1 U15712 ( .A1(n16552), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13669) );
  NOR2_X1 U15713 ( .A1(n13671), .A2(n13669), .ZN(n13674) );
  NAND2_X1 U15714 ( .A1(n13674), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13146) );
  INV_X1 U15715 ( .A(n13146), .ZN(n12526) );
  AND3_X1 U15716 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12552) );
  NAND3_X1 U15717 ( .A1(n12173), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n12530), .ZN(n12531) );
  NOR2_X1 U15718 ( .A1(n13890), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12529) );
  XNOR2_X1 U15719 ( .A(n12530), .B(n12529), .ZN(n13971) );
  NAND2_X1 U15720 ( .A1(n13971), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13973) );
  NAND2_X1 U15721 ( .A1(n12531), .A2(n13973), .ZN(n12534) );
  XNOR2_X1 U15722 ( .A(n13142), .B(n12534), .ZN(n14054) );
  OAI21_X1 U15723 ( .B1(n12533), .B2(n12563), .A(n12532), .ZN(n14053) );
  NAND2_X1 U15724 ( .A1(n14054), .A2(n14053), .ZN(n12536) );
  NAND2_X1 U15725 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12534), .ZN(
        n12535) );
  NAND2_X1 U15726 ( .A1(n12536), .A2(n12535), .ZN(n12537) );
  XNOR2_X1 U15727 ( .A(n12537), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16347) );
  NAND2_X1 U15728 ( .A1(n12537), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12538) );
  INV_X1 U15729 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12786) );
  INV_X1 U15730 ( .A(n12641), .ZN(n12539) );
  NAND2_X1 U15731 ( .A1(n16632), .A2(n16635), .ZN(n12543) );
  NAND3_X1 U15732 ( .A1(n16314), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12544) );
  NAND3_X1 U15733 ( .A1(n16632), .A2(n16635), .A3(n12547), .ZN(n12551) );
  INV_X1 U15734 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16401) );
  INV_X1 U15735 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16377) );
  INV_X1 U15736 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16376) );
  INV_X1 U15737 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16366) );
  NAND2_X1 U15738 ( .A1(n12553), .A2(n12566), .ZN(n12554) );
  NOR2_X1 U15739 ( .A1(n12569), .A2(n12554), .ZN(n12555) );
  NOR2_X1 U15740 ( .A1(n16800), .A2(n12555), .ZN(n12559) );
  AOI21_X1 U15741 ( .B1(n16693), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16803) );
  NAND2_X1 U15742 ( .A1(n12557), .A2(n16803), .ZN(n12558) );
  INV_X1 U15743 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13812) );
  NAND2_X1 U15744 ( .A1(n12558), .A2(n13812), .ZN(n20595) );
  MUX2_X1 U15745 ( .A(n12559), .B(n20595), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n20615) );
  INV_X1 U15746 ( .A(n16816), .ZN(n12560) );
  NAND2_X1 U15747 ( .A1(n12560), .A2(n9576), .ZN(n20614) );
  INV_X1 U15748 ( .A(n20614), .ZN(n12561) );
  NAND2_X1 U15749 ( .A1(n20615), .A2(n12561), .ZN(n12573) );
  INV_X1 U15750 ( .A(n14617), .ZN(n12562) );
  NAND2_X1 U15751 ( .A1(n14621), .A2(n12564), .ZN(n12565) );
  NAND2_X1 U15752 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  NAND2_X1 U15753 ( .A1(n12575), .A2(n12568), .ZN(n12571) );
  INV_X1 U15754 ( .A(n12569), .ZN(n12570) );
  NAND2_X1 U15755 ( .A1(n12571), .A2(n12570), .ZN(n20608) );
  NAND3_X1 U15756 ( .A1(n20609), .A2(n20608), .A3(n12572), .ZN(n13105) );
  NAND2_X1 U15757 ( .A1(n12573), .A2(n13105), .ZN(n12574) );
  INV_X1 U15758 ( .A(n13794), .ZN(n12778) );
  NAND2_X1 U15759 ( .A1(n9575), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n12578) );
  OAI21_X1 U15760 ( .B1(n12693), .B2(n12579), .A(n12578), .ZN(n12645) );
  INV_X1 U15761 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13908) );
  INV_X1 U15762 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14013) );
  NAND2_X1 U15763 ( .A1(n13908), .A2(n14013), .ZN(n12580) );
  NAND2_X1 U15764 ( .A1(n12583), .A2(n12582), .ZN(n12643) );
  NAND2_X1 U15765 ( .A1(n12693), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12584) );
  OAI21_X1 U15766 ( .B1(n12693), .B2(n12585), .A(n12584), .ZN(n12656) );
  NOR2_X2 U15767 ( .A1(n12643), .A2(n12656), .ZN(n12636) );
  INV_X1 U15768 ( .A(n12586), .ZN(n12587) );
  INV_X1 U15769 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14445) );
  MUX2_X1 U15770 ( .A(n12587), .B(n14445), .S(n12693), .Z(n12637) );
  INV_X1 U15771 ( .A(n12588), .ZN(n12589) );
  INV_X1 U15772 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n16001) );
  MUX2_X1 U15773 ( .A(n12589), .B(n16001), .S(n12693), .Z(n12610) );
  INV_X1 U15774 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14456) );
  MUX2_X1 U15775 ( .A(n12590), .B(n14456), .S(n12693), .Z(n12628) );
  INV_X1 U15776 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n15988) );
  NAND2_X1 U15777 ( .A1(n12625), .A2(n15988), .ZN(n12592) );
  NOR2_X2 U15778 ( .A1(n12632), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12620) );
  INV_X1 U15779 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n12593) );
  NAND2_X1 U15780 ( .A1(n12620), .A2(n12593), .ZN(n12685) );
  NAND2_X1 U15781 ( .A1(n12693), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12684) );
  OAI21_X1 U15782 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n12693), .ZN(n12594) );
  OAI21_X1 U15783 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(P2_EBX_REG_16__SCAN_IN), 
        .A(n12693), .ZN(n12595) );
  AND2_X2 U15784 ( .A1(n12698), .A2(n12595), .ZN(n12718) );
  OAI21_X1 U15785 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n12693), .ZN(n12596) );
  INV_X1 U15786 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n12597) );
  NAND2_X1 U15787 ( .A1(n12693), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U15788 ( .A1(n12693), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12745) );
  INV_X1 U15789 ( .A(n12745), .ZN(n12598) );
  NOR2_X2 U15790 ( .A1(n12762), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12755) );
  INV_X1 U15791 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15876) );
  NAND2_X1 U15792 ( .A1(n12755), .A2(n15876), .ZN(n12602) );
  NAND2_X1 U15793 ( .A1(n12602), .A2(n13087), .ZN(n12599) );
  NAND2_X1 U15794 ( .A1(n12693), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12603) );
  NAND2_X1 U15795 ( .A1(n12599), .A2(n12603), .ZN(n12601) );
  INV_X1 U15796 ( .A(n12601), .ZN(n12600) );
  NAND2_X1 U15797 ( .A1(n9575), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12771) );
  AOI21_X1 U15798 ( .B1(n15616), .B2(n12769), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16102) );
  INV_X1 U15799 ( .A(n16102), .ZN(n12607) );
  INV_X1 U15800 ( .A(n12603), .ZN(n12604) );
  NAND2_X1 U15801 ( .A1(n12602), .A2(n12604), .ZN(n12605) );
  NAND2_X1 U15802 ( .A1(n16115), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16100) );
  XNOR2_X1 U15803 ( .A(n12601), .B(n9725), .ZN(n15636) );
  NAND2_X1 U15804 ( .A1(n15636), .A2(n12769), .ZN(n16116) );
  NAND2_X1 U15805 ( .A1(n12607), .A2(n12606), .ZN(n12768) );
  NAND2_X1 U15806 ( .A1(n12609), .A2(n10320), .ZN(n12611) );
  NAND2_X1 U15807 ( .A1(n12608), .A2(n12611), .ZN(n19749) );
  OAI21_X1 U15808 ( .B1(n12615), .B2(n12614), .A(n19749), .ZN(n12612) );
  INV_X1 U15809 ( .A(n12612), .ZN(n12618) );
  INV_X1 U15810 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16624) );
  INV_X1 U15811 ( .A(n12619), .ZN(n12623) );
  NAND3_X1 U15812 ( .A1(n12621), .A2(n12693), .A3(P2_EBX_REG_11__SCAN_IN), 
        .ZN(n12622) );
  NAND2_X1 U15813 ( .A1(n12623), .A2(n12622), .ZN(n19706) );
  OAI21_X1 U15814 ( .B1(n19706), .B2(n12523), .A(n16551), .ZN(n16274) );
  INV_X1 U15815 ( .A(n12625), .ZN(n12626) );
  AND3_X1 U15816 ( .A1(n12626), .A2(n12693), .A3(P2_EBX_REG_8__SCAN_IN), .ZN(
        n12627) );
  NOR2_X1 U15817 ( .A1(n12624), .A2(n12627), .ZN(n19720) );
  NAND2_X1 U15818 ( .A1(n19720), .A2(n12769), .ZN(n12671) );
  NAND2_X1 U15819 ( .A1(n12671), .A2(n16593), .ZN(n16318) );
  XNOR2_X1 U15820 ( .A(n12608), .B(n12591), .ZN(n12673) );
  NAND2_X1 U15821 ( .A1(n12673), .A2(n16611), .ZN(n16330) );
  AND2_X1 U15822 ( .A1(n16318), .A2(n16330), .ZN(n16279) );
  NOR2_X1 U15823 ( .A1(n12624), .A2(n15973), .ZN(n12629) );
  MUX2_X1 U15824 ( .A(n12624), .B(n12629), .S(n12693), .Z(n12631) );
  INV_X1 U15825 ( .A(n12632), .ZN(n12630) );
  INV_X1 U15826 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16577) );
  OAI21_X1 U15827 ( .B1(n15803), .B2(n12523), .A(n16577), .ZN(n16303) );
  NAND2_X1 U15828 ( .A1(n12693), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12633) );
  MUX2_X1 U15829 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n12633), .S(n12632), .Z(
        n12634) );
  NAND2_X1 U15830 ( .A1(n12634), .A2(n12700), .ZN(n15788) );
  OR2_X1 U15831 ( .A1(n15788), .A2(n12523), .ZN(n12635) );
  INV_X1 U15832 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16563) );
  NAND2_X1 U15833 ( .A1(n12635), .A2(n16563), .ZN(n16291) );
  NAND4_X1 U15834 ( .A1(n16274), .A2(n16279), .A3(n16303), .A4(n16291), .ZN(
        n12680) );
  AOI21_X1 U15835 ( .B1(n16277), .B2(n16624), .A(n12680), .ZN(n12670) );
  INV_X1 U15836 ( .A(n12636), .ZN(n12639) );
  INV_X1 U15837 ( .A(n12637), .ZN(n12638) );
  NAND2_X1 U15838 ( .A1(n12639), .A2(n12638), .ZN(n12640) );
  NAND2_X1 U15839 ( .A1(n12609), .A2(n12640), .ZN(n19760) );
  OAI21_X1 U15840 ( .B1(n12641), .B2(n12769), .A(n19760), .ZN(n12642) );
  NAND2_X1 U15841 ( .A1(n12642), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12669) );
  OAI21_X1 U15842 ( .B1(n12644), .B2(n12649), .A(n12645), .ZN(n12646) );
  NAND2_X1 U15843 ( .A1(n12643), .A2(n12646), .ZN(n16349) );
  XNOR2_X1 U15844 ( .A(n12644), .B(n12649), .ZN(n15834) );
  XNOR2_X1 U15845 ( .A(n15834), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14060) );
  AND2_X1 U15846 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n12647) );
  NAND2_X1 U15847 ( .A1(n12693), .A2(n12647), .ZN(n12648) );
  NAND2_X1 U15848 ( .A1(n12649), .A2(n12648), .ZN(n15846) );
  NAND2_X1 U15849 ( .A1(n12721), .A2(n13890), .ZN(n12651) );
  NAND2_X1 U15850 ( .A1(n12693), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12650) );
  NAND2_X1 U15851 ( .A1(n12651), .A2(n12650), .ZN(n15852) );
  NAND2_X1 U15852 ( .A1(n15852), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13968) );
  OAI21_X1 U15853 ( .B1(n15846), .B2(n14633), .A(n13968), .ZN(n12653) );
  NAND2_X1 U15854 ( .A1(n15846), .A2(n14633), .ZN(n12652) );
  AND2_X1 U15855 ( .A1(n12653), .A2(n12652), .ZN(n14059) );
  NAND2_X1 U15856 ( .A1(n14060), .A2(n14059), .ZN(n19935) );
  INV_X1 U15857 ( .A(n15834), .ZN(n12654) );
  NAND2_X1 U15858 ( .A1(n12654), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12655) );
  NAND2_X1 U15859 ( .A1(n19935), .A2(n12655), .ZN(n19920) );
  INV_X1 U15860 ( .A(n12643), .ZN(n12658) );
  INV_X1 U15861 ( .A(n12656), .ZN(n12657) );
  XNOR2_X1 U15862 ( .A(n12658), .B(n12657), .ZN(n19925) );
  INV_X1 U15863 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19954) );
  NAND2_X1 U15864 ( .A1(n19925), .A2(n19954), .ZN(n12663) );
  AND2_X1 U15865 ( .A1(n12663), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12660) );
  INV_X1 U15866 ( .A(n19925), .ZN(n12659) );
  AOI22_X1 U15867 ( .A1(n19920), .A2(n12660), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n12659), .ZN(n12662) );
  AND2_X1 U15868 ( .A1(n16349), .A2(n12662), .ZN(n12661) );
  MUX2_X1 U15869 ( .A(n12786), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .S(
        n19760), .Z(n16629) );
  INV_X1 U15870 ( .A(n12662), .ZN(n12666) );
  OAI21_X1 U15871 ( .B1(n19920), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n12663), .ZN(n12664) );
  INV_X1 U15872 ( .A(n12664), .ZN(n12665) );
  OR2_X1 U15873 ( .A1(n12666), .A2(n12665), .ZN(n16627) );
  AND2_X1 U15874 ( .A1(n16629), .A2(n16627), .ZN(n12667) );
  NAND2_X1 U15875 ( .A1(n16628), .A2(n12667), .ZN(n12668) );
  NAND2_X1 U15876 ( .A1(n12669), .A2(n12668), .ZN(n16275) );
  NOR2_X1 U15877 ( .A1(n12680), .A2(n16624), .ZN(n12682) );
  INV_X1 U15878 ( .A(n12671), .ZN(n12672) );
  NAND2_X1 U15879 ( .A1(n12672), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16319) );
  INV_X1 U15880 ( .A(n12673), .ZN(n19737) );
  NAND2_X1 U15881 ( .A1(n19737), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16328) );
  AND2_X1 U15882 ( .A1(n16319), .A2(n16328), .ZN(n12679) );
  INV_X1 U15883 ( .A(n15803), .ZN(n12675) );
  AND2_X1 U15884 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12674) );
  NAND2_X1 U15885 ( .A1(n12675), .A2(n12674), .ZN(n16302) );
  NAND2_X1 U15886 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12676) );
  OR2_X1 U15887 ( .A1(n15788), .A2(n12676), .ZN(n16290) );
  AND2_X1 U15888 ( .A1(n16302), .A2(n16290), .ZN(n16280) );
  INV_X1 U15889 ( .A(n19706), .ZN(n12678) );
  AND2_X1 U15890 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12677) );
  NAND2_X1 U15891 ( .A1(n12678), .A2(n12677), .ZN(n16273) );
  OAI211_X1 U15892 ( .C1(n12680), .C2(n12679), .A(n16280), .B(n16273), .ZN(
        n12681) );
  NAND2_X1 U15893 ( .A1(n12685), .A2(n10044), .ZN(n12686) );
  NAND2_X1 U15894 ( .A1(n12683), .A2(n12686), .ZN(n12735) );
  NAND2_X1 U15895 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12687) );
  NOR2_X1 U15896 ( .A1(n12735), .A2(n12687), .ZN(n16264) );
  INV_X1 U15897 ( .A(n12688), .ZN(n12690) );
  NAND3_X1 U15898 ( .A1(n9609), .A2(n12693), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n12689) );
  AND2_X1 U15899 ( .A1(n12690), .A2(n12689), .ZN(n12691) );
  INV_X1 U15900 ( .A(n12691), .ZN(n15729) );
  NOR2_X1 U15901 ( .A1(n15729), .A2(n12523), .ZN(n13655) );
  NAND3_X1 U15902 ( .A1(n12691), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n12769), .ZN(n12716) );
  INV_X1 U15903 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n12692) );
  NAND2_X1 U15904 ( .A1(n12698), .A2(n12692), .ZN(n12705) );
  AND2_X1 U15905 ( .A1(n12693), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12694) );
  NAND2_X1 U15906 ( .A1(n12705), .A2(n12694), .ZN(n12695) );
  INV_X1 U15907 ( .A(n12718), .ZN(n12722) );
  NAND2_X1 U15908 ( .A1(n12695), .A2(n12722), .ZN(n15759) );
  NAND2_X1 U15909 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12696) );
  OR2_X1 U15910 ( .A1(n15759), .A2(n12696), .ZN(n13577) );
  INV_X1 U15911 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12697) );
  NAND2_X1 U15912 ( .A1(n12707), .A2(n12697), .ZN(n12713) );
  NAND3_X1 U15913 ( .A1(n12713), .A2(n12693), .A3(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n12699) );
  INV_X1 U15914 ( .A(n12698), .ZN(n12703) );
  NAND2_X1 U15915 ( .A1(n12731), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16232) );
  AND2_X1 U15916 ( .A1(n12693), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12702) );
  INV_X1 U15917 ( .A(n12700), .ZN(n12701) );
  AOI21_X1 U15918 ( .B1(n12703), .B2(n12702), .A(n12701), .ZN(n12704) );
  AND2_X1 U15919 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12706) );
  NAND2_X1 U15920 ( .A1(n19653), .A2(n12706), .ZN(n13575) );
  INV_X1 U15921 ( .A(n12707), .ZN(n12712) );
  NAND2_X1 U15922 ( .A1(n12683), .A2(n10437), .ZN(n12708) );
  NAND2_X1 U15923 ( .A1(n12712), .A2(n12708), .ZN(n15773) );
  NOR2_X1 U15924 ( .A1(n15773), .A2(n12523), .ZN(n12733) );
  NAND2_X1 U15925 ( .A1(n12733), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n16250) );
  AND4_X1 U15926 ( .A1(n13577), .A2(n16232), .A3(n13575), .A4(n16250), .ZN(
        n12715) );
  NAND2_X1 U15927 ( .A1(n12693), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12709) );
  XNOR2_X1 U15928 ( .A(n12719), .B(n12709), .ZN(n12741) );
  AND2_X1 U15929 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12710) );
  NAND2_X1 U15930 ( .A1(n12741), .A2(n12710), .ZN(n16192) );
  NAND2_X1 U15931 ( .A1(n12712), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12711) );
  MUX2_X1 U15932 ( .A(n12712), .B(n12711), .S(n12693), .Z(n12714) );
  NAND2_X1 U15933 ( .A1(n12714), .A2(n12713), .ZN(n19676) );
  NOR2_X1 U15934 ( .A1(n19676), .A2(n12523), .ZN(n12737) );
  NAND2_X1 U15935 ( .A1(n12737), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16238) );
  NAND4_X1 U15936 ( .A1(n12716), .A2(n12715), .A3(n16192), .A4(n16238), .ZN(
        n12728) );
  INV_X1 U15937 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15938 ( .A1(n12718), .A2(n12717), .ZN(n12724) );
  NAND3_X1 U15939 ( .A1(n12724), .A2(n12693), .A3(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n12720) );
  AND2_X1 U15940 ( .A1(n12720), .A2(n12719), .ZN(n19618) );
  NAND2_X1 U15941 ( .A1(n19618), .A2(n12769), .ZN(n13579) );
  INV_X1 U15942 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16474) );
  NAND2_X1 U15943 ( .A1(n12722), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12723) );
  MUX2_X1 U15944 ( .A(n12723), .B(n12722), .S(n12721), .Z(n12725) );
  INV_X1 U15945 ( .A(n19633), .ZN(n12727) );
  AND2_X1 U15946 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U15947 ( .A1(n12727), .A2(n12726), .ZN(n16202) );
  OAI21_X1 U15948 ( .B1(n13579), .B2(n16474), .A(n16202), .ZN(n13649) );
  NAND2_X1 U15949 ( .A1(n19653), .A2(n12769), .ZN(n12729) );
  INV_X1 U15950 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14547) );
  XNOR2_X1 U15951 ( .A(n12729), .B(n14547), .ZN(n16223) );
  INV_X1 U15952 ( .A(n15759), .ZN(n12730) );
  AOI21_X1 U15953 ( .B1(n12730), .B2(n12769), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13576) );
  INV_X1 U15954 ( .A(n12731), .ZN(n12732) );
  NAND2_X1 U15955 ( .A1(n12732), .A2(n14555), .ZN(n16231) );
  INV_X1 U15956 ( .A(n12733), .ZN(n12734) );
  INV_X1 U15957 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16254) );
  NAND2_X1 U15958 ( .A1(n12734), .A2(n16254), .ZN(n16249) );
  INV_X1 U15959 ( .A(n12735), .ZN(n19693) );
  NAND2_X1 U15960 ( .A1(n19693), .A2(n12769), .ZN(n12736) );
  INV_X1 U15961 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16526) );
  NAND2_X1 U15962 ( .A1(n12736), .A2(n16526), .ZN(n16263) );
  NAND4_X1 U15963 ( .A1(n16231), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16249), .A4(n16263), .ZN(n12739) );
  INV_X1 U15964 ( .A(n12737), .ZN(n12738) );
  INV_X1 U15965 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12832) );
  NOR4_X1 U15966 ( .A1(n16223), .A2(n13576), .A3(n12739), .A4(n13574), .ZN(
        n12742) );
  NAND2_X1 U15967 ( .A1(n13579), .A2(n16474), .ZN(n12740) );
  INV_X1 U15968 ( .A(n12741), .ZN(n15742) );
  INV_X1 U15969 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16457) );
  OAI21_X1 U15970 ( .B1(n15742), .B2(n12523), .A(n16457), .ZN(n16193) );
  AND2_X1 U15971 ( .A1(n12742), .A2(n13651), .ZN(n12743) );
  XNOR2_X1 U15972 ( .A(n12744), .B(n12745), .ZN(n15708) );
  NAND2_X1 U15973 ( .A1(n15708), .A2(n12769), .ZN(n12754) );
  XNOR2_X1 U15974 ( .A(n12754), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16173) );
  NAND2_X1 U15975 ( .A1(n12747), .A2(n10041), .ZN(n12748) );
  NAND2_X1 U15976 ( .A1(n12744), .A2(n12748), .ZN(n15717) );
  INV_X1 U15977 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16186) );
  NAND2_X1 U15978 ( .A1(n12753), .A2(n16186), .ZN(n16178) );
  AND2_X1 U15979 ( .A1(n16173), .A2(n16178), .ZN(n12749) );
  AND2_X1 U15980 ( .A1(n12693), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12750) );
  INV_X1 U15981 ( .A(n13087), .ZN(n12760) );
  AOI21_X1 U15982 ( .B1(n12751), .B2(n12750), .A(n12760), .ZN(n12752) );
  AND2_X1 U15983 ( .A1(n12752), .A2(n12762), .ZN(n15692) );
  NAND2_X1 U15984 ( .A1(n12764), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16157) );
  INV_X1 U15985 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21554) );
  OR2_X1 U15986 ( .A1(n12754), .A2(n21554), .ZN(n16137) );
  INV_X1 U15987 ( .A(n12755), .ZN(n12763) );
  NAND3_X1 U15988 ( .A1(n12763), .A2(n12693), .A3(P2_EBX_REG_26__SCAN_IN), 
        .ZN(n12756) );
  NAND3_X1 U15989 ( .A1(n12602), .A2(n12756), .A3(n13087), .ZN(n15654) );
  INV_X1 U15990 ( .A(n15654), .ZN(n12758) );
  INV_X1 U15991 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16399) );
  OAI21_X1 U15992 ( .B1(n15654), .B2(n12523), .A(n16399), .ZN(n12759) );
  AND2_X1 U15993 ( .A1(n12693), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12761) );
  NOR2_X1 U15994 ( .A1(n16139), .A2(n12765), .ZN(n12766) );
  NAND2_X1 U15995 ( .A1(n16376), .A2(n16377), .ZN(n16098) );
  INV_X1 U15996 ( .A(n16116), .ZN(n16097) );
  INV_X1 U15997 ( .A(n15671), .ZN(n12767) );
  NAND3_X1 U15998 ( .A1(n12767), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n12769), .ZN(n16148) );
  NAND2_X1 U15999 ( .A1(n16113), .A2(n16148), .ZN(n16099) );
  AND2_X1 U16000 ( .A1(n12769), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12770) );
  NAND2_X1 U16001 ( .A1(n15616), .A2(n12770), .ZN(n16101) );
  NAND2_X1 U16002 ( .A1(n13084), .A2(n16101), .ZN(n12777) );
  NAND2_X1 U16003 ( .A1(n12693), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12774) );
  INV_X1 U16004 ( .A(n12771), .ZN(n12772) );
  AOI21_X1 U16005 ( .B1(n14692), .B2(n12590), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13083) );
  INV_X1 U16006 ( .A(n13083), .ZN(n12775) );
  NAND3_X1 U16007 ( .A1(n14692), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12590), .ZN(n13079) );
  NAND2_X1 U16008 ( .A1(n12775), .A2(n13079), .ZN(n12776) );
  NAND2_X1 U16009 ( .A1(n9583), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12781) );
  NAND2_X1 U16010 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12780) );
  OAI211_X1 U16011 ( .C1(n12792), .C2(n20516), .A(n12781), .B(n12780), .ZN(
        n12782) );
  INV_X1 U16012 ( .A(n12782), .ZN(n12785) );
  OR2_X1 U16013 ( .A1(n12843), .A2(n16624), .ZN(n12784) );
  OR2_X1 U16014 ( .A1(n12843), .A2(n12786), .ZN(n12791) );
  INV_X1 U16015 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19759) );
  NAND2_X1 U16016 ( .A1(n9583), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U16017 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12787) );
  OAI211_X1 U16018 ( .C1(n12792), .C2(n19759), .A(n12788), .B(n12787), .ZN(
        n12789) );
  INV_X1 U16019 ( .A(n12789), .ZN(n12790) );
  OR2_X1 U16020 ( .A1(n12843), .A2(n16611), .ZN(n12794) );
  AOI22_X1 U16021 ( .A1(n12879), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12793) );
  OAI211_X1 U16022 ( .C1(n12792), .C2(n20518), .A(n12794), .B(n12793), .ZN(
        n14455) );
  OR2_X1 U16023 ( .A1(n12843), .A2(n16593), .ZN(n12797) );
  INV_X1 U16024 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n20520) );
  NAND2_X1 U16025 ( .A1(n9583), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12796) );
  NAND2_X1 U16026 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12795) );
  AND2_X1 U16027 ( .A1(n12797), .A2(n9684), .ZN(n15982) );
  INV_X1 U16028 ( .A(n15982), .ZN(n12798) );
  AND2_X2 U16029 ( .A1(n14454), .A2(n12798), .ZN(n15792) );
  OR2_X1 U16030 ( .A1(n12843), .A2(n16577), .ZN(n12803) );
  INV_X1 U16031 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n16306) );
  NAND2_X1 U16032 ( .A1(n12879), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12800) );
  NAND2_X1 U16033 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12799) );
  OAI211_X1 U16034 ( .C1(n12792), .C2(n16306), .A(n12800), .B(n12799), .ZN(
        n12801) );
  INV_X1 U16035 ( .A(n12801), .ZN(n12802) );
  AND2_X1 U16036 ( .A1(n12803), .A2(n12802), .ZN(n15793) );
  INV_X1 U16037 ( .A(n15793), .ZN(n12804) );
  INV_X1 U16038 ( .A(n12805), .ZN(n12807) );
  NAND2_X1 U16039 ( .A1(n12807), .A2(n12806), .ZN(n14375) );
  OR2_X1 U16040 ( .A1(n12843), .A2(n19954), .ZN(n12812) );
  INV_X1 U16041 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19915) );
  NAND2_X1 U16042 ( .A1(n9583), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U16043 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12808) );
  OAI211_X1 U16044 ( .C1(n12792), .C2(n19915), .A(n12809), .B(n12808), .ZN(
        n12810) );
  INV_X1 U16045 ( .A(n12810), .ZN(n12811) );
  OR2_X1 U16046 ( .A1(n12843), .A2(n16563), .ZN(n12817) );
  INV_X1 U16047 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n20523) );
  NAND2_X1 U16048 ( .A1(n9583), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U16049 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12813) );
  OAI211_X1 U16050 ( .C1(n12792), .C2(n20523), .A(n12814), .B(n12813), .ZN(
        n12815) );
  INV_X1 U16051 ( .A(n12815), .ZN(n12816) );
  AND2_X1 U16052 ( .A1(n12817), .A2(n12816), .ZN(n15778) );
  OR2_X1 U16053 ( .A1(n12843), .A2(n16551), .ZN(n12819) );
  AOI22_X1 U16054 ( .A1(n12879), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12818) );
  OAI211_X1 U16055 ( .C1(n12792), .C2(n19703), .A(n12819), .B(n12818), .ZN(
        n15962) );
  INV_X1 U16056 ( .A(n15948), .ZN(n12826) );
  OR2_X1 U16057 ( .A1(n12843), .A2(n16526), .ZN(n12824) );
  INV_X1 U16058 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n20526) );
  NAND2_X1 U16059 ( .A1(n9583), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12821) );
  NAND2_X1 U16060 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12820) );
  OAI211_X1 U16061 ( .C1(n12792), .C2(n20526), .A(n12821), .B(n12820), .ZN(
        n12822) );
  INV_X1 U16062 ( .A(n12822), .ZN(n12823) );
  NAND2_X1 U16063 ( .A1(n12826), .A2(n12825), .ZN(n15762) );
  OR2_X1 U16064 ( .A1(n12843), .A2(n16254), .ZN(n12831) );
  INV_X1 U16065 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15767) );
  NAND2_X1 U16066 ( .A1(n12879), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U16067 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12827) );
  OAI211_X1 U16068 ( .C1(n12792), .C2(n15767), .A(n12828), .B(n12827), .ZN(
        n12829) );
  INV_X1 U16069 ( .A(n12829), .ZN(n12830) );
  OR2_X1 U16070 ( .A1(n12843), .A2(n12832), .ZN(n12834) );
  AOI22_X1 U16071 ( .A1(n9583), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12833) );
  OAI211_X1 U16072 ( .C1(n12792), .C2(n20529), .A(n12834), .B(n12833), .ZN(
        n15938) );
  OR2_X1 U16073 ( .A1(n12843), .A2(n14555), .ZN(n12837) );
  INV_X1 U16074 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20531) );
  NAND2_X1 U16075 ( .A1(n9583), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12836) );
  NAND2_X1 U16076 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12835) );
  OR2_X1 U16077 ( .A1(n12843), .A2(n14547), .ZN(n12841) );
  INV_X1 U16078 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20533) );
  NAND2_X1 U16079 ( .A1(n9583), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U16080 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12839) );
  INV_X1 U16081 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12842) );
  OR2_X1 U16082 ( .A1(n12843), .A2(n12842), .ZN(n12845) );
  AOI22_X1 U16083 ( .A1(n12879), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12844) );
  OR2_X1 U16084 ( .A1(n12887), .A2(n16481), .ZN(n12847) );
  AOI22_X1 U16085 ( .A1(n9583), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n12846) );
  NAND2_X1 U16086 ( .A1(n14567), .A2(n15915), .ZN(n13587) );
  OR2_X1 U16087 ( .A1(n12887), .A2(n16474), .ZN(n12852) );
  INV_X1 U16088 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20538) );
  NAND2_X1 U16089 ( .A1(n12879), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12849) );
  NAND2_X1 U16090 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12848) );
  OAI211_X1 U16091 ( .C1(n12792), .C2(n20538), .A(n12849), .B(n12848), .ZN(
        n12850) );
  INV_X1 U16092 ( .A(n12850), .ZN(n12851) );
  NAND2_X1 U16093 ( .A1(n12854), .A2(n12853), .ZN(n13585) );
  OR2_X1 U16094 ( .A1(n12887), .A2(n16457), .ZN(n12857) );
  INV_X1 U16095 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20540) );
  NAND2_X1 U16096 ( .A1(n12879), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12856) );
  NAND2_X1 U16097 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12855) );
  INV_X1 U16098 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13672) );
  OR2_X1 U16099 ( .A1(n12887), .A2(n13672), .ZN(n12860) );
  INV_X1 U16100 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20542) );
  NAND2_X1 U16101 ( .A1(n12879), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U16102 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12858) );
  OR2_X1 U16103 ( .A1(n12887), .A2(n16186), .ZN(n12862) );
  AOI22_X1 U16104 ( .A1(n12879), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n12861) );
  OAI211_X1 U16105 ( .C1(n12792), .C2(n20544), .A(n12862), .B(n12861), .ZN(
        n15713) );
  INV_X1 U16106 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20546) );
  OR2_X1 U16107 ( .A1(n12887), .A2(n21554), .ZN(n12864) );
  AOI22_X1 U16108 ( .A1(n9583), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12863) );
  INV_X1 U16109 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16419) );
  OR2_X1 U16110 ( .A1(n12887), .A2(n16419), .ZN(n12869) );
  INV_X1 U16111 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20548) );
  NAND2_X1 U16112 ( .A1(n9583), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12866) );
  NAND2_X1 U16113 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12865) );
  INV_X1 U16114 ( .A(n12867), .ZN(n12868) );
  OR2_X1 U16115 ( .A1(n12887), .A2(n16401), .ZN(n12874) );
  NAND2_X1 U16116 ( .A1(n9582), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12871) );
  NAND2_X1 U16117 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12870) );
  INV_X1 U16118 ( .A(n12872), .ZN(n12873) );
  NOR2_X2 U16119 ( .A1(n15683), .A2(n15663), .ZN(n15649) );
  INV_X1 U16120 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n16142) );
  OR2_X1 U16121 ( .A1(n12887), .A2(n16399), .ZN(n12876) );
  AOI22_X1 U16122 ( .A1(n9582), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n12875) );
  OAI211_X1 U16123 ( .C1(n12792), .C2(n16142), .A(n12876), .B(n12875), .ZN(
        n15648) );
  INV_X1 U16124 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20554) );
  OR2_X1 U16125 ( .A1(n12887), .A2(n16377), .ZN(n12878) );
  AOI22_X1 U16126 ( .A1(n12879), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12877) );
  OR2_X1 U16127 ( .A1(n12887), .A2(n16376), .ZN(n12884) );
  NAND2_X1 U16128 ( .A1(n9583), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U16129 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12880) );
  INV_X1 U16130 ( .A(n12882), .ZN(n12883) );
  AOI22_X1 U16131 ( .A1(n12879), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n12885) );
  AOI21_X1 U16132 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n13070), .A(
        n12886), .ZN(n13682) );
  INV_X1 U16133 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20559) );
  INV_X1 U16134 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13635) );
  OR2_X1 U16135 ( .A1(n12887), .A2(n13635), .ZN(n12889) );
  AOI22_X1 U16136 ( .A1(n9583), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12888) );
  NOR2_X1 U16137 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20579) );
  OR2_X1 U16138 ( .A1(n20382), .A2(n20579), .ZN(n20600) );
  NAND2_X1 U16139 ( .A1(n20600), .A2(n16837), .ZN(n12890) );
  NOR2_X1 U16140 ( .A1(n13787), .A2(n19970), .ZN(n14146) );
  NOR2_X2 U16141 ( .A1(n14634), .A2(n19934), .ZN(n14637) );
  NOR2_X2 U16142 ( .A1(n14628), .A2(n16296), .ZN(n14627) );
  INV_X1 U16143 ( .A(n14627), .ZN(n14629) );
  NOR2_X2 U16144 ( .A1(n14644), .A2(n16257), .ZN(n14643) );
  AND2_X1 U16145 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12892) );
  NOR2_X2 U16146 ( .A1(n14664), .A2(n16169), .ZN(n14667) );
  INV_X1 U16147 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12893) );
  INV_X1 U16148 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15643) );
  AND2_X2 U16149 ( .A1(n14675), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14677) );
  XNOR2_X1 U16150 ( .A(n14677), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14701) );
  NAND2_X1 U16151 ( .A1(n19970), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14679) );
  NAND2_X1 U16152 ( .A1(n12894), .A2(n14679), .ZN(n13903) );
  INV_X2 U16153 ( .A(n16341), .ZN(n19701) );
  NOR2_X1 U16154 ( .A1(n19701), .A2(n20559), .ZN(n13158) );
  AOI21_X1 U16155 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n13158), .ZN(n12895) );
  OAI21_X1 U16156 ( .B1(n14701), .B2(n19939), .A(n12895), .ZN(n12896) );
  INV_X1 U16157 ( .A(n12896), .ZN(n12897) );
  INV_X1 U16158 ( .A(n13738), .ZN(n12899) );
  NAND3_X1 U16159 ( .A1(n14037), .A2(n15595), .A3(n20819), .ZN(n12914) );
  INV_X1 U16160 ( .A(n12901), .ZN(n13866) );
  NAND2_X1 U16161 ( .A1(n12902), .A2(n20819), .ZN(n13041) );
  AND2_X1 U16162 ( .A1(n13041), .A2(n14511), .ZN(n12903) );
  NAND2_X1 U16163 ( .A1(n12904), .A2(n12903), .ZN(n13033) );
  NAND2_X1 U16164 ( .A1(n9635), .A2(n13033), .ZN(n12905) );
  NAND2_X1 U16165 ( .A1(n13866), .A2(n12905), .ZN(n13941) );
  AND3_X1 U16166 ( .A1(n12909), .A2(n12908), .A3(n12907), .ZN(n12912) );
  AOI21_X1 U16167 ( .B1(n12912), .B2(n12911), .A(n12910), .ZN(n13867) );
  AND2_X1 U16168 ( .A1(n13867), .A2(n21419), .ZN(n13600) );
  OAI211_X1 U16169 ( .C1(n14140), .C2(n17186), .A(n20824), .B(n13600), .ZN(
        n12913) );
  NAND3_X1 U16170 ( .A1(n12914), .A2(n13941), .A3(n12913), .ZN(n12915) );
  NAND2_X1 U16171 ( .A1(n12915), .A2(n14043), .ZN(n12919) );
  INV_X1 U16172 ( .A(n13936), .ZN(n13915) );
  NOR2_X1 U16173 ( .A1(n13915), .A2(n21501), .ZN(n13597) );
  INV_X1 U16174 ( .A(n17186), .ZN(n21498) );
  NAND2_X1 U16175 ( .A1(n14140), .A2(n21498), .ZN(n13712) );
  NAND2_X1 U16176 ( .A1(n13028), .A2(n14511), .ZN(n12916) );
  AOI21_X1 U16177 ( .B1(n13597), .B2(n13712), .A(n12916), .ZN(n12917) );
  INV_X1 U16178 ( .A(n12921), .ZN(n17271) );
  NAND2_X1 U16179 ( .A1(n9635), .A2(n13862), .ZN(n13922) );
  AND2_X1 U16180 ( .A1(n13922), .A2(n12922), .ZN(n13864) );
  INV_X1 U16181 ( .A(n13023), .ZN(n12923) );
  NAND2_X1 U16182 ( .A1(n12923), .A2(n20833), .ZN(n12924) );
  NAND4_X1 U16183 ( .A1(n17271), .A2(n13864), .A3(n12925), .A4(n12924), .ZN(
        n12926) );
  OR2_X1 U16184 ( .A1(n14733), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12929) );
  INV_X1 U16185 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12930) );
  NAND2_X1 U16186 ( .A1(n12959), .A2(n12930), .ZN(n12928) );
  NAND2_X1 U16187 ( .A1(n12929), .A2(n12928), .ZN(n13698) );
  NAND2_X1 U16188 ( .A1(n12951), .A2(n12930), .ZN(n12931) );
  OAI21_X1 U16189 ( .B1(n13698), .B2(n12951), .A(n12931), .ZN(n13696) );
  INV_X1 U16190 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12933) );
  INV_X1 U16191 ( .A(n12969), .ZN(n12941) );
  NAND2_X1 U16192 ( .A1(n12941), .A2(n12933), .ZN(n12934) );
  OAI211_X1 U16193 ( .C1(n12932), .C2(n14473), .A(n12934), .B(n12999), .ZN(
        n12935) );
  NAND2_X1 U16194 ( .A1(n12936), .A2(n12935), .ZN(n12939) );
  INV_X1 U16195 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n12938) );
  NAND2_X1 U16196 ( .A1(n12932), .A2(n12938), .ZN(n12937) );
  OAI21_X1 U16197 ( .B1(n12999), .B2(n12938), .A(n12937), .ZN(n14035) );
  XNOR2_X1 U16198 ( .A(n12939), .B(n14035), .ZN(n14073) );
  INV_X1 U16199 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12940) );
  NAND2_X1 U16200 ( .A1(n12995), .A2(n12940), .ZN(n12944) );
  INV_X1 U16201 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20812) );
  NAND2_X1 U16202 ( .A1(n12941), .A2(n12940), .ZN(n12942) );
  OAI211_X1 U16203 ( .C1(n12951), .C2(n20812), .A(n12942), .B(n12999), .ZN(
        n12943) );
  AND2_X1 U16204 ( .A1(n12944), .A2(n12943), .ZN(n14255) );
  INV_X1 U16205 ( .A(n12945), .ZN(n13017) );
  MUX2_X1 U16206 ( .A(n12951), .B(n13017), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12948) );
  INV_X1 U16207 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12946) );
  NOR2_X1 U16208 ( .A1(n12959), .A2(n12946), .ZN(n12947) );
  NOR2_X1 U16209 ( .A1(n12948), .A2(n12947), .ZN(n14462) );
  MUX2_X1 U16210 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12949) );
  OAI21_X1 U16211 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n14733), .A(
        n12949), .ZN(n14461) );
  NOR2_X1 U16212 ( .A1(n14462), .A2(n14461), .ZN(n12950) );
  MUX2_X1 U16214 ( .A(n12951), .B(n13017), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n12953) );
  NOR2_X1 U16215 ( .A1(n12959), .A2(n13037), .ZN(n12952) );
  NOR2_X1 U16216 ( .A1(n12953), .A2(n12952), .ZN(n14479) );
  INV_X1 U16217 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n15103) );
  NAND2_X1 U16218 ( .A1(n12959), .A2(n15103), .ZN(n12956) );
  OAI211_X1 U16219 ( .C1(n12951), .C2(n17237), .A(n12956), .B(n12999), .ZN(
        n12957) );
  OAI21_X1 U16220 ( .B1(n13020), .B2(P1_EBX_REG_6__SCAN_IN), .A(n12957), .ZN(
        n15101) );
  INV_X1 U16221 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U16222 ( .A1(n12995), .A2(n15088), .ZN(n12962) );
  NAND2_X1 U16223 ( .A1(n12959), .A2(n15088), .ZN(n12960) );
  OAI211_X1 U16224 ( .C1(n12951), .C2(n11592), .A(n12960), .B(n12999), .ZN(
        n12961) );
  AND2_X1 U16225 ( .A1(n12962), .A2(n12961), .ZN(n14977) );
  MUX2_X1 U16226 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n12964) );
  NAND2_X1 U16227 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12963) );
  NAND2_X1 U16228 ( .A1(n12964), .A2(n12963), .ZN(n15095) );
  MUX2_X1 U16229 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12966) );
  NAND2_X1 U16230 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12965) );
  NAND2_X1 U16231 ( .A1(n12966), .A2(n12965), .ZN(n15083) );
  NAND2_X1 U16232 ( .A1(n15084), .A2(n15083), .ZN(n15086) );
  MUX2_X1 U16233 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n12967) );
  OAI21_X1 U16234 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n14733), .A(
        n12967), .ZN(n14962) );
  NAND2_X1 U16235 ( .A1(n12999), .A2(n15548), .ZN(n12971) );
  INV_X1 U16236 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n17215) );
  NAND2_X1 U16237 ( .A1(n12959), .A2(n17215), .ZN(n12970) );
  NAND3_X1 U16238 ( .A1(n12971), .A2(n14731), .A3(n12970), .ZN(n12973) );
  NAND2_X1 U16239 ( .A1(n12932), .A2(n17215), .ZN(n12972) );
  INV_X1 U16240 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15070) );
  NAND2_X1 U16241 ( .A1(n12995), .A2(n15070), .ZN(n12976) );
  NAND2_X1 U16242 ( .A1(n12959), .A2(n15070), .ZN(n12974) );
  OAI211_X1 U16243 ( .C1(n12951), .C2(n15531), .A(n12974), .B(n12999), .ZN(
        n12975) );
  MUX2_X1 U16244 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12978) );
  NAND2_X1 U16245 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12977) );
  NAND2_X1 U16246 ( .A1(n12978), .A2(n12977), .ZN(n14930) );
  INV_X1 U16247 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U16248 ( .A1(n12959), .A2(n17204), .ZN(n12979) );
  OAI211_X1 U16249 ( .C1(n12951), .C2(n15475), .A(n12979), .B(n12999), .ZN(
        n12980) );
  OAI21_X1 U16250 ( .B1(n13020), .B2(P1_EBX_REG_14__SCAN_IN), .A(n12980), .ZN(
        n15064) );
  MUX2_X1 U16251 ( .A(n12951), .B(n13017), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12982) );
  NOR2_X1 U16252 ( .A1(n12959), .A2(n15492), .ZN(n12981) );
  NOR2_X1 U16253 ( .A1(n12982), .A2(n12981), .ZN(n15052) );
  INV_X1 U16254 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n12983) );
  NAND2_X1 U16255 ( .A1(n12959), .A2(n12983), .ZN(n12984) );
  OAI211_X1 U16256 ( .C1(n12951), .C2(n15493), .A(n12984), .B(n12999), .ZN(
        n12985) );
  OAI21_X1 U16257 ( .B1(n13020), .B2(P1_EBX_REG_16__SCAN_IN), .A(n12985), .ZN(
        n14913) );
  MUX2_X1 U16258 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12988) );
  NAND2_X1 U16259 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12987) );
  NAND2_X1 U16260 ( .A1(n12988), .A2(n12987), .ZN(n14898) );
  MUX2_X1 U16261 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n12989) );
  OAI21_X1 U16262 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14733), .A(
        n12989), .ZN(n14891) );
  INV_X1 U16263 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15451) );
  NAND2_X1 U16264 ( .A1(n12999), .A2(n15451), .ZN(n12991) );
  INV_X1 U16265 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n12992) );
  NAND2_X1 U16266 ( .A1(n12959), .A2(n12992), .ZN(n12990) );
  NAND3_X1 U16267 ( .A1(n12991), .A2(n14731), .A3(n12990), .ZN(n12994) );
  NAND2_X1 U16268 ( .A1(n12932), .A2(n12992), .ZN(n12993) );
  INV_X1 U16269 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15045) );
  NAND2_X1 U16270 ( .A1(n12995), .A2(n15045), .ZN(n12998) );
  NAND2_X1 U16271 ( .A1(n12959), .A2(n15045), .ZN(n12996) );
  OAI211_X1 U16272 ( .C1(n12951), .C2(n10899), .A(n12996), .B(n12999), .ZN(
        n12997) );
  MUX2_X1 U16273 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13001) );
  NAND2_X1 U16274 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13000) );
  NAND2_X1 U16275 ( .A1(n13001), .A2(n13000), .ZN(n14844) );
  MUX2_X1 U16276 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13002) );
  OAI21_X1 U16277 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14733), .A(
        n13002), .ZN(n14828) );
  NAND2_X1 U16278 ( .A1(n12999), .A2(n15416), .ZN(n13004) );
  INV_X1 U16279 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n13005) );
  NAND2_X1 U16280 ( .A1(n12959), .A2(n13005), .ZN(n13003) );
  NAND3_X1 U16281 ( .A1(n13004), .A2(n14731), .A3(n13003), .ZN(n13007) );
  NAND2_X1 U16282 ( .A1(n12951), .A2(n13005), .ZN(n13006) );
  INV_X1 U16283 ( .A(n14816), .ZN(n13008) );
  MUX2_X1 U16284 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n13009) );
  OAI21_X1 U16285 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14733), .A(
        n13009), .ZN(n13010) );
  INV_X1 U16286 ( .A(n13010), .ZN(n14798) );
  MUX2_X1 U16287 ( .A(n14731), .B(n12999), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n13012) );
  NAND2_X1 U16288 ( .A1(n12969), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13011) );
  NAND2_X1 U16289 ( .A1(n13012), .A2(n13011), .ZN(n14794) );
  INV_X1 U16290 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n13013) );
  NAND2_X1 U16291 ( .A1(n12959), .A2(n13013), .ZN(n13014) );
  OAI211_X1 U16292 ( .C1(n12951), .C2(n13015), .A(n13014), .B(n12999), .ZN(
        n13016) );
  OAI21_X1 U16293 ( .B1(n13020), .B2(P1_EBX_REG_26__SCAN_IN), .A(n13016), .ZN(
        n14774) );
  MUX2_X1 U16294 ( .A(n12951), .B(n13017), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13019) );
  INV_X1 U16295 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15383) );
  NOR2_X1 U16296 ( .A1(n12959), .A2(n15383), .ZN(n13018) );
  NOR2_X1 U16297 ( .A1(n13019), .A2(n13018), .ZN(n14760) );
  MUX2_X1 U16298 ( .A(n13020), .B(n14731), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13021) );
  OAI21_X1 U16299 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14733), .A(
        n13021), .ZN(n13626) );
  XOR2_X1 U16300 ( .A(n13696), .B(n13697), .Z(n14724) );
  OAI22_X1 U16301 ( .A1(n13022), .A2(n20819), .B1(n13023), .B2(n20833), .ZN(
        n13024) );
  AND2_X2 U16302 ( .A1(n13044), .A2(n13024), .ZN(n20801) );
  AND2_X1 U16303 ( .A1(n12901), .A2(n20819), .ZN(n17140) );
  INV_X1 U16304 ( .A(n13862), .ZN(n14990) );
  INV_X1 U16305 ( .A(n13026), .ZN(n13032) );
  INV_X1 U16306 ( .A(n15003), .ZN(n13027) );
  OAI21_X1 U16307 ( .B1(n14039), .B2(n10602), .A(n13027), .ZN(n13030) );
  OAI21_X1 U16308 ( .B1(n13028), .B2(n14511), .A(n20824), .ZN(n13029) );
  AND2_X1 U16309 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  OAI211_X1 U16310 ( .C1(n13025), .C2(n14990), .A(n9669), .B(n13033), .ZN(
        n13917) );
  OAI21_X1 U16311 ( .B1(n13913), .B2(n14511), .A(n13034), .ZN(n13035) );
  OR2_X1 U16312 ( .A1(n13917), .A2(n13035), .ZN(n13036) );
  NAND2_X1 U16313 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20785) );
  OR2_X1 U16314 ( .A1(n13037), .A2(n20785), .ZN(n15529) );
  NOR3_X1 U16315 ( .A1(n20812), .A2(n14473), .A3(n15529), .ZN(n15553) );
  INV_X1 U16316 ( .A(n15553), .ZN(n13038) );
  AND2_X1 U16317 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15563) );
  NOR3_X1 U16318 ( .A1(n11592), .A2(n17251), .A3(n17237), .ZN(n15562) );
  NAND2_X1 U16319 ( .A1(n15563), .A2(n15562), .ZN(n15530) );
  NOR2_X1 U16320 ( .A1(n13038), .A2(n15530), .ZN(n15534) );
  AND2_X1 U16321 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13039) );
  NAND2_X1 U16322 ( .A1(n15534), .A2(n13039), .ZN(n15464) );
  AOI21_X1 U16323 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14472) );
  NOR2_X1 U16324 ( .A1(n14472), .A2(n15529), .ZN(n15554) );
  NOR2_X1 U16325 ( .A1(n15530), .A2(n15548), .ZN(n13042) );
  NAND2_X1 U16326 ( .A1(n15554), .A2(n13042), .ZN(n15532) );
  OR2_X1 U16327 ( .A1(n15532), .A2(n15531), .ZN(n13056) );
  NAND2_X1 U16328 ( .A1(n20805), .A2(n13056), .ZN(n13043) );
  NAND2_X1 U16329 ( .A1(n15428), .A2(n15426), .ZN(n13046) );
  OR2_X1 U16330 ( .A1(n13044), .A2(n20786), .ZN(n13045) );
  NAND2_X1 U16331 ( .A1(n13046), .A2(n13045), .ZN(n15533) );
  NOR2_X1 U16332 ( .A1(n13047), .A2(n15533), .ZN(n15521) );
  INV_X1 U16333 ( .A(n20805), .ZN(n15537) );
  NAND3_X1 U16334 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15477) );
  NAND2_X1 U16335 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n13048) );
  NOR2_X1 U16336 ( .A1(n15477), .A2(n13048), .ZN(n13060) );
  NAND2_X1 U16337 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n13060), .ZN(
        n15465) );
  NAND2_X1 U16338 ( .A1(n15580), .A2(n15465), .ZN(n13049) );
  NAND2_X1 U16339 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n13058) );
  AND2_X1 U16340 ( .A1(n15580), .A2(n13058), .ZN(n13050) );
  NOR2_X1 U16341 ( .A1(n15446), .A2(n13050), .ZN(n15417) );
  NAND2_X1 U16342 ( .A1(n20805), .A2(n15416), .ZN(n13051) );
  AOI22_X1 U16343 ( .A1(n20811), .A2(n15218), .B1(n20805), .B2(n13621), .ZN(
        n13052) );
  NAND2_X1 U16344 ( .A1(n15389), .A2(n17255), .ZN(n15368) );
  NAND2_X1 U16345 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15390) );
  NAND2_X1 U16346 ( .A1(n15580), .A2(n15390), .ZN(n13053) );
  NOR2_X1 U16347 ( .A1(n13742), .A2(n13054), .ZN(n13064) );
  NOR2_X1 U16348 ( .A1(n15464), .A2(n10879), .ZN(n13055) );
  NAND2_X1 U16349 ( .A1(n15539), .A2(n13055), .ZN(n15409) );
  INV_X1 U16350 ( .A(n13056), .ZN(n15425) );
  NAND3_X1 U16351 ( .A1(n20805), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15425), .ZN(n13057) );
  NAND2_X1 U16352 ( .A1(n15409), .A2(n13057), .ZN(n15513) );
  NOR2_X1 U16353 ( .A1(n15433), .A2(n13058), .ZN(n13059) );
  AND2_X1 U16354 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  NAND2_X1 U16355 ( .A1(n15513), .A2(n13061), .ZN(n15419) );
  NOR2_X1 U16356 ( .A1(n15400), .A2(n15390), .ZN(n15381) );
  INV_X1 U16357 ( .A(n13062), .ZN(n13627) );
  NAND2_X1 U16358 ( .A1(n15381), .A2(n13627), .ZN(n15374) );
  NAND2_X1 U16359 ( .A1(n20786), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n13751) );
  OAI21_X1 U16360 ( .B1(n15374), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13751), .ZN(n13063) );
  AOI211_X1 U16361 ( .C1(n14724), .C2(n20801), .A(n13064), .B(n13063), .ZN(
        n13065) );
  NAND2_X1 U16362 ( .A1(n13681), .A2(n13067), .ZN(n13072) );
  INV_X1 U16363 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20561) );
  AOI22_X1 U16364 ( .A1(n9582), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13068) );
  AOI21_X1 U16365 ( .B1(n13070), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13069), .ZN(n13071) );
  NAND2_X1 U16366 ( .A1(n14677), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13074) );
  INV_X1 U16367 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13073) );
  NOR2_X1 U16368 ( .A1(n19701), .A2(n20561), .ZN(n13637) );
  AOI21_X1 U16369 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13637), .ZN(n13075) );
  OAI21_X1 U16370 ( .B1(n14623), .B2(n19939), .A(n13075), .ZN(n13076) );
  INV_X1 U16371 ( .A(n13076), .ZN(n13077) );
  OAI21_X1 U16372 ( .B1(n14696), .B2(n19928), .A(n13077), .ZN(n13078) );
  INV_X1 U16373 ( .A(n13085), .ZN(n13086) );
  OAI21_X1 U16374 ( .B1(n13086), .B2(P2_EBX_REG_30__SCAN_IN), .A(n9575), .ZN(
        n13088) );
  NAND2_X1 U16375 ( .A1(n13088), .A2(n13087), .ZN(n14705) );
  NOR2_X1 U16376 ( .A1(n14705), .A2(n12523), .ZN(n13089) );
  XNOR2_X1 U16377 ( .A(n13089), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13090) );
  XNOR2_X1 U16378 ( .A(n13091), .B(n13090), .ZN(n13645) );
  OAI211_X1 U16379 ( .C1(n13648), .C2(n19941), .A(n13093), .B(n13092), .ZN(
        P2_U2983) );
  NOR2_X1 U16380 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20490) );
  INV_X1 U16381 ( .A(n20490), .ZN(n20501) );
  NAND2_X1 U16382 ( .A1(n20495), .A2(n20480), .ZN(n14616) );
  INV_X1 U16383 ( .A(n14616), .ZN(n13790) );
  NAND2_X1 U16384 ( .A1(n13123), .A2(n13790), .ZN(n13109) );
  AOI21_X1 U16385 ( .B1(n13094), .B2(n16815), .A(n20003), .ZN(n13107) );
  NAND2_X1 U16386 ( .A1(n13786), .A2(n13790), .ZN(n13097) );
  OAI21_X1 U16387 ( .B1(n13095), .B2(n13097), .A(n13096), .ZN(n13098) );
  NOR2_X1 U16388 ( .A1(n13099), .A2(n13098), .ZN(n13804) );
  NOR2_X1 U16389 ( .A1(n16816), .A2(n19985), .ZN(n13100) );
  NAND2_X1 U16390 ( .A1(n20615), .A2(n13100), .ZN(n13104) );
  NAND2_X1 U16391 ( .A1(n13095), .A2(n15871), .ZN(n13102) );
  NAND4_X1 U16392 ( .A1(n13102), .A2(n13786), .A3(n20480), .A4(n13101), .ZN(
        n13103) );
  NAND4_X1 U16393 ( .A1(n13804), .A2(n13105), .A3(n13104), .A4(n13103), .ZN(
        n13106) );
  AOI21_X1 U16394 ( .B1(n19836), .B2(n13107), .A(n13106), .ZN(n13108) );
  OAI21_X1 U16395 ( .B1(n19836), .B2(n13109), .A(n13108), .ZN(n13110) );
  NAND2_X1 U16396 ( .A1(n13141), .A2(n13112), .ZN(n16639) );
  AOI222_X1 U16397 ( .A1(n13640), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n12327), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n12216), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13114) );
  INV_X1 U16398 ( .A(n13114), .ZN(n13115) );
  NOR2_X2 U16399 ( .A1(n13642), .A2(n13117), .ZN(n14619) );
  INV_X1 U16400 ( .A(n12149), .ZN(n16799) );
  NAND2_X1 U16401 ( .A1(n16799), .A2(n15871), .ZN(n13121) );
  INV_X1 U16402 ( .A(n13118), .ZN(n13120) );
  NAND2_X1 U16403 ( .A1(n13120), .A2(n13119), .ZN(n16676) );
  NAND2_X1 U16404 ( .A1(n13121), .A2(n16676), .ZN(n13122) );
  NAND2_X1 U16405 ( .A1(n14619), .A2(n16645), .ZN(n13161) );
  NAND2_X1 U16406 ( .A1(n13141), .A2(n16798), .ZN(n14064) );
  AOI22_X1 U16407 ( .A1(n13799), .A2(n11699), .B1(n15607), .B2(n13123), .ZN(
        n13131) );
  NAND2_X1 U16408 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  NAND2_X1 U16409 ( .A1(n13128), .A2(n13127), .ZN(n13130) );
  AND4_X1 U16410 ( .A1(n13132), .A2(n13131), .A3(n13130), .A4(n13129), .ZN(
        n13138) );
  NAND2_X1 U16411 ( .A1(n13133), .A2(n15871), .ZN(n16650) );
  NAND2_X1 U16412 ( .A1(n16650), .A2(n13134), .ZN(n13136) );
  NAND2_X1 U16413 ( .A1(n13136), .A2(n13135), .ZN(n13137) );
  NAND2_X1 U16414 ( .A1(n16649), .A2(n16672), .ZN(n13140) );
  AND2_X1 U16415 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16362) );
  NAND2_X1 U16416 ( .A1(n16362), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13634) );
  NAND2_X1 U16417 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U16418 ( .A1(n13142), .A2(n14056), .ZN(n14065) );
  NAND2_X1 U16419 ( .A1(n13163), .A2(n19701), .ZN(n14046) );
  NOR2_X1 U16420 ( .A1(n13142), .A2(n14056), .ZN(n13151) );
  INV_X1 U16421 ( .A(n13151), .ZN(n14066) );
  NAND2_X1 U16422 ( .A1(n13143), .A2(n14066), .ZN(n14055) );
  AND3_X1 U16423 ( .A1(n14046), .A2(n14055), .A3(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13144) );
  OAI21_X1 U16424 ( .B1(n14064), .B2(n14065), .A(n13144), .ZN(n16636) );
  NAND2_X1 U16425 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16640) );
  NOR3_X1 U16426 ( .A1(n16624), .A2(n16636), .A3(n16640), .ZN(n16591) );
  NOR2_X1 U16427 ( .A1(n16611), .A2(n16593), .ZN(n16590) );
  INV_X1 U16428 ( .A(n14046), .ZN(n13145) );
  NOR2_X1 U16429 ( .A1(n16480), .A2(n13145), .ZN(n16637) );
  INV_X1 U16430 ( .A(n16637), .ZN(n16549) );
  NAND2_X1 U16431 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16432) );
  OR2_X1 U16432 ( .A1(n13146), .A2(n16432), .ZN(n13154) );
  NAND2_X1 U16433 ( .A1(n16480), .A2(n13154), .ZN(n13147) );
  AND2_X1 U16434 ( .A1(n16480), .A2(n16419), .ZN(n13148) );
  NAND2_X1 U16435 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n13149) );
  AND2_X1 U16436 ( .A1(n16480), .A2(n13149), .ZN(n13150) );
  OR2_X1 U16437 ( .A1(n16412), .A2(n13150), .ZN(n16388) );
  AOI21_X1 U16438 ( .B1(n16480), .B2(n13634), .A(n16388), .ZN(n13633) );
  INV_X1 U16439 ( .A(n13633), .ZN(n13159) );
  INV_X1 U16440 ( .A(n16640), .ZN(n13152) );
  INV_X1 U16441 ( .A(n14064), .ZN(n14549) );
  OAI211_X1 U16442 ( .C1(n14549), .C2(n13151), .A(n14065), .B(n16480), .ZN(
        n17305) );
  NOR2_X1 U16443 ( .A1(n17306), .A2(n17305), .ZN(n19955) );
  NAND2_X1 U16444 ( .A1(n13152), .A2(n19955), .ZN(n16589) );
  NAND2_X1 U16445 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16590), .ZN(
        n13153) );
  INV_X1 U16446 ( .A(n13154), .ZN(n13155) );
  AND2_X1 U16447 ( .A1(n16578), .A2(n13155), .ZN(n16420) );
  AND2_X1 U16448 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n13156) );
  AND2_X1 U16449 ( .A1(n16420), .A2(n13156), .ZN(n16400) );
  NAND2_X1 U16450 ( .A1(n16400), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16385) );
  NOR3_X1 U16451 ( .A1(n16385), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13634), .ZN(n13157) );
  AOI211_X1 U16452 ( .C1(n13159), .C2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13158), .B(n13157), .ZN(n13160) );
  OAI211_X1 U16453 ( .C1(n13111), .C2(n16639), .A(n13161), .B(n13160), .ZN(
        n13162) );
  INV_X1 U16454 ( .A(n13162), .ZN(n13166) );
  NAND2_X1 U16455 ( .A1(n13164), .A2(n19962), .ZN(n13165) );
  OAI211_X1 U16456 ( .C1(n13167), .C2(n19967), .A(n13166), .B(n13165), .ZN(
        P2_U3016) );
  INV_X2 U16457 ( .A(n13256), .ZN(n18067) );
  INV_X2 U16458 ( .A(n18067), .ZN(n18107) );
  NOR2_X2 U16459 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14393), .ZN(
        n13179) );
  AOI22_X1 U16460 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13176) );
  NAND2_X1 U16461 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13171) );
  NAND2_X1 U16462 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13170) );
  AND2_X2 U16463 ( .A1(n14215), .A2(n13182), .ZN(n13412) );
  NAND2_X1 U16464 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13169) );
  AND3_X1 U16465 ( .A1(n13171), .A2(n13170), .A3(n13169), .ZN(n13175) );
  AND2_X2 U16466 ( .A1(n13181), .A2(n14389), .ZN(n17109) );
  AOI22_X1 U16467 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13174) );
  INV_X1 U16468 ( .A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n18104) );
  OR2_X1 U16469 ( .A1(n18086), .A2(n18104), .ZN(n13173) );
  INV_X2 U16470 ( .A(n10442), .ZN(n18091) );
  AOI22_X1 U16471 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13186) );
  AND2_X2 U16472 ( .A1(n14215), .A2(n13181), .ZN(n13200) );
  AOI22_X1 U16473 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13184) );
  INV_X2 U16474 ( .A(n18030), .ZN(n18125) );
  AOI22_X1 U16475 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13183) );
  NAND4_X1 U16476 ( .A1(n13186), .A2(n13185), .A3(n13184), .A4(n13183), .ZN(
        n13187) );
  NAND2_X1 U16477 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13191) );
  INV_X2 U16478 ( .A(n10442), .ZN(n18122) );
  NAND2_X1 U16479 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n13190) );
  INV_X2 U16480 ( .A(n18030), .ZN(n18112) );
  NAND2_X1 U16481 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13189) );
  NAND2_X1 U16482 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n13188) );
  INV_X1 U16483 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17963) );
  OR2_X1 U16484 ( .A1(n18086), .A2(n17963), .ZN(n13195) );
  INV_X2 U16485 ( .A(n13297), .ZN(n17112) );
  NAND2_X1 U16486 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n13194) );
  NAND2_X1 U16487 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13193) );
  NAND2_X1 U16488 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n13192) );
  NAND2_X1 U16489 ( .A1(n13256), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n13199) );
  NAND2_X1 U16490 ( .A1(n13178), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n13198) );
  NAND2_X1 U16491 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n13197) );
  NAND2_X1 U16492 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n13196) );
  AND4_X1 U16493 ( .A1(n13199), .A2(n13198), .A3(n13197), .A4(n13196), .ZN(
        n13206) );
  INV_X4 U16494 ( .A(n9620), .ZN(n18106) );
  NAND2_X1 U16495 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13204) );
  NAND2_X1 U16496 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13203) );
  NAND2_X1 U16497 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n13202) );
  NAND2_X1 U16498 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13201) );
  NAND2_X1 U16499 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13212) );
  NAND2_X1 U16500 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13211) );
  INV_X4 U16501 ( .A(n17087), .ZN(n18123) );
  NAND2_X1 U16502 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13210) );
  NAND2_X1 U16503 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13209) );
  AND4_X1 U16504 ( .A1(n13212), .A2(n13211), .A3(n13210), .A4(n13209), .ZN(
        n13228) );
  NAND2_X1 U16505 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13216) );
  NAND2_X1 U16506 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13215) );
  NAND2_X1 U16507 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13214) );
  NAND2_X1 U16508 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13213) );
  AND4_X1 U16509 ( .A1(n13216), .A2(n13215), .A3(n13214), .A4(n13213), .ZN(
        n13227) );
  INV_X1 U16510 ( .A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17993) );
  OR2_X1 U16511 ( .A1(n18086), .A2(n17993), .ZN(n13220) );
  NAND2_X1 U16512 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13219) );
  NAND2_X1 U16513 ( .A1(n18131), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13218) );
  NAND2_X1 U16514 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13217) );
  AND4_X1 U16515 ( .A1(n13220), .A2(n13219), .A3(n13218), .A4(n13217), .ZN(
        n13226) );
  NAND2_X1 U16516 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13224) );
  NAND2_X1 U16517 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n13223) );
  NAND2_X1 U16518 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13222) );
  NAND2_X1 U16519 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13221) );
  AND4_X1 U16520 ( .A1(n13224), .A2(n13223), .A3(n13222), .A4(n13221), .ZN(
        n13225) );
  NAND4_X1 U16521 ( .A1(n13228), .A2(n13227), .A3(n13226), .A4(n13225), .ZN(
        n14270) );
  AND2_X1 U16522 ( .A1(n14270), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16933) );
  INV_X1 U16523 ( .A(n13528), .ZN(n14213) );
  NAND2_X1 U16524 ( .A1(n14213), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13229) );
  INV_X1 U16525 ( .A(n13230), .ZN(n13231) );
  NAND2_X1 U16526 ( .A1(n13231), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13232) );
  NAND2_X1 U16527 ( .A1(n13233), .A2(n13232), .ZN(n18710) );
  AOI22_X1 U16528 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13240) );
  NAND2_X1 U16529 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13236) );
  NAND2_X1 U16530 ( .A1(n18131), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16531 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n13234) );
  AND3_X1 U16532 ( .A1(n13236), .A2(n13235), .A3(n13234), .ZN(n13239) );
  AOI22_X1 U16533 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13238) );
  INV_X1 U16534 ( .A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13410) );
  OR2_X1 U16535 ( .A1(n18086), .A2(n13410), .ZN(n13237) );
  NAND4_X1 U16536 ( .A1(n13240), .A2(n13239), .A3(n13238), .A4(n13237), .ZN(
        n13246) );
  AOI22_X1 U16537 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18122), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U16538 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U16539 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16540 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13241) );
  NAND4_X1 U16541 ( .A1(n13244), .A2(n13243), .A3(n13242), .A4(n13241), .ZN(
        n13245) );
  XNOR2_X1 U16542 ( .A(n13249), .B(n13535), .ZN(n13247) );
  INV_X1 U16543 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18968) );
  XNOR2_X1 U16544 ( .A(n13247), .B(n18968), .ZN(n18709) );
  NAND2_X1 U16545 ( .A1(n13247), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13248) );
  INV_X1 U16546 ( .A(n13249), .ZN(n13250) );
  NAND2_X1 U16547 ( .A1(n13250), .A2(n13535), .ZN(n13270) );
  INV_X1 U16548 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13251) );
  OR2_X1 U16549 ( .A1(n18086), .A2(n13251), .ZN(n13255) );
  NAND2_X1 U16550 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n13254) );
  NAND2_X1 U16551 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13253) );
  NAND2_X1 U16552 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n13252) );
  AOI22_X1 U16553 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U16554 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13257) );
  NAND3_X1 U16555 ( .A1(n13259), .A2(n13258), .A3(n13257), .ZN(n13265) );
  AOI22_X1 U16556 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U16557 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U16558 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13261) );
  AOI22_X1 U16559 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13260) );
  NAND4_X1 U16560 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        n13264) );
  XNOR2_X1 U16561 ( .A(n13270), .B(n18317), .ZN(n13266) );
  INV_X1 U16562 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n16919) );
  INV_X1 U16563 ( .A(n13266), .ZN(n13267) );
  INV_X1 U16564 ( .A(n13270), .ZN(n13271) );
  NAND2_X1 U16565 ( .A1(n13271), .A2(n13532), .ZN(n13288) );
  AOI22_X1 U16566 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U16567 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13274) );
  NAND2_X1 U16568 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n13273) );
  NAND2_X1 U16569 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n13272) );
  AND3_X1 U16570 ( .A1(n13274), .A2(n13273), .A3(n13272), .ZN(n13277) );
  AOI22_X1 U16571 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13276) );
  OR2_X1 U16572 ( .A1(n18086), .A2(n17917), .ZN(n13275) );
  NAND4_X1 U16573 ( .A1(n13278), .A2(n13277), .A3(n13276), .A4(n13275), .ZN(
        n13284) );
  AOI22_X1 U16574 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18122), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U16575 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13281) );
  AOI22_X1 U16576 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13280) );
  INV_X1 U16577 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18156) );
  AOI22_X1 U16578 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13279) );
  NAND4_X1 U16579 ( .A1(n13282), .A2(n13281), .A3(n13280), .A4(n13279), .ZN(
        n13283) );
  XNOR2_X1 U16580 ( .A(n13288), .B(n18308), .ZN(n13285) );
  INV_X1 U16581 ( .A(n13288), .ZN(n13289) );
  NAND2_X1 U16582 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n13292) );
  NAND2_X1 U16583 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n13291) );
  NAND2_X1 U16584 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n13290) );
  AND3_X1 U16585 ( .A1(n13292), .A2(n13291), .A3(n13290), .ZN(n13296) );
  AOI22_X1 U16586 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16587 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13294) );
  INV_X1 U16588 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17893) );
  OR2_X1 U16589 ( .A1(n18086), .A2(n17893), .ZN(n13293) );
  NAND4_X1 U16590 ( .A1(n13296), .A2(n13295), .A3(n13294), .A4(n13293), .ZN(
        n13303) );
  AOI22_X1 U16591 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13301) );
  AOI22_X1 U16592 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9573), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13300) );
  AOI22_X1 U16593 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13299) );
  AOI22_X1 U16594 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13298) );
  NAND4_X1 U16595 ( .A1(n13301), .A2(n13300), .A3(n13299), .A4(n13298), .ZN(
        n13302) );
  XNOR2_X1 U16596 ( .A(n13306), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14296) );
  INV_X1 U16597 ( .A(n14296), .ZN(n13304) );
  XNOR2_X1 U16598 ( .A(n13305), .B(n13304), .ZN(n14301) );
  INV_X1 U16599 ( .A(n13305), .ZN(n13307) );
  OAI211_X1 U16600 ( .C1(n13307), .C2(n13306), .A(n13330), .B(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13308) );
  NAND2_X1 U16601 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n13312) );
  NAND2_X1 U16602 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16603 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n13310) );
  NAND2_X1 U16604 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n13309) );
  NAND2_X1 U16605 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n13316) );
  NAND2_X1 U16606 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n13315) );
  NAND2_X1 U16607 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13314) );
  NAND2_X1 U16608 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n13313) );
  INV_X1 U16609 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13317) );
  OR2_X1 U16610 ( .A1(n18086), .A2(n13317), .ZN(n13321) );
  NAND2_X1 U16611 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13320) );
  NAND2_X1 U16612 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n13319) );
  NAND2_X1 U16613 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n13318) );
  NAND2_X1 U16614 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13325) );
  NAND2_X1 U16615 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n13324) );
  NAND2_X1 U16616 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n13323) );
  INV_X1 U16617 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18151) );
  NAND2_X1 U16618 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13322) );
  NAND2_X1 U16619 ( .A1(n13330), .A2(n18302), .ZN(n13331) );
  NAND2_X1 U16620 ( .A1(n18565), .A2(n13331), .ZN(n13332) );
  NAND2_X1 U16621 ( .A1(n18567), .A2(n9838), .ZN(n13333) );
  INV_X1 U16622 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13336) );
  INV_X1 U16623 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18834) );
  INV_X1 U16624 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18868) );
  INV_X1 U16625 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18890) );
  NAND2_X1 U16626 ( .A1(n13338), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13339) );
  INV_X1 U16627 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18919) );
  NOR2_X1 U16628 ( .A1(n18931), .A2(n18919), .ZN(n18908) );
  NAND2_X1 U16629 ( .A1(n18908), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18889) );
  NAND2_X1 U16630 ( .A1(n18617), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n18861) );
  NAND2_X1 U16631 ( .A1(n18659), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13340) );
  INV_X1 U16632 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13341) );
  AND2_X1 U16633 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18813) );
  INV_X1 U16634 ( .A(n18813), .ZN(n18509) );
  OR2_X1 U16635 ( .A1(n18510), .A2(n18509), .ZN(n13342) );
  INV_X1 U16636 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21624) );
  NOR2_X1 U16637 ( .A1(n21624), .A2(n18800), .ZN(n18784) );
  NAND2_X1 U16638 ( .A1(n18784), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18766) );
  INV_X1 U16639 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18765) );
  NOR2_X1 U16640 ( .A1(n18766), .A2(n18765), .ZN(n16996) );
  AND2_X1 U16641 ( .A1(n16996), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13343) );
  NAND2_X1 U16642 ( .A1(n18813), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18757) );
  NOR2_X1 U16643 ( .A1(n18766), .A2(n18757), .ZN(n18772) );
  NAND2_X1 U16644 ( .A1(n18772), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18478) );
  INV_X1 U16645 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18750) );
  OR2_X1 U16646 ( .A1(n18478), .A2(n18750), .ZN(n16894) );
  INV_X1 U16647 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18818) );
  NAND2_X1 U16648 ( .A1(n18530), .A2(n18800), .ZN(n13344) );
  NOR2_X1 U16649 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n13344), .ZN(
        n18511) );
  INV_X1 U16650 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18770) );
  NAND2_X1 U16651 ( .A1(n18511), .A2(n18770), .ZN(n18489) );
  NAND2_X1 U16652 ( .A1(n18765), .A2(n18750), .ZN(n13345) );
  OAI22_X1 U16653 ( .A1(n18510), .A2(n16894), .B1(n18489), .B2(n13345), .ZN(
        n13346) );
  NAND2_X1 U16654 ( .A1(n13351), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13350) );
  INV_X1 U16655 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18743) );
  NAND2_X1 U16656 ( .A1(n18659), .A2(n18743), .ZN(n13348) );
  NAND2_X1 U16657 ( .A1(n13350), .A2(n13349), .ZN(n16878) );
  NAND2_X1 U16658 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U16659 ( .A1(n18659), .A2(n13554), .ZN(n13352) );
  NOR2_X2 U16660 ( .A1(n13354), .A2(n18565), .ZN(n18450) );
  NAND2_X1 U16661 ( .A1(n18450), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13359) );
  INV_X1 U16662 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n13355) );
  INV_X1 U16663 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n18438) );
  NAND2_X1 U16664 ( .A1(n18565), .A2(n18438), .ZN(n13357) );
  OR2_X1 U16665 ( .A1(n18446), .A2(n13357), .ZN(n13358) );
  NAND2_X1 U16666 ( .A1(n13359), .A2(n13358), .ZN(n13360) );
  XNOR2_X1 U16667 ( .A(n13360), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17139) );
  INV_X1 U16668 ( .A(n17139), .ZN(n13527) );
  INV_X1 U16669 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13361) );
  OR2_X1 U16670 ( .A1(n18086), .A2(n13361), .ZN(n13365) );
  NAND2_X1 U16671 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n13364) );
  NAND2_X1 U16672 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13363) );
  NAND2_X1 U16673 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13362) );
  NAND2_X1 U16674 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n13369) );
  NAND2_X1 U16675 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n13368) );
  NAND2_X1 U16676 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13367) );
  NAND2_X1 U16677 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13366) );
  NAND2_X1 U16678 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n13373) );
  NAND2_X1 U16679 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13372) );
  NAND2_X1 U16680 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n13371) );
  NAND2_X1 U16681 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13370) );
  NAND2_X1 U16682 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n13377) );
  NAND2_X1 U16683 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13376) );
  NAND2_X1 U16684 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n13375) );
  NAND2_X1 U16685 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13374) );
  NAND2_X1 U16686 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13385) );
  NAND2_X1 U16687 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n13384) );
  NAND2_X1 U16688 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13383) );
  NAND2_X1 U16689 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13382) );
  INV_X1 U16690 ( .A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n18136) );
  OR2_X1 U16691 ( .A1(n18086), .A2(n18136), .ZN(n13389) );
  NAND2_X1 U16692 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13388) );
  NAND2_X1 U16693 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n13387) );
  NAND2_X1 U16694 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13386) );
  NAND2_X1 U16695 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n13393) );
  NAND2_X1 U16696 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n13392) );
  NAND2_X1 U16697 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13391) );
  NAND2_X1 U16698 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n13390) );
  NAND2_X1 U16699 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n13397) );
  NAND2_X1 U16700 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n13396) );
  NAND2_X1 U16701 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13395) );
  NAND2_X1 U16702 ( .A1(n18112), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13394) );
  NOR2_X1 U16703 ( .A1(n14208), .A2(n17006), .ZN(n19587) );
  INV_X1 U16704 ( .A(n19587), .ZN(n19574) );
  INV_X1 U16705 ( .A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n18014) );
  AOI22_X1 U16706 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9573), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13402) );
  AOI22_X1 U16707 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13403) );
  AOI22_X1 U16708 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18080), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13407) );
  AOI22_X1 U16709 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13406) );
  AOI22_X1 U16710 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13405) );
  AOI22_X1 U16711 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17109), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n13404) );
  NAND4_X1 U16712 ( .A1(n13407), .A2(n13406), .A3(n13405), .A4(n13404), .ZN(
        n13408) );
  INV_X4 U16713 ( .A(n18120), .ZN(n19024) );
  NAND2_X1 U16714 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n13409) );
  INV_X1 U16715 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13411) );
  INV_X1 U16716 ( .A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17082) );
  OAI22_X1 U16717 ( .A1(n13423), .A2(n13411), .B1(n9626), .B2(n17082), .ZN(
        n13415) );
  INV_X1 U16718 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13413) );
  OAI22_X1 U16719 ( .A1(n18035), .A2(n17081), .B1(n18135), .B2(n13413), .ZN(
        n13414) );
  AOI22_X1 U16720 ( .A1(n18091), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13419) );
  AOI22_X1 U16721 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13418) );
  AOI22_X1 U16722 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U16723 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13416) );
  INV_X1 U16724 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17919) );
  AOI22_X1 U16725 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13421) );
  NAND2_X1 U16726 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n13420) );
  OAI211_X1 U16727 ( .C1(n17919), .C2(n18135), .A(n13421), .B(n13420), .ZN(
        n13422) );
  INV_X1 U16728 ( .A(n13422), .ZN(n13428) );
  INV_X1 U16729 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17107) );
  INV_X1 U16730 ( .A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17110) );
  OAI22_X1 U16731 ( .A1(n13423), .A2(n17107), .B1(n9626), .B2(n17110), .ZN(
        n13424) );
  INV_X1 U16732 ( .A(n13424), .ZN(n13427) );
  INV_X1 U16733 ( .A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17111) );
  OAI22_X1 U16734 ( .A1(n18141), .A2(n17111), .B1(n18030), .B2(n17917), .ZN(
        n13425) );
  INV_X1 U16735 ( .A(n13425), .ZN(n13426) );
  NAND3_X1 U16736 ( .A1(n13428), .A2(n13427), .A3(n13426), .ZN(n13434) );
  AOI22_X1 U16737 ( .A1(n18091), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U16738 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13431) );
  AOI22_X1 U16739 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13430) );
  AOI22_X1 U16740 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13429) );
  NAND4_X1 U16741 ( .A1(n13432), .A2(n13431), .A3(n13430), .A4(n13429), .ZN(
        n13433) );
  AOI22_X1 U16742 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13442) );
  NAND2_X1 U16743 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13437) );
  NAND2_X1 U16744 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13436) );
  NAND2_X1 U16745 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13435) );
  AOI22_X1 U16746 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13440) );
  INV_X1 U16747 ( .A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13438) );
  OR2_X1 U16748 ( .A1(n18086), .A2(n13438), .ZN(n13439) );
  NAND4_X1 U16749 ( .A1(n13442), .A2(n13441), .A3(n13440), .A4(n13439), .ZN(
        n13448) );
  AOI22_X1 U16750 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U16751 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U16752 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U16753 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13443) );
  NAND4_X1 U16754 ( .A1(n13446), .A2(n13445), .A3(n13444), .A4(n13443), .ZN(
        n13447) );
  NAND2_X1 U16755 ( .A1(n19016), .A2(n14104), .ZN(n14103) );
  INV_X1 U16756 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n18051) );
  AOI22_X1 U16757 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13450) );
  NAND2_X1 U16758 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n13449) );
  OAI211_X1 U16759 ( .C1(n18051), .C2(n18086), .A(n13450), .B(n13449), .ZN(
        n13451) );
  INV_X1 U16760 ( .A(n13451), .ZN(n13454) );
  AOI22_X1 U16761 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U16762 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13452) );
  NAND3_X1 U16763 ( .A1(n13454), .A2(n13453), .A3(n13452), .ZN(n13460) );
  AOI22_X1 U16764 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U16765 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13457) );
  AOI22_X1 U16766 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18081), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13456) );
  AOI22_X1 U16767 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13455) );
  NAND4_X1 U16768 ( .A1(n13458), .A2(n13457), .A3(n13456), .A4(n13455), .ZN(
        n13459) );
  INV_X1 U16769 ( .A(n14205), .ZN(n19012) );
  AOI22_X1 U16770 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13466) );
  NAND2_X1 U16771 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13463) );
  NAND2_X1 U16772 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n13462) );
  NAND2_X1 U16773 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13461) );
  AOI22_X1 U16774 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13465) );
  INV_X1 U16775 ( .A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17846) );
  OR2_X1 U16776 ( .A1(n18086), .A2(n17846), .ZN(n13464) );
  NAND4_X1 U16777 ( .A1(n13466), .A2(n9668), .A3(n13465), .A4(n13464), .ZN(
        n13472) );
  AOI22_X1 U16778 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U16779 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13469) );
  AOI22_X1 U16780 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13468) );
  AOI22_X1 U16781 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13467) );
  NAND4_X1 U16782 ( .A1(n13470), .A2(n13469), .A3(n13468), .A4(n13467), .ZN(
        n13471) );
  NAND2_X1 U16783 ( .A1(n19012), .A2(n18186), .ZN(n14171) );
  NOR3_X2 U16784 ( .A1(n14096), .A2(n14103), .A3(n14171), .ZN(n14162) );
  NAND2_X1 U16785 ( .A1(n14205), .A2(n18186), .ZN(n13480) );
  NOR4_X4 U16786 ( .A1(n14096), .A2(n19016), .A3(n13478), .A4(n14214), .ZN(
        n18379) );
  NOR3_X1 U16787 ( .A1(n18120), .A2(n18992), .A3(n19008), .ZN(n13475) );
  NAND2_X1 U16788 ( .A1(n19004), .A2(n14175), .ZN(n17421) );
  NOR2_X1 U16789 ( .A1(n13481), .A2(n19019), .ZN(n14354) );
  NOR3_X1 U16790 ( .A1(n14214), .A2(n14210), .A3(n19001), .ZN(n14099) );
  AOI211_X1 U16791 ( .C1(n14103), .C2(n13478), .A(n13474), .B(n14099), .ZN(
        n13476) );
  INV_X1 U16792 ( .A(n13483), .ZN(n13477) );
  AOI21_X1 U16793 ( .B1(n19024), .B2(n13477), .A(n14205), .ZN(n13486) );
  NAND2_X1 U16794 ( .A1(n14104), .A2(n13483), .ZN(n14105) );
  AOI21_X1 U16795 ( .B1(n13478), .B2(n14105), .A(n18992), .ZN(n13485) );
  NOR2_X1 U16796 ( .A1(n13479), .A2(n19004), .ZN(n14094) );
  NOR2_X1 U16797 ( .A1(n13481), .A2(n13480), .ZN(n14097) );
  OAI21_X1 U16798 ( .B1(n14094), .B2(n13483), .A(n13482), .ZN(n13484) );
  NAND2_X1 U16799 ( .A1(n14175), .A2(n13489), .ZN(n13768) );
  NAND3_X1 U16800 ( .A1(n14096), .A2(n14160), .A3(n19001), .ZN(n13490) );
  NAND2_X1 U16801 ( .A1(n13490), .A2(n13489), .ZN(n14172) );
  AOI21_X4 U16802 ( .B1(n14173), .B2(n14388), .A(n14172), .ZN(n18926) );
  NOR2_X4 U16803 ( .A1(n18836), .A2(n19001), .ZN(n19399) );
  MUX2_X1 U16804 ( .A(n13491), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n13514) );
  NAND2_X1 U16805 ( .A1(n13514), .A2(n13515), .ZN(n13493) );
  NAND2_X1 U16806 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n13491), .ZN(
        n13492) );
  NAND2_X1 U16807 ( .A1(n13493), .A2(n13492), .ZN(n13502) );
  MUX2_X1 U16808 ( .A(n19430), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13501) );
  NAND2_X1 U16809 ( .A1(n13502), .A2(n13501), .ZN(n13500) );
  NAND2_X1 U16810 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19430), .ZN(
        n13494) );
  NAND2_X1 U16811 ( .A1(n13500), .A2(n13494), .ZN(n13495) );
  NAND2_X1 U16812 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n19410), .ZN(
        n13496) );
  OAI21_X1 U16813 ( .B1(n13495), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13496), .ZN(n13503) );
  NAND2_X1 U16814 ( .A1(n13503), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13499) );
  NAND2_X1 U16815 ( .A1(n13495), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13504) );
  INV_X1 U16816 ( .A(n13496), .ZN(n13497) );
  NAND2_X1 U16817 ( .A1(n13504), .A2(n13497), .ZN(n13498) );
  NAND2_X1 U16818 ( .A1(n13499), .A2(n13498), .ZN(n13511) );
  OAI21_X1 U16819 ( .B1(n13502), .B2(n13501), .A(n13500), .ZN(n13521) );
  INV_X1 U16820 ( .A(n13518), .ZN(n13513) );
  INV_X1 U16821 ( .A(n13503), .ZN(n13507) );
  NAND2_X1 U16822 ( .A1(n13504), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13506) );
  INV_X1 U16823 ( .A(n13515), .ZN(n13508) );
  OAI21_X1 U16824 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13509), .A(
        n13508), .ZN(n13510) );
  NOR2_X1 U16825 ( .A1(n13511), .A2(n13510), .ZN(n13523) );
  NAND2_X1 U16826 ( .A1(n13523), .A2(n13514), .ZN(n13512) );
  NAND2_X1 U16827 ( .A1(n19399), .A2(n19401), .ZN(n13526) );
  XNOR2_X1 U16828 ( .A(n19570), .B(n14104), .ZN(n14102) );
  INV_X1 U16829 ( .A(n13514), .ZN(n13516) );
  XNOR2_X1 U16830 ( .A(n13516), .B(n13515), .ZN(n13517) );
  NAND2_X1 U16831 ( .A1(n13518), .A2(n13517), .ZN(n13520) );
  INV_X1 U16832 ( .A(n13521), .ZN(n13522) );
  NAND2_X1 U16833 ( .A1(n13523), .A2(n13522), .ZN(n13524) );
  NAND2_X1 U16834 ( .A1(n16961), .A2(n19405), .ZN(n13525) );
  NOR2_X2 U16835 ( .A1(n17423), .A2(n19570), .ZN(n16923) );
  NOR2_X1 U16836 ( .A1(n13355), .A2(n18438), .ZN(n17136) );
  NAND2_X1 U16837 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18737) );
  NOR2_X1 U16838 ( .A1(n18478), .A2(n18737), .ZN(n18741) );
  NAND2_X1 U16839 ( .A1(n13528), .A2(n14270), .ZN(n13539) );
  INV_X1 U16840 ( .A(n14281), .ZN(n13538) );
  NAND2_X1 U16841 ( .A1(n13539), .A2(n13538), .ZN(n13537) );
  NAND2_X1 U16842 ( .A1(n13537), .A2(n13535), .ZN(n13533) );
  NAND2_X1 U16843 ( .A1(n13529), .A2(n18308), .ZN(n14292) );
  NOR2_X1 U16844 ( .A1(n18305), .A2(n14292), .ZN(n13547) );
  NAND2_X1 U16845 ( .A1(n13547), .A2(n17130), .ZN(n13548) );
  INV_X1 U16846 ( .A(n14292), .ZN(n14294) );
  XNOR2_X1 U16847 ( .A(n18305), .B(n14294), .ZN(n13546) );
  INV_X1 U16848 ( .A(n18308), .ZN(n13530) );
  XNOR2_X1 U16849 ( .A(n13530), .B(n13529), .ZN(n13531) );
  NAND2_X1 U16850 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13531), .ZN(
        n13545) );
  INV_X1 U16851 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18942) );
  XNOR2_X1 U16852 ( .A(n18942), .B(n13531), .ZN(n18696) );
  XNOR2_X1 U16853 ( .A(n13533), .B(n13532), .ZN(n13534) );
  NAND2_X1 U16854 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13534), .ZN(
        n13544) );
  XOR2_X1 U16855 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n13534), .Z(
        n16926) );
  INV_X1 U16856 ( .A(n13535), .ZN(n14288) );
  XNOR2_X1 U16857 ( .A(n13537), .B(n14288), .ZN(n13536) );
  NAND2_X1 U16858 ( .A1(n13536), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13543) );
  XNOR2_X1 U16859 ( .A(n13536), .B(n18968), .ZN(n18705) );
  OAI21_X1 U16860 ( .B1(n13539), .B2(n13538), .A(n13537), .ZN(n13541) );
  NAND2_X1 U16861 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13541), .ZN(
        n13542) );
  INV_X1 U16862 ( .A(n13539), .ZN(n13540) );
  OR2_X1 U16863 ( .A1(n14270), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16935) );
  NOR2_X1 U16864 ( .A1(n16936), .A2(n16935), .ZN(n16934) );
  AOI211_X1 U16865 ( .C1(n14213), .C2(n9830), .A(n13540), .B(n16934), .ZN(
        n14089) );
  NAND2_X1 U16866 ( .A1(n13543), .A2(n18706), .ZN(n16925) );
  NAND2_X1 U16867 ( .A1(n16926), .A2(n16925), .ZN(n16924) );
  XOR2_X1 U16868 ( .A(n18302), .B(n13547), .Z(n14197) );
  NAND2_X1 U16869 ( .A1(n14196), .A2(n14197), .ZN(n14195) );
  NAND2_X1 U16870 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n14195), .ZN(
        n13551) );
  NOR2_X1 U16871 ( .A1(n13548), .A2(n13551), .ZN(n13553) );
  INV_X1 U16872 ( .A(n13548), .ZN(n13552) );
  NOR2_X1 U16873 ( .A1(n14196), .A2(n14197), .ZN(n13550) );
  NOR2_X1 U16874 ( .A1(n13552), .A2(n13551), .ZN(n13549) );
  AOI211_X1 U16875 ( .C1(n13552), .C2(n13551), .A(n13550), .B(n13549), .ZN(
        n14260) );
  NAND2_X1 U16876 ( .A1(n17136), .A2(n16978), .ZN(n16963) );
  INV_X1 U16877 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n17135) );
  NAND2_X1 U16878 ( .A1(n16963), .A2(n17135), .ZN(n13571) );
  NOR2_X4 U16879 ( .A1(n17423), .A2(n19001), .ZN(n18647) );
  INV_X1 U16880 ( .A(n13554), .ZN(n16977) );
  NAND2_X1 U16881 ( .A1(n18741), .A2(n16977), .ZN(n18437) );
  NAND2_X1 U16882 ( .A1(n17136), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n17179) );
  NOR2_X1 U16883 ( .A1(n18437), .A2(n17179), .ZN(n17177) );
  NAND2_X1 U16884 ( .A1(n17177), .A2(n13555), .ZN(n17133) );
  NAND2_X1 U16885 ( .A1(n18647), .A2(n17133), .ZN(n17313) );
  INV_X1 U16886 ( .A(n17313), .ZN(n13570) );
  AND2_X2 U16887 ( .A1(n13556), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18901) );
  NAND2_X1 U16888 ( .A1(n18901), .A2(n18858), .ZN(n18601) );
  NOR2_X2 U16889 ( .A1(n18868), .A2(n18601), .ZN(n18845) );
  NAND2_X1 U16890 ( .A1(n18845), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18844) );
  NOR2_X1 U16891 ( .A1(n18844), .A2(n18437), .ZN(n16979) );
  NAND2_X1 U16892 ( .A1(n17136), .A2(n16979), .ZN(n16962) );
  INV_X1 U16893 ( .A(n17177), .ZN(n13557) );
  NOR2_X1 U16894 ( .A1(n18844), .A2(n13557), .ZN(n17315) );
  AND2_X2 U16895 ( .A1(n16923), .A2(n18302), .ZN(n18645) );
  INV_X1 U16896 ( .A(n18645), .ZN(n17314) );
  AOI211_X1 U16897 ( .C1(n17135), .C2(n16962), .A(n17315), .B(n17314), .ZN(
        n13568) );
  INV_X1 U16898 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19571) );
  INV_X1 U16899 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17761) );
  NAND4_X1 U16900 ( .A1(n18637), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17636) );
  INV_X1 U16901 ( .A(n17636), .ZN(n13558) );
  NAND2_X1 U16902 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18572) );
  NAND2_X1 U16903 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18538) );
  NAND2_X1 U16904 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n18498) );
  NAND2_X1 U16905 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18465) );
  INV_X1 U16906 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13559) );
  NOR2_X1 U16907 ( .A1(n18465), .A2(n13559), .ZN(n16881) );
  INV_X1 U16908 ( .A(n18433), .ZN(n13560) );
  NAND2_X1 U16909 ( .A1(n13560), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13565) );
  NOR2_X1 U16910 ( .A1(n17474), .A2(n13565), .ZN(n16863) );
  OR2_X1 U16911 ( .A1(n19180), .A2(n16863), .ZN(n13566) );
  NOR2_X1 U16912 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n13561) );
  NAND2_X2 U16913 ( .A1(n19584), .A2(n13561), .ZN(n18981) );
  INV_X2 U16914 ( .A(n18981), .ZN(n18954) );
  INV_X1 U16915 ( .A(n17439), .ZN(n13562) );
  NOR2_X1 U16916 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21628), .ZN(n16883) );
  INV_X1 U16917 ( .A(n16883), .ZN(n18608) );
  INV_X1 U16918 ( .A(n19584), .ZN(n17817) );
  NAND2_X1 U16919 ( .A1(n21628), .A2(n19552), .ZN(n17417) );
  NAND2_X1 U16920 ( .A1(n17817), .A2(n17417), .ZN(n18983) );
  OAI211_X1 U16921 ( .C1(n13562), .C2(n18608), .A(n18708), .B(n13566), .ZN(
        n16867) );
  AOI22_X1 U16922 ( .A1(n18954), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16867), .ZN(n13564) );
  NOR2_X1 U16923 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18495), .ZN(
        n16868) );
  NAND2_X1 U16924 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16928) );
  AOI21_X1 U16925 ( .B1(n17474), .B2(n17439), .A(n17308), .ZN(n17473) );
  OAI21_X1 U16926 ( .B1(n16868), .B2(n18529), .A(n17473), .ZN(n13563) );
  OAI211_X1 U16927 ( .C1(n13566), .C2(n13565), .A(n13564), .B(n13563), .ZN(
        n13567) );
  INV_X1 U16928 ( .A(n13576), .ZN(n13578) );
  NAND2_X1 U16929 ( .A1(n13578), .A2(n13577), .ZN(n14561) );
  INV_X1 U16930 ( .A(n13582), .ZN(n14553) );
  NAND2_X1 U16931 ( .A1(n16207), .A2(n16474), .ZN(n13584) );
  NAND2_X1 U16932 ( .A1(n13587), .A2(n13588), .ZN(n13589) );
  NAND2_X1 U16933 ( .A1(n19621), .A2(n19946), .ZN(n13596) );
  INV_X1 U16934 ( .A(n14660), .ZN(n13592) );
  INV_X1 U16935 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n13590) );
  NAND2_X1 U16936 ( .A1(n9691), .A2(n13590), .ZN(n13591) );
  NAND2_X1 U16937 ( .A1(n13592), .A2(n13591), .ZN(n19625) );
  NOR2_X1 U16938 ( .A1(n19701), .A2(n20538), .ZN(n16468) );
  AOI21_X1 U16939 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16468), .ZN(n13593) );
  OAI21_X1 U16940 ( .B1(n19939), .B2(n19625), .A(n13593), .ZN(n13594) );
  NAND2_X1 U16941 ( .A1(n13597), .A2(n12959), .ZN(n13598) );
  INV_X1 U16942 ( .A(n10599), .ZN(n14045) );
  NAND2_X1 U16943 ( .A1(n12921), .A2(n13600), .ZN(n13940) );
  OAI21_X1 U16944 ( .B1(n13914), .B2(n14038), .A(n13940), .ZN(n13601) );
  NAND2_X1 U16945 ( .A1(n13601), .A2(n14043), .ZN(n13602) );
  AND2_X1 U16946 ( .A1(n17230), .A2(n14045), .ZN(n13604) );
  NOR4_X1 U16947 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n13608) );
  NOR4_X1 U16948 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13607) );
  NOR4_X1 U16949 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(
        P1_ADDRESS_REG_6__SCAN_IN), .A3(P1_ADDRESS_REG_5__SCAN_IN), .A4(
        P1_ADDRESS_REG_4__SCAN_IN), .ZN(n13606) );
  NOR4_X1 U16950 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13605) );
  AND4_X1 U16951 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13613) );
  NOR4_X1 U16952 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_3__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13611) );
  NOR4_X1 U16953 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13610) );
  NOR4_X1 U16954 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13609) );
  AND4_X1 U16955 ( .A1(n13611), .A2(n13610), .A3(n13609), .A4(n21428), .ZN(
        n13612) );
  NAND2_X1 U16956 ( .A1(n13613), .A2(n13612), .ZN(n13614) );
  AOI22_X1 U16957 ( .A1(n13615), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15123), .ZN(n13616) );
  INV_X1 U16958 ( .A(n13616), .ZN(n13618) );
  INV_X1 U16959 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n17324) );
  NOR2_X1 U16960 ( .A1(n13618), .A2(n13617), .ZN(n13619) );
  NAND2_X1 U16961 ( .A1(n13620), .A2(n13619), .ZN(P1_U2873) );
  AND3_X1 U16962 ( .A1(n15353), .A2(n15416), .A3(n13621), .ZN(n15220) );
  NOR2_X1 U16963 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15391) );
  NAND3_X1 U16964 ( .A1(n15220), .A2(n15391), .A3(n15383), .ZN(n13623) );
  NOR2_X1 U16965 ( .A1(n15353), .A2(n13622), .ZN(n15211) );
  INV_X1 U16966 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13624) );
  AOI21_X1 U16967 ( .B1(n14758), .B2(n13626), .A(n13697), .ZN(n15035) );
  NAND2_X1 U16968 ( .A1(n15035), .A2(n20801), .ZN(n13631) );
  INV_X1 U16969 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21471) );
  NOR2_X1 U16970 ( .A1(n15360), .A2(n21471), .ZN(n15196) );
  INV_X1 U16971 ( .A(n15381), .ZN(n13628) );
  NOR3_X1 U16972 ( .A1(n13628), .A2(n13627), .A3(n13735), .ZN(n13629) );
  AOI211_X1 U16973 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15379), .A(
        n15196), .B(n13629), .ZN(n13630) );
  OAI21_X1 U16974 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14559), .A(
        n13633), .ZN(n13638) );
  NOR4_X1 U16975 ( .A1(n16385), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13635), .A4(n13634), .ZN(n13636) );
  AOI211_X1 U16976 ( .C1(n13638), .C2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n13637), .B(n13636), .ZN(n13639) );
  OAI21_X1 U16977 ( .B1(n14696), .B2(n16639), .A(n13639), .ZN(n13644) );
  AOI222_X1 U16978 ( .A1(n13640), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12327), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12216), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13641) );
  NOR2_X1 U16979 ( .A1(n14695), .A2(n19959), .ZN(n13643) );
  NAND2_X1 U16980 ( .A1(n13645), .A2(n19962), .ZN(n13646) );
  OAI211_X1 U16981 ( .C1(n13648), .C2(n19967), .A(n13647), .B(n13646), .ZN(
        P2_U3015) );
  XNOR2_X1 U16982 ( .A(n13655), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13652) );
  INV_X1 U16983 ( .A(n13652), .ZN(n13650) );
  AND2_X1 U16984 ( .A1(n13650), .A2(n16192), .ZN(n13659) );
  INV_X1 U16985 ( .A(n13659), .ZN(n13662) );
  INV_X1 U16986 ( .A(n16190), .ZN(n13658) );
  INV_X1 U16987 ( .A(n13655), .ZN(n13654) );
  OAI21_X1 U16988 ( .B1(n16193), .B2(n13672), .A(n13654), .ZN(n13657) );
  OAI21_X1 U16989 ( .B1(n13672), .B2(n16192), .A(n13655), .ZN(n13656) );
  AOI22_X1 U16990 ( .A1(n13659), .A2(n13658), .B1(n13657), .B2(n13656), .ZN(
        n13660) );
  AND2_X1 U16991 ( .A1(n15739), .A2(n13666), .ZN(n13667) );
  NOR2_X1 U16992 ( .A1(n13665), .A2(n13667), .ZN(n16044) );
  AOI21_X1 U16993 ( .B1(n13668), .B2(n15740), .A(n15714), .ZN(n13691) );
  INV_X1 U16994 ( .A(n13691), .ZN(n15903) );
  NAND2_X1 U16995 ( .A1(n16341), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n13688) );
  INV_X1 U16996 ( .A(n13669), .ZN(n13670) );
  NOR2_X1 U16997 ( .A1(n16543), .A2(n13671), .ZN(n16431) );
  NAND2_X1 U16998 ( .A1(n16431), .A2(n13672), .ZN(n13673) );
  OAI211_X1 U16999 ( .C1(n13674), .C2(n14559), .A(n13673), .B(n16576), .ZN(
        n16447) );
  OAI21_X1 U17000 ( .B1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n16431), .A(
        n16447), .ZN(n13675) );
  OAI211_X1 U17001 ( .C1(n15903), .C2(n16639), .A(n13688), .B(n13675), .ZN(
        n13676) );
  AOI21_X1 U17002 ( .B1(n16645), .B2(n16044), .A(n13676), .ZN(n13677) );
  AOI21_X1 U17003 ( .B1(n13682), .B2(n15633), .A(n13681), .ZN(n16369) );
  INV_X1 U17004 ( .A(n16369), .ZN(n13684) );
  NAND2_X1 U17005 ( .A1(n9574), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13683) );
  OAI21_X1 U17006 ( .B1(n13684), .B2(n9574), .A(n13683), .ZN(n13685) );
  NAND2_X1 U17007 ( .A1(n13687), .A2(n19936), .ZN(n13695) );
  AOI21_X1 U17008 ( .B1(n15728), .B2(n14659), .A(n14663), .ZN(n15733) );
  NAND2_X1 U17009 ( .A1(n19917), .A2(n15733), .ZN(n13689) );
  OAI211_X1 U17010 ( .C1(n15728), .C2(n19950), .A(n13689), .B(n13688), .ZN(
        n13690) );
  AOI21_X1 U17011 ( .B1(n13691), .B2(n19946), .A(n13690), .ZN(n13692) );
  NAND2_X1 U17012 ( .A1(n13695), .A2(n13694), .ZN(P2_U2993) );
  NAND2_X1 U17013 ( .A1(n13697), .A2(n13696), .ZN(n14730) );
  NAND2_X1 U17014 ( .A1(n14730), .A2(n12951), .ZN(n13699) );
  NAND2_X1 U17015 ( .A1(n13699), .A2(n13698), .ZN(n13701) );
  OR2_X1 U17016 ( .A1(n13697), .A2(n12932), .ZN(n13700) );
  NAND2_X1 U17017 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  AOI22_X1 U17018 ( .A1(n14733), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n12969), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14732) );
  XNOR2_X1 U17019 ( .A(n13702), .B(n14732), .ZN(n15033) );
  INV_X1 U17020 ( .A(n15033), .ZN(n13747) );
  AND2_X1 U17021 ( .A1(n12901), .A2(n14043), .ZN(n13703) );
  NAND2_X1 U17022 ( .A1(n13867), .A2(n13703), .ZN(n13802) );
  NAND2_X1 U17023 ( .A1(n11005), .A2(n21403), .ZN(n21503) );
  NAND2_X1 U17024 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n17172), .ZN(n17281) );
  NOR2_X1 U17025 ( .A1(n17281), .A2(n10276), .ZN(n13706) );
  NAND2_X1 U17026 ( .A1(n11431), .A2(n21508), .ZN(n13704) );
  NAND2_X1 U17027 ( .A1(n15360), .A2(n13704), .ZN(n13705) );
  AND2_X1 U17028 ( .A1(n20819), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13713) );
  INV_X1 U17029 ( .A(n13713), .ZN(n13708) );
  NAND2_X1 U17030 ( .A1(n21419), .A2(n21497), .ZN(n17165) );
  INV_X1 U17031 ( .A(n17165), .ZN(n13711) );
  NOR2_X1 U17032 ( .A1(n13708), .A2(n13711), .ZN(n13709) );
  INV_X1 U17033 ( .A(n13730), .ZN(n13710) );
  AND2_X1 U17034 ( .A1(n13712), .A2(n13711), .ZN(n13715) );
  NOR2_X1 U17035 ( .A1(n13715), .A2(n13713), .ZN(n13714) );
  AND2_X2 U17036 ( .A1(n13716), .A2(n13714), .ZN(n20685) );
  AND2_X2 U17037 ( .A1(n15001), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20698) );
  AOI22_X1 U17038 ( .A1(n20685), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20698), .ZN(n13725) );
  INV_X1 U17039 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n21465) );
  INV_X1 U17040 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21435) );
  INV_X1 U17041 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21431) );
  NAND4_X1 U17042 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14992)
         );
  NOR2_X1 U17043 ( .A1(n21431), .A2(n14992), .ZN(n20670) );
  NAND2_X1 U17044 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20670), .ZN(n20671) );
  NOR2_X1 U17045 ( .A1(n21435), .A2(n20671), .ZN(n14984) );
  NAND2_X1 U17046 ( .A1(n14984), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n14869) );
  NAND2_X1 U17047 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14935) );
  AND2_X1 U17048 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14933) );
  NAND2_X1 U17049 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14933), .ZN(n13717) );
  NOR2_X1 U17050 ( .A1(n14935), .A2(n13717), .ZN(n17202) );
  NAND2_X1 U17051 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n17202), .ZN(n14871) );
  NAND3_X1 U17052 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14874) );
  NOR3_X1 U17053 ( .A1(n14869), .A2(n14871), .A3(n14874), .ZN(n13718) );
  NAND3_X1 U17054 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n13718), .ZN(n14854) );
  INV_X1 U17055 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21454) );
  NOR2_X1 U17056 ( .A1(n14854), .A2(n21454), .ZN(n14839) );
  NAND2_X1 U17057 ( .A1(n14839), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14817) );
  NAND2_X1 U17058 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n13719) );
  OR2_X1 U17059 ( .A1(n14817), .A2(n13719), .ZN(n14806) );
  INV_X1 U17060 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21461) );
  NOR2_X1 U17061 ( .A1(n14806), .A2(n21461), .ZN(n14790) );
  NAND2_X1 U17062 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n14790), .ZN(n14775) );
  NOR2_X1 U17063 ( .A1(n21465), .A2(n14775), .ZN(n14765) );
  NAND2_X1 U17064 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(n14765), .ZN(n14747) );
  NOR2_X1 U17065 ( .A1(n21471), .A2(n14747), .ZN(n14718) );
  NAND2_X1 U17066 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(n14718), .ZN(n13720) );
  NOR2_X1 U17067 ( .A1(n20687), .A2(n13720), .ZN(n14737) );
  AND2_X1 U17068 ( .A1(n20687), .A2(n15001), .ZN(n14981) );
  AND2_X1 U17069 ( .A1(n15001), .A2(n14718), .ZN(n13721) );
  NOR2_X1 U17070 ( .A1(n14981), .A2(n13721), .ZN(n14749) );
  AOI21_X1 U17071 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(P1_REIP_REG_30__SCAN_IN), 
        .A(n20687), .ZN(n13722) );
  NOR2_X1 U17072 ( .A1(n14749), .A2(n13722), .ZN(n14741) );
  INV_X1 U17073 ( .A(n14741), .ZN(n13723) );
  OAI21_X1 U17074 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14737), .A(n13723), 
        .ZN(n13724) );
  OAI211_X1 U17075 ( .C1(n20691), .C2(n14522), .A(n13725), .B(n13724), .ZN(
        n13726) );
  AOI21_X1 U17076 ( .B1(n13747), .B2(n20705), .A(n13726), .ZN(n13734) );
  NAND2_X1 U17077 ( .A1(n15032), .A2(n13732), .ZN(n13733) );
  NAND2_X1 U17078 ( .A1(n13734), .A2(n13733), .ZN(P1_U2810) );
  INV_X1 U17079 ( .A(n13735), .ZN(n13736) );
  NOR2_X1 U17080 ( .A1(n13737), .A2(n13736), .ZN(n13740) );
  AOI22_X1 U17081 ( .A1(n15203), .A2(n13740), .B1(n13739), .B2(n13738), .ZN(
        n13741) );
  XNOR2_X1 U17082 ( .A(n13741), .B(n10909), .ZN(n14525) );
  OAI211_X1 U17083 ( .C1(n17255), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n13742), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15369) );
  INV_X1 U17084 ( .A(n15369), .ZN(n13745) );
  INV_X1 U17085 ( .A(n15374), .ZN(n13743) );
  AOI21_X1 U17086 ( .B1(n13743), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13744) );
  NAND2_X1 U17087 ( .A1(n20786), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14521) );
  OAI21_X1 U17088 ( .B1(n13745), .B2(n13744), .A(n14521), .ZN(n13746) );
  OAI21_X1 U17089 ( .B1(n14525), .B2(n20807), .A(n13748), .ZN(P1_U3001) );
  OR2_X1 U17090 ( .A1(n14745), .A2(n13749), .ZN(n13750) );
  NOR2_X1 U17091 ( .A1(n14710), .A2(n17244), .ZN(n13756) );
  NAND2_X1 U17092 ( .A1(n14723), .A2(n15274), .ZN(n13754) );
  OAI21_X1 U17093 ( .B1(n15271), .B2(n9914), .A(n13751), .ZN(n13752) );
  INV_X1 U17094 ( .A(n13752), .ZN(n13753) );
  NAND2_X1 U17095 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  OAI21_X1 U17096 ( .B1(n13758), .B2(n20631), .A(n13757), .ZN(P1_U2970) );
  NOR2_X1 U17097 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13760) );
  NOR4_X1 U17098 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13759) );
  NAND4_X1 U17099 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13760), .A4(n13759), .ZN(n13763) );
  INV_X1 U17100 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21496) );
  NOR3_X1 U17101 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n21496), .ZN(n13762) );
  NOR4_X1 U17102 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_2__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13761) );
  NAND4_X1 U17103 ( .A1(n15135), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13762), .A4(
        n13761), .ZN(U214) );
  NOR2_X1 U17104 ( .A1(n16714), .A2(n13763), .ZN(n17323) );
  NAND2_X1 U17105 ( .A1(n17323), .A2(U214), .ZN(U212) );
  NOR2_X1 U17106 ( .A1(n16927), .A2(n9624), .ZN(n18493) );
  NAND2_X1 U17107 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18493), .ZN(
        n17448) );
  OAI21_X1 U17108 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18493), .A(
        n17448), .ZN(n13764) );
  INV_X1 U17109 ( .A(n13764), .ZN(n18519) );
  NAND2_X1 U17110 ( .A1(n17308), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13765) );
  XNOR2_X2 U17111 ( .A(n13765), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14217) );
  INV_X1 U17112 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17634) );
  NAND2_X1 U17113 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18596), .ZN(
        n17647) );
  NOR2_X1 U17114 ( .A1(n17634), .A2(n17647), .ZN(n18570) );
  NAND2_X1 U17115 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18570), .ZN(
        n17618) );
  NOR2_X1 U17116 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17618), .ZN(
        n17597) );
  AND2_X1 U17117 ( .A1(n17597), .A2(n18493), .ZN(n13766) );
  NAND3_X1 U17118 ( .A1(n21628), .A2(n19452), .A3(n19571), .ZN(n19461) );
  NOR2_X2 U17119 ( .A1(n19451), .A2(n19461), .ZN(n17784) );
  AOI211_X1 U17120 ( .C1(n18519), .C2(n13767), .A(n17446), .B(n19459), .ZN(
        n13784) );
  NAND2_X1 U17121 ( .A1(n17792), .A2(n17787), .ZN(n17785) );
  NAND2_X1 U17122 ( .A1(n17759), .A2(n17754), .ZN(n17753) );
  NAND2_X1 U17123 ( .A1(n17735), .A2(n17734), .ZN(n17731) );
  NOR2_X2 U17124 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17731), .ZN(n17710) );
  NAND2_X1 U17125 ( .A1(n17710), .A2(n17705), .ZN(n17685) );
  NOR2_X2 U17126 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17685), .ZN(n17684) );
  NAND2_X1 U17127 ( .A1(n17684), .A2(n17675), .ZN(n17674) );
  NOR2_X2 U17128 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17674), .ZN(n17661) );
  NAND2_X1 U17129 ( .A1(n17661), .A2(n17653), .ZN(n17650) );
  INV_X1 U17130 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17627) );
  NAND2_X1 U17131 ( .A1(n17632), .A2(n17627), .ZN(n17626) );
  NAND2_X1 U17132 ( .A1(n17609), .A2(n17605), .ZN(n17604) );
  NOR2_X2 U17133 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17604), .ZN(n17588) );
  INV_X1 U17134 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17581) );
  NAND2_X1 U17135 ( .A1(n17588), .A2(n17581), .ZN(n17580) );
  NOR2_X2 U17136 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17580), .ZN(n17568) );
  INV_X1 U17137 ( .A(n13768), .ZN(n13769) );
  NAND2_X1 U17138 ( .A1(n19001), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n13775) );
  AOI211_X4 U17139 ( .C1(n19571), .C2(n19572), .A(n13778), .B(n13775), .ZN(
        n17786) );
  AOI211_X1 U17140 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17580), .A(n17568), .B(
        n17811), .ZN(n13783) );
  INV_X1 U17141 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n18517) );
  INV_X1 U17142 ( .A(n19456), .ZN(n17416) );
  NOR2_X1 U17143 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19552), .ZN(n19318) );
  NOR2_X1 U17144 ( .A1(n17416), .A2(n19454), .ZN(n19440) );
  OR2_X1 U17145 ( .A1(n17784), .A2(n18954), .ZN(n13771) );
  OR2_X1 U17146 ( .A1(n19440), .A2(n13771), .ZN(n13772) );
  NAND2_X2 U17147 ( .A1(n19583), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19538) );
  NOR2_X1 U17148 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19463) );
  INV_X1 U17149 ( .A(n19463), .ZN(n13773) );
  NAND3_X1 U17150 ( .A1(n19479), .A2(n19538), .A3(n13773), .ZN(n19569) );
  INV_X1 U17151 ( .A(n19572), .ZN(n19467) );
  AOI211_X1 U17152 ( .C1(n19569), .C2(n19570), .A(n19467), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13777) );
  INV_X1 U17153 ( .A(n13778), .ZN(n13774) );
  NAND2_X1 U17154 ( .A1(n13775), .A2(n13774), .ZN(n13776) );
  INV_X1 U17155 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17821) );
  OAI22_X1 U17156 ( .A1(n18517), .A2(n17791), .B1(n17812), .B2(n17821), .ZN(
        n13782) );
  NAND2_X1 U17157 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n13779) );
  INV_X1 U17158 ( .A(n13777), .ZN(n19441) );
  INV_X1 U17159 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19504) );
  INV_X1 U17160 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19488) );
  INV_X1 U17161 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19485) );
  NAND3_X1 U17162 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17758) );
  NOR3_X1 U17163 ( .A1(n19488), .A2(n19485), .A3(n17758), .ZN(n17711) );
  NAND4_X1 U17164 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17711), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n17690) );
  NAND3_X1 U17165 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(P3_REIP_REG_10__SCAN_IN), 
        .A3(P3_REIP_REG_9__SCAN_IN), .ZN(n17644) );
  NOR2_X1 U17166 ( .A1(n17690), .A2(n17644), .ZN(n17664) );
  NAND2_X1 U17167 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17664), .ZN(n17631) );
  NOR2_X1 U17168 ( .A1(n17712), .A2(n17608), .ZN(n17625) );
  NAND4_X1 U17169 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .A4(n17625), .ZN(n17594) );
  NOR2_X1 U17170 ( .A1(n13779), .A2(n17594), .ZN(n13780) );
  INV_X1 U17171 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19510) );
  INV_X1 U17172 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19507) );
  INV_X1 U17173 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19505) );
  NOR4_X1 U17174 ( .A1(n17608), .A2(n19510), .A3(n19507), .A4(n19505), .ZN(
        n17572) );
  INV_X1 U17175 ( .A(n13779), .ZN(n17573) );
  AND3_X1 U17176 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n17572), .A3(n17573), 
        .ZN(n17549) );
  OAI21_X1 U17177 ( .B1(n17712), .B2(n17549), .A(n17816), .ZN(n17566) );
  MUX2_X1 U17178 ( .A(n13780), .B(n17566), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n13781) );
  AND2_X1 U17179 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14151), .ZN(n16842) );
  NAND2_X1 U17180 ( .A1(n20392), .A2(n13787), .ZN(n16835) );
  INV_X1 U17181 ( .A(n16835), .ZN(n14680) );
  NAND2_X1 U17182 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20392), .ZN(n20484) );
  NOR2_X1 U17183 ( .A1(n20480), .A2(n20484), .ZN(n16840) );
  NOR3_X1 U17184 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n13785) );
  NOR4_X1 U17185 ( .A1(n16842), .A2(n14680), .A3(n16840), .A4(n13785), .ZN(
        P2_U3178) );
  OR2_X1 U17186 ( .A1(n13795), .A2(n19833), .ZN(n19787) );
  AND2_X1 U17187 ( .A1(n20382), .A2(n13787), .ZN(n13796) );
  AOI211_X1 U17188 ( .C1(P2_MEMORYFETCH_REG_SCAN_IN), .C2(n19787), .A(n13796), 
        .B(n14684), .ZN(n13789) );
  INV_X1 U17189 ( .A(n13789), .ZN(P2_U2814) );
  NOR2_X1 U17190 ( .A1(n13791), .A2(n13790), .ZN(n13792) );
  NAND2_X1 U17191 ( .A1(n13793), .A2(n13792), .ZN(n16822) );
  AND2_X1 U17192 ( .A1(n16822), .A2(n13810), .ZN(n20616) );
  OAI21_X1 U17193 ( .B1(n20616), .B2(n13812), .A(n13794), .ZN(P2_U2819) );
  INV_X1 U17194 ( .A(n19594), .ZN(n13798) );
  OAI21_X1 U17195 ( .B1(n13796), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n13798), 
        .ZN(n13797) );
  OAI21_X1 U17196 ( .B1(n13799), .B2(n13798), .A(n13797), .ZN(P2_U3612) );
  AOI22_X1 U17197 ( .A1(P2_EAX_REG_6__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13801) );
  NAND3_X1 U17198 ( .A1(n14684), .A2(n20480), .A3(n15871), .ZN(n13876) );
  NAND2_X1 U17199 ( .A1(n16713), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13800) );
  OAI21_X1 U17200 ( .B1(n16713), .B2(n19020), .A(n13800), .ZN(n16734) );
  NAND2_X1 U17201 ( .A1(n19909), .A2(n16734), .ZN(n13856) );
  NAND2_X1 U17202 ( .A1(n13801), .A2(n13856), .ZN(P2_U2973) );
  AND2_X1 U17203 ( .A1(n21349), .A2(n21403), .ZN(n14878) );
  AOI21_X1 U17204 ( .B1(n13802), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n14878), 
        .ZN(n13803) );
  NAND2_X1 U17205 ( .A1(n14139), .A2(n13803), .ZN(P1_U2801) );
  OR2_X1 U17206 ( .A1(n19833), .A2(n14616), .ZN(n13809) );
  INV_X1 U17207 ( .A(n13804), .ZN(n13805) );
  NOR2_X1 U17208 ( .A1(n13806), .A2(n13805), .ZN(n13807) );
  OAI211_X1 U17209 ( .C1(n19836), .C2(n13809), .A(n13808), .B(n13807), .ZN(
        n16825) );
  NAND2_X1 U17210 ( .A1(n16825), .A2(n13810), .ZN(n13816) );
  INV_X1 U17211 ( .A(n16842), .ZN(n13811) );
  NAND2_X1 U17212 ( .A1(n9587), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13813) );
  NAND2_X1 U17213 ( .A1(n13811), .A2(n13813), .ZN(n16846) );
  NAND2_X1 U17214 ( .A1(n13813), .A2(n13812), .ZN(n13814) );
  NAND2_X1 U17215 ( .A1(n16846), .A2(n13814), .ZN(n13815) );
  NAND2_X1 U17216 ( .A1(n13816), .A2(n13815), .ZN(n16707) );
  NOR2_X1 U17217 ( .A1(n19833), .A2(n15871), .ZN(n16819) );
  INV_X1 U17218 ( .A(n20579), .ZN(n16705) );
  NOR2_X1 U17219 ( .A1(n16803), .A2(n16705), .ZN(n13817) );
  NAND3_X1 U17220 ( .A1(n16707), .A2(n16819), .A3(n13817), .ZN(n13818) );
  OAI21_X1 U17221 ( .B1(n16707), .B2(n12127), .A(n13818), .ZN(P2_U3595) );
  AOI22_X1 U17222 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13821) );
  INV_X1 U17223 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n13820) );
  NAND2_X1 U17224 ( .A1(n16713), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13819) );
  OAI21_X1 U17225 ( .B1(n16713), .B2(n13820), .A(n13819), .ZN(n16016) );
  NAND2_X1 U17226 ( .A1(n19909), .A2(n16016), .ZN(n13844) );
  NAND2_X1 U17227 ( .A1(n13821), .A2(n13844), .ZN(P2_U2961) );
  AOI22_X1 U17228 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13824) );
  INV_X1 U17229 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n13823) );
  NAND2_X1 U17230 ( .A1(n16713), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13822) );
  OAI21_X1 U17231 ( .B1(n16713), .B2(n13823), .A(n13822), .ZN(n16003) );
  NAND2_X1 U17232 ( .A1(n19909), .A2(n16003), .ZN(n13955) );
  NAND2_X1 U17233 ( .A1(n13824), .A2(n13955), .ZN(P2_U2979) );
  AOI22_X1 U17234 ( .A1(P2_EAX_REG_21__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13827) );
  INV_X1 U17235 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n13826) );
  NAND2_X1 U17236 ( .A1(n16713), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13825) );
  OAI21_X1 U17237 ( .B1(n16713), .B2(n13826), .A(n13825), .ZN(n16784) );
  NAND2_X1 U17238 ( .A1(n19909), .A2(n16784), .ZN(n13833) );
  NAND2_X1 U17239 ( .A1(n13827), .A2(n13833), .ZN(P2_U2957) );
  AOI22_X1 U17240 ( .A1(P2_EAX_REG_24__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13830) );
  INV_X1 U17241 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n13829) );
  NAND2_X1 U17242 ( .A1(n16713), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13828) );
  OAI21_X1 U17243 ( .B1(n16713), .B2(n13829), .A(n13828), .ZN(n16023) );
  NAND2_X1 U17244 ( .A1(n19909), .A2(n16023), .ZN(n13831) );
  NAND2_X1 U17245 ( .A1(n13830), .A2(n13831), .ZN(P2_U2960) );
  AOI22_X1 U17246 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_8__SCAN_IN), .ZN(n13832) );
  NAND2_X1 U17247 ( .A1(n13832), .A2(n13831), .ZN(P2_U2975) );
  AOI22_X1 U17248 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13834) );
  NAND2_X1 U17249 ( .A1(n13834), .A2(n13833), .ZN(P2_U2972) );
  AOI22_X1 U17250 ( .A1(P2_EAX_REG_23__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13837) );
  INV_X1 U17251 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n13836) );
  NAND2_X1 U17252 ( .A1(n16713), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13835) );
  OAI21_X1 U17253 ( .B1(n16713), .B2(n13836), .A(n13835), .ZN(n16739) );
  NAND2_X1 U17254 ( .A1(n19909), .A2(n16739), .ZN(n13846) );
  NAND2_X1 U17255 ( .A1(n13837), .A2(n13846), .ZN(P2_U2959) );
  AOI22_X1 U17256 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13840) );
  NAND2_X1 U17257 ( .A1(n16714), .A2(BUF2_REG_3__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U17258 ( .A1(n16713), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13838) );
  AND2_X1 U17259 ( .A1(n13839), .A2(n13838), .ZN(n19822) );
  NAND2_X1 U17260 ( .A1(n19909), .A2(n19995), .ZN(n13952) );
  NAND2_X1 U17261 ( .A1(n13840), .A2(n13952), .ZN(P2_U2970) );
  AOI22_X1 U17262 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13843) );
  INV_X1 U17263 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n13842) );
  NAND2_X1 U17264 ( .A1(n16713), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13841) );
  OAI21_X1 U17265 ( .B1(n16713), .B2(n13842), .A(n13841), .ZN(n14533) );
  NAND2_X1 U17266 ( .A1(n19909), .A2(n14533), .ZN(n13848) );
  NAND2_X1 U17267 ( .A1(n13843), .A2(n13848), .ZN(P2_U2963) );
  AOI22_X1 U17268 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13845) );
  NAND2_X1 U17269 ( .A1(n13845), .A2(n13844), .ZN(P2_U2976) );
  AOI22_X1 U17270 ( .A1(P2_EAX_REG_7__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13847) );
  NAND2_X1 U17271 ( .A1(n13847), .A2(n13846), .ZN(P2_U2974) );
  AOI22_X1 U17272 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U17273 ( .A1(n13849), .A2(n13848), .ZN(P2_U2978) );
  INV_X1 U17274 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19864) );
  INV_X1 U17275 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n19013) );
  NAND2_X1 U17276 ( .A1(n16713), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13851) );
  OAI21_X1 U17277 ( .B1(n16713), .B2(n19013), .A(n13851), .ZN(n20001) );
  NAND2_X1 U17278 ( .A1(n19909), .A2(n20001), .ZN(n13859) );
  NAND2_X1 U17279 ( .A1(n13961), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13852) );
  OAI211_X1 U17280 ( .C1(n19834), .C2(n19864), .A(n13859), .B(n13852), .ZN(
        P2_U2956) );
  INV_X1 U17281 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n21632) );
  INV_X1 U17282 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n19005) );
  NAND2_X1 U17283 ( .A1(n16713), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13853) );
  OAI21_X1 U17284 ( .B1(n16713), .B2(n19005), .A(n13853), .ZN(n19989) );
  NAND2_X1 U17285 ( .A1(n19909), .A2(n19989), .ZN(n13962) );
  NAND2_X1 U17286 ( .A1(n13961), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13854) );
  OAI211_X1 U17287 ( .C1(n19834), .C2(n21632), .A(n13962), .B(n13854), .ZN(
        P2_U2954) );
  INV_X1 U17288 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19860) );
  NAND2_X1 U17289 ( .A1(n13961), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13855) );
  OAI211_X1 U17290 ( .C1(n19834), .C2(n19860), .A(n13856), .B(n13855), .ZN(
        P2_U2958) );
  INV_X1 U17291 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n21566) );
  MUX2_X1 U17292 ( .A(BUF2_REG_0__SCAN_IN), .B(BUF1_REG_0__SCAN_IN), .S(n16713), .Z(n19797) );
  NAND2_X1 U17293 ( .A1(n19909), .A2(n19797), .ZN(n13861) );
  NAND2_X1 U17294 ( .A1(n13961), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13857) );
  OAI211_X1 U17295 ( .C1(n19834), .C2(n21566), .A(n13861), .B(n13857), .ZN(
        P2_U2952) );
  INV_X1 U17296 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19895) );
  NAND2_X1 U17297 ( .A1(n13961), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13858) );
  OAI211_X1 U17298 ( .C1(n19834), .C2(n19895), .A(n13859), .B(n13858), .ZN(
        P2_U2971) );
  NAND2_X1 U17299 ( .A1(n13961), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13860) );
  OAI211_X1 U17300 ( .C1(n19834), .C2(n12181), .A(n13861), .B(n13860), .ZN(
        P2_U2967) );
  NOR3_X1 U17301 ( .A1(n13862), .A2(n12959), .A3(n17186), .ZN(n21500) );
  NAND2_X1 U17302 ( .A1(n13867), .A2(n12901), .ZN(n13863) );
  AOI22_X1 U17303 ( .A1(n14037), .A2(n14990), .B1(n13022), .B2(n13863), .ZN(
        n20625) );
  OAI21_X1 U17304 ( .B1(n21500), .B2(n21501), .A(n20625), .ZN(n17156) );
  AND2_X1 U17305 ( .A1(n17156), .A2(n14043), .ZN(n20632) );
  INV_X1 U17306 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17157) );
  INV_X1 U17307 ( .A(n14036), .ZN(n13865) );
  MUX2_X1 U17308 ( .A(n13865), .B(n13864), .S(n14037), .Z(n13871) );
  INV_X1 U17309 ( .A(n13022), .ZN(n13869) );
  NOR2_X1 U17310 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  AOI21_X1 U17311 ( .B1(n14037), .B2(n13869), .A(n13868), .ZN(n13870) );
  NAND2_X1 U17312 ( .A1(n13871), .A2(n13870), .ZN(n17158) );
  NAND2_X1 U17313 ( .A1(n20632), .A2(n17158), .ZN(n13872) );
  OAI21_X1 U17314 ( .B1(n20632), .B2(n17157), .A(n13872), .ZN(P1_U3484) );
  INV_X1 U17315 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14181) );
  NOR2_X1 U17316 ( .A1(n16714), .A2(n14181), .ZN(n13873) );
  AOI21_X1 U17317 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n16714), .A(n13873), .ZN(
        n14325) );
  INV_X1 U17318 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13875) );
  OAI222_X1 U17319 ( .A1(n19834), .A2(n19873), .B1(n13876), .B2(n14325), .C1(
        n13875), .C2(n13874), .ZN(P2_U2982) );
  XNOR2_X1 U17320 ( .A(n13877), .B(n13878), .ZN(n19752) );
  INV_X1 U17321 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19891) );
  INV_X1 U17322 ( .A(n19798), .ZN(n13880) );
  INV_X1 U17323 ( .A(n16734), .ZN(n13881) );
  OAI222_X1 U17324 ( .A1(n19752), .A2(n16096), .B1(n19891), .B2(n19832), .C1(
        n19821), .C2(n13881), .ZN(P2_U2913) );
  NAND2_X1 U17325 ( .A1(n13883), .A2(n13884), .ZN(n13885) );
  NAND2_X1 U17326 ( .A1(n13882), .A2(n13885), .ZN(n19725) );
  INV_X1 U17327 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19887) );
  INV_X1 U17328 ( .A(n16023), .ZN(n13886) );
  OAI222_X1 U17329 ( .A1(n19725), .A2(n16096), .B1(n19832), .B2(n19887), .C1(
        n19821), .C2(n13886), .ZN(P2_U2911) );
  OAI21_X1 U17330 ( .B1(n13888), .B2(n13887), .A(n13883), .ZN(n19739) );
  INV_X1 U17331 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19889) );
  INV_X1 U17332 ( .A(n16739), .ZN(n13889) );
  OAI222_X1 U17333 ( .A1(n19739), .A2(n16096), .B1(n19889), .B2(n19832), .C1(
        n19821), .C2(n13889), .ZN(P2_U2912) );
  XNOR2_X1 U17334 ( .A(n13890), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13902) );
  INV_X1 U17335 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19606) );
  OR2_X1 U17336 ( .A1(n19701), .A2(n19606), .ZN(n13898) );
  OAI21_X1 U17337 ( .B1(n16639), .B2(n13909), .A(n13898), .ZN(n13895) );
  OR2_X1 U17338 ( .A1(n15852), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13891) );
  NAND2_X1 U17339 ( .A1(n13968), .A2(n13891), .ZN(n13899) );
  XNOR2_X1 U17340 ( .A(n13893), .B(n13892), .ZN(n15851) );
  OAI22_X1 U17341 ( .A1(n16648), .A2(n13899), .B1(n19959), .B2(n15851), .ZN(
        n13894) );
  AOI211_X1 U17342 ( .C1(n16603), .C2(n13902), .A(n13895), .B(n13894), .ZN(
        n13897) );
  MUX2_X1 U17343 ( .A(n14559), .B(n14046), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13896) );
  NAND2_X1 U17344 ( .A1(n13897), .A2(n13896), .ZN(P2_U3046) );
  INV_X1 U17345 ( .A(n13898), .ZN(n13901) );
  NOR2_X1 U17346 ( .A1(n17292), .A2(n13899), .ZN(n13900) );
  AOI211_X1 U17347 ( .C1(n13902), .C2(n16335), .A(n13901), .B(n13900), .ZN(
        n13905) );
  OAI21_X1 U17348 ( .B1(n17289), .B2(n13903), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13904) );
  OAI211_X1 U17349 ( .C1(n19928), .C2(n13909), .A(n13905), .B(n13904), .ZN(
        P2_U3014) );
  NAND2_X1 U17350 ( .A1(n15871), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13906) );
  AND4_X1 U17351 ( .A1(n13906), .A2(n16735), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n20581), .ZN(n13907) );
  MUX2_X1 U17352 ( .A(n13909), .B(n13908), .S(n9574), .Z(n13910) );
  OAI21_X1 U17353 ( .B1(n16745), .B2(n15975), .A(n13910), .ZN(P2_U2887) );
  INV_X1 U17354 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19885) );
  XNOR2_X1 U17355 ( .A(n13882), .B(n13911), .ZN(n16583) );
  INV_X1 U17356 ( .A(n16016), .ZN(n13912) );
  OAI222_X1 U17357 ( .A1(n19832), .A2(n19885), .B1(n16583), .B2(n16096), .C1(
        n13912), .C2(n19821), .ZN(P2_U2910) );
  NAND3_X1 U17358 ( .A1(n13915), .A2(n13914), .A3(n13913), .ZN(n13916) );
  NOR2_X1 U17359 ( .A1(n13917), .A2(n13916), .ZN(n13918) );
  NAND2_X1 U17360 ( .A1(n17271), .A2(n13918), .ZN(n15591) );
  NAND2_X1 U17361 ( .A1(n21088), .A2(n15591), .ZN(n13934) );
  NAND2_X1 U17362 ( .A1(n15593), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13919) );
  NAND2_X1 U17363 ( .A1(n13919), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13920) );
  NAND2_X1 U17364 ( .A1(n13921), .A2(n13920), .ZN(n13935) );
  NAND2_X1 U17365 ( .A1(n14039), .A2(n13935), .ZN(n13931) );
  INV_X1 U17366 ( .A(n13922), .ZN(n13923) );
  NOR2_X1 U17367 ( .A1(n14036), .A2(n13923), .ZN(n13991) );
  OR3_X1 U17368 ( .A1(n13991), .A2(n13925), .A3(n13924), .ZN(n13930) );
  NAND2_X1 U17369 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13926) );
  NAND2_X1 U17370 ( .A1(n10948), .A2(n13926), .ZN(n13927) );
  NAND3_X1 U17371 ( .A1(n17140), .A2(n13928), .A3(n13927), .ZN(n13929) );
  OAI211_X1 U17372 ( .C1(n15591), .C2(n13931), .A(n13930), .B(n13929), .ZN(
        n13932) );
  INV_X1 U17373 ( .A(n13932), .ZN(n13933) );
  NAND2_X1 U17374 ( .A1(n13934), .A2(n13933), .ZN(n14406) );
  AOI22_X1 U17375 ( .A1(n14406), .A2(n20624), .B1(n17173), .B2(n13935), .ZN(
        n13947) );
  OAI211_X1 U17376 ( .C1(n17140), .C2(n13936), .A(n17186), .B(n21419), .ZN(
        n13938) );
  NAND2_X1 U17377 ( .A1(n13938), .A2(n13937), .ZN(n13939) );
  MUX2_X1 U17378 ( .A(n13939), .B(n14036), .S(n14037), .Z(n13944) );
  INV_X1 U17379 ( .A(n13940), .ZN(n13943) );
  OAI21_X1 U17380 ( .B1(n20824), .B2(n15003), .A(n13941), .ZN(n13942) );
  INV_X1 U17381 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21646) );
  NAND2_X1 U17382 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n17280), .ZN(n17285) );
  NOR2_X1 U17383 ( .A1(n21646), .A2(n17285), .ZN(n13945) );
  AOI21_X1 U17384 ( .B1(n17143), .B2(n14043), .A(n13945), .ZN(n17273) );
  NAND2_X1 U17385 ( .A1(n10276), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13946) );
  NAND2_X1 U17386 ( .A1(n17273), .A2(n13946), .ZN(n17276) );
  MUX2_X1 U17387 ( .A(n10948), .B(n13947), .S(n17276), .Z(n13948) );
  INV_X1 U17388 ( .A(n13948), .ZN(P1_U3469) );
  AOI22_X1 U17389 ( .A1(P2_EAX_REG_17__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13951) );
  INV_X1 U17390 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n13950) );
  NAND2_X1 U17391 ( .A1(n16713), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13949) );
  OAI21_X1 U17392 ( .B1(n16713), .B2(n13950), .A(n13949), .ZN(n19983) );
  NAND2_X1 U17393 ( .A1(n19909), .A2(n19983), .ZN(n13959) );
  NAND2_X1 U17394 ( .A1(n13951), .A2(n13959), .ZN(P2_U2953) );
  AOI22_X1 U17395 ( .A1(P2_EAX_REG_19__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13953) );
  NAND2_X1 U17396 ( .A1(n13953), .A2(n13952), .ZN(P2_U2955) );
  AOI22_X1 U17397 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13954) );
  NAND2_X1 U17398 ( .A1(n19909), .A2(n14186), .ZN(n13957) );
  NAND2_X1 U17399 ( .A1(n13954), .A2(n13957), .ZN(P2_U2965) );
  AOI22_X1 U17400 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13956) );
  NAND2_X1 U17401 ( .A1(n13956), .A2(n13955), .ZN(P2_U2964) );
  AOI22_X1 U17402 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13958) );
  NAND2_X1 U17403 ( .A1(n13958), .A2(n13957), .ZN(P2_U2980) );
  AOI22_X1 U17404 ( .A1(P2_EAX_REG_1__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13960) );
  NAND2_X1 U17405 ( .A1(n13960), .A2(n13959), .ZN(P2_U2968) );
  AOI22_X1 U17406 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(n13850), .B1(n13961), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13963) );
  NAND2_X1 U17407 ( .A1(n13963), .A2(n13962), .ZN(P2_U2969) );
  INV_X1 U17408 ( .A(n14056), .ZN(n14047) );
  AOI211_X1 U17409 ( .C1(n14632), .C2(n14633), .A(n14047), .B(n14559), .ZN(
        n13976) );
  OR2_X1 U17410 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  NAND2_X1 U17411 ( .A1(n13967), .A2(n13966), .ZN(n16086) );
  XNOR2_X1 U17412 ( .A(n13968), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13969) );
  XNOR2_X1 U17413 ( .A(n13969), .B(n15846), .ZN(n14019) );
  AOI22_X1 U17414 ( .A1(n16645), .A2(n16086), .B1(n19962), .B2(n14019), .ZN(
        n13970) );
  NAND2_X1 U17415 ( .A1(n16341), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14015) );
  OAI211_X1 U17416 ( .C1(n16639), .C2(n15847), .A(n13970), .B(n14015), .ZN(
        n13975) );
  OR2_X1 U17417 ( .A1(n13971), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13972) );
  NAND2_X1 U17418 ( .A1(n13973), .A2(n13972), .ZN(n14016) );
  OAI22_X1 U17419 ( .A1(n19967), .A2(n14016), .B1(n14633), .B2(n14046), .ZN(
        n13974) );
  OR3_X1 U17420 ( .A1(n13976), .A2(n13975), .A3(n13974), .ZN(P2_U3045) );
  INV_X1 U17421 ( .A(n13977), .ZN(n13981) );
  NAND2_X1 U17422 ( .A1(n13979), .A2(n13978), .ZN(n13980) );
  NAND2_X1 U17423 ( .A1(n13981), .A2(n13980), .ZN(n16570) );
  INV_X1 U17424 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n21539) );
  NAND2_X1 U17425 ( .A1(n16713), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13982) );
  OAI21_X1 U17426 ( .B1(n16713), .B2(n21539), .A(n13982), .ZN(n19906) );
  AOI22_X1 U17427 ( .A1(n19824), .A2(n19906), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19813), .ZN(n13983) );
  OAI21_X1 U17428 ( .B1(n16570), .B2(n16096), .A(n13983), .ZN(P2_U2909) );
  XNOR2_X1 U17429 ( .A(n15593), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13985) );
  INV_X1 U17430 ( .A(n13985), .ZN(n13993) );
  INV_X1 U17431 ( .A(n13984), .ZN(n15005) );
  NAND2_X1 U17432 ( .A1(n15005), .A2(n15591), .ZN(n13990) );
  XNOR2_X1 U17433 ( .A(n10934), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13988) );
  NOR3_X1 U17434 ( .A1(n15591), .A2(n13986), .A3(n13985), .ZN(n13987) );
  AOI21_X1 U17435 ( .B1(n17140), .B2(n13988), .A(n13987), .ZN(n13989) );
  OAI211_X1 U17436 ( .C1(n13993), .C2(n13991), .A(n13990), .B(n13989), .ZN(
        n14405) );
  INV_X1 U17437 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15426) );
  NOR2_X1 U17438 ( .A1(n21403), .A2(n15426), .ZN(n15601) );
  INV_X1 U17439 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13992) );
  AOI22_X1 U17440 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14473), .B2(n13992), .ZN(
        n15599) );
  AOI222_X1 U17441 ( .A1(n14405), .A2(n20624), .B1(n15601), .B2(n15599), .C1(
        n13993), .C2(n17173), .ZN(n13994) );
  MUX2_X1 U17442 ( .A(n10934), .B(n13994), .S(n17276), .Z(n13995) );
  INV_X1 U17443 ( .A(n13995), .ZN(P1_U3472) );
  INV_X1 U17444 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14001) );
  NAND2_X1 U17445 ( .A1(n14140), .A2(n17186), .ZN(n13996) );
  OR2_X1 U17446 ( .A1(n13022), .A2(n13996), .ZN(n17166) );
  INV_X1 U17447 ( .A(n17166), .ZN(n13997) );
  AOI21_X1 U17448 ( .B1(n17140), .B2(n17186), .A(n13997), .ZN(n13998) );
  NAND2_X1 U17449 ( .A1(n10276), .A2(n17280), .ZN(n20720) );
  INV_X2 U17450 ( .A(n20720), .ZN(n20738) );
  NOR2_X4 U17451 ( .A1(n20718), .A2(n20738), .ZN(n20737) );
  AOI22_X1 U17452 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n14000) );
  OAI21_X1 U17453 ( .B1(n14001), .B2(n14248), .A(n14000), .ZN(P1_U2908) );
  AOI22_X1 U17454 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14002) );
  OAI21_X1 U17455 ( .B1(n15138), .B2(n14248), .A(n14002), .ZN(P1_U2911) );
  AOI22_X1 U17456 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14003) );
  OAI21_X1 U17457 ( .B1(n15142), .B2(n14248), .A(n14003), .ZN(P1_U2912) );
  INV_X1 U17458 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17459 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n14004) );
  OAI21_X1 U17460 ( .B1(n14005), .B2(n14248), .A(n14004), .ZN(P1_U2909) );
  INV_X1 U17461 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17462 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14006) );
  OAI21_X1 U17463 ( .B1(n14007), .B2(n14248), .A(n14006), .ZN(P1_U2910) );
  AOI22_X1 U17464 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n14008) );
  OAI21_X1 U17465 ( .B1(n14714), .B2(n14248), .A(n14008), .ZN(P1_U2907) );
  INV_X1 U17466 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n14010) );
  AOI22_X1 U17467 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n14009) );
  OAI21_X1 U17468 ( .B1(n14010), .B2(n14248), .A(n14009), .ZN(P1_U2906) );
  MUX2_X1 U17469 ( .A(n14013), .B(n15847), .S(n16002), .Z(n14014) );
  OAI21_X1 U17470 ( .B1(n19968), .B2(n15975), .A(n14014), .ZN(P2_U2886) );
  OAI21_X1 U17471 ( .B1(n19941), .B2(n14016), .A(n14015), .ZN(n14018) );
  MUX2_X1 U17472 ( .A(n19917), .B(n17289), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n14017) );
  AOI211_X1 U17473 ( .C1(n14019), .C2(n19936), .A(n14018), .B(n14017), .ZN(
        n14020) );
  OAI21_X1 U17474 ( .B1(n15847), .B2(n19928), .A(n14020), .ZN(P2_U3013) );
  OAI21_X1 U17475 ( .B1(n13977), .B2(n14023), .A(n14022), .ZN(n19707) );
  INV_X1 U17476 ( .A(n14533), .ZN(n14024) );
  INV_X1 U17477 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U17478 ( .A1(n19707), .A2(n16096), .B1(n14024), .B2(n19821), .C1(
        n19881), .C2(n19832), .ZN(P2_U2908) );
  INV_X1 U17479 ( .A(n14025), .ZN(n14028) );
  OAI21_X1 U17480 ( .B1(n14028), .B2(n14027), .A(n14026), .ZN(n15030) );
  NOR2_X1 U17481 ( .A1(n14030), .A2(n10601), .ZN(n14029) );
  NAND2_X1 U17482 ( .A1(n14030), .A2(n17230), .ZN(n15177) );
  NAND2_X1 U17483 ( .A1(n14509), .A2(DATAI_0_), .ZN(n14033) );
  NAND2_X1 U17484 ( .A1(n15135), .A2(BUF1_REG_0__SCAN_IN), .ZN(n14032) );
  AND2_X1 U17485 ( .A1(n14033), .A2(n14032), .ZN(n15176) );
  INV_X1 U17486 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U17487 ( .A1(n15030), .A2(n15195), .B1(n17225), .B2(n15176), .C1(
        n17230), .C2(n20741), .ZN(P1_U2904) );
  NOR2_X1 U17488 ( .A1(n14733), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14034) );
  OR2_X1 U17489 ( .A1(n14035), .A2(n14034), .ZN(n15023) );
  NAND2_X1 U17490 ( .A1(n14037), .A2(n14036), .ZN(n14042) );
  INV_X1 U17491 ( .A(n14038), .ZN(n14040) );
  NAND4_X1 U17492 ( .A1(n14040), .A2(n10916), .A3(n12959), .A4(n14039), .ZN(
        n14041) );
  OAI222_X1 U17493 ( .A1(n15023), .A2(n15105), .B1(n12938), .B2(n15104), .C1(
        n15030), .C2(n15079), .ZN(P1_U2872) );
  OAI21_X1 U17494 ( .B1(n14554), .B2(n14047), .A(n14046), .ZN(n14069) );
  OR2_X1 U17495 ( .A1(n14051), .A2(n14050), .ZN(n14052) );
  NAND2_X1 U17496 ( .A1(n14049), .A2(n14052), .ZN(n20592) );
  XNOR2_X1 U17497 ( .A(n14054), .B(n14053), .ZN(n19942) );
  OAI22_X1 U17498 ( .A1(n19967), .A2(n19942), .B1(n14056), .B2(n14055), .ZN(
        n14058) );
  NAND2_X1 U17499 ( .A1(n16341), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19947) );
  INV_X1 U17500 ( .A(n19947), .ZN(n14057) );
  AOI211_X1 U17501 ( .C1(n16645), .C2(n20592), .A(n14058), .B(n14057), .ZN(
        n14062) );
  OR2_X1 U17502 ( .A1(n14060), .A2(n14059), .ZN(n19937) );
  NAND3_X1 U17503 ( .A1(n19962), .A2(n19935), .A3(n19937), .ZN(n14061) );
  OAI211_X1 U17504 ( .C1(n16639), .C2(n14063), .A(n14062), .B(n14061), .ZN(
        n14068) );
  AOI21_X1 U17505 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n14067) );
  AOI211_X1 U17506 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n14069), .A(
        n14068), .B(n14067), .ZN(n14070) );
  INV_X1 U17507 ( .A(n14070), .ZN(P2_U3044) );
  OAI21_X1 U17508 ( .B1(n14072), .B2(n14071), .A(n14250), .ZN(n15022) );
  XNOR2_X1 U17509 ( .A(n14073), .B(n12959), .ZN(n15583) );
  AOI22_X1 U17510 ( .A1(n15097), .A2(n15583), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15096), .ZN(n14074) );
  OAI21_X1 U17511 ( .B1(n15022), .B2(n15099), .A(n14074), .ZN(P1_U2871) );
  NAND3_X1 U17512 ( .A1(n14076), .A2(n14075), .A3(n15426), .ZN(n14077) );
  AOI21_X1 U17513 ( .B1(n14502), .B2(n14078), .A(n14077), .ZN(n14080) );
  INV_X1 U17514 ( .A(n14079), .ZN(n14436) );
  NOR2_X1 U17515 ( .A1(n14080), .A2(n14436), .ZN(n14129) );
  AND2_X1 U17516 ( .A1(n20786), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n14133) );
  INV_X1 U17517 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14081) );
  AOI21_X1 U17518 ( .B1(n15271), .B2(n14082), .A(n14081), .ZN(n14083) );
  AOI211_X1 U17519 ( .C1(n14129), .C2(n20780), .A(n14133), .B(n14083), .ZN(
        n14084) );
  OAI21_X1 U17520 ( .B1(n17244), .B2(n15030), .A(n14084), .ZN(P1_U2999) );
  NAND2_X1 U17521 ( .A1(n14509), .A2(DATAI_1_), .ZN(n14086) );
  NAND2_X1 U17522 ( .A1(n15135), .A2(BUF1_REG_1__SCAN_IN), .ZN(n14085) );
  AND2_X1 U17523 ( .A1(n14086), .A2(n14085), .ZN(n20821) );
  OAI222_X1 U17524 ( .A1(n15022), .A2(n15195), .B1(n17225), .B2(n20821), .C1(
        n17230), .C2(n10980), .ZN(P1_U2903) );
  INV_X1 U17525 ( .A(n19399), .ZN(n16991) );
  OAI21_X1 U17526 ( .B1(n14089), .B2(n14088), .A(n14087), .ZN(n18726) );
  INV_X1 U17527 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14356) );
  NOR2_X1 U17528 ( .A1(n9877), .A2(n9830), .ZN(n16943) );
  INV_X1 U17529 ( .A(n16943), .ZN(n14192) );
  OAI21_X1 U17530 ( .B1(n9830), .B2(n14356), .A(n9877), .ZN(n16941) );
  OAI21_X1 U17531 ( .B1(n14356), .B2(n14192), .A(n16941), .ZN(n14092) );
  OAI21_X1 U17532 ( .B1(n18926), .B2(n14356), .A(n18927), .ZN(n16950) );
  INV_X1 U17533 ( .A(n16950), .ZN(n14193) );
  NOR3_X1 U17534 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n9830), .A3(
        n14193), .ZN(n14091) );
  NOR2_X1 U17535 ( .A1(n18926), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16976) );
  INV_X1 U17536 ( .A(n16976), .ZN(n14190) );
  INV_X1 U17537 ( .A(n18926), .ZN(n18905) );
  NOR2_X1 U17538 ( .A1(n18978), .A2(n18905), .ZN(n18817) );
  AOI211_X1 U17539 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n14190), .A(
        n18817), .B(n9877), .ZN(n14090) );
  AOI211_X1 U17540 ( .C1(n19400), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14093) );
  OAI21_X1 U17541 ( .B1(n16991), .B2(n18726), .A(n14093), .ZN(n14116) );
  OAI221_X1 U17542 ( .B1(n14354), .B2(n14205), .C1(n14354), .C2(n18992), .A(
        n14094), .ZN(n14095) );
  NOR4_X1 U17543 ( .A1(n14098), .A2(n14097), .A3(n14096), .A4(n14095), .ZN(
        n14101) );
  INV_X1 U17544 ( .A(n14099), .ZN(n14100) );
  OAI21_X1 U17545 ( .B1(n17413), .B2(n14101), .A(n14100), .ZN(n14161) );
  AOI21_X1 U17546 ( .B1(n19569), .B2(n14102), .A(n19467), .ZN(n17420) );
  NAND4_X1 U17547 ( .A1(n19405), .A2(n14104), .A3(n19001), .A4(n19019), .ZN(
        n14108) );
  NAND2_X1 U17548 ( .A1(n14205), .A2(n14105), .ZN(n14106) );
  NAND2_X1 U17549 ( .A1(n19401), .A2(n14106), .ZN(n14107) );
  NAND3_X1 U17550 ( .A1(n10432), .A2(n14108), .A3(n14107), .ZN(n14109) );
  XNOR2_X1 U17551 ( .A(n14112), .B(n14111), .ZN(n18718) );
  INV_X1 U17552 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n14113) );
  OR2_X1 U17553 ( .A1(n18981), .A2(n14113), .ZN(n18724) );
  NOR2_X2 U17554 ( .A1(n18954), .A2(n18958), .ZN(n18976) );
  NAND2_X1 U17555 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18976), .ZN(
        n14114) );
  OAI211_X1 U17556 ( .C1(n18971), .C2(n18718), .A(n18724), .B(n14114), .ZN(
        n14115) );
  AOI21_X1 U17557 ( .B1(n14116), .B2(n18958), .A(n14115), .ZN(n14117) );
  INV_X1 U17558 ( .A(n14117), .ZN(P3_U2860) );
  AOI21_X1 U17559 ( .B1(n14119), .B2(n14022), .A(n10383), .ZN(n19696) );
  INV_X1 U17560 ( .A(n19696), .ZN(n14121) );
  INV_X1 U17561 ( .A(n16003), .ZN(n14120) );
  INV_X1 U17562 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19879) );
  OAI222_X1 U17563 ( .A1(n14121), .A2(n16096), .B1(n14120), .B2(n19821), .C1(
        n19879), .C2(n19832), .ZN(P2_U2907) );
  INV_X1 U17564 ( .A(n16933), .ZN(n14122) );
  AND2_X1 U17565 ( .A1(n14122), .A2(n16935), .ZN(n14277) );
  INV_X1 U17566 ( .A(n14277), .ZN(n14128) );
  AOI21_X1 U17567 ( .B1(n18927), .B2(n18958), .A(n14356), .ZN(n14125) );
  INV_X1 U17568 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n14123) );
  NOR2_X1 U17569 ( .A1(n18981), .A2(n14123), .ZN(n14273) );
  NOR2_X1 U17570 ( .A1(n18973), .A2(n14277), .ZN(n14124) );
  AOI211_X1 U17571 ( .C1(n14125), .C2(n18981), .A(n14273), .B(n14124), .ZN(
        n14127) );
  NOR2_X1 U17572 ( .A1(n19400), .A2(n18905), .ZN(n18857) );
  NOR3_X1 U17573 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18857), .A3(
        n18888), .ZN(n18975) );
  INV_X1 U17574 ( .A(n18975), .ZN(n14126) );
  OAI211_X1 U17575 ( .C1(n14128), .C2(n18971), .A(n14127), .B(n14126), .ZN(
        P3_U2862) );
  INV_X1 U17576 ( .A(n14129), .ZN(n14136) );
  INV_X1 U17577 ( .A(n15023), .ZN(n14134) );
  AOI21_X1 U17578 ( .B1(n20805), .B2(n15426), .A(n15533), .ZN(n15581) );
  INV_X1 U17579 ( .A(n14130), .ZN(n15452) );
  NOR3_X1 U17580 ( .A1(n20805), .A2(n15428), .A3(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14131) );
  AOI21_X1 U17581 ( .B1(n15581), .B2(n15452), .A(n14131), .ZN(n14132) );
  AOI211_X1 U17582 ( .C1(n14134), .C2(n20801), .A(n14133), .B(n14132), .ZN(
        n14135) );
  OAI21_X1 U17583 ( .B1(n20807), .B2(n14136), .A(n14135), .ZN(P1_U3031) );
  NAND2_X1 U17584 ( .A1(n20765), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n14143) );
  NOR2_X2 U17585 ( .A1(n20765), .A2(n14140), .ZN(n20757) );
  INV_X1 U17586 ( .A(DATAI_8_), .ZN(n14141) );
  MUX2_X1 U17587 ( .A(n14141), .B(n17354), .S(n15135), .Z(n15193) );
  INV_X1 U17588 ( .A(n15193), .ZN(n14142) );
  NAND2_X1 U17589 ( .A1(n20757), .A2(n14142), .ZN(n14144) );
  OAI211_X1 U17590 ( .C1(n14326), .C2(n15142), .A(n14143), .B(n14144), .ZN(
        P1_U2945) );
  INV_X1 U17591 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20728) );
  NAND2_X1 U17592 ( .A1(n20765), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n14145) );
  OAI211_X1 U17593 ( .C1(n14326), .C2(n20728), .A(n14145), .B(n14144), .ZN(
        P1_U2960) );
  NAND2_X1 U17594 ( .A1(n20382), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20589) );
  INV_X1 U17595 ( .A(n20589), .ZN(n14149) );
  INV_X1 U17596 ( .A(n20600), .ZN(n14147) );
  NOR2_X1 U17597 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  MUX2_X1 U17598 ( .A(n14149), .B(n14148), .S(n16744), .Z(n14150) );
  AOI21_X1 U17599 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n16086), .A(n14150), 
        .ZN(n14156) );
  NAND2_X1 U17600 ( .A1(n16835), .A2(n20597), .ZN(n14152) );
  NAND2_X1 U17601 ( .A1(n20615), .A2(n13812), .ZN(n14153) );
  NAND2_X1 U17602 ( .A1(n14153), .A2(n16842), .ZN(n14154) );
  NAND2_X1 U17603 ( .A1(n20183), .A2(n14154), .ZN(n20602) );
  INV_X1 U17604 ( .A(n20602), .ZN(n20605) );
  NAND2_X1 U17605 ( .A1(n20605), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14155) );
  OAI21_X1 U17606 ( .B1(n14156), .B2(n20605), .A(n14155), .ZN(P2_U3604) );
  NOR2_X1 U17607 ( .A1(n16745), .A2(n15851), .ZN(n16087) );
  XNOR2_X1 U17608 ( .A(n16744), .B(n16086), .ZN(n16088) );
  XOR2_X1 U17609 ( .A(n16087), .B(n16088), .Z(n14159) );
  AOI22_X1 U17610 ( .A1(n19823), .A2(n16086), .B1(n19813), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n14158) );
  NAND2_X1 U17611 ( .A1(n19824), .A2(n19983), .ZN(n14157) );
  OAI211_X1 U17612 ( .C1(n14159), .C2(n16062), .A(n14158), .B(n14157), .ZN(
        P2_U2918) );
  NAND2_X1 U17613 ( .A1(n19404), .A2(n19572), .ZN(n14165) );
  NAND2_X1 U17614 ( .A1(n19570), .A2(n18379), .ZN(n19442) );
  INV_X1 U17615 ( .A(n18322), .ZN(n14164) );
  NOR2_X1 U17616 ( .A1(n14209), .A2(n14161), .ZN(n14163) );
  NAND2_X1 U17617 ( .A1(n19401), .A2(n14162), .ZN(n14207) );
  INV_X1 U17618 ( .A(n19418), .ZN(n19427) );
  INV_X1 U17619 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n17424) );
  NAND3_X1 U17620 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_1__SCAN_IN), .ZN(n19551)
         );
  OAI22_X1 U17621 ( .A1(n19427), .A2(n19449), .B1(n17424), .B2(n19551), .ZN(
        n14166) );
  NOR2_X1 U17622 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18978), .ZN(
        n14355) );
  NAND2_X1 U17623 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14397) );
  OR2_X1 U17624 ( .A1(n14355), .A2(n14397), .ZN(n14169) );
  INV_X1 U17625 ( .A(n14389), .ZN(n14394) );
  NAND2_X1 U17626 ( .A1(n14394), .A2(n14167), .ZN(n14382) );
  NAND2_X1 U17627 ( .A1(n19400), .A2(n14382), .ZN(n14168) );
  AOI21_X1 U17628 ( .B1(n14169), .B2(n14168), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19414) );
  INV_X1 U17629 ( .A(n14397), .ZN(n14170) );
  AND2_X1 U17630 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n14170), .ZN(
        n14380) );
  OAI21_X1 U17631 ( .B1(n14380), .B2(n19412), .A(n18035), .ZN(n17779) );
  AOI22_X1 U17632 ( .A1(n19414), .A2(n19584), .B1(n19444), .B2(n17779), .ZN(
        n14180) );
  INV_X1 U17633 ( .A(n14171), .ZN(n14174) );
  AOI21_X1 U17634 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14391) );
  OR2_X1 U17635 ( .A1(n14391), .A2(n14380), .ZN(n14178) );
  OAI21_X1 U17636 ( .B1(n14175), .B2(n14392), .A(n14397), .ZN(n14176) );
  AND2_X1 U17637 ( .A1(n14176), .A2(n14382), .ZN(n14177) );
  NAND2_X1 U17638 ( .A1(n14178), .A2(n14177), .ZN(n19411) );
  AOI21_X1 U17639 ( .B1(n19584), .B2(n19411), .A(n14404), .ZN(n14179) );
  OAI22_X1 U17640 ( .A1(n14404), .A2(n14180), .B1(n14179), .B2(n19412), .ZN(
        P3_U3285) );
  INV_X1 U17641 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n15182) );
  INV_X1 U17642 ( .A(n20757), .ZN(n14183) );
  NOR2_X1 U17643 ( .A1(n14509), .A2(n14181), .ZN(n14182) );
  AOI21_X1 U17644 ( .B1(DATAI_15_), .B2(n14509), .A(n14182), .ZN(n15183) );
  INV_X1 U17645 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n21615) );
  OAI222_X1 U17646 ( .A1(n14326), .A2(n15182), .B1(n14183), .B2(n15183), .C1(
        n14327), .C2(n21615), .ZN(P1_U2967) );
  AOI21_X1 U17647 ( .B1(n14185), .B2(n14118), .A(n14184), .ZN(n16528) );
  INV_X1 U17648 ( .A(n16528), .ZN(n15776) );
  INV_X1 U17649 ( .A(n14186), .ZN(n14187) );
  INV_X1 U17650 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19877) );
  OAI222_X1 U17651 ( .A1(n15776), .A2(n16096), .B1(n14187), .B2(n19821), .C1(
        n19877), .C2(n19832), .ZN(P2_U2906) );
  INV_X1 U17652 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14189) );
  XNOR2_X1 U17653 ( .A(n14188), .B(n14189), .ZN(n16913) );
  INV_X1 U17654 ( .A(n16913), .ZN(n14203) );
  INV_X1 U17655 ( .A(n18836), .ZN(n16999) );
  INV_X1 U17656 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14299) );
  NAND3_X1 U17657 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14300) );
  NOR2_X1 U17658 ( .A1(n14299), .A2(n14300), .ZN(n16944) );
  INV_X1 U17659 ( .A(n16941), .ZN(n14194) );
  AOI21_X1 U17660 ( .B1(n16943), .B2(n14190), .A(n18817), .ZN(n14191) );
  AOI21_X1 U17661 ( .B1(n14194), .B2(n19400), .A(n14191), .ZN(n18961) );
  OAI211_X1 U17662 ( .C1(n16999), .C2(n16944), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n18961), .ZN(n14263) );
  OAI22_X1 U17663 ( .A1(n14194), .A2(n18762), .B1(n14193), .B2(n14192), .ZN(
        n18940) );
  NAND2_X1 U17664 ( .A1(n16944), .A2(n18940), .ZN(n18806) );
  AOI21_X1 U17665 ( .B1(n14189), .B2(n18806), .A(n18888), .ZN(n14201) );
  OAI21_X1 U17666 ( .B1(n14197), .B2(n14196), .A(n14195), .ZN(n14198) );
  XOR2_X1 U17667 ( .A(n14198), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n16918) );
  INV_X1 U17668 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19490) );
  NOR2_X1 U17669 ( .A1(n18981), .A2(n19490), .ZN(n16914) );
  AOI21_X1 U17670 ( .B1(n18976), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16914), .ZN(n14199) );
  OAI21_X1 U17671 ( .B1(n18973), .B2(n16918), .A(n14199), .ZN(n14200) );
  AOI21_X1 U17672 ( .B1(n14263), .B2(n14201), .A(n14200), .ZN(n14202) );
  OAI21_X1 U17673 ( .B1(n14203), .B2(n18971), .A(n14202), .ZN(P3_U2855) );
  NAND3_X1 U17674 ( .A1(n18120), .A2(n14205), .A3(n14204), .ZN(n14206) );
  NAND2_X1 U17675 ( .A1(n18120), .A2(n14279), .ZN(n18300) );
  INV_X1 U17676 ( .A(n18300), .ZN(n14280) );
  INV_X1 U17677 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n18403) );
  INV_X1 U17678 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n18377) );
  NOR2_X1 U17679 ( .A1(n18403), .A2(n18377), .ZN(n18182) );
  INV_X1 U17680 ( .A(n18182), .ZN(n14278) );
  OAI211_X1 U17681 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n14280), .B(n14278), .ZN(n14212) );
  NAND2_X1 U17682 ( .A1(n14210), .A2(n14279), .ZN(n18321) );
  AOI22_X1 U17683 ( .A1(n18183), .A2(P3_EAX_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n18310), .ZN(n14211) );
  OAI211_X1 U17684 ( .C1(n14213), .C2(n18318), .A(n14212), .B(n14211), .ZN(
        P3_U2734) );
  AND2_X1 U17685 ( .A1(n19586), .A2(n14214), .ZN(n19588) );
  INV_X1 U17686 ( .A(n19588), .ZN(n17820) );
  INV_X1 U17687 ( .A(n14215), .ZN(n14216) );
  NAND2_X1 U17688 ( .A1(n14216), .A2(n14394), .ZN(n14359) );
  INV_X1 U17689 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17635) );
  NAND2_X1 U17690 ( .A1(n14217), .A2(n17784), .ZN(n17738) );
  OAI21_X1 U17691 ( .B1(n17635), .B2(n17738), .A(n17791), .ZN(n14219) );
  OAI21_X1 U17692 ( .B1(n17775), .B2(n17635), .A(n17784), .ZN(n17649) );
  INV_X1 U17693 ( .A(n17649), .ZN(n17740) );
  INV_X1 U17694 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n18173) );
  OAI22_X1 U17695 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17712), .B1(n17812), 
        .B2(n18173), .ZN(n14218) );
  AOI221_X1 U17696 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n14219), .C1(
        n16927), .C2(n17740), .A(n14218), .ZN(n14222) );
  INV_X1 U17697 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n18179) );
  NAND2_X1 U17698 ( .A1(n18179), .A2(n18173), .ZN(n17793) );
  OAI21_X1 U17699 ( .B1(n18173), .B2(n18179), .A(n17793), .ZN(n18175) );
  INV_X1 U17700 ( .A(n18175), .ZN(n14220) );
  AOI22_X1 U17701 ( .A1(n17786), .A2(n14220), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n17796), .ZN(n14221) );
  OAI211_X1 U17702 ( .C1(n17820), .C2(n14359), .A(n14222), .B(n14221), .ZN(
        P3_U2670) );
  OAI21_X1 U17703 ( .B1(n14184), .B2(n14224), .A(n14223), .ZN(n19680) );
  INV_X1 U17704 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U17705 ( .A1(n16713), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14225) );
  OAI21_X1 U17706 ( .B1(n16713), .B2(n14226), .A(n14225), .ZN(n19908) );
  AOI22_X1 U17707 ( .A1(n19824), .A2(n19908), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19813), .ZN(n14227) );
  OAI21_X1 U17708 ( .B1(n19680), .B2(n16096), .A(n14227), .ZN(P2_U2905) );
  XNOR2_X2 U17709 ( .A(n14228), .B(n14229), .ZN(n20590) );
  INV_X1 U17710 ( .A(n20590), .ZN(n16683) );
  MUX2_X1 U17711 ( .A(P2_EBX_REG_2__SCAN_IN), .B(n19945), .S(n16002), .Z(
        n14230) );
  AOI21_X1 U17712 ( .B1(n16683), .B2(n15992), .A(n14230), .ZN(n14231) );
  INV_X1 U17713 ( .A(n14231), .ZN(P2_U2885) );
  NOR2_X1 U17714 ( .A1(n14236), .A2(n9574), .ZN(n14237) );
  AOI21_X1 U17715 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n9574), .A(n14237), .ZN(
        n14238) );
  OAI21_X1 U17716 ( .B1(n20582), .B2(n15975), .A(n14238), .ZN(P2_U2884) );
  AOI22_X1 U17717 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n14239) );
  OAI21_X1 U17718 ( .B1(n15155), .B2(n14248), .A(n14239), .ZN(P1_U2915) );
  INV_X1 U17719 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15165) );
  AOI22_X1 U17720 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n14240) );
  OAI21_X1 U17721 ( .B1(n15165), .B2(n14248), .A(n14240), .ZN(P1_U2918) );
  INV_X1 U17722 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U17723 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n14241) );
  OAI21_X1 U17724 ( .B1(n14242), .B2(n14248), .A(n14241), .ZN(P1_U2917) );
  AOI22_X1 U17725 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14243) );
  OAI21_X1 U17726 ( .B1(n15150), .B2(n14248), .A(n14243), .ZN(P1_U2914) );
  AOI22_X1 U17727 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n14244) );
  OAI21_X1 U17728 ( .B1(n15169), .B2(n14248), .A(n14244), .ZN(P1_U2919) );
  AOI22_X1 U17729 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n14245) );
  OAI21_X1 U17730 ( .B1(n15175), .B2(n14248), .A(n14245), .ZN(P1_U2920) );
  INV_X1 U17731 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21555) );
  AOI22_X1 U17732 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14246) );
  OAI21_X1 U17733 ( .B1(n21555), .B2(n14248), .A(n14246), .ZN(P1_U2913) );
  INV_X1 U17734 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14249) );
  AOI22_X1 U17735 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n14247) );
  OAI21_X1 U17736 ( .B1(n14249), .B2(n14248), .A(n14247), .ZN(P1_U2916) );
  NAND2_X1 U17737 ( .A1(n14251), .A2(n14250), .ZN(n14252) );
  NAND2_X1 U17738 ( .A1(n14253), .A2(n14252), .ZN(n15013) );
  NOR2_X1 U17739 ( .A1(n14256), .A2(n14255), .ZN(n14257) );
  AOI22_X1 U17740 ( .A1(n15097), .A2(n10433), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15096), .ZN(n14258) );
  OAI21_X1 U17741 ( .B1(n15013), .B2(n15099), .A(n14258), .ZN(P1_U2870) );
  XNOR2_X1 U17742 ( .A(n16907), .B(n18565), .ZN(n16910) );
  AOI21_X1 U17743 ( .B1(n14260), .B2(n13334), .A(n14259), .ZN(n16906) );
  INV_X1 U17744 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n14261) );
  INV_X1 U17745 ( .A(n18976), .ZN(n18969) );
  OAI22_X1 U17746 ( .A1(n18981), .A2(n14261), .B1(n13334), .B2(n18969), .ZN(
        n14262) );
  AOI21_X1 U17747 ( .B1(n16906), .B2(n18870), .A(n14262), .ZN(n14269) );
  INV_X1 U17748 ( .A(n18878), .ZN(n18902) );
  INV_X1 U17749 ( .A(n16907), .ZN(n14266) );
  NAND4_X1 U17750 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16944), .A3(
        n13334), .A4(n18940), .ZN(n14265) );
  NAND3_X1 U17751 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18836), .A3(
        n14263), .ZN(n14264) );
  OAI211_X1 U17752 ( .C1(n18902), .C2(n14266), .A(n14265), .B(n14264), .ZN(
        n14267) );
  NAND2_X1 U17753 ( .A1(n14267), .A2(n18958), .ZN(n14268) );
  OAI211_X1 U17754 ( .C1(n16910), .C2(n18913), .A(n14269), .B(n14268), .ZN(
        P3_U2854) );
  NAND2_X1 U17755 ( .A1(n18309), .A2(n14270), .ZN(n14272) );
  AOI22_X1 U17756 ( .A1(n18183), .A2(P3_EAX_REG_0__SCAN_IN), .B1(n18310), .B2(
        BUF2_REG_0__SCAN_IN), .ZN(n14271) );
  OAI211_X1 U17757 ( .C1(n18300), .C2(P3_EAX_REG_0__SCAN_IN), .A(n14272), .B(
        n14271), .ZN(P3_U2735) );
  INV_X2 U17758 ( .A(n18647), .ZN(n18727) );
  AOI21_X1 U17759 ( .B1(n16923), .B2(n14277), .A(n14273), .ZN(n14276) );
  NAND3_X1 U17760 ( .A1(n19451), .A2(n18608), .A3(n18708), .ZN(n14274) );
  NAND2_X1 U17761 ( .A1(n14274), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14275) );
  OAI211_X1 U17762 ( .C1(n18727), .C2(n14277), .A(n14276), .B(n14275), .ZN(
        P3_U2830) );
  INV_X1 U17763 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n18372) );
  NAND2_X2 U17764 ( .A1(n19024), .A2(n14279), .ZN(n18316) );
  AOI22_X1 U17765 ( .A1(n14280), .A2(n18182), .B1(P3_EAX_REG_2__SCAN_IN), .B2(
        n18316), .ZN(n14284) );
  NAND2_X1 U17766 ( .A1(n18310), .A2(BUF2_REG_2__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U17767 ( .A1(n18309), .A2(n14281), .ZN(n14282) );
  OAI211_X1 U17768 ( .C1(n14287), .C2(n14284), .A(n14283), .B(n14282), .ZN(
        P3_U2733) );
  NAND2_X1 U17769 ( .A1(n14509), .A2(DATAI_2_), .ZN(n14286) );
  NAND2_X1 U17770 ( .A1(n15135), .A2(BUF1_REG_2__SCAN_IN), .ZN(n14285) );
  AND2_X1 U17771 ( .A1(n14286), .A2(n14285), .ZN(n20826) );
  OAI222_X1 U17772 ( .A1(n15013), .A2(n15195), .B1(n17225), .B2(n20826), .C1(
        n17230), .C2(n10972), .ZN(P1_U2902) );
  AOI21_X1 U17773 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n18316), .A(n14287), .ZN(
        n14291) );
  INV_X1 U17774 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n19009) );
  OAI22_X1 U17775 ( .A1(n18321), .A2(n19009), .B1(n18318), .B2(n14288), .ZN(
        n14289) );
  INV_X1 U17776 ( .A(n14289), .ZN(n14290) );
  OAI21_X1 U17777 ( .B1(n14291), .B2(n18315), .A(n14290), .ZN(P3_U2732) );
  AOI22_X1 U17778 ( .A1(n14294), .A2(n18694), .B1(n14293), .B2(n14292), .ZN(
        n14295) );
  XNOR2_X1 U17779 ( .A(n14296), .B(n14295), .ZN(n18693) );
  INV_X1 U17780 ( .A(n14300), .ZN(n14297) );
  OAI21_X1 U17781 ( .B1(n16999), .B2(n14297), .A(n18961), .ZN(n14298) );
  AOI21_X1 U17782 ( .B1(n14298), .B2(n18958), .A(n18976), .ZN(n18943) );
  OAI22_X1 U17783 ( .A1(n18693), .A2(n18973), .B1(n18943), .B2(n14299), .ZN(
        n14306) );
  NAND2_X1 U17784 ( .A1(n18958), .A2(n18940), .ZN(n18960) );
  NOR3_X1 U17785 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14300), .A3(
        n18960), .ZN(n14305) );
  XNOR2_X1 U17786 ( .A(n14302), .B(n14301), .ZN(n18688) );
  INV_X1 U17787 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n14303) );
  OAI22_X1 U17788 ( .A1(n18971), .A2(n18688), .B1(n18981), .B2(n14303), .ZN(
        n14304) );
  OR3_X1 U17789 ( .A1(n14306), .A2(n14305), .A3(n14304), .ZN(P3_U2856) );
  AOI22_X1 U17790 ( .A1(n20770), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20765), .ZN(n14310) );
  NAND2_X1 U17791 ( .A1(n14509), .A2(DATAI_4_), .ZN(n14308) );
  NAND2_X1 U17792 ( .A1(n15135), .A2(BUF1_REG_4__SCAN_IN), .ZN(n14307) );
  AND2_X1 U17793 ( .A1(n14308), .A2(n14307), .ZN(n20835) );
  INV_X1 U17794 ( .A(n20835), .ZN(n14309) );
  NAND2_X1 U17795 ( .A1(n20757), .A2(n14309), .ZN(n14336) );
  NAND2_X1 U17796 ( .A1(n14310), .A2(n14336), .ZN(P1_U2956) );
  AOI22_X1 U17797 ( .A1(n20770), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20765), .ZN(n14314) );
  NAND2_X1 U17798 ( .A1(n14509), .A2(DATAI_7_), .ZN(n14312) );
  NAND2_X1 U17799 ( .A1(n15135), .A2(BUF1_REG_7__SCAN_IN), .ZN(n14311) );
  INV_X1 U17800 ( .A(n20857), .ZN(n14313) );
  NAND2_X1 U17801 ( .A1(n20757), .A2(n14313), .ZN(n14344) );
  NAND2_X1 U17802 ( .A1(n14314), .A2(n14344), .ZN(P1_U2959) );
  AOI22_X1 U17803 ( .A1(n20770), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20765), .ZN(n14318) );
  NAND2_X1 U17804 ( .A1(n14509), .A2(DATAI_5_), .ZN(n14316) );
  NAND2_X1 U17805 ( .A1(n15135), .A2(BUF1_REG_5__SCAN_IN), .ZN(n14315) );
  AND2_X1 U17806 ( .A1(n14316), .A2(n14315), .ZN(n20840) );
  INV_X1 U17807 ( .A(n20840), .ZN(n14317) );
  NAND2_X1 U17808 ( .A1(n20757), .A2(n14317), .ZN(n14348) );
  NAND2_X1 U17809 ( .A1(n14318), .A2(n14348), .ZN(P1_U2957) );
  AOI22_X1 U17810 ( .A1(n20770), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20765), .ZN(n14322) );
  NAND2_X1 U17811 ( .A1(n14509), .A2(DATAI_6_), .ZN(n14320) );
  NAND2_X1 U17812 ( .A1(n15135), .A2(BUF1_REG_6__SCAN_IN), .ZN(n14319) );
  AND2_X1 U17813 ( .A1(n14320), .A2(n14319), .ZN(n20844) );
  INV_X1 U17814 ( .A(n20844), .ZN(n14321) );
  NAND2_X1 U17815 ( .A1(n20757), .A2(n14321), .ZN(n14350) );
  NAND2_X1 U17816 ( .A1(n14322), .A2(n14350), .ZN(P1_U2958) );
  INV_X1 U17817 ( .A(n14223), .ZN(n14324) );
  OAI21_X1 U17818 ( .B1(n14324), .B2(n10450), .A(n16496), .ZN(n19665) );
  INV_X1 U17819 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19873) );
  OAI222_X1 U17820 ( .A1(n19665), .A2(n16096), .B1(n19832), .B2(n19873), .C1(
        n14325), .C2(n19821), .ZN(P2_U2904) );
  AOI22_X1 U17821 ( .A1(n20770), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20765), .ZN(n14329) );
  INV_X1 U17822 ( .A(n20821), .ZN(n14328) );
  NAND2_X1 U17823 ( .A1(n20757), .A2(n14328), .ZN(n14346) );
  NAND2_X1 U17824 ( .A1(n14329), .A2(n14346), .ZN(P1_U2938) );
  AOI22_X1 U17825 ( .A1(n20770), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20765), .ZN(n14331) );
  INV_X1 U17826 ( .A(n15176), .ZN(n14330) );
  NAND2_X1 U17827 ( .A1(n20757), .A2(n14330), .ZN(n14334) );
  NAND2_X1 U17828 ( .A1(n14331), .A2(n14334), .ZN(P1_U2937) );
  AOI22_X1 U17829 ( .A1(n20770), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20765), .ZN(n14333) );
  INV_X1 U17830 ( .A(n20826), .ZN(n14332) );
  NAND2_X1 U17831 ( .A1(n20757), .A2(n14332), .ZN(n14342) );
  NAND2_X1 U17832 ( .A1(n14333), .A2(n14342), .ZN(P1_U2954) );
  AOI22_X1 U17833 ( .A1(n20770), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20765), .ZN(n14335) );
  NAND2_X1 U17834 ( .A1(n14335), .A2(n14334), .ZN(P1_U2952) );
  AOI22_X1 U17835 ( .A1(n20770), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20765), .ZN(n14337) );
  NAND2_X1 U17836 ( .A1(n14337), .A2(n14336), .ZN(P1_U2941) );
  AOI22_X1 U17837 ( .A1(n20770), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20765), .ZN(n14341) );
  NAND2_X1 U17838 ( .A1(n14509), .A2(DATAI_3_), .ZN(n14339) );
  NAND2_X1 U17839 ( .A1(n15135), .A2(BUF1_REG_3__SCAN_IN), .ZN(n14338) );
  AND2_X1 U17840 ( .A1(n14339), .A2(n14338), .ZN(n20830) );
  INV_X1 U17841 ( .A(n20830), .ZN(n14340) );
  NAND2_X1 U17842 ( .A1(n20757), .A2(n14340), .ZN(n14352) );
  NAND2_X1 U17843 ( .A1(n14341), .A2(n14352), .ZN(P1_U2955) );
  AOI22_X1 U17844 ( .A1(n20770), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20765), .ZN(n14343) );
  NAND2_X1 U17845 ( .A1(n14343), .A2(n14342), .ZN(P1_U2939) );
  AOI22_X1 U17846 ( .A1(n20770), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20765), .ZN(n14345) );
  NAND2_X1 U17847 ( .A1(n14345), .A2(n14344), .ZN(P1_U2944) );
  AOI22_X1 U17848 ( .A1(n20770), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20765), .ZN(n14347) );
  NAND2_X1 U17849 ( .A1(n14347), .A2(n14346), .ZN(P1_U2953) );
  AOI22_X1 U17850 ( .A1(n20770), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20765), .ZN(n14349) );
  NAND2_X1 U17851 ( .A1(n14349), .A2(n14348), .ZN(P1_U2942) );
  AOI22_X1 U17852 ( .A1(n20770), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20765), .ZN(n14351) );
  NAND2_X1 U17853 ( .A1(n14351), .A2(n14350), .ZN(P1_U2943) );
  AOI22_X1 U17854 ( .A1(n20770), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20765), .ZN(n14353) );
  NAND2_X1 U17855 ( .A1(n14353), .A2(n14352), .ZN(P1_U2940) );
  NOR2_X1 U17856 ( .A1(n14354), .A2(n18905), .ZN(n14363) );
  OAI22_X1 U17857 ( .A1(n14363), .A2(n14359), .B1(n14355), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19424) );
  INV_X1 U17858 ( .A(n19444), .ZN(n14384) );
  NOR2_X1 U17859 ( .A1(n19451), .A2(n14356), .ZN(n14387) );
  INV_X1 U17860 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U17861 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n9830), .B2(n16873), .ZN(
        n14386) );
  INV_X1 U17862 ( .A(n14386), .ZN(n14357) );
  NAND2_X1 U17863 ( .A1(n14387), .A2(n14357), .ZN(n14358) );
  OAI211_X1 U17864 ( .C1(n14384), .C2(n14359), .A(n17129), .B(n14358), .ZN(
        n14360) );
  AOI21_X1 U17865 ( .B1(n19424), .B2(n19584), .A(n14360), .ZN(n14361) );
  AOI21_X1 U17866 ( .B1(n14404), .B2(n14393), .A(n14361), .ZN(P3_U3289) );
  NAND2_X1 U17867 ( .A1(n19444), .A2(n14362), .ZN(n14367) );
  MUX2_X1 U17868 ( .A(n14363), .B(n18927), .S(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n19421) );
  NOR2_X1 U17869 ( .A1(n19421), .A2(n17817), .ZN(n14365) );
  OAI21_X1 U17870 ( .B1(n19451), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17129), .ZN(n14364) );
  OAI22_X1 U17871 ( .A1(n17129), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n14365), .B2(n14364), .ZN(n14366) );
  OAI21_X1 U17872 ( .B1(n14404), .B2(n14367), .A(n14366), .ZN(P3_U3290) );
  AND2_X1 U17873 ( .A1(n14368), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14371) );
  INV_X1 U17874 ( .A(n14370), .ZN(n14372) );
  OR3_X1 U17875 ( .A1(n14373), .A2(n14372), .A3(n14371), .ZN(n14374) );
  NAND2_X1 U17876 ( .A1(n15990), .A2(n14374), .ZN(n19808) );
  INV_X1 U17877 ( .A(n14452), .ZN(n14443) );
  NAND2_X1 U17878 ( .A1(n14375), .A2(n14376), .ZN(n14377) );
  NAND2_X1 U17879 ( .A1(n14443), .A2(n14377), .ZN(n19951) );
  NOR2_X1 U17880 ( .A1(n19951), .A2(n9574), .ZN(n14378) );
  AOI21_X1 U17881 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n9574), .A(n14378), .ZN(
        n14379) );
  OAI21_X1 U17882 ( .B1(n19808), .B2(n15975), .A(n14379), .ZN(P2_U2883) );
  INV_X1 U17883 ( .A(n14380), .ZN(n14381) );
  AND2_X1 U17884 ( .A1(n14382), .A2(n14381), .ZN(n17795) );
  INV_X1 U17885 ( .A(n17795), .ZN(n14383) );
  NOR2_X1 U17886 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  AOI211_X1 U17887 ( .C1(n14387), .C2(n14386), .A(n14404), .B(n14385), .ZN(
        n14403) );
  OR2_X1 U17888 ( .A1(n14388), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14390) );
  AOI21_X1 U17889 ( .B1(n14391), .B2(n14390), .A(n14389), .ZN(n14396) );
  OAI22_X1 U17890 ( .A1(n18926), .A2(n14394), .B1(n14393), .B2(n14388), .ZN(
        n14395) );
  MUX2_X1 U17891 ( .A(n14396), .B(n14395), .S(n14167), .Z(n14401) );
  OAI211_X1 U17892 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n14398), .B(n14397), .ZN(
        n14399) );
  OAI21_X1 U17893 ( .B1(n18762), .B2(n17795), .A(n14399), .ZN(n14400) );
  NOR2_X1 U17894 ( .A1(n14401), .A2(n14400), .ZN(n19417) );
  OR2_X1 U17895 ( .A1(n19417), .A2(n17817), .ZN(n14402) );
  AOI22_X1 U17896 ( .A1(n14404), .A2(n14167), .B1(n14403), .B2(n14402), .ZN(
        P3_U3288) );
  MUX2_X1 U17897 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14405), .S(
        n17143), .Z(n17149) );
  NOR2_X1 U17898 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21403), .ZN(n14413) );
  AOI22_X1 U17899 ( .A1(n17149), .A2(n21403), .B1(n14413), .B2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14408) );
  MUX2_X1 U17900 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14406), .S(
        n17143), .Z(n17154) );
  AOI22_X1 U17901 ( .A1(n14413), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21403), .B2(n17154), .ZN(n14407) );
  NOR2_X1 U17902 ( .A1(n14408), .A2(n14407), .ZN(n17161) );
  INV_X1 U17903 ( .A(n14409), .ZN(n14410) );
  NAND2_X1 U17904 ( .A1(n17161), .A2(n14410), .ZN(n14424) );
  NOR2_X1 U17905 ( .A1(n9642), .A2(n9872), .ZN(n14411) );
  XNOR2_X1 U17906 ( .A(n14411), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20690) );
  OAI21_X1 U17907 ( .B1(n20690), .B2(n17271), .A(n17143), .ZN(n14415) );
  INV_X1 U17908 ( .A(n17143), .ZN(n14412) );
  AOI21_X1 U17909 ( .B1(n14412), .B2(n17275), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n14414) );
  AOI22_X1 U17910 ( .A1(n14415), .A2(n14414), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n14413), .ZN(n17163) );
  AND3_X1 U17911 ( .A1(n14424), .A2(n21646), .A3(n17163), .ZN(n14416) );
  AND2_X1 U17912 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21222), .ZN(n15589) );
  NOR2_X1 U17913 ( .A1(n13984), .A2(n15589), .ZN(n14422) );
  INV_X1 U17914 ( .A(n14417), .ZN(n14418) );
  NOR2_X1 U17915 ( .A1(n14418), .A2(n21497), .ZN(n14419) );
  INV_X1 U17916 ( .A(n14419), .ZN(n21346) );
  NOR2_X1 U17917 ( .A1(n21346), .A2(n21341), .ZN(n14420) );
  NOR2_X1 U17918 ( .A1(n14419), .A2(n21341), .ZN(n20929) );
  INV_X1 U17919 ( .A(n10975), .ZN(n14500) );
  MUX2_X1 U17920 ( .A(n14420), .B(n20929), .S(n14500), .Z(n14421) );
  OAI21_X1 U17921 ( .B1(n14422), .B2(n14421), .A(n20817), .ZN(n14423) );
  OAI21_X1 U17922 ( .B1(n20817), .B2(n21143), .A(n14423), .ZN(P1_U3476) );
  AND3_X1 U17923 ( .A1(n14424), .A2(n17163), .A3(n17280), .ZN(n17168) );
  INV_X1 U17924 ( .A(n10986), .ZN(n15024) );
  OAI22_X1 U17925 ( .A1(n20889), .A2(n21341), .B1(n15024), .B2(n15589), .ZN(
        n14425) );
  OAI21_X1 U17926 ( .B1(n17168), .B2(n14425), .A(n20817), .ZN(n14426) );
  OAI21_X1 U17927 ( .B1(n20817), .B2(n21264), .A(n14426), .ZN(P1_U3478) );
  INV_X1 U17928 ( .A(n14428), .ZN(n14427) );
  MUX2_X1 U17929 ( .A(n21345), .B(n21064), .S(n14417), .Z(n14430) );
  AOI211_X1 U17930 ( .C1(n14430), .C2(n21193), .A(P1_STATE2_REG_3__SCAN_IN), 
        .B(n14429), .ZN(n14433) );
  INV_X1 U17931 ( .A(n14501), .ZN(n14431) );
  NAND2_X1 U17932 ( .A1(n21349), .A2(n21497), .ZN(n21219) );
  INV_X1 U17933 ( .A(n21088), .ZN(n20702) );
  OAI22_X1 U17934 ( .A1(n14431), .A2(n21219), .B1(n20702), .B2(n15589), .ZN(
        n14432) );
  OAI21_X1 U17935 ( .B1(n14433), .B2(n14432), .A(n20817), .ZN(n14434) );
  OAI21_X1 U17936 ( .B1(n20817), .B2(n21184), .A(n14434), .ZN(P1_U3475) );
  NAND2_X1 U17937 ( .A1(n20786), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15586) );
  OAI21_X1 U17938 ( .B1(n15271), .B2(n15020), .A(n15586), .ZN(n14435) );
  AOI21_X1 U17939 ( .B1(n15274), .B2(n15020), .A(n14435), .ZN(n14441) );
  XNOR2_X1 U17940 ( .A(n14437), .B(n14436), .ZN(n14438) );
  NAND2_X1 U17941 ( .A1(n14438), .A2(n14473), .ZN(n15579) );
  INV_X1 U17942 ( .A(n14438), .ZN(n14439) );
  NAND2_X1 U17943 ( .A1(n14439), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15578) );
  NAND3_X1 U17944 ( .A1(n15579), .A2(n15578), .A3(n20780), .ZN(n14440) );
  OAI211_X1 U17945 ( .C1(n15022), .C2(n17244), .A(n14441), .B(n14440), .ZN(
        P1_U2998) );
  XOR2_X1 U17946 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n15990), .Z(n14447)
         );
  OR2_X1 U17947 ( .A1(n14443), .A2(n14442), .ZN(n15996) );
  NAND2_X1 U17948 ( .A1(n14443), .A2(n14442), .ZN(n14444) );
  NAND2_X1 U17949 ( .A1(n15996), .A2(n14444), .ZN(n19769) );
  MUX2_X1 U17950 ( .A(n19769), .B(n14445), .S(n9574), .Z(n14446) );
  OAI21_X1 U17951 ( .B1(n14447), .B2(n15975), .A(n14446), .ZN(P2_U2882) );
  OAI21_X1 U17952 ( .B1(n14450), .B2(n14449), .A(n14448), .ZN(n20706) );
  OAI222_X1 U17953 ( .A1(n20706), .A2(n15195), .B1(n17225), .B2(n20830), .C1(
        n17230), .C2(n11000), .ZN(P1_U2901) );
  XNOR2_X1 U17954 ( .A(n15991), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14458) );
  AND2_X1 U17955 ( .A1(n14452), .A2(n14453), .ZN(n15998) );
  NAND2_X1 U17956 ( .A1(n14452), .A2(n14454), .ZN(n15983) );
  OAI21_X1 U17957 ( .B1(n15998), .B2(n14455), .A(n15983), .ZN(n19740) );
  MUX2_X1 U17958 ( .A(n14456), .B(n19740), .S(n16002), .Z(n14457) );
  OAI21_X1 U17959 ( .B1(n14458), .B2(n15975), .A(n14457), .ZN(P2_U2880) );
  XNOR2_X1 U17960 ( .A(n14448), .B(n14459), .ZN(n20778) );
  INV_X1 U17961 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U17962 ( .A1(n15195), .A2(n20778), .B1(n17230), .B2(n20733), .C1(
        n17225), .C2(n20835), .ZN(P1_U2900) );
  INV_X1 U17963 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14460) );
  INV_X1 U17964 ( .A(n14254), .ZN(n14463) );
  XNOR2_X1 U17965 ( .A(n14463), .B(n14462), .ZN(n20704) );
  OAI222_X1 U17966 ( .A1(n15079), .A2(n20706), .B1(n14460), .B2(n15104), .C1(
        n15105), .C2(n20704), .ZN(P1_U2869) );
  OAI21_X1 U17967 ( .B1(n14463), .B2(n14462), .A(n14461), .ZN(n14465) );
  NAND2_X1 U17968 ( .A1(n14465), .A2(n14464), .ZN(n20684) );
  INV_X1 U17969 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14466) );
  OAI222_X1 U17970 ( .A1(n20684), .A2(n15105), .B1(n14466), .B2(n15104), .C1(
        n15079), .C2(n20778), .ZN(P1_U2868) );
  OAI21_X1 U17971 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n17246) );
  NOR2_X1 U17972 ( .A1(n20812), .A2(n14473), .ZN(n14471) );
  INV_X1 U17973 ( .A(n14472), .ZN(n14470) );
  NOR2_X1 U17974 ( .A1(n20799), .A2(n20785), .ZN(n14475) );
  NAND2_X1 U17975 ( .A1(n20805), .A2(n14472), .ZN(n20814) );
  AOI21_X1 U17976 ( .B1(n14473), .B2(n20811), .A(n15533), .ZN(n20802) );
  OAI211_X1 U17977 ( .C1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n15555), .A(
        n20814), .B(n20802), .ZN(n20794) );
  AOI21_X1 U17978 ( .B1(n15580), .B2(n15529), .A(n20794), .ZN(n17270) );
  INV_X1 U17979 ( .A(n17270), .ZN(n14474) );
  MUX2_X1 U17980 ( .A(n14475), .B(n14474), .S(
        P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n14476) );
  INV_X1 U17981 ( .A(n14476), .ZN(n14481) );
  INV_X1 U17982 ( .A(n14477), .ZN(n14478) );
  AOI21_X1 U17983 ( .B1(n14479), .B2(n14464), .A(n14478), .ZN(n14998) );
  AOI22_X1 U17984 ( .A1(n20801), .A2(n14998), .B1(n20786), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n14480) );
  OAI211_X1 U17985 ( .C1(n17246), .C2(n20807), .A(n14481), .B(n14480), .ZN(
        P1_U3026) );
  OAI21_X1 U17986 ( .B1(n14484), .B2(n14483), .A(n14482), .ZN(n20808) );
  INV_X1 U17987 ( .A(n20808), .ZN(n14488) );
  INV_X1 U17988 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n14485) );
  NOR2_X1 U17989 ( .A1(n15360), .A2(n14485), .ZN(n20800) );
  AOI21_X1 U17990 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20800), .ZN(n14486) );
  OAI21_X1 U17991 ( .B1(n20784), .B2(n15009), .A(n14486), .ZN(n14487) );
  AOI21_X1 U17992 ( .B1(n14488), .B2(n20780), .A(n14487), .ZN(n14489) );
  OAI21_X1 U17993 ( .B1(n17244), .B2(n15013), .A(n14489), .ZN(P1_U2997) );
  XNOR2_X1 U17994 ( .A(n20775), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14492) );
  INV_X1 U17995 ( .A(n14490), .ZN(n14491) );
  NOR2_X1 U17996 ( .A1(n14492), .A2(n14491), .ZN(n20774) );
  AOI21_X1 U17997 ( .B1(n14492), .B2(n14491), .A(n20774), .ZN(n20796) );
  NAND2_X1 U17998 ( .A1(n20796), .A2(n20780), .ZN(n14496) );
  INV_X1 U17999 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14493) );
  NOR2_X1 U18000 ( .A1(n15360), .A2(n14493), .ZN(n20792) );
  NOR2_X1 U18001 ( .A1(n20784), .A2(n20707), .ZN(n14494) );
  AOI211_X1 U18002 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20792), .B(n14494), .ZN(n14495) );
  OAI211_X1 U18003 ( .C1(n17244), .C2(n20706), .A(n14496), .B(n14495), .ZN(
        P1_U2996) );
  OAI222_X1 U18004 ( .A1(n17245), .A2(n15195), .B1(n20840), .B2(n17225), .C1(
        n17230), .C2(n11024), .ZN(P1_U2899) );
  INV_X1 U18005 ( .A(n14998), .ZN(n14499) );
  INV_X1 U18006 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n14995) );
  OAI222_X1 U18007 ( .A1(n14499), .A2(n15105), .B1(n14995), .B2(n15104), .C1(
        n17245), .C2(n15079), .ZN(P1_U2867) );
  INV_X1 U18008 ( .A(n21401), .ZN(n21388) );
  OAI21_X1 U18009 ( .B1(n20876), .B2(n21388), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14503) );
  NAND2_X1 U18010 ( .A1(n14503), .A2(n21349), .ZN(n14516) );
  INV_X1 U18011 ( .A(n14516), .ZN(n14508) );
  OR2_X1 U18012 ( .A1(n21088), .A2(n15005), .ZN(n20933) );
  NAND2_X1 U18013 ( .A1(n14514), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21293) );
  INV_X1 U18014 ( .A(n21293), .ZN(n14505) );
  INV_X1 U18015 ( .A(n21149), .ZN(n20894) );
  NAND2_X1 U18016 ( .A1(n21089), .A2(n21148), .ZN(n20970) );
  INV_X1 U18017 ( .A(n20970), .ZN(n14506) );
  NAND3_X1 U18018 ( .A1(n21184), .A2(n21143), .A3(n21216), .ZN(n20864) );
  NOR2_X1 U18019 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20864), .ZN(
        n14512) );
  OAI22_X1 U18020 ( .A1(n14506), .A2(n11005), .B1(n14512), .B2(n21222), .ZN(
        n14507) );
  INV_X1 U18021 ( .A(n21354), .ZN(n21303) );
  AOI22_X1 U18022 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20852), .B1(DATAI_24_), 
        .B2(n20853), .ZN(n21306) );
  NAND2_X1 U18023 ( .A1(n20854), .A2(n14511), .ZN(n21217) );
  INV_X1 U18024 ( .A(n14512), .ZN(n20855) );
  OAI22_X1 U18025 ( .A1(n21401), .A2(n21306), .B1(n21217), .B2(n20855), .ZN(
        n14513) );
  AOI21_X1 U18026 ( .B1(n20876), .B2(n21303), .A(n14513), .ZN(n14518) );
  NOR2_X1 U18027 ( .A1(n14514), .A2(n11005), .ZN(n20974) );
  INV_X1 U18028 ( .A(n20974), .ZN(n21154) );
  NOR2_X2 U18029 ( .A1(n20973), .A2(n15176), .ZN(n21342) );
  NAND2_X1 U18030 ( .A1(n20858), .A2(n21342), .ZN(n14517) );
  OAI211_X1 U18031 ( .C1(n20851), .C2(n14519), .A(n14518), .B(n14517), .ZN(
        P1_U3033) );
  NAND2_X1 U18032 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14520) );
  OAI211_X1 U18033 ( .C1(n14522), .C2(n20784), .A(n14521), .B(n14520), .ZN(
        n14523) );
  AOI21_X1 U18034 ( .B1(n15032), .B2(n20779), .A(n14523), .ZN(n14524) );
  OAI21_X1 U18035 ( .B1(n14525), .B2(n20631), .A(n14524), .ZN(P1_U2969) );
  OAI21_X1 U18036 ( .B1(n14528), .B2(n14527), .A(n14526), .ZN(n14543) );
  AOI21_X1 U18037 ( .B1(n14532), .B2(n15659), .A(n14531), .ZN(n16389) );
  INV_X1 U18038 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U18039 ( .A1(n19798), .A2(n14533), .B1(n19813), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n14535) );
  NAND2_X1 U18040 ( .A1(n19800), .A2(BUF1_REG_27__SCAN_IN), .ZN(n14534) );
  OAI211_X1 U18041 ( .C1(n16077), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        n14537) );
  AOI21_X1 U18042 ( .B1(n16389), .B2(n19823), .A(n14537), .ZN(n14538) );
  OAI21_X1 U18043 ( .B1(n14543), .B2(n16062), .A(n14538), .ZN(P2_U2892) );
  NOR2_X1 U18044 ( .A1(n16392), .A2(n9574), .ZN(n14541) );
  AOI21_X1 U18045 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n9574), .A(n14541), .ZN(
        n14542) );
  OAI21_X1 U18046 ( .B1(n14543), .B2(n15975), .A(n14542), .ZN(P2_U2860) );
  AOI211_X1 U18047 ( .C1(n16745), .C2(n15851), .A(n16062), .B(n16087), .ZN(
        n14544) );
  AOI21_X1 U18048 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19813), .A(n14544), .ZN(
        n14546) );
  NAND2_X1 U18049 ( .A1(n19824), .A2(n19797), .ZN(n14545) );
  OAI211_X1 U18050 ( .C1(n15851), .C2(n16081), .A(n14546), .B(n14545), .ZN(
        P2_U2919) );
  OR2_X1 U18051 ( .A1(n16543), .A2(n14553), .ZN(n16485) );
  AOI22_X1 U18052 ( .A1(n16206), .A2(n16603), .B1(n14548), .B2(n16512), .ZN(
        n14575) );
  NOR2_X1 U18053 ( .A1(n16603), .A2(n14549), .ZN(n14550) );
  NAND2_X1 U18054 ( .A1(n16576), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16562) );
  NAND2_X1 U18055 ( .A1(n16576), .A2(n14559), .ZN(n14551) );
  AOI21_X1 U18056 ( .B1(n14553), .B2(n16480), .A(n16545), .ZN(n16509) );
  NAND2_X1 U18057 ( .A1(n13143), .A2(n14555), .ZN(n14556) );
  AND2_X1 U18058 ( .A1(n16509), .A2(n14556), .ZN(n14557) );
  NAND2_X1 U18059 ( .A1(n14558), .A2(n14557), .ZN(n16495) );
  NOR2_X1 U18060 ( .A1(n14559), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14560) );
  OAI21_X1 U18061 ( .B1(n16495), .B2(n14560), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14574) );
  XNOR2_X1 U18062 ( .A(n14562), .B(n14561), .ZN(n16213) );
  INV_X1 U18063 ( .A(n14564), .ZN(n14565) );
  OAI21_X1 U18064 ( .B1(n14563), .B2(n14566), .A(n14565), .ZN(n16082) );
  NOR2_X1 U18065 ( .A1(n16082), .A2(n19959), .ZN(n14572) );
  NOR2_X1 U18066 ( .A1(n14568), .A2(n14569), .ZN(n14570) );
  OR2_X1 U18067 ( .A1(n14567), .A2(n14570), .ZN(n15923) );
  NAND2_X1 U18068 ( .A1(n16341), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n16216) );
  OAI21_X1 U18069 ( .B1(n15923), .B2(n16639), .A(n16216), .ZN(n14571) );
  AOI211_X1 U18070 ( .C1(n16213), .C2(n19962), .A(n14572), .B(n14571), .ZN(
        n14573) );
  OAI211_X1 U18071 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n14575), .A(
        n14574), .B(n14573), .ZN(P2_U3029) );
  INV_X1 U18072 ( .A(n17276), .ZN(n14582) );
  AOI21_X1 U18073 ( .B1(n17140), .B2(n20624), .A(n14582), .ZN(n14584) );
  NOR2_X1 U18074 ( .A1(n14576), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14577) );
  AOI21_X1 U18075 ( .B1(n10986), .B2(n15591), .A(n14577), .ZN(n17142) );
  INV_X1 U18076 ( .A(n17142), .ZN(n14580) );
  OAI22_X1 U18077 ( .A1(n14578), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21403), .ZN(n14579) );
  AOI21_X1 U18078 ( .B1(n20624), .B2(n14580), .A(n14579), .ZN(n14581) );
  OAI22_X1 U18079 ( .A1(n14584), .A2(n14583), .B1(n14582), .B2(n14581), .ZN(
        P1_U3474) );
  AOI22_X1 U18080 ( .A1(n11970), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11784), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14589) );
  AOI22_X1 U18081 ( .A1(n14592), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14588) );
  NAND3_X1 U18082 ( .A1(n14589), .A2(n14588), .A3(n14587), .ZN(n14605) );
  AOI22_X1 U18083 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14591) );
  AOI22_X1 U18084 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14590) );
  NAND2_X1 U18085 ( .A1(n14591), .A2(n14590), .ZN(n14604) );
  AOI22_X1 U18086 ( .A1(n9584), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14592), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14596) );
  AOI22_X1 U18087 ( .A1(n9579), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14593), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14594) );
  NAND3_X1 U18088 ( .A1(n14596), .A2(n14595), .A3(n14594), .ZN(n14603) );
  AOI22_X1 U18089 ( .A1(n14598), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14597), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14601) );
  AOI22_X1 U18090 ( .A1(n16692), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14599), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14600) );
  NAND2_X1 U18091 ( .A1(n14601), .A2(n14600), .ZN(n14602) );
  OAI22_X1 U18092 ( .A1(n14605), .A2(n14604), .B1(n14603), .B2(n14602), .ZN(
        n14606) );
  INV_X1 U18093 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14609) );
  AOI22_X1 U18094 ( .A1(n19798), .A2(n19908), .B1(n19813), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14608) );
  NAND2_X1 U18095 ( .A1(n19800), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14607) );
  OAI211_X1 U18096 ( .C1(n16077), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        n14610) );
  AOI21_X1 U18097 ( .B1(n14619), .B2(n19823), .A(n14610), .ZN(n14611) );
  OAI21_X1 U18098 ( .B1(n14614), .B2(n16062), .A(n14611), .ZN(P2_U2889) );
  OAI21_X1 U18099 ( .B1(n14614), .B2(n15975), .A(n14613), .ZN(P2_U2857) );
  NAND2_X1 U18100 ( .A1(n20480), .A2(n19970), .ZN(n14682) );
  NOR2_X1 U18101 ( .A1(n14621), .A2(n14682), .ZN(n14615) );
  NOR2_X1 U18102 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n14616), .ZN(n16829) );
  AND2_X1 U18103 ( .A1(n14617), .A2(n16829), .ZN(n14618) );
  NAND2_X1 U18104 ( .A1(n14619), .A2(n19785), .ZN(n14694) );
  NAND2_X1 U18105 ( .A1(n14682), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14620) );
  NOR2_X1 U18106 ( .A1(n14621), .A2(n14620), .ZN(n14622) );
  INV_X2 U18107 ( .A(n14700), .ZN(n19790) );
  NAND2_X1 U18108 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n14624), .ZN(
        n14651) );
  OAI21_X1 U18109 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14624), .A(
        n14651), .ZN(n19647) );
  INV_X1 U18110 ( .A(n19647), .ZN(n14649) );
  OAI21_X1 U18111 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14643), .A(
        n14646), .ZN(n16242) );
  INV_X1 U18112 ( .A(n16242), .ZN(n19686) );
  OAI21_X1 U18113 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n14625), .A(
        n14644), .ZN(n19690) );
  INV_X1 U18114 ( .A(n19690), .ZN(n14642) );
  INV_X1 U18115 ( .A(n14625), .ZN(n14626) );
  OAI21_X1 U18116 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n14627), .A(
        n14626), .ZN(n19715) );
  NAND2_X1 U18117 ( .A1(n16296), .A2(n14640), .ZN(n14630) );
  AND2_X1 U18118 ( .A1(n14630), .A2(n14629), .ZN(n16298) );
  AOI21_X1 U18119 ( .B1(n14638), .B2(n19721), .A(n14641), .ZN(n19719) );
  AOI21_X1 U18120 ( .B1(n19748), .B2(n14636), .A(n14639), .ZN(n19747) );
  AOI21_X1 U18121 ( .B1(n19934), .B2(n14634), .A(n14637), .ZN(n19916) );
  AOI21_X1 U18122 ( .B1(n19949), .B2(n15842), .A(n14635), .ZN(n19938) );
  INV_X1 U18123 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14631) );
  MUX2_X1 U18124 ( .A(n14632), .B(n14631), .S(n9587), .Z(n15853) );
  MUX2_X1 U18125 ( .A(n14633), .B(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .S(n16837), .Z(n15838) );
  NAND2_X1 U18126 ( .A1(n15853), .A2(n15838), .ZN(n15837) );
  OAI21_X1 U18127 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n14635), .A(
        n14634), .ZN(n16354) );
  NAND2_X1 U18128 ( .A1(n15813), .A2(n16354), .ZN(n19789) );
  OAI21_X1 U18129 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n14637), .A(
        n14636), .ZN(n19766) );
  NAND2_X1 U18130 ( .A1(n19763), .A2(n19766), .ZN(n19745) );
  NOR2_X1 U18131 ( .A1(n19747), .A2(n19745), .ZN(n19731) );
  OAI21_X1 U18132 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n14639), .A(
        n14638), .ZN(n19733) );
  NAND2_X1 U18133 ( .A1(n19731), .A2(n19733), .ZN(n19717) );
  OAI21_X1 U18134 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n14641), .A(
        n14640), .ZN(n16307) );
  NAND2_X1 U18135 ( .A1(n15795), .A2(n16307), .ZN(n15783) );
  NAND2_X1 U18136 ( .A1(n19715), .A2(n19712), .ZN(n19687) );
  AOI21_X1 U18137 ( .B1(n16257), .B2(n14644), .A(n14643), .ZN(n16255) );
  INV_X1 U18138 ( .A(n16255), .ZN(n14645) );
  NAND2_X1 U18139 ( .A1(n15768), .A2(n14645), .ZN(n19672) );
  NOR2_X1 U18140 ( .A1(n19686), .A2(n19672), .ZN(n19661) );
  INV_X1 U18141 ( .A(n14646), .ZN(n14648) );
  INV_X1 U18142 ( .A(n14624), .ZN(n14647) );
  OAI21_X1 U18143 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n14648), .A(
        n14647), .ZN(n19663) );
  NAND2_X1 U18144 ( .A1(n19661), .A2(n19663), .ZN(n19645) );
  INV_X1 U18145 ( .A(n14651), .ZN(n14650) );
  NAND2_X1 U18146 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n14650), .ZN(
        n14655) );
  INV_X1 U18147 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14652) );
  NAND2_X1 U18148 ( .A1(n14652), .A2(n14651), .ZN(n14653) );
  NAND2_X1 U18149 ( .A1(n14655), .A2(n14653), .ZN(n16217) );
  NAND2_X1 U18150 ( .A1(n15755), .A2(n16217), .ZN(n19638) );
  INV_X1 U18151 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14654) );
  NAND2_X1 U18152 ( .A1(n14655), .A2(n14654), .ZN(n14656) );
  NAND2_X1 U18153 ( .A1(n9691), .A2(n14656), .ZN(n19641) );
  INV_X1 U18154 ( .A(n19641), .ZN(n14657) );
  NOR2_X1 U18155 ( .A1(n19638), .A2(n14657), .ZN(n19622) );
  NAND2_X1 U18156 ( .A1(n19622), .A2(n19625), .ZN(n14658) );
  OAI21_X1 U18157 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14660), .A(
        n14659), .ZN(n16199) );
  INV_X1 U18158 ( .A(n15733), .ZN(n14661) );
  NAND2_X1 U18159 ( .A1(n14662), .A2(n19790), .ZN(n15718) );
  OAI21_X1 U18160 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n14663), .A(
        n14664), .ZN(n16182) );
  NAND2_X1 U18161 ( .A1(n15718), .A2(n16182), .ZN(n15701) );
  AOI21_X1 U18162 ( .B1(n16169), .B2(n14664), .A(n14667), .ZN(n16172) );
  OAI21_X1 U18163 ( .B1(n15701), .B2(n16172), .A(n19790), .ZN(n15686) );
  INV_X1 U18164 ( .A(n14665), .ZN(n14666) );
  OAI21_X1 U18165 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n14667), .A(
        n14666), .ZN(n16165) );
  NAND2_X1 U18166 ( .A1(n15686), .A2(n16165), .ZN(n15667) );
  NOR2_X1 U18167 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n14665), .ZN(
        n14668) );
  NOR2_X1 U18168 ( .A1(n14669), .A2(n14668), .ZN(n16154) );
  OAI21_X1 U18169 ( .B1(n15667), .B2(n16154), .A(n19790), .ZN(n15651) );
  OAI21_X1 U18170 ( .B1(n14669), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14670), .ZN(n16144) );
  AND2_X1 U18171 ( .A1(n14670), .A2(n15643), .ZN(n14671) );
  NOR2_X1 U18172 ( .A1(n14670), .A2(n15643), .ZN(n14673) );
  OR2_X1 U18173 ( .A1(n14671), .A2(n14673), .ZN(n16133) );
  NAND2_X1 U18174 ( .A1(n15638), .A2(n16133), .ZN(n14672) );
  NAND2_X1 U18175 ( .A1(n14672), .A2(n19790), .ZN(n15626) );
  NOR2_X1 U18176 ( .A1(n14673), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14674) );
  OR2_X1 U18177 ( .A1(n14675), .A2(n14674), .ZN(n16120) );
  NAND2_X1 U18178 ( .A1(n15626), .A2(n16120), .ZN(n15617) );
  NOR2_X1 U18179 ( .A1(n14675), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14676) );
  OR2_X1 U18180 ( .A1(n14677), .A2(n14676), .ZN(n16104) );
  INV_X1 U18181 ( .A(n16104), .ZN(n15622) );
  XNOR2_X1 U18182 ( .A(n14702), .B(n14701), .ZN(n14690) );
  NAND2_X1 U18183 ( .A1(n20392), .A2(n16837), .ZN(n14678) );
  NAND3_X1 U18184 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .A3(n14680), .ZN(n16839) );
  NAND2_X1 U18185 ( .A1(n19701), .A2(n16839), .ZN(n14681) );
  INV_X1 U18186 ( .A(n19778), .ZN(n19613) );
  INV_X1 U18187 ( .A(n16829), .ZN(n14697) );
  NAND2_X1 U18188 ( .A1(n13850), .A2(n14697), .ZN(n14686) );
  INV_X1 U18189 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n14683) );
  NAND3_X1 U18190 ( .A1(n14684), .A2(n14683), .A3(n14682), .ZN(n14685) );
  INV_X2 U18191 ( .A(n19651), .ZN(n19784) );
  AOI22_X1 U18192 ( .A1(n19613), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_30__SCAN_IN), .ZN(n14687) );
  INV_X1 U18193 ( .A(n14687), .ZN(n14688) );
  OAI21_X1 U18194 ( .B1(n14690), .B2(n20488), .A(n14689), .ZN(n14691) );
  AOI21_X1 U18195 ( .B1(n14692), .B2(n19736), .A(n14691), .ZN(n14693) );
  OAI211_X1 U18196 ( .C1(n13111), .C2(n19786), .A(n14694), .B(n14693), .ZN(
        P2_U2825) );
  INV_X1 U18197 ( .A(n14696), .ZN(n15862) );
  NAND3_X1 U18198 ( .A1(n13850), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n14697), 
        .ZN(n14698) );
  OAI21_X1 U18199 ( .B1(n19778), .B2(n20561), .A(n14698), .ZN(n14699) );
  AOI21_X1 U18200 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19777), .A(
        n14699), .ZN(n14704) );
  NAND3_X1 U18201 ( .A1(n14702), .A2(n15855), .A3(n14701), .ZN(n14703) );
  OAI211_X1 U18202 ( .C1(n14705), .C2(n19782), .A(n14704), .B(n14703), .ZN(
        n14706) );
  AOI21_X1 U18203 ( .B1(n15862), .B2(n19754), .A(n14706), .ZN(n14707) );
  OAI21_X1 U18204 ( .B1(n14695), .B2(n19767), .A(n14707), .ZN(P2_U2824) );
  AOI22_X1 U18205 ( .A1(n19800), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19813), .ZN(n14709) );
  NAND2_X1 U18206 ( .A1(n19799), .A2(BUF2_REG_31__SCAN_IN), .ZN(n14708) );
  OAI211_X1 U18207 ( .C1(n14695), .C2(n16081), .A(n14709), .B(n14708), .ZN(
        P2_U2888) );
  AOI22_X1 U18208 ( .A1(n14724), .A2(n15097), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n15096), .ZN(n14711) );
  OAI21_X1 U18209 ( .B1(n14710), .B2(n15079), .A(n14711), .ZN(P1_U2843) );
  INV_X1 U18210 ( .A(DATAI_13_), .ZN(n14713) );
  INV_X1 U18211 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14712) );
  MUX2_X1 U18212 ( .A(n14713), .B(n14712), .S(n15135), .Z(n20753) );
  OAI22_X1 U18213 ( .A1(n15177), .A2(n20753), .B1(n14714), .B2(n17230), .ZN(
        n14715) );
  AOI21_X1 U18214 ( .B1(n13615), .B2(DATAI_29_), .A(n14715), .ZN(n14717) );
  NAND2_X1 U18215 ( .A1(n15171), .A2(BUF1_REG_29__SCAN_IN), .ZN(n14716) );
  OAI211_X1 U18216 ( .C1(n14710), .C2(n15195), .A(n14717), .B(n14716), .ZN(
        P1_U2875) );
  INV_X1 U18217 ( .A(n14749), .ZN(n14721) );
  INV_X1 U18218 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21469) );
  AOI22_X1 U18219 ( .A1(n20685), .A2(P1_EBX_REG_29__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20698), .ZN(n14720) );
  NAND3_X1 U18220 ( .A1(n20672), .A2(n14718), .A3(n21469), .ZN(n14719) );
  OAI211_X1 U18221 ( .C1(n14721), .C2(n21469), .A(n14720), .B(n14719), .ZN(
        n14722) );
  AOI21_X1 U18222 ( .B1(n20709), .B2(n14723), .A(n14722), .ZN(n14726) );
  NAND2_X1 U18223 ( .A1(n14724), .A2(n20705), .ZN(n14725) );
  OAI211_X1 U18224 ( .C1(n14710), .C2(n20677), .A(n14726), .B(n14725), .ZN(
        P1_U2811) );
  OR2_X1 U18225 ( .A1(n14878), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n14728) );
  NAND2_X1 U18226 ( .A1(n14731), .A2(n14990), .ZN(n14727) );
  MUX2_X1 U18227 ( .A(n14728), .B(n14727), .S(n21505), .Z(P1_U3487) );
  INV_X1 U18228 ( .A(n14729), .ZN(n14744) );
  MUX2_X1 U18229 ( .A(n14732), .B(n14731), .S(n14730), .Z(n14736) );
  AOI22_X1 U18230 ( .A1(n14733), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n12969), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14734) );
  INV_X1 U18231 ( .A(n14734), .ZN(n14735) );
  AOI22_X1 U18232 ( .A1(n20685), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20698), .ZN(n14739) );
  NAND3_X1 U18233 ( .A1(n14737), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n14740), 
        .ZN(n14738) );
  OAI211_X1 U18234 ( .C1(n14741), .C2(n14740), .A(n14739), .B(n14738), .ZN(
        n14742) );
  OAI21_X1 U18235 ( .B1(n14744), .B2(n20677), .A(n14743), .ZN(P1_U2809) );
  AOI21_X1 U18236 ( .B1(n14755), .B2(n14746), .A(n14745), .ZN(n15200) );
  INV_X1 U18237 ( .A(n15200), .ZN(n15120) );
  AOI22_X1 U18238 ( .A1(n20685), .A2(P1_EBX_REG_28__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20698), .ZN(n14751) );
  OAI21_X1 U18239 ( .B1(n20687), .B2(n14747), .A(n21471), .ZN(n14748) );
  NAND2_X1 U18240 ( .A1(n14749), .A2(n14748), .ZN(n14750) );
  OAI211_X1 U18241 ( .C1(n20691), .C2(n15198), .A(n14751), .B(n14750), .ZN(
        n14752) );
  AOI21_X1 U18242 ( .B1(n15035), .B2(n20705), .A(n14752), .ZN(n14753) );
  OAI21_X1 U18243 ( .B1(n15120), .B2(n20677), .A(n14753), .ZN(P1_U2812) );
  INV_X1 U18244 ( .A(n14755), .ZN(n14756) );
  AOI21_X1 U18245 ( .B1(n14757), .B2(n14754), .A(n14756), .ZN(n15208) );
  INV_X1 U18246 ( .A(n15208), .ZN(n15130) );
  INV_X1 U18247 ( .A(n14758), .ZN(n14759) );
  AOI21_X1 U18248 ( .B1(n14760), .B2(n14772), .A(n14759), .ZN(n15386) );
  INV_X1 U18249 ( .A(n14761), .ZN(n15206) );
  INV_X1 U18250 ( .A(n15001), .ZN(n20660) );
  NOR2_X1 U18251 ( .A1(n14765), .A2(n20687), .ZN(n14762) );
  NOR2_X1 U18252 ( .A1(n20660), .A2(n14762), .ZN(n14776) );
  INV_X1 U18253 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21467) );
  INV_X1 U18254 ( .A(n20698), .ZN(n20646) );
  OAI22_X1 U18255 ( .A1(n14776), .A2(n21467), .B1(n20646), .B2(n14763), .ZN(
        n14764) );
  AOI21_X1 U18256 ( .B1(n20685), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14764), .ZN(
        n14767) );
  NAND3_X1 U18257 ( .A1(n20672), .A2(n14765), .A3(n21467), .ZN(n14766) );
  OAI211_X1 U18258 ( .C1(n20691), .C2(n15206), .A(n14767), .B(n14766), .ZN(
        n14768) );
  AOI21_X1 U18259 ( .B1(n15386), .B2(n20705), .A(n14768), .ZN(n14769) );
  OAI21_X1 U18260 ( .B1(n15130), .B2(n20677), .A(n14769), .ZN(P1_U2813) );
  AOI21_X1 U18261 ( .B1(n14771), .B2(n14770), .A(n11489), .ZN(n15216) );
  INV_X1 U18262 ( .A(n15216), .ZN(n15039) );
  INV_X1 U18263 ( .A(n14772), .ZN(n14773) );
  AOI21_X1 U18264 ( .B1(n14774), .B2(n14793), .A(n14773), .ZN(n15395) );
  AOI22_X1 U18265 ( .A1(n20685), .A2(P1_EBX_REG_26__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20698), .ZN(n14780) );
  NOR2_X1 U18266 ( .A1(n20687), .A2(n14775), .ZN(n14778) );
  INV_X1 U18267 ( .A(n14776), .ZN(n14777) );
  OAI21_X1 U18268 ( .B1(n14778), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14777), 
        .ZN(n14779) );
  OAI211_X1 U18269 ( .C1(n20691), .C2(n15214), .A(n14780), .B(n14779), .ZN(
        n14781) );
  AOI21_X1 U18270 ( .B1(n15395), .B2(n20705), .A(n14781), .ZN(n14782) );
  OAI21_X1 U18271 ( .B1(n15039), .B2(n20677), .A(n14782), .ZN(P1_U2814) );
  AND2_X1 U18272 ( .A1(n14783), .A2(n14838), .ZN(n14785) );
  OAI21_X1 U18273 ( .B1(n14802), .B2(n14786), .A(n14770), .ZN(n15226) );
  INV_X1 U18274 ( .A(n14806), .ZN(n14787) );
  OR2_X1 U18275 ( .A1(n20687), .A2(n14787), .ZN(n14788) );
  AND2_X1 U18276 ( .A1(n14788), .A2(n15001), .ZN(n14821) );
  INV_X1 U18277 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21462) );
  AOI22_X1 U18278 ( .A1(n20685), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20698), .ZN(n14792) );
  NAND2_X1 U18279 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_24__SCAN_IN), 
        .ZN(n14789) );
  OAI211_X1 U18280 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14790), .A(n20672), 
        .B(n14789), .ZN(n14791) );
  OAI211_X1 U18281 ( .C1(n14821), .C2(n21462), .A(n14792), .B(n14791), .ZN(
        n14796) );
  OAI21_X1 U18282 ( .B1(n14800), .B2(n14794), .A(n14793), .ZN(n15406) );
  NOR2_X1 U18283 ( .A1(n15406), .A2(n20650), .ZN(n14795) );
  AOI211_X1 U18284 ( .C1(n20709), .C2(n15223), .A(n14796), .B(n14795), .ZN(
        n14797) );
  OAI21_X1 U18285 ( .B1(n15226), .B2(n20677), .A(n14797), .ZN(P1_U2815) );
  NOR2_X1 U18286 ( .A1(n14815), .A2(n14798), .ZN(n14799) );
  OR2_X1 U18287 ( .A1(n14800), .A2(n14799), .ZN(n15415) );
  NAND2_X1 U18288 ( .A1(n14783), .A2(n14838), .ZN(n14837) );
  NOR2_X1 U18289 ( .A1(n14837), .A2(n14801), .ZN(n14812) );
  INV_X1 U18290 ( .A(n14802), .ZN(n14803) );
  OAI21_X1 U18291 ( .B1(n14804), .B2(n14812), .A(n14803), .ZN(n15233) );
  INV_X1 U18292 ( .A(n15233), .ZN(n14805) );
  NAND2_X1 U18293 ( .A1(n14805), .A2(n13732), .ZN(n14811) );
  AOI22_X1 U18294 ( .A1(n20685), .A2(P1_EBX_REG_24__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n20698), .ZN(n14808) );
  OR3_X1 U18295 ( .A1(n20687), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14806), .ZN(
        n14807) );
  OAI211_X1 U18296 ( .C1(n14821), .C2(n21461), .A(n14808), .B(n14807), .ZN(
        n14809) );
  AOI21_X1 U18297 ( .B1(n20709), .B2(n15230), .A(n14809), .ZN(n14810) );
  OAI211_X1 U18298 ( .C1(n15415), .C2(n20650), .A(n14811), .B(n14810), .ZN(
        P1_U2816) );
  OR2_X1 U18299 ( .A1(n14837), .A2(n14826), .ZN(n14824) );
  AOI21_X1 U18300 ( .B1(n14813), .B2(n14824), .A(n14812), .ZN(n15241) );
  INV_X1 U18301 ( .A(n15241), .ZN(n15149) );
  INV_X1 U18302 ( .A(n14814), .ZN(n14827) );
  AOI21_X1 U18303 ( .B1(n14816), .B2(n14827), .A(n14815), .ZN(n15422) );
  NOR2_X1 U18304 ( .A1(n20687), .A2(n14817), .ZN(n14829) );
  AOI21_X1 U18305 ( .B1(n14829), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n14820) );
  NAND2_X1 U18306 ( .A1(n20709), .A2(n15238), .ZN(n14819) );
  AOI22_X1 U18307 ( .A1(n20685), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20698), .ZN(n14818) );
  OAI211_X1 U18308 ( .C1(n14821), .C2(n14820), .A(n14819), .B(n14818), .ZN(
        n14822) );
  AOI21_X1 U18309 ( .B1(n15422), .B2(n20705), .A(n14822), .ZN(n14823) );
  OAI21_X1 U18310 ( .B1(n15149), .B2(n20677), .A(n14823), .ZN(P1_U2817) );
  INV_X1 U18311 ( .A(n14824), .ZN(n14825) );
  AOI21_X1 U18312 ( .B1(n14826), .B2(n14837), .A(n14825), .ZN(n15249) );
  INV_X1 U18313 ( .A(n15249), .ZN(n15154) );
  AOI21_X1 U18314 ( .B1(n14828), .B2(n9600), .A(n14814), .ZN(n15438) );
  NOR2_X1 U18315 ( .A1(n20691), .A2(n15247), .ZN(n14835) );
  INV_X1 U18316 ( .A(n14829), .ZN(n14833) );
  OAI21_X1 U18317 ( .B1(n20687), .B2(n14839), .A(n15001), .ZN(n14855) );
  NOR2_X1 U18318 ( .A1(n20687), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14830) );
  OAI21_X1 U18319 ( .B1(n14855), .B2(n14830), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14832) );
  AOI22_X1 U18320 ( .A1(n20685), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20698), .ZN(n14831) );
  OAI211_X1 U18321 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n14833), .A(n14832), 
        .B(n14831), .ZN(n14834) );
  AOI211_X1 U18322 ( .C1(n15438), .C2(n20705), .A(n14835), .B(n14834), .ZN(
        n14836) );
  OAI21_X1 U18323 ( .B1(n15154), .B2(n20677), .A(n14836), .ZN(P1_U2818) );
  OAI21_X1 U18324 ( .B1(n14783), .B2(n14838), .A(n14837), .ZN(n15258) );
  INV_X1 U18325 ( .A(n14855), .ZN(n14842) );
  INV_X1 U18326 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n21456) );
  AOI22_X1 U18327 ( .A1(n20685), .A2(P1_EBX_REG_21__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20698), .ZN(n14841) );
  NAND3_X1 U18328 ( .A1(n20672), .A2(n14839), .A3(n21456), .ZN(n14840) );
  OAI211_X1 U18329 ( .C1(n14842), .C2(n21456), .A(n14841), .B(n14840), .ZN(
        n14846) );
  OAI21_X1 U18330 ( .B1(n14843), .B2(n14844), .A(n9600), .ZN(n15449) );
  NOR2_X1 U18331 ( .A1(n15449), .A2(n20650), .ZN(n14845) );
  AOI211_X1 U18332 ( .C1(n20709), .C2(n15255), .A(n14846), .B(n14845), .ZN(
        n14847) );
  OAI21_X1 U18333 ( .B1(n15258), .B2(n20677), .A(n14847), .ZN(P1_U2819) );
  NOR2_X1 U18334 ( .A1(n14848), .A2(n14849), .ZN(n14850) );
  INV_X1 U18335 ( .A(n15262), .ZN(n14860) );
  NOR2_X1 U18336 ( .A1(n14851), .A2(n14852), .ZN(n14853) );
  OR2_X1 U18337 ( .A1(n14843), .A2(n14853), .ZN(n15461) );
  AOI22_X1 U18338 ( .A1(n20685), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20698), .ZN(n14858) );
  NOR2_X1 U18339 ( .A1(n20687), .A2(n14854), .ZN(n14856) );
  OAI21_X1 U18340 ( .B1(n14856), .B2(P1_REIP_REG_20__SCAN_IN), .A(n14855), 
        .ZN(n14857) );
  OAI211_X1 U18341 ( .C1(n15461), .C2(n20650), .A(n14858), .B(n14857), .ZN(
        n14859) );
  AOI21_X1 U18342 ( .B1(n14860), .B2(n20709), .A(n14859), .ZN(n14861) );
  OAI21_X1 U18343 ( .B1(n15266), .B2(n20677), .A(n14861), .ZN(P1_U2820) );
  AND2_X1 U18344 ( .A1(n14862), .A2(n14863), .ZN(n14864) );
  OR2_X1 U18345 ( .A1(n14864), .A2(n14848), .ZN(n15277) );
  AND2_X1 U18346 ( .A1(n9619), .A2(n14865), .ZN(n14866) );
  NOR2_X1 U18347 ( .A1(n14851), .A2(n14866), .ZN(n15469) );
  AND2_X1 U18348 ( .A1(n17202), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n14867) );
  NAND2_X1 U18349 ( .A1(n20652), .A2(n14867), .ZN(n17201) );
  INV_X1 U18350 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15290) );
  INV_X1 U18351 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21447) );
  OR3_X1 U18352 ( .A1(n17201), .A2(n15290), .A3(n21447), .ZN(n14903) );
  INV_X1 U18353 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15269) );
  NAND3_X1 U18354 ( .A1(n15269), .A2(P1_REIP_REG_17__SCAN_IN), .A3(
        P1_REIP_REG_18__SCAN_IN), .ZN(n14883) );
  INV_X1 U18355 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21451) );
  NAND2_X1 U18356 ( .A1(n21451), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n14868) );
  OR2_X1 U18357 ( .A1(n14903), .A2(n14868), .ZN(n14888) );
  INV_X1 U18358 ( .A(n14869), .ZN(n14870) );
  AND2_X1 U18359 ( .A1(n15001), .A2(n14870), .ZN(n14980) );
  INV_X1 U18360 ( .A(n14871), .ZN(n14872) );
  AND2_X1 U18361 ( .A1(n14980), .A2(n14872), .ZN(n14873) );
  OR2_X1 U18362 ( .A1(n14981), .A2(n14873), .ZN(n17212) );
  INV_X1 U18363 ( .A(n14874), .ZN(n14875) );
  OR2_X1 U18364 ( .A1(n14981), .A2(n14875), .ZN(n14876) );
  AND2_X1 U18365 ( .A1(n17212), .A2(n14876), .ZN(n14902) );
  NAND2_X1 U18366 ( .A1(n14888), .A2(n14902), .ZN(n14877) );
  NAND2_X1 U18367 ( .A1(n14877), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14882) );
  NAND2_X1 U18368 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14879) );
  NAND2_X1 U18369 ( .A1(n15001), .A2(n14878), .ZN(n20688) );
  NAND2_X1 U18370 ( .A1(n14879), .A2(n20688), .ZN(n14880) );
  AOI21_X1 U18371 ( .B1(n20685), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14880), .ZN(
        n14881) );
  OAI211_X1 U18372 ( .C1(n14903), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n14884) );
  AOI21_X1 U18373 ( .B1(n15469), .B2(n20705), .A(n14884), .ZN(n14886) );
  NAND2_X1 U18374 ( .A1(n20709), .A2(n15273), .ZN(n14885) );
  OAI211_X1 U18375 ( .C1(n15277), .C2(n20677), .A(n14886), .B(n14885), .ZN(
        P1_U2821) );
  OAI21_X1 U18376 ( .B1(n11262), .B2(n10423), .A(n14862), .ZN(n15284) );
  INV_X1 U18377 ( .A(n15278), .ZN(n14895) );
  INV_X1 U18378 ( .A(n20688), .ZN(n20662) );
  INV_X1 U18379 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15047) );
  NOR2_X1 U18380 ( .A1(n17214), .A2(n15047), .ZN(n14887) );
  AOI211_X1 U18381 ( .C1(n20698), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20662), .B(n14887), .ZN(n14889) );
  OAI211_X1 U18382 ( .C1(n14902), .C2(n21451), .A(n14889), .B(n14888), .ZN(
        n14894) );
  INV_X1 U18383 ( .A(n14891), .ZN(n14892) );
  OAI21_X1 U18384 ( .B1(n10321), .B2(n14892), .A(n9619), .ZN(n15484) );
  NOR2_X1 U18385 ( .A1(n15484), .A2(n20650), .ZN(n14893) );
  AOI211_X1 U18386 ( .C1(n20709), .C2(n14895), .A(n14894), .B(n14893), .ZN(
        n14896) );
  OAI21_X1 U18387 ( .B1(n15284), .B2(n20677), .A(n14896), .ZN(P1_U2822) );
  NAND2_X1 U18388 ( .A1(n14897), .A2(n13732), .ZN(n14908) );
  OR2_X1 U18389 ( .A1(n10434), .A2(n14898), .ZN(n14899) );
  AND2_X1 U18390 ( .A1(n14890), .A2(n14899), .ZN(n15489) );
  NAND2_X1 U18391 ( .A1(n20685), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14900) );
  OAI211_X1 U18392 ( .C1(n20646), .C2(n14901), .A(n14900), .B(n20688), .ZN(
        n14906) );
  AOI21_X1 U18393 ( .B1(n14904), .B2(n14903), .A(n14902), .ZN(n14905) );
  AOI211_X1 U18394 ( .C1(n15489), .C2(n20705), .A(n14906), .B(n14905), .ZN(
        n14907) );
  OAI211_X1 U18395 ( .C1(n20691), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        P1_U2823) );
  AOI21_X1 U18396 ( .B1(n14912), .B2(n14910), .A(n14911), .ZN(n15294) );
  NAND2_X1 U18397 ( .A1(n15294), .A2(n13732), .ZN(n14921) );
  AOI21_X1 U18398 ( .B1(n14913), .B2(n9695), .A(n10434), .ZN(n15499) );
  OAI21_X1 U18399 ( .B1(n20646), .B2(n14914), .A(n20688), .ZN(n14917) );
  XNOR2_X1 U18400 ( .A(P1_REIP_REG_16__SCAN_IN), .B(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n14915) );
  NOR2_X1 U18401 ( .A1(n17201), .A2(n14915), .ZN(n14916) );
  AOI211_X1 U18402 ( .C1(P1_EBX_REG_16__SCAN_IN), .C2(n20685), .A(n14917), .B(
        n14916), .ZN(n14918) );
  OAI21_X1 U18403 ( .B1(n15290), .B2(n17212), .A(n14918), .ZN(n14919) );
  AOI21_X1 U18404 ( .B1(n20705), .B2(n15499), .A(n14919), .ZN(n14920) );
  OAI211_X1 U18405 ( .C1(n20691), .C2(n15292), .A(n14921), .B(n14920), .ZN(
        P1_U2824) );
  INV_X1 U18406 ( .A(n14922), .ZN(n14960) );
  NAND2_X1 U18407 ( .A1(n14960), .A2(n14923), .ZN(n14924) );
  OAI21_X1 U18408 ( .B1(n14960), .B2(n14923), .A(n14924), .ZN(n15072) );
  INV_X1 U18409 ( .A(n15071), .ZN(n14925) );
  OAI21_X1 U18410 ( .B1(n15072), .B2(n14925), .A(n14924), .ZN(n14944) );
  NAND2_X1 U18411 ( .A1(n14944), .A2(n14943), .ZN(n14942) );
  INV_X1 U18412 ( .A(n14926), .ZN(n14928) );
  OAI21_X1 U18413 ( .B1(n14925), .B2(n14922), .A(n14924), .ZN(n14927) );
  AOI21_X1 U18414 ( .B1(n14942), .B2(n14928), .A(n15054), .ZN(n15322) );
  INV_X1 U18415 ( .A(n15322), .ZN(n15185) );
  INV_X1 U18416 ( .A(n15320), .ZN(n14940) );
  OAI21_X1 U18417 ( .B1(n14929), .B2(n14930), .A(n15063), .ZN(n15067) );
  INV_X1 U18418 ( .A(n15067), .ZN(n15523) );
  AOI22_X1 U18419 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n20685), .B1(n20705), 
        .B2(n15523), .ZN(n14931) );
  OAI211_X1 U18420 ( .C1(n20646), .C2(n14932), .A(n14931), .B(n20688), .ZN(
        n14939) );
  NAND2_X1 U18421 ( .A1(n20652), .A2(n14933), .ZN(n14950) );
  NOR2_X1 U18422 ( .A1(n14935), .A2(n14950), .ZN(n14937) );
  INV_X1 U18423 ( .A(n14981), .ZN(n15027) );
  AND2_X1 U18424 ( .A1(n14980), .A2(n14933), .ZN(n14934) );
  NOR2_X1 U18425 ( .A1(n14981), .A2(n14934), .ZN(n17218) );
  AOI21_X1 U18426 ( .B1(n15027), .B2(n14935), .A(n17218), .ZN(n14952) );
  INV_X1 U18427 ( .A(n14952), .ZN(n14936) );
  MUX2_X1 U18428 ( .A(n14937), .B(n14936), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14938) );
  AOI211_X1 U18429 ( .C1(n20709), .C2(n14940), .A(n14939), .B(n14938), .ZN(
        n14941) );
  OAI21_X1 U18430 ( .B1(n15185), .B2(n20677), .A(n14941), .ZN(P1_U2827) );
  OAI21_X1 U18431 ( .B1(n14944), .B2(n14943), .A(n14942), .ZN(n15332) );
  INV_X1 U18432 ( .A(n15332), .ZN(n14945) );
  NAND2_X1 U18433 ( .A1(n14945), .A2(n13732), .ZN(n14956) );
  NOR2_X1 U18434 ( .A1(n14946), .A2(n14947), .ZN(n14948) );
  OR2_X1 U18435 ( .A1(n14929), .A2(n14948), .ZN(n15069) );
  INV_X1 U18436 ( .A(n15069), .ZN(n15528) );
  AOI21_X1 U18437 ( .B1(n20698), .B2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n20662), .ZN(n14949) );
  OAI21_X1 U18438 ( .B1(n17214), .B2(n15070), .A(n14949), .ZN(n14954) );
  INV_X1 U18439 ( .A(n14950), .ZN(n17219) );
  AOI21_X1 U18440 ( .B1(n17219), .B2(P1_REIP_REG_11__SCAN_IN), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14951) );
  NOR2_X1 U18441 ( .A1(n14952), .A2(n14951), .ZN(n14953) );
  AOI211_X1 U18442 ( .C1(n15528), .C2(n20705), .A(n14954), .B(n14953), .ZN(
        n14955) );
  OAI211_X1 U18443 ( .C1(n20691), .C2(n15328), .A(n14956), .B(n14955), .ZN(
        P1_U2828) );
  INV_X1 U18444 ( .A(n14957), .ZN(n15091) );
  INV_X1 U18445 ( .A(n14974), .ZN(n14958) );
  NAND2_X1 U18446 ( .A1(n15082), .A2(n15081), .ZN(n15080) );
  INV_X1 U18447 ( .A(n14959), .ZN(n14961) );
  AOI21_X1 U18448 ( .B1(n15080), .B2(n14961), .A(n14960), .ZN(n15351) );
  INV_X1 U18449 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21439) );
  NOR2_X1 U18450 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n21439), .ZN(n14968) );
  NAND2_X1 U18451 ( .A1(n15086), .A2(n14962), .ZN(n14963) );
  NAND2_X1 U18452 ( .A1(n15074), .A2(n14963), .ZN(n15561) );
  INV_X1 U18453 ( .A(n15561), .ZN(n14964) );
  AOI22_X1 U18454 ( .A1(n20705), .A2(n14964), .B1(n20685), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n14965) );
  OAI211_X1 U18455 ( .C1(n20646), .C2(n14966), .A(n14965), .B(n20688), .ZN(
        n14967) );
  AOI21_X1 U18456 ( .B1(n20652), .B2(n14968), .A(n14967), .ZN(n14970) );
  NAND2_X1 U18457 ( .A1(n17218), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U18458 ( .C1(n20691), .C2(n15349), .A(n14970), .B(n14969), .ZN(
        n14971) );
  AOI21_X1 U18459 ( .B1(n15351), .B2(n13732), .A(n14971), .ZN(n14972) );
  INV_X1 U18460 ( .A(n14972), .ZN(P1_U2830) );
  INV_X1 U18461 ( .A(n15094), .ZN(n14975) );
  INV_X1 U18462 ( .A(n15082), .ZN(n14973) );
  INV_X1 U18463 ( .A(n15361), .ZN(n14988) );
  INV_X1 U18464 ( .A(n14976), .ZN(n14978) );
  AOI21_X1 U18465 ( .B1(n14978), .B2(n15095), .A(n14977), .ZN(n14979) );
  OR2_X1 U18466 ( .A1(n14979), .A2(n15084), .ZN(n17252) );
  NOR2_X1 U18467 ( .A1(n14981), .A2(n14980), .ZN(n20653) );
  AOI21_X1 U18468 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20653), .A(n20662), .ZN(
        n14983) );
  NAND2_X1 U18469 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14982) );
  OAI211_X1 U18470 ( .C1(n20650), .C2(n17252), .A(n14983), .B(n14982), .ZN(
        n14987) );
  INV_X1 U18471 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21436) );
  NAND3_X1 U18472 ( .A1(n20672), .A2(n14984), .A3(n21436), .ZN(n14985) );
  OAI21_X1 U18473 ( .B1(n17214), .B2(n15088), .A(n14985), .ZN(n14986) );
  AOI211_X1 U18474 ( .C1(n20709), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        n14989) );
  OAI21_X1 U18475 ( .B1(n15365), .B2(n20677), .A(n14989), .ZN(P1_U2832) );
  INV_X1 U18476 ( .A(n17245), .ZN(n14991) );
  NAND2_X1 U18477 ( .A1(n14991), .A2(n20710), .ZN(n15000) );
  NOR3_X1 U18478 ( .A1(n20687), .A2(P1_REIP_REG_5__SCAN_IN), .A3(n14992), .ZN(
        n14997) );
  AOI21_X1 U18479 ( .B1(n20672), .B2(n14992), .A(n20660), .ZN(n20696) );
  OAI21_X1 U18480 ( .B1(n20696), .B2(n21431), .A(n20688), .ZN(n14993) );
  AOI21_X1 U18481 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n20698), .A(
        n14993), .ZN(n14994) );
  OAI21_X1 U18482 ( .B1(n17214), .B2(n14995), .A(n14994), .ZN(n14996) );
  AOI211_X1 U18483 ( .C1(n14998), .C2(n20705), .A(n14997), .B(n14996), .ZN(
        n14999) );
  OAI211_X1 U18484 ( .C1(n20691), .C2(n17250), .A(n15000), .B(n14999), .ZN(
        P1_U2835) );
  OR2_X1 U18485 ( .A1(n20687), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15002) );
  NAND2_X1 U18486 ( .A1(n15002), .A2(n15001), .ZN(n20712) );
  NOR2_X1 U18487 ( .A1(n20687), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20713) );
  NAND2_X1 U18488 ( .A1(n20713), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n15008) );
  NOR2_X1 U18489 ( .A1(n15004), .A2(n15003), .ZN(n15014) );
  AOI22_X1 U18490 ( .A1(n15014), .A2(n15005), .B1(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20698), .ZN(n15007) );
  AOI22_X1 U18491 ( .A1(n10433), .A2(n20705), .B1(n20685), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n15006) );
  NAND3_X1 U18492 ( .A1(n15008), .A2(n15007), .A3(n15006), .ZN(n15011) );
  NOR2_X1 U18493 ( .A1(n20691), .A2(n15009), .ZN(n15010) );
  AOI211_X1 U18494 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n20712), .A(n15011), .B(
        n15010), .ZN(n15012) );
  OAI21_X1 U18495 ( .B1(n20692), .B2(n15013), .A(n15012), .ZN(P1_U2838) );
  INV_X1 U18496 ( .A(n15014), .ZN(n20701) );
  NAND2_X1 U18497 ( .A1(n20685), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n15016) );
  AOI22_X1 U18498 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20660), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n15015) );
  OAI211_X1 U18499 ( .C1(n20701), .C2(n14504), .A(n15016), .B(n15015), .ZN(
        n15019) );
  INV_X1 U18500 ( .A(n14073), .ZN(n15017) );
  OAI22_X1 U18501 ( .A1(n20650), .A2(n15017), .B1(P1_REIP_REG_1__SCAN_IN), 
        .B2(n20687), .ZN(n15018) );
  AOI211_X1 U18502 ( .C1(n20709), .C2(n15020), .A(n15019), .B(n15018), .ZN(
        n15021) );
  OAI21_X1 U18503 ( .B1(n20692), .B2(n15022), .A(n15021), .ZN(P1_U2839) );
  NOR2_X1 U18504 ( .A1(n20650), .A2(n15023), .ZN(n15026) );
  OAI22_X1 U18505 ( .A1(n17214), .A2(n12938), .B1(n15024), .B2(n20701), .ZN(
        n15025) );
  AOI211_X1 U18506 ( .C1(P1_REIP_REG_0__SCAN_IN), .C2(n15027), .A(n15026), .B(
        n15025), .ZN(n15029) );
  OAI21_X1 U18507 ( .B1(n20709), .B2(n20698), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15028) );
  OAI211_X1 U18508 ( .C1(n20692), .C2(n15030), .A(n15029), .B(n15028), .ZN(
        P1_U2840) );
  INV_X1 U18509 ( .A(n15376), .ZN(n15031) );
  INV_X1 U18510 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n21572) );
  OAI22_X1 U18511 ( .A1(n15031), .A2(n15105), .B1(n15104), .B2(n21572), .ZN(
        P1_U2841) );
  INV_X1 U18512 ( .A(n15032), .ZN(n15114) );
  INV_X1 U18513 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15034) );
  OAI222_X1 U18514 ( .A1(n15079), .A2(n15114), .B1(n15034), .B2(n15104), .C1(
        n15105), .C2(n15033), .ZN(P1_U2842) );
  AOI22_X1 U18515 ( .A1(n15035), .A2(n15097), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15096), .ZN(n15036) );
  OAI21_X1 U18516 ( .B1(n15120), .B2(n15099), .A(n15036), .ZN(P1_U2844) );
  AOI22_X1 U18517 ( .A1(n15386), .A2(n15097), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15096), .ZN(n15037) );
  OAI21_X1 U18518 ( .B1(n15130), .B2(n15099), .A(n15037), .ZN(P1_U2845) );
  AOI22_X1 U18519 ( .A1(n15395), .A2(n15097), .B1(P1_EBX_REG_26__SCAN_IN), 
        .B2(n15096), .ZN(n15038) );
  OAI21_X1 U18520 ( .B1(n15039), .B2(n15099), .A(n15038), .ZN(P1_U2846) );
  INV_X1 U18521 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15040) );
  OAI222_X1 U18522 ( .A1(n15079), .A2(n15226), .B1(n15040), .B2(n15104), .C1(
        n15406), .C2(n15105), .ZN(P1_U2847) );
  INV_X1 U18523 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15041) );
  OAI222_X1 U18524 ( .A1(n15079), .A2(n15233), .B1(n15041), .B2(n15104), .C1(
        n15415), .C2(n15105), .ZN(P1_U2848) );
  AOI22_X1 U18525 ( .A1(n15422), .A2(n15097), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n15096), .ZN(n15042) );
  OAI21_X1 U18526 ( .B1(n15149), .B2(n15099), .A(n15042), .ZN(P1_U2849) );
  AOI22_X1 U18527 ( .A1(n15438), .A2(n15097), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n15096), .ZN(n15043) );
  OAI21_X1 U18528 ( .B1(n15154), .B2(n15099), .A(n15043), .ZN(P1_U2850) );
  INV_X1 U18529 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15044) );
  OAI222_X1 U18530 ( .A1(n15258), .A2(n15099), .B1(n15044), .B2(n15104), .C1(
        n15449), .C2(n15105), .ZN(P1_U2851) );
  OAI222_X1 U18531 ( .A1(n15266), .A2(n15099), .B1(n15045), .B2(n15104), .C1(
        n15461), .C2(n15105), .ZN(P1_U2852) );
  AOI22_X1 U18532 ( .A1(n15469), .A2(n15097), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15096), .ZN(n15046) );
  OAI21_X1 U18533 ( .B1(n15277), .B2(n15099), .A(n15046), .ZN(P1_U2853) );
  OAI222_X1 U18534 ( .A1(n15284), .A2(n15079), .B1(n15047), .B2(n15104), .C1(
        n15484), .C2(n15105), .ZN(P1_U2854) );
  INV_X1 U18535 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15049) );
  INV_X1 U18536 ( .A(n15489), .ZN(n15048) );
  OAI222_X1 U18537 ( .A1(n15079), .A2(n15174), .B1(n15104), .B2(n15049), .C1(
        n15048), .C2(n15105), .ZN(P1_U2855) );
  INV_X1 U18538 ( .A(n15294), .ZN(n15051) );
  AOI22_X1 U18539 ( .A1(n15499), .A2(n15097), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n15096), .ZN(n15050) );
  OAI21_X1 U18540 ( .B1(n15051), .B2(n15079), .A(n15050), .ZN(P1_U2856) );
  NAND2_X1 U18541 ( .A1(n15061), .A2(n15052), .ZN(n15053) );
  AND2_X1 U18542 ( .A1(n9695), .A2(n15053), .ZN(n17195) );
  INV_X1 U18543 ( .A(n17195), .ZN(n15057) );
  INV_X1 U18544 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15056) );
  NOR2_X1 U18545 ( .A1(n15059), .A2(n15060), .ZN(n15058) );
  OAI21_X1 U18546 ( .B1(n15058), .B2(n15055), .A(n14910), .ZN(n17190) );
  OAI222_X1 U18547 ( .A1(n15057), .A2(n15105), .B1(n15104), .B2(n15056), .C1(
        n17190), .C2(n15079), .ZN(P1_U2857) );
  AOI21_X1 U18548 ( .B1(n15060), .B2(n15059), .A(n15058), .ZN(n17228) );
  INV_X1 U18549 ( .A(n17228), .ZN(n15066) );
  INV_X1 U18550 ( .A(n15061), .ZN(n15062) );
  AOI21_X1 U18551 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n17206) );
  AOI22_X1 U18552 ( .A1(n17206), .A2(n15097), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n15096), .ZN(n15065) );
  OAI21_X1 U18553 ( .B1(n15066), .B2(n15079), .A(n15065), .ZN(P1_U2858) );
  INV_X1 U18554 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n15068) );
  OAI222_X1 U18555 ( .A1(n15185), .A2(n15079), .B1(n15104), .B2(n15068), .C1(
        n15067), .C2(n15105), .ZN(P1_U2859) );
  OAI222_X1 U18556 ( .A1(n15332), .A2(n15099), .B1(n15070), .B2(n15104), .C1(
        n15069), .C2(n15105), .ZN(P1_U2860) );
  XNOR2_X1 U18557 ( .A(n15072), .B(n15071), .ZN(n17220) );
  AND2_X1 U18558 ( .A1(n15074), .A2(n15073), .ZN(n15075) );
  OR2_X1 U18559 ( .A1(n15075), .A2(n14946), .ZN(n17213) );
  OAI22_X1 U18560 ( .A1(n17213), .A2(n15105), .B1(n17215), .B2(n15104), .ZN(
        n15076) );
  AOI21_X1 U18561 ( .B1(n17220), .B2(n15107), .A(n15076), .ZN(n15077) );
  INV_X1 U18562 ( .A(n15077), .ZN(P1_U2861) );
  INV_X1 U18563 ( .A(n15351), .ZN(n15191) );
  INV_X1 U18564 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15078) );
  OAI222_X1 U18565 ( .A1(n15191), .A2(n15079), .B1(n15078), .B2(n15104), .C1(
        n15561), .C2(n15105), .ZN(P1_U2862) );
  OAI21_X1 U18566 ( .B1(n15082), .B2(n15081), .A(n15080), .ZN(n20654) );
  INV_X1 U18567 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n15087) );
  OR2_X1 U18568 ( .A1(n15084), .A2(n15083), .ZN(n15085) );
  NAND2_X1 U18569 ( .A1(n15086), .A2(n15085), .ZN(n20649) );
  OAI222_X1 U18570 ( .A1(n20654), .A2(n15099), .B1(n15087), .B2(n15104), .C1(
        n20649), .C2(n15105), .ZN(P1_U2863) );
  OAI22_X1 U18571 ( .A1(n17252), .A2(n15105), .B1(n15088), .B2(n15104), .ZN(
        n15089) );
  INV_X1 U18572 ( .A(n15089), .ZN(n15090) );
  OAI21_X1 U18573 ( .B1(n15365), .B2(n15099), .A(n15090), .ZN(P1_U2864) );
  NAND2_X1 U18574 ( .A1(n15092), .A2(n15091), .ZN(n15093) );
  INV_X1 U18575 ( .A(n20668), .ZN(n15194) );
  XNOR2_X1 U18576 ( .A(n14976), .B(n15095), .ZN(n20663) );
  AOI22_X1 U18577 ( .A1(n15097), .A2(n20663), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n15096), .ZN(n15098) );
  OAI21_X1 U18578 ( .B1(n15194), .B2(n15099), .A(n15098), .ZN(P1_U2865) );
  NAND2_X1 U18579 ( .A1(n14477), .A2(n15101), .ZN(n15102) );
  NAND2_X1 U18580 ( .A1(n14976), .A2(n15102), .ZN(n17265) );
  OAI22_X1 U18581 ( .A1(n17265), .A2(n15105), .B1(n15104), .B2(n15103), .ZN(
        n15106) );
  AOI21_X1 U18582 ( .B1(n17241), .B2(n15107), .A(n15106), .ZN(n15108) );
  INV_X1 U18583 ( .A(n15108), .ZN(P1_U2866) );
  INV_X1 U18584 ( .A(DATAI_14_), .ZN(n15110) );
  INV_X1 U18585 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n15109) );
  MUX2_X1 U18586 ( .A(n15110), .B(n15109), .S(n15135), .Z(n17224) );
  OAI22_X1 U18587 ( .A1(n15177), .A2(n17224), .B1(n14010), .B2(n17230), .ZN(
        n15111) );
  AOI21_X1 U18588 ( .B1(n13615), .B2(DATAI_30_), .A(n15111), .ZN(n15113) );
  NAND2_X1 U18589 ( .A1(n15171), .A2(BUF1_REG_30__SCAN_IN), .ZN(n15112) );
  OAI211_X1 U18590 ( .C1(n15114), .C2(n15195), .A(n15113), .B(n15112), .ZN(
        P1_U2874) );
  INV_X1 U18591 ( .A(DATAI_12_), .ZN(n15116) );
  INV_X1 U18592 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n15115) );
  MUX2_X1 U18593 ( .A(n15116), .B(n15115), .S(n15135), .Z(n20750) );
  OAI22_X1 U18594 ( .A1(n15177), .A2(n20750), .B1(n14001), .B2(n17230), .ZN(
        n15117) );
  AOI21_X1 U18595 ( .B1(n13615), .B2(DATAI_28_), .A(n15117), .ZN(n15119) );
  NAND2_X1 U18596 ( .A1(n15171), .A2(BUF1_REG_28__SCAN_IN), .ZN(n15118) );
  OAI211_X1 U18597 ( .C1(n15120), .C2(n15195), .A(n15119), .B(n15118), .ZN(
        P1_U2876) );
  INV_X1 U18598 ( .A(n13615), .ZN(n15127) );
  INV_X1 U18599 ( .A(DATAI_27_), .ZN(n15126) );
  INV_X1 U18600 ( .A(n15177), .ZN(n15124) );
  INV_X1 U18601 ( .A(DATAI_11_), .ZN(n15122) );
  NAND2_X1 U18602 ( .A1(n15135), .A2(BUF1_REG_11__SCAN_IN), .ZN(n15121) );
  OAI21_X1 U18603 ( .B1(n15135), .B2(n15122), .A(n15121), .ZN(n20748) );
  AOI22_X1 U18604 ( .A1(n15124), .A2(n20748), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15123), .ZN(n15125) );
  OAI21_X1 U18605 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15128) );
  AOI21_X1 U18606 ( .B1(n15171), .B2(BUF1_REG_27__SCAN_IN), .A(n15128), .ZN(
        n15129) );
  OAI21_X1 U18607 ( .B1(n15130), .B2(n15195), .A(n15129), .ZN(P1_U2877) );
  INV_X1 U18608 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n19991) );
  INV_X1 U18609 ( .A(n15195), .ZN(n17227) );
  NAND2_X1 U18610 ( .A1(n15216), .A2(n17227), .ZN(n15134) );
  INV_X1 U18611 ( .A(DATAI_10_), .ZN(n15131) );
  INV_X1 U18612 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n21596) );
  MUX2_X1 U18613 ( .A(n15131), .B(n21596), .S(n15135), .Z(n20745) );
  OAI22_X1 U18614 ( .A1(n15177), .A2(n20745), .B1(n14007), .B2(n17230), .ZN(
        n15132) );
  AOI21_X1 U18615 ( .B1(n13615), .B2(DATAI_26_), .A(n15132), .ZN(n15133) );
  OAI211_X1 U18616 ( .C1(n19991), .C2(n15181), .A(n15134), .B(n15133), .ZN(
        P1_U2878) );
  INV_X1 U18617 ( .A(DATAI_9_), .ZN(n15137) );
  INV_X1 U18618 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n15136) );
  MUX2_X1 U18619 ( .A(n15137), .B(n15136), .S(n15135), .Z(n20742) );
  OAI22_X1 U18620 ( .A1(n15177), .A2(n20742), .B1(n15138), .B2(n17230), .ZN(
        n15139) );
  AOI21_X1 U18621 ( .B1(n13615), .B2(DATAI_25_), .A(n15139), .ZN(n15141) );
  NAND2_X1 U18622 ( .A1(n15171), .A2(BUF1_REG_25__SCAN_IN), .ZN(n15140) );
  OAI211_X1 U18623 ( .C1(n15226), .C2(n15195), .A(n15141), .B(n15140), .ZN(
        P1_U2879) );
  OAI22_X1 U18624 ( .A1(n15177), .A2(n15193), .B1(n15142), .B2(n17230), .ZN(
        n15143) );
  AOI21_X1 U18625 ( .B1(n15171), .B2(BUF1_REG_24__SCAN_IN), .A(n15143), .ZN(
        n15145) );
  NAND2_X1 U18626 ( .A1(n13615), .A2(DATAI_24_), .ZN(n15144) );
  OAI211_X1 U18627 ( .C1(n15233), .C2(n15195), .A(n15145), .B(n15144), .ZN(
        P1_U2880) );
  OAI22_X1 U18628 ( .A1(n15177), .A2(n20857), .B1(n21555), .B2(n17230), .ZN(
        n15146) );
  AOI21_X1 U18629 ( .B1(n13615), .B2(DATAI_23_), .A(n15146), .ZN(n15148) );
  NAND2_X1 U18630 ( .A1(n15171), .A2(BUF1_REG_23__SCAN_IN), .ZN(n15147) );
  OAI211_X1 U18631 ( .C1(n15149), .C2(n15195), .A(n15148), .B(n15147), .ZN(
        P1_U2881) );
  OAI22_X1 U18632 ( .A1(n15177), .A2(n20844), .B1(n15150), .B2(n17230), .ZN(
        n15151) );
  AOI21_X1 U18633 ( .B1(n13615), .B2(DATAI_22_), .A(n15151), .ZN(n15153) );
  NAND2_X1 U18634 ( .A1(n15171), .A2(BUF1_REG_22__SCAN_IN), .ZN(n15152) );
  OAI211_X1 U18635 ( .C1(n15154), .C2(n15195), .A(n15153), .B(n15152), .ZN(
        P1_U2882) );
  OAI22_X1 U18636 ( .A1(n15177), .A2(n20840), .B1(n15155), .B2(n17230), .ZN(
        n15156) );
  AOI21_X1 U18637 ( .B1(n13615), .B2(DATAI_21_), .A(n15156), .ZN(n15158) );
  NAND2_X1 U18638 ( .A1(n15171), .A2(BUF1_REG_21__SCAN_IN), .ZN(n15157) );
  OAI211_X1 U18639 ( .C1(n15258), .C2(n15195), .A(n15158), .B(n15157), .ZN(
        P1_U2883) );
  OAI22_X1 U18640 ( .A1(n15177), .A2(n20835), .B1(n14249), .B2(n17230), .ZN(
        n15159) );
  AOI21_X1 U18641 ( .B1(n13615), .B2(DATAI_20_), .A(n15159), .ZN(n15161) );
  NAND2_X1 U18642 ( .A1(n15171), .A2(BUF1_REG_20__SCAN_IN), .ZN(n15160) );
  OAI211_X1 U18643 ( .C1(n15266), .C2(n15195), .A(n15161), .B(n15160), .ZN(
        P1_U2884) );
  OAI22_X1 U18644 ( .A1(n15177), .A2(n20830), .B1(n14242), .B2(n17230), .ZN(
        n15162) );
  AOI21_X1 U18645 ( .B1(n13615), .B2(DATAI_19_), .A(n15162), .ZN(n15164) );
  NAND2_X1 U18646 ( .A1(n15171), .A2(BUF1_REG_19__SCAN_IN), .ZN(n15163) );
  OAI211_X1 U18647 ( .C1(n15277), .C2(n15195), .A(n15164), .B(n15163), .ZN(
        P1_U2885) );
  OAI22_X1 U18648 ( .A1(n15177), .A2(n20826), .B1(n15165), .B2(n17230), .ZN(
        n15166) );
  AOI21_X1 U18649 ( .B1(n13615), .B2(DATAI_18_), .A(n15166), .ZN(n15168) );
  NAND2_X1 U18650 ( .A1(n15171), .A2(BUF1_REG_18__SCAN_IN), .ZN(n15167) );
  OAI211_X1 U18651 ( .C1(n15284), .C2(n15195), .A(n15168), .B(n15167), .ZN(
        P1_U2886) );
  OAI22_X1 U18652 ( .A1(n15177), .A2(n20821), .B1(n15169), .B2(n17230), .ZN(
        n15170) );
  AOI21_X1 U18653 ( .B1(n13615), .B2(DATAI_17_), .A(n15170), .ZN(n15173) );
  NAND2_X1 U18654 ( .A1(n15171), .A2(BUF1_REG_17__SCAN_IN), .ZN(n15172) );
  OAI211_X1 U18655 ( .C1(n15174), .C2(n15195), .A(n15173), .B(n15172), .ZN(
        P1_U2887) );
  INV_X1 U18656 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n17344) );
  NAND2_X1 U18657 ( .A1(n15294), .A2(n17227), .ZN(n15180) );
  OAI22_X1 U18658 ( .A1(n15177), .A2(n15176), .B1(n15175), .B2(n17230), .ZN(
        n15178) );
  AOI21_X1 U18659 ( .B1(n13615), .B2(DATAI_16_), .A(n15178), .ZN(n15179) );
  OAI211_X1 U18660 ( .C1(n15181), .C2(n17344), .A(n15180), .B(n15179), .ZN(
        P1_U2888) );
  OAI222_X1 U18661 ( .A1(n17190), .A2(n15195), .B1(n17225), .B2(n15183), .C1(
        n17230), .C2(n15182), .ZN(P1_U2889) );
  OAI222_X1 U18662 ( .A1(n15185), .A2(n15195), .B1(n20753), .B2(n17225), .C1(
        n15184), .C2(n17230), .ZN(P1_U2891) );
  OAI222_X1 U18663 ( .A1(n15332), .A2(n15195), .B1(n20750), .B2(n17225), .C1(
        n15186), .C2(n17230), .ZN(P1_U2892) );
  INV_X1 U18664 ( .A(n17220), .ZN(n15189) );
  INV_X1 U18665 ( .A(n20748), .ZN(n15188) );
  OAI222_X1 U18666 ( .A1(n15189), .A2(n15195), .B1(n15188), .B2(n17225), .C1(
        n15187), .C2(n17230), .ZN(P1_U2893) );
  OAI222_X1 U18667 ( .A1(n15191), .A2(n15195), .B1(n20745), .B2(n17225), .C1(
        n15190), .C2(n17230), .ZN(P1_U2894) );
  OAI222_X1 U18668 ( .A1(n20654), .A2(n15195), .B1(n20742), .B2(n17225), .C1(
        n15192), .C2(n17230), .ZN(P1_U2895) );
  OAI222_X1 U18669 ( .A1(n15365), .A2(n15195), .B1(n15193), .B2(n17225), .C1(
        n20728), .C2(n17230), .ZN(P1_U2896) );
  OAI222_X1 U18670 ( .A1(n15194), .A2(n15195), .B1(n20857), .B2(n17225), .C1(
        n17230), .C2(n11031), .ZN(P1_U2897) );
  INV_X1 U18671 ( .A(n17241), .ZN(n20678) );
  OAI222_X1 U18672 ( .A1(n15195), .A2(n20678), .B1(n17230), .B2(n11039), .C1(
        n17225), .C2(n20844), .ZN(P1_U2898) );
  AOI21_X1 U18673 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15196), .ZN(n15197) );
  OAI21_X1 U18674 ( .B1(n15198), .B2(n20784), .A(n15197), .ZN(n15199) );
  AOI21_X1 U18675 ( .B1(n15200), .B2(n20779), .A(n15199), .ZN(n15201) );
  OAI21_X1 U18676 ( .B1(n15202), .B2(n20631), .A(n15201), .ZN(P1_U2971) );
  NOR2_X1 U18677 ( .A1(n15360), .A2(n21467), .ZN(n15380) );
  AOI21_X1 U18678 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15380), .ZN(n15205) );
  OAI21_X1 U18679 ( .B1(n15206), .B2(n20784), .A(n15205), .ZN(n15207) );
  AOI21_X1 U18680 ( .B1(n15208), .B2(n20779), .A(n15207), .ZN(n15209) );
  OAI21_X1 U18681 ( .B1(n15388), .B2(n20631), .A(n15209), .ZN(P1_U2972) );
  XNOR2_X1 U18682 ( .A(n15212), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15398) );
  NOR2_X1 U18683 ( .A1(n15360), .A2(n21465), .ZN(n15394) );
  AOI21_X1 U18684 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15394), .ZN(n15213) );
  OAI21_X1 U18685 ( .B1(n15214), .B2(n20784), .A(n15213), .ZN(n15215) );
  AOI21_X1 U18686 ( .B1(n15216), .B2(n20779), .A(n15215), .ZN(n15217) );
  OAI21_X1 U18687 ( .B1(n15398), .B2(n20631), .A(n15217), .ZN(P1_U2973) );
  INV_X1 U18688 ( .A(n15218), .ZN(n15219) );
  NAND2_X1 U18689 ( .A1(n15399), .A2(n20780), .ZN(n15225) );
  NOR2_X1 U18690 ( .A1(n15360), .A2(n21462), .ZN(n15402) );
  NOR2_X1 U18691 ( .A1(n15271), .A2(n9909), .ZN(n15222) );
  AOI211_X1 U18692 ( .C1(n15223), .C2(n15274), .A(n15402), .B(n15222), .ZN(
        n15224) );
  NAND2_X1 U18693 ( .A1(n15353), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15227) );
  AOI22_X1 U18694 ( .A1(n15237), .A2(n15227), .B1(n15333), .B2(n15416), .ZN(
        n15229) );
  XNOR2_X1 U18695 ( .A(n15353), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15228) );
  XNOR2_X1 U18696 ( .A(n15229), .B(n15228), .ZN(n15407) );
  NOR2_X1 U18697 ( .A1(n15360), .A2(n21461), .ZN(n15411) );
  AOI21_X1 U18698 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15411), .ZN(n15232) );
  NAND2_X1 U18699 ( .A1(n15230), .A2(n15274), .ZN(n15231) );
  OAI211_X1 U18700 ( .C1(n15233), .C2(n17244), .A(n15232), .B(n15231), .ZN(
        n15234) );
  AOI21_X1 U18701 ( .B1(n15407), .B2(n20780), .A(n15234), .ZN(n15235) );
  INV_X1 U18702 ( .A(n15235), .ZN(P1_U2975) );
  XNOR2_X1 U18703 ( .A(n15353), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15236) );
  XNOR2_X1 U18704 ( .A(n15237), .B(n15236), .ZN(n15424) );
  NAND2_X1 U18705 ( .A1(n15238), .A2(n15274), .ZN(n15239) );
  NAND2_X1 U18706 ( .A1(n20786), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15418) );
  OAI211_X1 U18707 ( .C1(n15271), .C2(n9908), .A(n15239), .B(n15418), .ZN(
        n15240) );
  AOI21_X1 U18708 ( .B1(n15241), .B2(n20779), .A(n15240), .ZN(n15242) );
  OAI21_X1 U18709 ( .B1(n15424), .B2(n20631), .A(n15242), .ZN(P1_U2976) );
  NOR2_X1 U18710 ( .A1(n15243), .A2(n15244), .ZN(n15245) );
  XNOR2_X1 U18711 ( .A(n15245), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15441) );
  INV_X1 U18712 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21458) );
  NOR2_X1 U18713 ( .A1(n15360), .A2(n21458), .ZN(n15437) );
  AOI21_X1 U18714 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15437), .ZN(n15246) );
  OAI21_X1 U18715 ( .B1(n15247), .B2(n20784), .A(n15246), .ZN(n15248) );
  AOI21_X1 U18716 ( .B1(n15249), .B2(n20779), .A(n15248), .ZN(n15250) );
  OAI21_X1 U18717 ( .B1(n20631), .B2(n15441), .A(n15250), .ZN(P1_U2977) );
  NOR3_X1 U18718 ( .A1(n15251), .A2(n15353), .A3(n15451), .ZN(n15260) );
  NOR2_X1 U18719 ( .A1(n15252), .A2(n15333), .ZN(n15259) );
  AOI22_X1 U18720 ( .A1(n15260), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15259), .B2(n10899), .ZN(n15253) );
  XNOR2_X1 U18721 ( .A(n15253), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15442) );
  NAND2_X1 U18722 ( .A1(n15442), .A2(n20780), .ZN(n15257) );
  NOR2_X1 U18723 ( .A1(n15360), .A2(n21456), .ZN(n15445) );
  NOR2_X1 U18724 ( .A1(n15271), .A2(n9912), .ZN(n15254) );
  AOI211_X1 U18725 ( .C1(n15274), .C2(n15255), .A(n15445), .B(n15254), .ZN(
        n15256) );
  OAI211_X1 U18726 ( .C1(n17244), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        P1_U2978) );
  NOR2_X1 U18727 ( .A1(n15260), .A2(n15259), .ZN(n15261) );
  XNOR2_X1 U18728 ( .A(n15261), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15450) );
  NAND2_X1 U18729 ( .A1(n15450), .A2(n20780), .ZN(n15265) );
  NOR2_X1 U18730 ( .A1(n15360), .A2(n21454), .ZN(n15456) );
  NOR2_X1 U18731 ( .A1(n20784), .A2(n15262), .ZN(n15263) );
  AOI211_X1 U18732 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15456), .B(n15263), .ZN(n15264) );
  OAI211_X1 U18733 ( .C1(n17244), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        P1_U2979) );
  NOR2_X1 U18734 ( .A1(n15333), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15267) );
  MUX2_X1 U18735 ( .A(n15333), .B(n15267), .S(n15251), .Z(n15268) );
  XNOR2_X1 U18736 ( .A(n15268), .B(n15451), .ZN(n15462) );
  NAND2_X1 U18737 ( .A1(n15462), .A2(n20780), .ZN(n15276) );
  NOR2_X1 U18738 ( .A1(n15360), .A2(n15269), .ZN(n15466) );
  INV_X1 U18739 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15270) );
  NOR2_X1 U18740 ( .A1(n15271), .A2(n15270), .ZN(n15272) );
  AOI211_X1 U18741 ( .C1(n15274), .C2(n15273), .A(n15466), .B(n15272), .ZN(
        n15275) );
  OAI211_X1 U18742 ( .C1(n17244), .C2(n15277), .A(n15276), .B(n15275), .ZN(
        P1_U2980) );
  NOR2_X1 U18743 ( .A1(n15360), .A2(n21451), .ZN(n15480) );
  NOR2_X1 U18744 ( .A1(n20784), .A2(n15278), .ZN(n15279) );
  AOI211_X1 U18745 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15480), .B(n15279), .ZN(n15283) );
  OR2_X1 U18746 ( .A1(n15281), .A2(n15280), .ZN(n15474) );
  NAND3_X1 U18747 ( .A1(n15474), .A2(n15251), .A3(n20780), .ZN(n15282) );
  OAI211_X1 U18748 ( .C1(n15284), .C2(n17244), .A(n15283), .B(n15282), .ZN(
        P1_U2981) );
  OAI21_X1 U18749 ( .B1(n15296), .B2(n15287), .A(n15297), .ZN(n15288) );
  XOR2_X1 U18750 ( .A(n15289), .B(n15288), .Z(n15502) );
  NOR2_X1 U18751 ( .A1(n15360), .A2(n15290), .ZN(n15496) );
  AOI21_X1 U18752 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15496), .ZN(n15291) );
  OAI21_X1 U18753 ( .B1(n20784), .B2(n15292), .A(n15291), .ZN(n15293) );
  AOI21_X1 U18754 ( .B1(n15294), .B2(n20779), .A(n15293), .ZN(n15295) );
  OAI21_X1 U18755 ( .B1(n15502), .B2(n20631), .A(n15295), .ZN(P1_U2983) );
  NAND2_X1 U18756 ( .A1(n15503), .A2(n20780), .ZN(n15301) );
  NOR2_X1 U18757 ( .A1(n15360), .A2(n21447), .ZN(n15504) );
  NOR2_X1 U18758 ( .A1(n20784), .A2(n17197), .ZN(n15299) );
  AOI211_X1 U18759 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15504), .B(n15299), .ZN(n15300) );
  OAI211_X1 U18760 ( .C1(n17244), .C2(n17190), .A(n15301), .B(n15300), .ZN(
        P1_U2984) );
  INV_X1 U18761 ( .A(n15302), .ZN(n15303) );
  AOI21_X1 U18762 ( .B1(n15305), .B2(n15304), .A(n15303), .ZN(n15307) );
  XNOR2_X1 U18763 ( .A(n15353), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15306) );
  XNOR2_X1 U18764 ( .A(n15307), .B(n15306), .ZN(n15516) );
  AND2_X1 U18765 ( .A1(n20786), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n15511) );
  AOI21_X1 U18766 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n15511), .ZN(n15308) );
  OAI21_X1 U18767 ( .B1(n20784), .B2(n17207), .A(n15308), .ZN(n15309) );
  AOI21_X1 U18768 ( .B1(n17228), .B2(n20779), .A(n15309), .ZN(n15310) );
  OAI21_X1 U18769 ( .B1(n15516), .B2(n20631), .A(n15310), .ZN(P1_U2985) );
  INV_X1 U18770 ( .A(n15341), .ZN(n15314) );
  INV_X1 U18771 ( .A(n15311), .ZN(n15312) );
  AOI21_X1 U18772 ( .B1(n15314), .B2(n15313), .A(n15312), .ZN(n15326) );
  AND2_X1 U18773 ( .A1(n15315), .A2(n15316), .ZN(n15325) );
  NAND2_X1 U18774 ( .A1(n15326), .A2(n15325), .ZN(n15324) );
  NAND2_X1 U18775 ( .A1(n15324), .A2(n15316), .ZN(n15317) );
  XNOR2_X1 U18776 ( .A(n15318), .B(n15317), .ZN(n15525) );
  INV_X1 U18777 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21444) );
  OR2_X1 U18778 ( .A1(n15360), .A2(n21444), .ZN(n15520) );
  NAND2_X1 U18779 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15319) );
  OAI211_X1 U18780 ( .C1(n20784), .C2(n15320), .A(n15520), .B(n15319), .ZN(
        n15321) );
  AOI21_X1 U18781 ( .B1(n15322), .B2(n20779), .A(n15321), .ZN(n15323) );
  OAI21_X1 U18782 ( .B1(n15525), .B2(n20631), .A(n15323), .ZN(P1_U2986) );
  OAI21_X1 U18783 ( .B1(n15326), .B2(n15325), .A(n15324), .ZN(n15526) );
  NAND2_X1 U18784 ( .A1(n15526), .A2(n20780), .ZN(n15331) );
  INV_X1 U18785 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15327) );
  NOR2_X1 U18786 ( .A1(n15360), .A2(n15327), .ZN(n15527) );
  NOR2_X1 U18787 ( .A1(n20784), .A2(n15328), .ZN(n15329) );
  AOI211_X1 U18788 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n15527), .B(n15329), .ZN(n15330) );
  OAI211_X1 U18789 ( .C1(n17244), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        P1_U2987) );
  NOR3_X1 U18790 ( .A1(n15341), .A2(n15353), .A3(n15564), .ZN(n15334) );
  NOR3_X1 U18791 ( .A1(n15340), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n15333), .ZN(n15345) );
  NOR2_X1 U18792 ( .A1(n15334), .A2(n15345), .ZN(n15335) );
  XNOR2_X1 U18793 ( .A(n15335), .B(n15548), .ZN(n15552) );
  INV_X1 U18794 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15336) );
  NOR2_X1 U18795 ( .A1(n15360), .A2(n15336), .ZN(n15546) );
  AOI21_X1 U18796 ( .B1(n20773), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15546), .ZN(n15337) );
  OAI21_X1 U18797 ( .B1(n20784), .B2(n17223), .A(n15337), .ZN(n15338) );
  AOI21_X1 U18798 ( .B1(n17220), .B2(n20779), .A(n15338), .ZN(n15339) );
  OAI21_X1 U18799 ( .B1(n15552), .B2(n20631), .A(n15339), .ZN(P1_U2988) );
  AND2_X1 U18800 ( .A1(n15340), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15344) );
  XNOR2_X1 U18801 ( .A(n15341), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15343) );
  MUX2_X1 U18802 ( .A(n15344), .B(n15343), .S(n15342), .Z(n15346) );
  NOR2_X1 U18803 ( .A1(n15346), .A2(n15345), .ZN(n15569) );
  INV_X1 U18804 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15347) );
  OR2_X1 U18805 ( .A1(n15360), .A2(n15347), .ZN(n15560) );
  NAND2_X1 U18806 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15348) );
  OAI211_X1 U18807 ( .C1(n20784), .C2(n15349), .A(n15560), .B(n15348), .ZN(
        n15350) );
  AOI21_X1 U18808 ( .B1(n15351), .B2(n20779), .A(n15350), .ZN(n15352) );
  OAI21_X1 U18809 ( .B1(n15569), .B2(n20631), .A(n15352), .ZN(P1_U2989) );
  INV_X1 U18810 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15565) );
  NAND2_X1 U18811 ( .A1(n15570), .A2(n20780), .ZN(n15356) );
  NOR2_X1 U18812 ( .A1(n15360), .A2(n21439), .ZN(n15573) );
  NOR2_X1 U18813 ( .A1(n20784), .A2(n20655), .ZN(n15354) );
  AOI211_X1 U18814 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15573), .B(n15354), .ZN(n15355) );
  OAI211_X1 U18815 ( .C1(n17244), .C2(n20654), .A(n15356), .B(n15355), .ZN(
        P1_U2990) );
  XNOR2_X1 U18816 ( .A(n15357), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15358) );
  XNOR2_X1 U18817 ( .A(n15359), .B(n15358), .ZN(n17256) );
  NAND2_X1 U18818 ( .A1(n17256), .A2(n20780), .ZN(n15364) );
  NOR2_X1 U18819 ( .A1(n15360), .A2(n21436), .ZN(n17253) );
  NOR2_X1 U18820 ( .A1(n20784), .A2(n15361), .ZN(n15362) );
  AOI211_X1 U18821 ( .C1(n20773), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n17253), .B(n15362), .ZN(n15363) );
  OAI211_X1 U18822 ( .C1(n17244), .C2(n15365), .A(n15364), .B(n15363), .ZN(
        P1_U2991) );
  INV_X1 U18823 ( .A(n15366), .ZN(n15378) );
  NAND2_X1 U18824 ( .A1(n15367), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15373) );
  NAND3_X1 U18825 ( .A1(n15369), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15368), .ZN(n15372) );
  INV_X1 U18826 ( .A(n15370), .ZN(n15371) );
  OAI211_X1 U18827 ( .C1(n15374), .C2(n15373), .A(n15372), .B(n15371), .ZN(
        n15375) );
  AOI21_X1 U18828 ( .B1(n15376), .B2(n20801), .A(n15375), .ZN(n15377) );
  OAI21_X1 U18829 ( .B1(n15378), .B2(n20807), .A(n15377), .ZN(P1_U3000) );
  INV_X1 U18830 ( .A(n15379), .ZN(n15384) );
  AOI21_X1 U18831 ( .B1(n15381), .B2(n15383), .A(n15380), .ZN(n15382) );
  OAI21_X1 U18832 ( .B1(n15384), .B2(n15383), .A(n15382), .ZN(n15385) );
  AOI21_X1 U18833 ( .B1(n15386), .B2(n20801), .A(n15385), .ZN(n15387) );
  INV_X1 U18834 ( .A(n15389), .ZN(n15403) );
  INV_X1 U18835 ( .A(n15390), .ZN(n15392) );
  NOR3_X1 U18836 ( .A1(n15400), .A2(n15392), .A3(n15391), .ZN(n15393) );
  AOI211_X1 U18837 ( .C1(n15403), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15394), .B(n15393), .ZN(n15397) );
  NAND2_X1 U18838 ( .A1(n15395), .A2(n20801), .ZN(n15396) );
  OAI211_X1 U18839 ( .C1(n15398), .C2(n20807), .A(n15397), .B(n15396), .ZN(
        P1_U3005) );
  NAND2_X1 U18840 ( .A1(n15399), .A2(n20795), .ZN(n15405) );
  NOR2_X1 U18841 ( .A1(n15400), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15401) );
  AOI211_X1 U18842 ( .C1(n15403), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15402), .B(n15401), .ZN(n15404) );
  NAND2_X1 U18843 ( .A1(n15407), .A2(n20795), .ZN(n15414) );
  OAI21_X1 U18844 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15409), .A(
        n15408), .ZN(n15412) );
  NOR3_X1 U18845 ( .A1(n15419), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15416), .ZN(n15410) );
  AOI211_X1 U18846 ( .C1(n15412), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15411), .B(n15410), .ZN(n15413) );
  OAI211_X1 U18847 ( .C1(n15571), .C2(n15415), .A(n15414), .B(n15413), .ZN(
        P1_U3007) );
  NOR2_X1 U18848 ( .A1(n15417), .A2(n15416), .ZN(n15421) );
  OAI21_X1 U18849 ( .B1(n15419), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15418), .ZN(n15420) );
  AOI211_X1 U18850 ( .C1(n15422), .C2(n20801), .A(n15421), .B(n15420), .ZN(
        n15423) );
  OAI21_X1 U18851 ( .B1(n15424), .B2(n20807), .A(n15423), .ZN(P1_U3008) );
  NOR2_X1 U18852 ( .A1(n15452), .A2(n15464), .ZN(n15518) );
  INV_X1 U18853 ( .A(n15518), .ZN(n15432) );
  NAND2_X1 U18854 ( .A1(n20805), .A2(n15425), .ZN(n15430) );
  NOR2_X1 U18855 ( .A1(n15464), .A2(n15426), .ZN(n15427) );
  NAND2_X1 U18856 ( .A1(n15428), .A2(n15427), .ZN(n15429) );
  NAND2_X1 U18857 ( .A1(n15430), .A2(n15429), .ZN(n15517) );
  INV_X1 U18858 ( .A(n15465), .ZN(n15431) );
  NAND2_X1 U18859 ( .A1(n15517), .A2(n15431), .ZN(n15463) );
  OAI21_X1 U18860 ( .B1(n15432), .B2(n15465), .A(n15463), .ZN(n15457) );
  INV_X1 U18861 ( .A(n15433), .ZN(n15434) );
  NAND2_X1 U18862 ( .A1(n15457), .A2(n15434), .ZN(n15443) );
  XNOR2_X1 U18863 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15435) );
  NOR2_X1 U18864 ( .A1(n15443), .A2(n15435), .ZN(n15436) );
  AOI211_X1 U18865 ( .C1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n15446), .A(
        n15437), .B(n15436), .ZN(n15440) );
  NAND2_X1 U18866 ( .A1(n15438), .A2(n20801), .ZN(n15439) );
  OAI211_X1 U18867 ( .C1(n15441), .C2(n20807), .A(n15440), .B(n15439), .ZN(
        P1_U3009) );
  NAND2_X1 U18868 ( .A1(n15442), .A2(n20795), .ZN(n15448) );
  NOR2_X1 U18869 ( .A1(n15443), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15444) );
  AOI211_X1 U18870 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15446), .A(
        n15445), .B(n15444), .ZN(n15447) );
  OAI211_X1 U18871 ( .C1(n15571), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        P1_U3010) );
  NAND2_X1 U18872 ( .A1(n15450), .A2(n20795), .ZN(n15460) );
  NOR2_X1 U18873 ( .A1(n15451), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15458) );
  AOI21_X1 U18874 ( .B1(n15463), .B2(n15452), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15468) );
  INV_X1 U18875 ( .A(n15468), .ZN(n15453) );
  AOI21_X1 U18876 ( .B1(n15454), .B2(n15453), .A(n10899), .ZN(n15455) );
  AOI211_X1 U18877 ( .C1(n15458), .C2(n15457), .A(n15456), .B(n15455), .ZN(
        n15459) );
  OAI211_X1 U18878 ( .C1(n15571), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        P1_U3011) );
  NAND2_X1 U18879 ( .A1(n15462), .A2(n20795), .ZN(n15473) );
  OAI21_X1 U18880 ( .B1(n15465), .B2(n15464), .A(n15463), .ZN(n15467) );
  AOI21_X1 U18881 ( .B1(n15468), .B2(n15467), .A(n15466), .ZN(n15472) );
  NAND2_X1 U18882 ( .A1(n15469), .A2(n20801), .ZN(n15471) );
  NAND4_X1 U18883 ( .A1(n15473), .A2(n15472), .A3(n15471), .A4(n15470), .ZN(
        P1_U3012) );
  NAND3_X1 U18884 ( .A1(n15251), .A2(n15474), .A3(n20795), .ZN(n15483) );
  NAND2_X1 U18885 ( .A1(n15513), .A2(n15475), .ZN(n15476) );
  OAI211_X1 U18886 ( .C1(n17255), .C2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15521), .B(n15476), .ZN(n15512) );
  AOI21_X1 U18887 ( .B1(n15580), .B2(n15477), .A(n15512), .ZN(n15485) );
  INV_X1 U18888 ( .A(n15485), .ZN(n15481) );
  AND2_X1 U18889 ( .A1(n15513), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15498) );
  INV_X1 U18890 ( .A(n15498), .ZN(n15478) );
  NOR3_X1 U18891 ( .A1(n15478), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15477), .ZN(n15479) );
  AOI211_X1 U18892 ( .C1(n15481), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15480), .B(n15479), .ZN(n15482) );
  OAI211_X1 U18893 ( .C1(n15571), .C2(n15484), .A(n15483), .B(n15482), .ZN(
        P1_U3013) );
  NAND3_X1 U18894 ( .A1(n15498), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15486) );
  AOI21_X1 U18895 ( .B1(n11597), .B2(n15486), .A(n15485), .ZN(n15487) );
  AOI211_X1 U18896 ( .C1(n15489), .C2(n20801), .A(n15488), .B(n15487), .ZN(
        n15490) );
  OAI21_X1 U18897 ( .B1(n15491), .B2(n20807), .A(n15490), .ZN(P1_U3014) );
  NOR2_X1 U18898 ( .A1(n15492), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15497) );
  INV_X1 U18899 ( .A(n15512), .ZN(n15494) );
  NAND2_X1 U18900 ( .A1(n15498), .A2(n15492), .ZN(n15506) );
  AOI21_X1 U18901 ( .B1(n15494), .B2(n15506), .A(n15493), .ZN(n15495) );
  AOI211_X1 U18902 ( .C1(n15498), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15501) );
  NAND2_X1 U18903 ( .A1(n15499), .A2(n20801), .ZN(n15500) );
  OAI211_X1 U18904 ( .C1(n15502), .C2(n20807), .A(n15501), .B(n15500), .ZN(
        P1_U3015) );
  INV_X1 U18905 ( .A(n15503), .ZN(n15510) );
  NAND2_X1 U18906 ( .A1(n15512), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15507) );
  INV_X1 U18907 ( .A(n15504), .ZN(n15505) );
  NAND3_X1 U18908 ( .A1(n15507), .A2(n15506), .A3(n15505), .ZN(n15508) );
  AOI21_X1 U18909 ( .B1(n20801), .B2(n17195), .A(n15508), .ZN(n15509) );
  OAI21_X1 U18910 ( .B1(n15510), .B2(n20807), .A(n15509), .ZN(P1_U3016) );
  AOI21_X1 U18911 ( .B1(n17206), .B2(n20801), .A(n15511), .ZN(n15515) );
  OAI21_X1 U18912 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15513), .A(
        n15512), .ZN(n15514) );
  OAI211_X1 U18913 ( .C1(n15516), .C2(n20807), .A(n15515), .B(n15514), .ZN(
        P1_U3017) );
  OAI21_X1 U18914 ( .B1(n15518), .B2(n15517), .A(n10879), .ZN(n15519) );
  OAI211_X1 U18915 ( .C1(n15521), .C2(n10879), .A(n15520), .B(n15519), .ZN(
        n15522) );
  AOI21_X1 U18916 ( .B1(n20801), .B2(n15523), .A(n15522), .ZN(n15524) );
  OAI21_X1 U18917 ( .B1(n15525), .B2(n20807), .A(n15524), .ZN(P1_U3018) );
  NAND2_X1 U18918 ( .A1(n15526), .A2(n20795), .ZN(n15544) );
  AOI21_X1 U18919 ( .B1(n15528), .B2(n20801), .A(n15527), .ZN(n15543) );
  INV_X1 U18920 ( .A(n15530), .ZN(n15549) );
  NAND4_X1 U18921 ( .A1(n17266), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        n15549), .A4(n15531), .ZN(n15542) );
  INV_X1 U18922 ( .A(n15532), .ZN(n15538) );
  INV_X1 U18923 ( .A(n15533), .ZN(n15558) );
  INV_X1 U18924 ( .A(n15534), .ZN(n15535) );
  NAND2_X1 U18925 ( .A1(n20811), .A2(n15535), .ZN(n15536) );
  OAI211_X1 U18926 ( .C1(n15538), .C2(n15537), .A(n15558), .B(n15536), .ZN(
        n15547) );
  AND2_X1 U18927 ( .A1(n15539), .A2(n15548), .ZN(n15540) );
  OAI21_X1 U18928 ( .B1(n15547), .B2(n15540), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15541) );
  NAND4_X1 U18929 ( .A1(n15544), .A2(n15543), .A3(n15542), .A4(n15541), .ZN(
        P1_U3019) );
  NOR2_X1 U18930 ( .A1(n17213), .A2(n15571), .ZN(n15545) );
  AOI211_X1 U18931 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15547), .A(
        n15546), .B(n15545), .ZN(n15551) );
  NAND3_X1 U18932 ( .A1(n17266), .A2(n15549), .A3(n15548), .ZN(n15550) );
  OAI211_X1 U18933 ( .C1(n15552), .C2(n20807), .A(n15551), .B(n15550), .ZN(
        P1_U3020) );
  AOI21_X1 U18934 ( .B1(n15555), .B2(n15554), .A(n15553), .ZN(n15557) );
  INV_X1 U18935 ( .A(n15562), .ZN(n15556) );
  OAI21_X1 U18936 ( .B1(n15557), .B2(n15556), .A(n15580), .ZN(n15559) );
  NAND2_X1 U18937 ( .A1(n15559), .A2(n15558), .ZN(n15574) );
  OAI21_X1 U18938 ( .B1(n15561), .B2(n15571), .A(n15560), .ZN(n15567) );
  NAND2_X1 U18939 ( .A1(n17266), .A2(n15562), .ZN(n15577) );
  AOI211_X1 U18940 ( .C1(n15565), .C2(n15564), .A(n15563), .B(n15577), .ZN(
        n15566) );
  AOI211_X1 U18941 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15574), .A(
        n15567), .B(n15566), .ZN(n15568) );
  OAI21_X1 U18942 ( .B1(n15569), .B2(n20807), .A(n15568), .ZN(P1_U3021) );
  NAND2_X1 U18943 ( .A1(n15570), .A2(n20795), .ZN(n15576) );
  NOR2_X1 U18944 ( .A1(n15571), .A2(n20649), .ZN(n15572) );
  AOI211_X1 U18945 ( .C1(n15574), .C2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15573), .B(n15572), .ZN(n15575) );
  OAI211_X1 U18946 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15577), .A(
        n15576), .B(n15575), .ZN(P1_U3022) );
  NAND3_X1 U18947 ( .A1(n15579), .A2(n15578), .A3(n20795), .ZN(n15587) );
  NAND2_X1 U18948 ( .A1(n15580), .A2(n20810), .ZN(n15582) );
  MUX2_X1 U18949 ( .A(n15582), .B(n15581), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n15585) );
  NAND2_X1 U18950 ( .A1(n20801), .A2(n15583), .ZN(n15584) );
  NAND4_X1 U18951 ( .A1(n15587), .A2(n15586), .A3(n15585), .A4(n15584), .ZN(
        P1_U3030) );
  OAI21_X1 U18952 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14417), .A(n20929), 
        .ZN(n15588) );
  OAI21_X1 U18953 ( .B1(n15589), .B2(n14504), .A(n15588), .ZN(n15590) );
  MUX2_X1 U18954 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15590), .S(
        n20817), .Z(P1_U3477) );
  INV_X1 U18955 ( .A(n15591), .ZN(n15592) );
  OR2_X1 U18956 ( .A1(n14504), .A2(n15592), .ZN(n15598) );
  NOR2_X1 U18957 ( .A1(n14409), .A2(n15593), .ZN(n15602) );
  AOI22_X1 U18958 ( .A1(n17140), .A2(n15596), .B1(n15602), .B2(n15595), .ZN(
        n15597) );
  NAND2_X1 U18959 ( .A1(n15598), .A2(n15597), .ZN(n17144) );
  INV_X1 U18960 ( .A(n17144), .ZN(n15604) );
  INV_X1 U18961 ( .A(n20624), .ZN(n17272) );
  INV_X1 U18962 ( .A(n15599), .ZN(n15600) );
  AOI22_X1 U18963 ( .A1(n17173), .A2(n15602), .B1(n15601), .B2(n15600), .ZN(
        n15603) );
  OAI21_X1 U18964 ( .B1(n15604), .B2(n17272), .A(n15603), .ZN(n15605) );
  MUX2_X1 U18965 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15605), .S(
        n17276), .Z(P1_U3473) );
  AOI21_X1 U18966 ( .B1(n20495), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n15606), 
        .ZN(n15609) );
  NOR3_X1 U18967 ( .A1(n20495), .A2(n15607), .A3(n16837), .ZN(n15608) );
  MUX2_X1 U18968 ( .A(n15609), .B(n15608), .S(n15871), .Z(n15611) );
  AOI22_X1 U18969 ( .A1(n20480), .A2(P2_STATE2_REG_2__SCAN_IN), .B1(n16835), 
        .B2(n16837), .ZN(n15610) );
  OR2_X1 U18970 ( .A1(n15611), .A2(n15610), .ZN(n15615) );
  INV_X2 U18971 ( .A(n19841), .ZN(n19902) );
  OAI21_X1 U18972 ( .B1(n15612), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n20575), 
        .ZN(n15613) );
  AOI211_X1 U18973 ( .C1(n20480), .C2(n19902), .A(n15613), .B(n19594), .ZN(
        n15614) );
  MUX2_X1 U18974 ( .A(n15615), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n15614), 
        .Z(P2_U3610) );
  OAI21_X1 U18975 ( .B1(n15617), .B2(n20488), .A(n19716), .ZN(n15621) );
  INV_X1 U18976 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16105) );
  NAND3_X1 U18977 ( .A1(n15617), .A2(n15855), .A3(n16104), .ZN(n15619) );
  AOI22_X1 U18978 ( .A1(n19613), .A2(P2_REIP_REG_29__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_29__SCAN_IN), .ZN(n15618) );
  OAI211_X1 U18979 ( .C1(n19775), .C2(n16105), .A(n15619), .B(n15618), .ZN(
        n15620) );
  NOR2_X1 U18980 ( .A1(n14531), .A2(n15623), .ZN(n15624) );
  XNOR2_X1 U18981 ( .A(n15626), .B(n16120), .ZN(n15629) );
  AOI22_X1 U18982 ( .A1(n19613), .A2(P2_REIP_REG_28__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_28__SCAN_IN), .ZN(n15628) );
  NAND2_X1 U18983 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15627) );
  OAI211_X1 U18984 ( .C1(n15629), .C2(n20488), .A(n15628), .B(n15627), .ZN(
        n15635) );
  NAND2_X1 U18985 ( .A1(n15631), .A2(n15630), .ZN(n15632) );
  NAND2_X1 U18986 ( .A1(n15633), .A2(n15632), .ZN(n16380) );
  NOR2_X1 U18987 ( .A1(n16380), .A2(n19786), .ZN(n15634) );
  AOI211_X1 U18988 ( .C1(n19736), .C2(n15636), .A(n15635), .B(n15634), .ZN(
        n15637) );
  OAI21_X1 U18989 ( .B1(n16374), .B2(n19767), .A(n15637), .ZN(P2_U2827) );
  NAND2_X1 U18990 ( .A1(n15638), .A2(n19771), .ZN(n15639) );
  AOI21_X1 U18991 ( .B1(n15639), .B2(n19716), .A(n16133), .ZN(n15645) );
  INV_X1 U18992 ( .A(n15638), .ZN(n15640) );
  NAND3_X1 U18993 ( .A1(n15640), .A2(n15855), .A3(n16133), .ZN(n15642) );
  AOI22_X1 U18994 ( .A1(n19613), .A2(P2_REIP_REG_27__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_27__SCAN_IN), .ZN(n15641) );
  OAI211_X1 U18995 ( .C1(n19775), .C2(n15643), .A(n15642), .B(n15641), .ZN(
        n15644) );
  AOI211_X1 U18996 ( .C1(n9607), .C2(n19736), .A(n15645), .B(n15644), .ZN(
        n15647) );
  NAND2_X1 U18997 ( .A1(n16389), .A2(n19785), .ZN(n15646) );
  OAI211_X1 U18998 ( .C1(n16392), .C2(n19786), .A(n15647), .B(n15646), .ZN(
        P2_U2828) );
  INV_X1 U18999 ( .A(n15648), .ZN(n15650) );
  INV_X1 U19000 ( .A(n15649), .ZN(n15664) );
  AOI21_X1 U19001 ( .B1(n15650), .B2(n15664), .A(n14539), .ZN(n16146) );
  INV_X1 U19002 ( .A(n16146), .ZN(n16405) );
  XOR2_X1 U19003 ( .A(n16144), .B(n15651), .Z(n15657) );
  INV_X1 U19004 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15653) );
  AOI22_X1 U19005 ( .A1(n19613), .A2(P2_REIP_REG_26__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n15652) );
  OAI21_X1 U19006 ( .B1(n19775), .B2(n15653), .A(n15652), .ZN(n15656) );
  NOR2_X1 U19007 ( .A1(n15654), .A2(n19782), .ZN(n15655) );
  AOI211_X1 U19008 ( .C1(n19771), .C2(n15657), .A(n15656), .B(n15655), .ZN(
        n15662) );
  AOI21_X1 U19009 ( .B1(n15660), .B2(n15678), .A(n14530), .ZN(n16407) );
  NAND2_X1 U19010 ( .A1(n16407), .A2(n19785), .ZN(n15661) );
  OAI211_X1 U19011 ( .C1(n16405), .C2(n19786), .A(n15662), .B(n15661), .ZN(
        P2_U2829) );
  INV_X1 U19012 ( .A(n15683), .ZN(n15666) );
  INV_X1 U19013 ( .A(n15663), .ZN(n15665) );
  OAI21_X1 U19014 ( .B1(n15667), .B2(n20488), .A(n19716), .ZN(n15674) );
  INV_X1 U19015 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16151) );
  INV_X1 U19016 ( .A(n16154), .ZN(n15668) );
  NAND3_X1 U19017 ( .A1(n15667), .A2(n15855), .A3(n15668), .ZN(n15670) );
  AOI22_X1 U19018 ( .A1(n19613), .A2(P2_REIP_REG_25__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_25__SCAN_IN), .ZN(n15669) );
  OAI211_X1 U19019 ( .C1(n19775), .C2(n16151), .A(n15670), .B(n15669), .ZN(
        n15673) );
  NOR2_X1 U19020 ( .A1(n15671), .A2(n19782), .ZN(n15672) );
  AOI211_X1 U19021 ( .C1(n16154), .C2(n15674), .A(n15673), .B(n15672), .ZN(
        n15680) );
  OR2_X1 U19022 ( .A1(n15675), .A2(n15676), .ZN(n15677) );
  AND2_X1 U19023 ( .A1(n15678), .A2(n15677), .ZN(n16416) );
  NAND2_X1 U19024 ( .A1(n16416), .A2(n19785), .ZN(n15679) );
  OAI211_X1 U19025 ( .C1(n16414), .C2(n19786), .A(n15680), .B(n15679), .ZN(
        P2_U2830) );
  NAND2_X1 U19026 ( .A1(n9621), .A2(n15681), .ZN(n15682) );
  NAND2_X1 U19027 ( .A1(n15683), .A2(n15682), .ZN(n16424) );
  AOI21_X1 U19028 ( .B1(n15685), .B2(n15684), .A(n15675), .ZN(n16426) );
  NAND2_X1 U19029 ( .A1(n16426), .A2(n19785), .ZN(n15694) );
  INV_X1 U19030 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15690) );
  XOR2_X1 U19031 ( .A(n16165), .B(n15686), .Z(n15687) );
  NAND2_X1 U19032 ( .A1(n15687), .A2(n19771), .ZN(n15689) );
  AOI22_X1 U19033 ( .A1(n19613), .A2(P2_REIP_REG_24__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_24__SCAN_IN), .ZN(n15688) );
  OAI211_X1 U19034 ( .C1(n15690), .C2(n19775), .A(n15689), .B(n15688), .ZN(
        n15691) );
  AOI21_X1 U19035 ( .B1(n15692), .B2(n19736), .A(n15691), .ZN(n15693) );
  OAI211_X1 U19036 ( .C1(n19786), .C2(n16424), .A(n15694), .B(n15693), .ZN(
        P2_U2831) );
  OR2_X1 U19037 ( .A1(n15695), .A2(n15696), .ZN(n15697) );
  NAND2_X1 U19038 ( .A1(n9621), .A2(n15697), .ZN(n16437) );
  INV_X1 U19039 ( .A(n15684), .ZN(n15699) );
  AOI21_X1 U19040 ( .B1(n15700), .B2(n15698), .A(n15699), .ZN(n16439) );
  NAND2_X1 U19041 ( .A1(n16439), .A2(n19785), .ZN(n15710) );
  OAI21_X1 U19042 ( .B1(n15701), .B2(n20488), .A(n19716), .ZN(n15702) );
  AND2_X1 U19043 ( .A1(n15702), .A2(n16172), .ZN(n15707) );
  INV_X1 U19044 ( .A(n16172), .ZN(n15703) );
  NAND3_X1 U19045 ( .A1(n15701), .A2(n15855), .A3(n15703), .ZN(n15705) );
  AOI22_X1 U19046 ( .A1(n19613), .A2(P2_REIP_REG_23__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_23__SCAN_IN), .ZN(n15704) );
  OAI211_X1 U19047 ( .C1(n19775), .C2(n16169), .A(n15705), .B(n15704), .ZN(
        n15706) );
  AOI211_X1 U19048 ( .C1(n15708), .C2(n19736), .A(n15707), .B(n15706), .ZN(
        n15709) );
  OAI211_X1 U19049 ( .C1(n19786), .C2(n16437), .A(n15710), .B(n15709), .ZN(
        P2_U2832) );
  OR2_X1 U19050 ( .A1(n13665), .A2(n15711), .ZN(n15712) );
  AND2_X1 U19051 ( .A1(n15698), .A2(n15712), .ZN(n16451) );
  INV_X1 U19052 ( .A(n16451), .ZN(n16043) );
  INV_X1 U19053 ( .A(n15713), .ZN(n15716) );
  INV_X1 U19054 ( .A(n15714), .ZN(n15715) );
  AOI21_X1 U19055 ( .B1(n15716), .B2(n15715), .A(n15695), .ZN(n16184) );
  NOR2_X1 U19056 ( .A1(n15717), .A2(n19782), .ZN(n15723) );
  XNOR2_X1 U19057 ( .A(n15718), .B(n16182), .ZN(n15721) );
  AOI22_X1 U19058 ( .A1(n19613), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n15720) );
  NAND2_X1 U19059 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15719) );
  OAI211_X1 U19060 ( .C1(n15721), .C2(n20488), .A(n15720), .B(n15719), .ZN(
        n15722) );
  AOI211_X1 U19061 ( .C1(n16184), .C2(n19754), .A(n15723), .B(n15722), .ZN(
        n15724) );
  OAI21_X1 U19062 ( .B1(n16043), .B2(n19767), .A(n15724), .ZN(P2_U2833) );
  OAI21_X1 U19063 ( .B1(n15725), .B2(n20488), .A(n19716), .ZN(n15732) );
  NAND3_X1 U19064 ( .A1(n15725), .A2(n15855), .A3(n14661), .ZN(n15727) );
  AOI22_X1 U19065 ( .A1(n19613), .A2(P2_REIP_REG_21__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_21__SCAN_IN), .ZN(n15726) );
  OAI211_X1 U19066 ( .C1(n19775), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15731) );
  NOR2_X1 U19067 ( .A1(n15729), .A2(n19782), .ZN(n15730) );
  AOI211_X1 U19068 ( .C1(n15733), .C2(n15732), .A(n15731), .B(n15730), .ZN(
        n15735) );
  NAND2_X1 U19069 ( .A1(n16044), .A2(n19785), .ZN(n15734) );
  OAI211_X1 U19070 ( .C1(n15903), .C2(n19786), .A(n15735), .B(n15734), .ZN(
        P2_U2834) );
  NAND2_X1 U19071 ( .A1(n15737), .A2(n15736), .ZN(n15738) );
  NAND2_X1 U19072 ( .A1(n15739), .A2(n15738), .ZN(n16463) );
  AOI21_X1 U19073 ( .B1(n15741), .B2(n13586), .A(n10415), .ZN(n16461) );
  NOR2_X1 U19074 ( .A1(n15742), .A2(n19782), .ZN(n15748) );
  XNOR2_X1 U19075 ( .A(n15743), .B(n16199), .ZN(n15746) );
  AOI22_X1 U19076 ( .A1(n19613), .A2(P2_REIP_REG_20__SCAN_IN), .B1(n19784), 
        .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n15745) );
  NAND2_X1 U19077 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15744) );
  OAI211_X1 U19078 ( .C1(n15746), .C2(n20488), .A(n15745), .B(n15744), .ZN(
        n15747) );
  AOI211_X1 U19079 ( .C1(n16461), .C2(n19754), .A(n15748), .B(n15747), .ZN(
        n15749) );
  OAI21_X1 U19080 ( .B1(n16463), .B2(n19767), .A(n15749), .ZN(P2_U2835) );
  INV_X1 U19081 ( .A(n15923), .ZN(n16219) );
  NAND2_X1 U19082 ( .A1(n15755), .A2(n19771), .ZN(n15750) );
  AOI21_X1 U19083 ( .B1(n15750), .B2(n19716), .A(n16217), .ZN(n15757) );
  NAND2_X1 U19084 ( .A1(n15855), .A2(n16217), .ZN(n15754) );
  NAND2_X1 U19085 ( .A1(n19784), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n15751) );
  OAI211_X1 U19086 ( .C1(n20535), .C2(n19778), .A(n15751), .B(n19701), .ZN(
        n15752) );
  AOI21_X1 U19087 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19777), .A(
        n15752), .ZN(n15753) );
  OAI21_X1 U19088 ( .B1(n15755), .B2(n15754), .A(n15753), .ZN(n15756) );
  NOR2_X1 U19089 ( .A1(n15757), .A2(n15756), .ZN(n15758) );
  OAI21_X1 U19090 ( .B1(n15759), .B2(n19782), .A(n15758), .ZN(n15760) );
  AOI21_X1 U19091 ( .B1(n16219), .B2(n19754), .A(n15760), .ZN(n15761) );
  OAI21_X1 U19092 ( .B1(n16082), .B2(n19767), .A(n15761), .ZN(P2_U2838) );
  AOI21_X1 U19093 ( .B1(n15764), .B2(n15762), .A(n15763), .ZN(n16259) );
  NAND2_X1 U19094 ( .A1(n19784), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n15766) );
  INV_X1 U19095 ( .A(n19716), .ZN(n15843) );
  AOI21_X1 U19096 ( .B1(n15843), .B2(n16255), .A(n16341), .ZN(n15765) );
  OAI211_X1 U19097 ( .C1(n19778), .C2(n15767), .A(n15766), .B(n15765), .ZN(
        n15771) );
  INV_X1 U19098 ( .A(n15768), .ZN(n15769) );
  NAND2_X1 U19099 ( .A1(n15855), .A2(n19672), .ZN(n19685) );
  AOI21_X1 U19100 ( .B1(n15769), .B2(n16255), .A(n19685), .ZN(n15770) );
  AOI211_X1 U19101 ( .C1(n19777), .C2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15771), .B(n15770), .ZN(n15772) );
  OAI21_X1 U19102 ( .B1(n15773), .B2(n19782), .A(n15772), .ZN(n15774) );
  AOI21_X1 U19103 ( .B1(n16259), .B2(n19754), .A(n15774), .ZN(n15775) );
  OAI21_X1 U19104 ( .B1(n15776), .B2(n19767), .A(n15775), .ZN(P2_U2842) );
  AND2_X1 U19105 ( .A1(n15777), .A2(n15778), .ZN(n15780) );
  OR2_X1 U19106 ( .A1(n15780), .A2(n15779), .ZN(n16566) );
  INV_X1 U19107 ( .A(n16566), .ZN(n15790) );
  NAND2_X1 U19108 ( .A1(n19784), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15781) );
  OAI211_X1 U19109 ( .C1(n20523), .C2(n19778), .A(n15781), .B(n19701), .ZN(
        n15782) );
  AOI21_X1 U19110 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19777), .A(
        n15782), .ZN(n15787) );
  NAND2_X1 U19111 ( .A1(n15783), .A2(n19790), .ZN(n15784) );
  XNOR2_X1 U19112 ( .A(n15784), .B(n16298), .ZN(n15785) );
  NAND2_X1 U19113 ( .A1(n15785), .A2(n19771), .ZN(n15786) );
  OAI211_X1 U19114 ( .C1(n15788), .C2(n19782), .A(n15787), .B(n15786), .ZN(
        n15789) );
  AOI21_X1 U19115 ( .B1(n15790), .B2(n19754), .A(n15789), .ZN(n15791) );
  OAI21_X1 U19116 ( .B1(n16570), .B2(n19767), .A(n15791), .ZN(P2_U2845) );
  NAND2_X1 U19117 ( .A1(n14452), .A2(n15792), .ZN(n15985) );
  NAND2_X1 U19118 ( .A1(n15985), .A2(n15793), .ZN(n15794) );
  NAND2_X1 U19119 ( .A1(n15777), .A2(n15794), .ZN(n16310) );
  INV_X1 U19120 ( .A(n16310), .ZN(n16580) );
  AOI21_X1 U19121 ( .B1(n15795), .B2(n19771), .A(n15843), .ZN(n15798) );
  NAND3_X1 U19122 ( .A1(n15855), .A2(n16307), .A3(n15796), .ZN(n15797) );
  OAI211_X1 U19123 ( .C1(n15798), .C2(n16307), .A(n19701), .B(n15797), .ZN(
        n15800) );
  NOR2_X1 U19124 ( .A1(n19778), .A2(n16306), .ZN(n15799) );
  AOI211_X1 U19125 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19784), .A(n15800), .B(
        n15799), .ZN(n15802) );
  NAND2_X1 U19126 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15801) );
  OAI211_X1 U19127 ( .C1(n15803), .C2(n19782), .A(n15802), .B(n15801), .ZN(
        n15804) );
  AOI21_X1 U19128 ( .B1(n16580), .B2(n19754), .A(n15804), .ZN(n15805) );
  OAI21_X1 U19129 ( .B1(n16583), .B2(n19767), .A(n15805), .ZN(P2_U2846) );
  NAND2_X1 U19130 ( .A1(n14049), .A2(n15806), .ZN(n16090) );
  NAND2_X1 U19131 ( .A1(n15808), .A2(n15807), .ZN(n15809) );
  NAND2_X1 U19132 ( .A1(n14049), .A2(n15809), .ZN(n15811) );
  NAND2_X1 U19133 ( .A1(n15811), .A2(n15810), .ZN(n15812) );
  NAND2_X1 U19134 ( .A1(n16090), .A2(n15812), .ZN(n20580) );
  INV_X1 U19135 ( .A(n20580), .ZN(n19814) );
  NOR2_X1 U19136 ( .A1(n19782), .A2(n16349), .ZN(n15821) );
  INV_X1 U19137 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16355) );
  AOI21_X1 U19138 ( .B1(n19771), .B2(n15813), .A(n15843), .ZN(n15816) );
  NAND3_X1 U19139 ( .A1(n15855), .A2(n16354), .A3(n15814), .ZN(n15815) );
  OAI21_X1 U19140 ( .B1(n15816), .B2(n16354), .A(n15815), .ZN(n15818) );
  INV_X1 U19141 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n20513) );
  NOR2_X1 U19142 ( .A1(n19778), .A2(n20513), .ZN(n15817) );
  AOI211_X1 U19143 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19784), .A(n15818), .B(
        n15817), .ZN(n15819) );
  OAI21_X1 U19144 ( .B1(n16355), .B2(n19775), .A(n15819), .ZN(n15820) );
  AOI211_X1 U19145 ( .C1(n19814), .C2(n19785), .A(n15821), .B(n15820), .ZN(
        n15824) );
  NAND2_X1 U19146 ( .A1(n15822), .A2(n19754), .ZN(n15823) );
  OAI211_X1 U19147 ( .C1(n20582), .C2(n19787), .A(n15824), .B(n15823), .ZN(
        P2_U2852) );
  OAI21_X1 U19148 ( .B1(n20488), .B2(n15837), .A(n19716), .ZN(n15828) );
  INV_X1 U19149 ( .A(n15837), .ZN(n15825) );
  NOR3_X1 U19150 ( .A1(n15826), .A2(n15825), .A3(n19938), .ZN(n15827) );
  AOI21_X1 U19151 ( .B1(n19938), .B2(n15828), .A(n15827), .ZN(n15829) );
  OAI21_X1 U19152 ( .B1(n19778), .B2(n20511), .A(n15829), .ZN(n15831) );
  NOR2_X1 U19153 ( .A1(n19775), .A2(n19949), .ZN(n15830) );
  AOI211_X1 U19154 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n19784), .A(n15831), .B(
        n15830), .ZN(n15833) );
  NAND2_X1 U19155 ( .A1(n20592), .A2(n19785), .ZN(n15832) );
  OAI211_X1 U19156 ( .C1(n19782), .C2(n15834), .A(n15833), .B(n15832), .ZN(
        n15835) );
  AOI21_X1 U19157 ( .B1(n19945), .B2(n19754), .A(n15835), .ZN(n15836) );
  OAI21_X1 U19158 ( .B1(n20590), .B2(n19787), .A(n15836), .ZN(P2_U2853) );
  NAND2_X1 U19159 ( .A1(n19784), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n15845) );
  OAI22_X1 U19160 ( .A1(n15842), .A2(n19775), .B1(n20509), .B2(n19778), .ZN(
        n15841) );
  OAI21_X1 U19161 ( .B1(n15838), .B2(n15853), .A(n15837), .ZN(n15839) );
  OR2_X1 U19162 ( .A1(n19764), .A2(n15839), .ZN(n16667) );
  NOR2_X1 U19163 ( .A1(n16667), .A2(n20488), .ZN(n15840) );
  AOI211_X1 U19164 ( .C1(n15843), .C2(n15842), .A(n15841), .B(n15840), .ZN(
        n15844) );
  OAI211_X1 U19165 ( .C1(n19782), .C2(n15846), .A(n15845), .B(n15844), .ZN(
        n15849) );
  NOR2_X1 U19166 ( .A1(n15847), .A2(n19786), .ZN(n15848) );
  AOI211_X1 U19167 ( .C1(n19785), .C2(n16086), .A(n15849), .B(n15848), .ZN(
        n15850) );
  OAI21_X1 U19168 ( .B1(n19968), .B2(n19787), .A(n15850), .ZN(P2_U2854) );
  OAI22_X1 U19169 ( .A1(n19606), .A2(n19778), .B1(n19767), .B2(n15851), .ZN(
        n15860) );
  INV_X1 U19170 ( .A(n15852), .ZN(n15858) );
  NAND2_X1 U19171 ( .A1(n19784), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n15857) );
  INV_X1 U19172 ( .A(n15853), .ZN(n16653) );
  NAND2_X1 U19173 ( .A1(n19775), .A2(n19716), .ZN(n15854) );
  AOI22_X1 U19174 ( .A1(n15855), .A2(n16653), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n15854), .ZN(n15856) );
  OAI211_X1 U19175 ( .C1(n15858), .C2(n19782), .A(n15857), .B(n15856), .ZN(
        n15859) );
  AOI211_X1 U19176 ( .C1(n16652), .C2(n19754), .A(n15860), .B(n15859), .ZN(
        n15861) );
  OAI21_X1 U19177 ( .B1(n16745), .B2(n19787), .A(n15861), .ZN(P2_U2855) );
  MUX2_X1 U19178 ( .A(n15862), .B(P2_EBX_REG_31__SCAN_IN), .S(n9574), .Z(
        P2_U2856) );
  NAND2_X1 U19179 ( .A1(n10031), .A2(n15863), .ZN(n15864) );
  XOR2_X1 U19180 ( .A(n15865), .B(n15864), .Z(n16009) );
  NOR2_X1 U19181 ( .A1(n16380), .A2(n9574), .ZN(n15866) );
  AOI21_X1 U19182 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9574), .A(n15866), .ZN(
        n15867) );
  OAI21_X1 U19183 ( .B1(n16009), .B2(n15975), .A(n15867), .ZN(P2_U2859) );
  NOR2_X1 U19184 ( .A1(n15868), .A2(n15879), .ZN(n15878) );
  NOR2_X1 U19185 ( .A1(n15878), .A2(n15869), .ZN(n15875) );
  NOR2_X1 U19186 ( .A1(n15871), .A2(n15870), .ZN(n15872) );
  XNOR2_X1 U19187 ( .A(n15873), .B(n15872), .ZN(n15874) );
  XNOR2_X1 U19188 ( .A(n15875), .B(n15874), .ZN(n16014) );
  MUX2_X1 U19189 ( .A(n15876), .B(n16405), .S(n16002), .Z(n15877) );
  OAI21_X1 U19190 ( .B1(n16014), .B2(n15975), .A(n15877), .ZN(P2_U2861) );
  AOI21_X1 U19191 ( .B1(n15868), .B2(n15879), .A(n15878), .ZN(n16015) );
  NAND2_X1 U19192 ( .A1(n16015), .A2(n15992), .ZN(n15881) );
  NAND2_X1 U19193 ( .A1(n9574), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15880) );
  OAI211_X1 U19194 ( .C1(n16414), .C2(n9574), .A(n15881), .B(n15880), .ZN(
        P2_U2862) );
  AOI21_X1 U19195 ( .B1(n15884), .B2(n15883), .A(n15882), .ZN(n15885) );
  XOR2_X1 U19196 ( .A(n15886), .B(n15885), .Z(n16029) );
  NOR2_X1 U19197 ( .A1(n16424), .A2(n9574), .ZN(n15887) );
  AOI21_X1 U19198 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n9574), .A(n15887), .ZN(
        n15888) );
  OAI21_X1 U19199 ( .B1(n16029), .B2(n15975), .A(n15888), .ZN(P2_U2863) );
  AOI21_X1 U19200 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(n16033) );
  NAND2_X1 U19201 ( .A1(n16033), .A2(n15992), .ZN(n15893) );
  NAND2_X1 U19202 ( .A1(n9574), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15892) );
  OAI211_X1 U19203 ( .C1(n16437), .C2(n9574), .A(n15893), .B(n15892), .ZN(
        P2_U2864) );
  INV_X1 U19204 ( .A(n16184), .ZN(n16449) );
  NAND2_X1 U19205 ( .A1(n15912), .A2(n15895), .ZN(n15899) );
  AOI21_X1 U19206 ( .B1(n15897), .B2(n15899), .A(n15896), .ZN(n16041) );
  AOI22_X1 U19207 ( .A1(n16041), .A2(n15992), .B1(P2_EBX_REG_22__SCAN_IN), 
        .B2(n9574), .ZN(n15898) );
  OAI21_X1 U19208 ( .B1(n16449), .B2(n9574), .A(n15898), .ZN(P2_U2865) );
  AND2_X1 U19209 ( .A1(n15912), .A2(n15904), .ZN(n15905) );
  OAI21_X1 U19210 ( .B1(n15905), .B2(n15900), .A(n15899), .ZN(n16050) );
  INV_X1 U19211 ( .A(n16050), .ZN(n15901) );
  AOI22_X1 U19212 ( .A1(n15901), .A2(n15992), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n9574), .ZN(n15902) );
  OAI21_X1 U19213 ( .B1(n15903), .B2(n9574), .A(n15902), .ZN(P2_U2866) );
  INV_X1 U19214 ( .A(n16461), .ZN(n15909) );
  INV_X1 U19215 ( .A(n15904), .ZN(n15907) );
  INV_X1 U19216 ( .A(n15912), .ZN(n15906) );
  AOI21_X1 U19217 ( .B1(n15907), .B2(n15906), .A(n15905), .ZN(n16056) );
  AOI22_X1 U19218 ( .A1(n16056), .A2(n15992), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n9574), .ZN(n15908) );
  OAI21_X1 U19219 ( .B1(n15909), .B2(n9574), .A(n15908), .ZN(P2_U2867) );
  NOR2_X1 U19220 ( .A1(n15894), .A2(n15910), .ZN(n15911) );
  OR2_X1 U19221 ( .A1(n15912), .A2(n15911), .ZN(n16063) );
  NAND2_X1 U19222 ( .A1(n19621), .A2(n16002), .ZN(n15914) );
  NAND2_X1 U19223 ( .A1(n9574), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15913) );
  OAI211_X1 U19224 ( .C1(n16063), .C2(n15975), .A(n15914), .B(n15913), .ZN(
        P2_U2868) );
  OAI21_X1 U19225 ( .B1(n14567), .B2(n15915), .A(n13587), .ZN(n16483) );
  AOI21_X1 U19226 ( .B1(n15917), .B2(n15916), .A(n15894), .ZN(n16072) );
  AOI22_X1 U19227 ( .A1(n16072), .A2(n15992), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n9574), .ZN(n15918) );
  OAI21_X1 U19228 ( .B1(n16483), .B2(n9574), .A(n15918), .ZN(P2_U2869) );
  INV_X1 U19229 ( .A(n15916), .ZN(n15920) );
  AOI21_X1 U19230 ( .B1(n15921), .B2(n15919), .A(n15920), .ZN(n16079) );
  AOI22_X1 U19231 ( .A1(n16079), .A2(n15992), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n9574), .ZN(n15922) );
  OAI21_X1 U19232 ( .B1(n15923), .B2(n9574), .A(n15922), .ZN(P2_U2870) );
  NOR2_X1 U19233 ( .A1(n15955), .A2(n15944), .ZN(n15941) );
  NAND2_X1 U19234 ( .A1(n15941), .A2(n15940), .ZN(n15939) );
  NOR2_X1 U19235 ( .A1(n15939), .A2(n15931), .ZN(n15926) );
  OAI21_X1 U19236 ( .B1(n15926), .B2(n15925), .A(n15919), .ZN(n19801) );
  AND2_X1 U19237 ( .A1(n15927), .A2(n15928), .ZN(n15929) );
  OR2_X1 U19238 ( .A1(n15929), .A2(n14568), .ZN(n16500) );
  MUX2_X1 U19239 ( .A(n16500), .B(n12692), .S(n9574), .Z(n15930) );
  OAI21_X1 U19240 ( .B1(n15975), .B2(n19801), .A(n15930), .ZN(P2_U2871) );
  XNOR2_X1 U19241 ( .A(n15939), .B(n15931), .ZN(n15937) );
  INV_X1 U19242 ( .A(n15927), .ZN(n15933) );
  AOI21_X1 U19243 ( .B1(n15934), .B2(n15932), .A(n15933), .ZN(n19664) );
  NAND2_X1 U19244 ( .A1(n19664), .A2(n16002), .ZN(n15936) );
  NAND2_X1 U19245 ( .A1(n9574), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n15935) );
  OAI211_X1 U19246 ( .C1(n15937), .C2(n15975), .A(n15936), .B(n15935), .ZN(
        P2_U2872) );
  OAI21_X1 U19247 ( .B1(n15763), .B2(n15938), .A(n15932), .ZN(n16245) );
  INV_X1 U19248 ( .A(n16245), .ZN(n19682) );
  NAND2_X1 U19249 ( .A1(n19682), .A2(n16002), .ZN(n15943) );
  OAI211_X1 U19250 ( .C1(n15941), .C2(n15940), .A(n15939), .B(n15992), .ZN(
        n15942) );
  OAI211_X1 U19251 ( .C1(n16002), .C2(n12697), .A(n15943), .B(n15942), .ZN(
        P2_U2873) );
  XNOR2_X1 U19252 ( .A(n15955), .B(n15944), .ZN(n15947) );
  INV_X1 U19253 ( .A(n16259), .ZN(n16531) );
  NOR2_X1 U19254 ( .A1(n16531), .A2(n9574), .ZN(n15945) );
  AOI21_X1 U19255 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n9574), .A(n15945), .ZN(
        n15946) );
  OAI21_X1 U19256 ( .B1(n15947), .B2(n15975), .A(n15946), .ZN(P2_U2874) );
  INV_X1 U19257 ( .A(n15762), .ZN(n15949) );
  AOI21_X1 U19258 ( .B1(n15950), .B2(n15948), .A(n15949), .ZN(n19697) );
  INV_X1 U19259 ( .A(n19697), .ZN(n15959) );
  NAND2_X1 U19260 ( .A1(n15991), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n15977) );
  NAND2_X1 U19261 ( .A1(n15978), .A2(n15972), .ZN(n15966) );
  NOR2_X1 U19262 ( .A1(n15966), .A2(n15952), .ZN(n15961) );
  INV_X1 U19263 ( .A(n15961), .ZN(n15967) );
  OAI21_X1 U19264 ( .B1(n15967), .B2(n15954), .A(n15953), .ZN(n15956) );
  NAND3_X1 U19265 ( .A1(n15956), .A2(n15992), .A3(n15955), .ZN(n15958) );
  NAND2_X1 U19266 ( .A1(n9574), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15957) );
  OAI211_X1 U19267 ( .C1(n15959), .C2(n9574), .A(n15958), .B(n15957), .ZN(
        P2_U2875) );
  XNOR2_X1 U19268 ( .A(n15961), .B(n15960), .ZN(n15965) );
  OAI21_X1 U19269 ( .B1(n15779), .B2(n15962), .A(n15948), .ZN(n16553) );
  NOR2_X1 U19270 ( .A1(n16553), .A2(n9574), .ZN(n15963) );
  AOI21_X1 U19271 ( .B1(P2_EBX_REG_11__SCAN_IN), .B2(n9574), .A(n15963), .ZN(
        n15964) );
  OAI21_X1 U19272 ( .B1(n15965), .B2(n15975), .A(n15964), .ZN(P2_U2876) );
  INV_X1 U19273 ( .A(n15966), .ZN(n15969) );
  OAI211_X1 U19274 ( .C1(n15969), .C2(n15968), .A(n15967), .B(n15992), .ZN(
        n15971) );
  NAND2_X1 U19275 ( .A1(n9574), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15970) );
  OAI211_X1 U19276 ( .C1(n16566), .C2(n9574), .A(n15971), .B(n15970), .ZN(
        P2_U2877) );
  XNOR2_X1 U19277 ( .A(n15978), .B(n15972), .ZN(n15976) );
  MUX2_X1 U19278 ( .A(n16310), .B(n15973), .S(n9574), .Z(n15974) );
  OAI21_X1 U19279 ( .B1(n15976), .B2(n15975), .A(n15974), .ZN(P2_U2878) );
  INV_X1 U19280 ( .A(n15977), .ZN(n15981) );
  INV_X1 U19281 ( .A(n15978), .ZN(n15979) );
  OAI211_X1 U19282 ( .C1(n15981), .C2(n15980), .A(n15979), .B(n15992), .ZN(
        n15987) );
  NAND2_X1 U19283 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  NAND2_X1 U19284 ( .A1(n15985), .A2(n15984), .ZN(n19726) );
  INV_X1 U19285 ( .A(n19726), .ZN(n16595) );
  NAND2_X1 U19286 ( .A1(n16595), .A2(n16002), .ZN(n15986) );
  OAI211_X1 U19287 ( .C1(n16002), .C2(n15988), .A(n15987), .B(n15986), .ZN(
        P2_U2879) );
  NOR2_X1 U19288 ( .A1(n15990), .A2(n15989), .ZN(n15994) );
  INV_X1 U19289 ( .A(n15991), .ZN(n15993) );
  OAI211_X1 U19290 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n15994), .A(
        n15993), .B(n15992), .ZN(n16000) );
  AND2_X1 U19291 ( .A1(n15996), .A2(n15995), .ZN(n15997) );
  NOR2_X1 U19292 ( .A1(n15998), .A2(n15997), .ZN(n19755) );
  NAND2_X1 U19293 ( .A1(n19755), .A2(n16002), .ZN(n15999) );
  OAI211_X1 U19294 ( .C1(n16002), .C2(n16001), .A(n16000), .B(n15999), .ZN(
        P2_U2881) );
  INV_X1 U19295 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19296 ( .A1(n19798), .A2(n16003), .B1(n19813), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n16004) );
  OAI21_X1 U19297 ( .B1(n16077), .B2(n16005), .A(n16004), .ZN(n16007) );
  NOR2_X1 U19298 ( .A1(n16374), .A2(n16081), .ZN(n16006) );
  AOI211_X1 U19299 ( .C1(n19800), .C2(BUF1_REG_28__SCAN_IN), .A(n16007), .B(
        n16006), .ZN(n16008) );
  OAI21_X1 U19300 ( .B1(n16009), .B2(n16062), .A(n16008), .ZN(P2_U2891) );
  INV_X1 U19301 ( .A(n19800), .ZN(n16054) );
  AOI22_X1 U19302 ( .A1(n19798), .A2(n19906), .B1(n19813), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n16011) );
  NAND2_X1 U19303 ( .A1(n19799), .A2(BUF2_REG_26__SCAN_IN), .ZN(n16010) );
  OAI211_X1 U19304 ( .C1(n16054), .C2(n19991), .A(n16011), .B(n16010), .ZN(
        n16012) );
  AOI21_X1 U19305 ( .B1(n16407), .B2(n19823), .A(n16012), .ZN(n16013) );
  OAI21_X1 U19306 ( .B1(n16014), .B2(n16062), .A(n16013), .ZN(P2_U2893) );
  INV_X1 U19307 ( .A(n16416), .ZN(n16022) );
  NAND2_X1 U19308 ( .A1(n16015), .A2(n19828), .ZN(n16021) );
  INV_X1 U19309 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n16018) );
  AOI22_X1 U19310 ( .A1(n19798), .A2(n16016), .B1(n19813), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16017) );
  OAI21_X1 U19311 ( .B1(n16077), .B2(n16018), .A(n16017), .ZN(n16019) );
  AOI21_X1 U19312 ( .B1(n19800), .B2(BUF1_REG_25__SCAN_IN), .A(n16019), .ZN(
        n16020) );
  OAI211_X1 U19313 ( .C1(n16022), .C2(n16081), .A(n16021), .B(n16020), .ZN(
        P2_U2894) );
  INV_X1 U19314 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n16026) );
  AOI22_X1 U19315 ( .A1(n19798), .A2(n16023), .B1(n19813), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16025) );
  NAND2_X1 U19316 ( .A1(n19800), .A2(BUF1_REG_24__SCAN_IN), .ZN(n16024) );
  OAI211_X1 U19317 ( .C1(n16077), .C2(n16026), .A(n16025), .B(n16024), .ZN(
        n16027) );
  AOI21_X1 U19318 ( .B1(n16426), .B2(n19823), .A(n16027), .ZN(n16028) );
  OAI21_X1 U19319 ( .B1(n16029), .B2(n16062), .A(n16028), .ZN(P2_U2895) );
  INV_X1 U19320 ( .A(n16439), .ZN(n16036) );
  INV_X1 U19321 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n16031) );
  AOI22_X1 U19322 ( .A1(n19798), .A2(n16739), .B1(n19813), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16030) );
  OAI21_X1 U19323 ( .B1(n16077), .B2(n16031), .A(n16030), .ZN(n16032) );
  AOI21_X1 U19324 ( .B1(n19800), .B2(BUF1_REG_23__SCAN_IN), .A(n16032), .ZN(
        n16035) );
  NAND2_X1 U19325 ( .A1(n16033), .A2(n19828), .ZN(n16034) );
  OAI211_X1 U19326 ( .C1(n16036), .C2(n16081), .A(n16035), .B(n16034), .ZN(
        P2_U2896) );
  INV_X1 U19327 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16039) );
  AOI22_X1 U19328 ( .A1(n19798), .A2(n16734), .B1(n19813), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U19329 ( .A1(n19799), .A2(BUF2_REG_22__SCAN_IN), .ZN(n16037) );
  OAI211_X1 U19330 ( .C1(n16054), .C2(n16039), .A(n16038), .B(n16037), .ZN(
        n16040) );
  AOI21_X1 U19331 ( .B1(n16041), .B2(n19828), .A(n16040), .ZN(n16042) );
  OAI21_X1 U19332 ( .B1(n16043), .B2(n16081), .A(n16042), .ZN(P2_U2897) );
  NAND2_X1 U19333 ( .A1(n16044), .A2(n19823), .ZN(n16049) );
  INV_X1 U19334 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n16046) );
  AOI22_X1 U19335 ( .A1(n19798), .A2(n16784), .B1(n19813), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n16045) );
  OAI21_X1 U19336 ( .B1(n16077), .B2(n16046), .A(n16045), .ZN(n16047) );
  AOI21_X1 U19337 ( .B1(n19800), .B2(BUF1_REG_21__SCAN_IN), .A(n16047), .ZN(
        n16048) );
  OAI211_X1 U19338 ( .C1(n16062), .C2(n16050), .A(n16049), .B(n16048), .ZN(
        P2_U2898) );
  INV_X1 U19339 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16053) );
  AOI22_X1 U19340 ( .A1(n19798), .A2(n20001), .B1(n19813), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16052) );
  NAND2_X1 U19341 ( .A1(n19799), .A2(BUF2_REG_20__SCAN_IN), .ZN(n16051) );
  OAI211_X1 U19342 ( .C1(n16054), .C2(n16053), .A(n16052), .B(n16051), .ZN(
        n16055) );
  AOI21_X1 U19343 ( .B1(n16056), .B2(n19828), .A(n16055), .ZN(n16057) );
  OAI21_X1 U19344 ( .B1(n16463), .B2(n16081), .A(n16057), .ZN(P2_U2899) );
  XNOR2_X1 U19345 ( .A(n16058), .B(n16059), .ZN(n19619) );
  INV_X1 U19346 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U19347 ( .A1(n19798), .A2(n19995), .B1(n19813), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n16060) );
  OAI21_X1 U19348 ( .B1(n16077), .B2(n16061), .A(n16060), .ZN(n16065) );
  NOR2_X1 U19349 ( .A1(n16063), .A2(n16062), .ZN(n16064) );
  AOI211_X1 U19350 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n19800), .A(n16065), .B(
        n16064), .ZN(n16066) );
  OAI21_X1 U19351 ( .B1(n19619), .B2(n16081), .A(n16066), .ZN(P2_U2900) );
  OAI21_X1 U19352 ( .B1(n14564), .B2(n16067), .A(n16058), .ZN(n19635) );
  INV_X1 U19353 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n16070) );
  AOI22_X1 U19354 ( .A1(n19798), .A2(n19989), .B1(n19813), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16069) );
  NAND2_X1 U19355 ( .A1(n19800), .A2(BUF1_REG_18__SCAN_IN), .ZN(n16068) );
  OAI211_X1 U19356 ( .C1(n16077), .C2(n16070), .A(n16069), .B(n16068), .ZN(
        n16071) );
  AOI21_X1 U19357 ( .B1(n16072), .B2(n19828), .A(n16071), .ZN(n16073) );
  OAI21_X1 U19358 ( .B1(n19635), .B2(n16081), .A(n16073), .ZN(P2_U2901) );
  INV_X1 U19359 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19360 ( .A1(n19798), .A2(n19983), .B1(n19813), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16075) );
  NAND2_X1 U19361 ( .A1(n19800), .A2(BUF1_REG_17__SCAN_IN), .ZN(n16074) );
  OAI211_X1 U19362 ( .C1(n16077), .C2(n16076), .A(n16075), .B(n16074), .ZN(
        n16078) );
  AOI21_X1 U19363 ( .B1(n16079), .B2(n19828), .A(n16078), .ZN(n16080) );
  OAI21_X1 U19364 ( .B1(n16082), .B2(n16081), .A(n16080), .ZN(P2_U2902) );
  INV_X1 U19365 ( .A(n16084), .ZN(n16085) );
  XNOR2_X1 U19366 ( .A(n16083), .B(n16085), .ZN(n16644) );
  INV_X1 U19367 ( .A(n16644), .ZN(n19768) );
  XNOR2_X1 U19368 ( .A(n20590), .B(n20592), .ZN(n19827) );
  OAI22_X1 U19369 ( .A1(n16088), .A2(n16087), .B1(n16744), .B2(n16086), .ZN(
        n19826) );
  NAND2_X1 U19370 ( .A1(n19827), .A2(n19826), .ZN(n19825) );
  OAI21_X1 U19371 ( .B1(n16683), .B2(n20592), .A(n19825), .ZN(n19816) );
  XNOR2_X1 U19372 ( .A(n16746), .B(n20580), .ZN(n19817) );
  NAND2_X1 U19373 ( .A1(n19816), .A2(n19817), .ZN(n19815) );
  OAI21_X1 U19374 ( .B1(n19814), .B2(n16746), .A(n19815), .ZN(n16092) );
  NAND2_X1 U19375 ( .A1(n16090), .A2(n16089), .ZN(n16091) );
  NAND2_X1 U19376 ( .A1(n16083), .A2(n16091), .ZN(n19960) );
  NAND2_X1 U19377 ( .A1(n16092), .A2(n19960), .ZN(n19809) );
  INV_X1 U19378 ( .A(n19808), .ZN(n16093) );
  NAND3_X1 U19379 ( .A1(n19809), .A2(n19828), .A3(n16093), .ZN(n16095) );
  AOI22_X1 U19380 ( .A1(n19824), .A2(n16784), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19813), .ZN(n16094) );
  OAI211_X1 U19381 ( .C1(n19768), .C2(n16096), .A(n16095), .B(n16094), .ZN(
        P2_U2914) );
  INV_X1 U19382 ( .A(n16099), .ZN(n16125) );
  NOR2_X1 U19383 ( .A1(n16102), .A2(n13080), .ZN(n16103) );
  NOR2_X1 U19384 ( .A1(n19939), .A2(n16104), .ZN(n16107) );
  OR2_X1 U19385 ( .A1(n19701), .A2(n20556), .ZN(n16365) );
  OAI21_X1 U19386 ( .B1(n19950), .B2(n16105), .A(n16365), .ZN(n16106) );
  AOI211_X1 U19387 ( .C1(n16369), .C2(n19946), .A(n16107), .B(n16106), .ZN(
        n16109) );
  NAND2_X1 U19388 ( .A1(n16370), .A2(n16335), .ZN(n16108) );
  INV_X1 U19389 ( .A(n16110), .ZN(n16112) );
  OAI21_X1 U19390 ( .B1(n16112), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16111), .ZN(n16384) );
  OAI211_X1 U19391 ( .C1(n12523), .C2(n16377), .A(n16113), .B(n16148), .ZN(
        n16114) );
  NAND2_X1 U19392 ( .A1(n9777), .A2(n19946), .ZN(n16119) );
  NOR2_X1 U19393 ( .A1(n19701), .A2(n16117), .ZN(n16378) );
  AOI21_X1 U19394 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16378), .ZN(n16118) );
  OAI211_X1 U19395 ( .C1(n19939), .C2(n16120), .A(n16119), .B(n16118), .ZN(
        n16121) );
  AOI21_X1 U19396 ( .B1(n19936), .B2(n16382), .A(n16121), .ZN(n16122) );
  OAI21_X1 U19397 ( .B1(n19941), .B2(n16384), .A(n16122), .ZN(P2_U2986) );
  INV_X1 U19398 ( .A(n16123), .ZN(n16124) );
  OAI21_X1 U19399 ( .B1(n16124), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16110), .ZN(n16396) );
  NAND2_X1 U19400 ( .A1(n16126), .A2(n16125), .ZN(n16129) );
  XNOR2_X1 U19401 ( .A(n16127), .B(n16377), .ZN(n16128) );
  XNOR2_X1 U19402 ( .A(n16129), .B(n16128), .ZN(n16394) );
  INV_X1 U19403 ( .A(n16392), .ZN(n16130) );
  NAND2_X1 U19404 ( .A1(n16130), .A2(n19946), .ZN(n16132) );
  NOR2_X1 U19405 ( .A1(n19701), .A2(n20554), .ZN(n16387) );
  AOI21_X1 U19406 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16387), .ZN(n16131) );
  OAI211_X1 U19407 ( .C1(n19939), .C2(n16133), .A(n16132), .B(n16131), .ZN(
        n16134) );
  AOI21_X1 U19408 ( .B1(n19936), .B2(n16394), .A(n16134), .ZN(n16135) );
  OAI21_X1 U19409 ( .B1(n19941), .B2(n16396), .A(n16135), .ZN(P2_U2987) );
  INV_X1 U19410 ( .A(n16178), .ZN(n16136) );
  INV_X1 U19411 ( .A(n16157), .ZN(n16138) );
  INV_X1 U19412 ( .A(n16139), .ZN(n16140) );
  NOR2_X1 U19413 ( .A1(n19701), .A2(n16142), .ZN(n16398) );
  AOI21_X1 U19414 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16398), .ZN(n16143) );
  OAI21_X1 U19415 ( .B1(n19939), .B2(n16144), .A(n16143), .ZN(n16145) );
  NAND2_X1 U19416 ( .A1(n16148), .A2(n16147), .ZN(n16149) );
  NOR2_X1 U19417 ( .A1(n19701), .A2(n20550), .ZN(n16411) );
  INV_X1 U19418 ( .A(n16411), .ZN(n16150) );
  OAI21_X1 U19419 ( .B1(n19950), .B2(n16151), .A(n16150), .ZN(n16153) );
  NOR2_X1 U19420 ( .A1(n16414), .A2(n19928), .ZN(n16152) );
  AOI211_X1 U19421 ( .C1(n19917), .C2(n16154), .A(n16153), .B(n16152), .ZN(
        n16156) );
  OR3_X1 U19422 ( .A1(n16409), .A2(n16141), .A3(n19941), .ZN(n16155) );
  OAI211_X1 U19423 ( .C1(n16417), .C2(n17292), .A(n16156), .B(n16155), .ZN(
        P2_U2989) );
  NAND2_X1 U19424 ( .A1(n16158), .A2(n16157), .ZN(n16160) );
  XOR2_X1 U19425 ( .A(n16160), .B(n16159), .Z(n16430) );
  INV_X1 U19426 ( .A(n16424), .ZN(n16162) );
  NAND2_X1 U19427 ( .A1(n16162), .A2(n19946), .ZN(n16164) );
  NOR2_X1 U19428 ( .A1(n19701), .A2(n20548), .ZN(n16418) );
  AOI21_X1 U19429 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16418), .ZN(n16163) );
  OAI211_X1 U19430 ( .C1(n16165), .C2(n19939), .A(n16164), .B(n16163), .ZN(
        n16166) );
  OAI21_X1 U19431 ( .B1(n16430), .B2(n17292), .A(n16167), .ZN(P2_U2990) );
  OAI21_X1 U19432 ( .B1(n16185), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16168), .ZN(n16443) );
  NAND2_X1 U19433 ( .A1(n16341), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n16433) );
  OAI21_X1 U19434 ( .B1(n19950), .B2(n16169), .A(n16433), .ZN(n16171) );
  NOR2_X1 U19435 ( .A1(n16437), .A2(n19928), .ZN(n16170) );
  AOI211_X1 U19436 ( .C1(n19917), .C2(n16172), .A(n16171), .B(n16170), .ZN(
        n16177) );
  OR2_X1 U19437 ( .A1(n16174), .A2(n16173), .ZN(n16440) );
  NAND3_X1 U19438 ( .A1(n16440), .A2(n16175), .A3(n19936), .ZN(n16176) );
  OAI211_X1 U19439 ( .C1(n16443), .C2(n19941), .A(n16177), .B(n16176), .ZN(
        P2_U2991) );
  NAND2_X1 U19440 ( .A1(n16179), .A2(n16178), .ZN(n16180) );
  XNOR2_X1 U19441 ( .A(n9681), .B(n16180), .ZN(n16456) );
  NOR2_X1 U19442 ( .A1(n19701), .A2(n20544), .ZN(n16446) );
  AOI21_X1 U19443 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n16446), .ZN(n16181) );
  OAI21_X1 U19444 ( .B1(n16182), .B2(n19939), .A(n16181), .ZN(n16183) );
  AOI21_X1 U19445 ( .B1(n16184), .B2(n19946), .A(n16183), .ZN(n16189) );
  INV_X1 U19446 ( .A(n16185), .ZN(n16453) );
  NAND2_X1 U19447 ( .A1(n16187), .A2(n16186), .ZN(n16452) );
  NAND3_X1 U19448 ( .A1(n16453), .A2(n16335), .A3(n16452), .ZN(n16188) );
  OAI211_X1 U19449 ( .C1(n16456), .C2(n17292), .A(n16189), .B(n16188), .ZN(
        P2_U2992) );
  NAND2_X1 U19450 ( .A1(n16191), .A2(n16190), .ZN(n16195) );
  NAND2_X1 U19451 ( .A1(n16193), .A2(n16192), .ZN(n16194) );
  NAND2_X1 U19452 ( .A1(n16461), .A2(n19946), .ZN(n16198) );
  NOR2_X1 U19453 ( .A1(n19701), .A2(n20540), .ZN(n16460) );
  AOI21_X1 U19454 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16460), .ZN(n16197) );
  OAI211_X1 U19455 ( .C1(n16199), .C2(n19939), .A(n16198), .B(n16197), .ZN(
        n16200) );
  AOI21_X1 U19456 ( .B1(n16466), .B2(n16335), .A(n16200), .ZN(n16201) );
  NAND2_X1 U19457 ( .A1(n16203), .A2(n16202), .ZN(n16204) );
  XNOR2_X1 U19458 ( .A(n16205), .B(n16204), .ZN(n16493) );
  NAND2_X1 U19459 ( .A1(n16206), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16214) );
  INV_X1 U19460 ( .A(n16207), .ZN(n16208) );
  AOI21_X2 U19461 ( .B1(n16214), .B2(n16481), .A(n16208), .ZN(n16491) );
  NOR2_X1 U19462 ( .A1(n19701), .A2(n19630), .ZN(n16487) );
  NOR2_X1 U19463 ( .A1(n19939), .A2(n19641), .ZN(n16209) );
  AOI211_X1 U19464 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17289), .A(
        n16487), .B(n16209), .ZN(n16210) );
  OAI21_X1 U19465 ( .B1(n16483), .B2(n19928), .A(n16210), .ZN(n16211) );
  AOI21_X1 U19466 ( .B1(n16491), .B2(n16335), .A(n16211), .ZN(n16212) );
  OAI21_X1 U19467 ( .B1(n17292), .B2(n16493), .A(n16212), .ZN(P2_U2996) );
  INV_X1 U19468 ( .A(n16213), .ZN(n16222) );
  OAI211_X1 U19469 ( .C1(n16206), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16214), .B(n16335), .ZN(n16221) );
  NAND2_X1 U19470 ( .A1(n17289), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n16215) );
  OAI211_X1 U19471 ( .C1(n19939), .C2(n16217), .A(n16216), .B(n16215), .ZN(
        n16218) );
  AOI21_X1 U19472 ( .B1(n16219), .B2(n19946), .A(n16218), .ZN(n16220) );
  OAI211_X1 U19473 ( .C1(n16222), .C2(n17292), .A(n16221), .B(n16220), .ZN(
        P2_U2997) );
  INV_X1 U19474 ( .A(n16502), .ZN(n16229) );
  INV_X1 U19475 ( .A(n16224), .ZN(n16494) );
  OAI211_X1 U19476 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16494), .A(
        n9932), .B(n16335), .ZN(n16228) );
  INV_X1 U19477 ( .A(n16500), .ZN(n19654) );
  NAND2_X1 U19478 ( .A1(n16341), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n16499) );
  NAND2_X1 U19479 ( .A1(n17289), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16225) );
  OAI211_X1 U19480 ( .C1(n19939), .C2(n19647), .A(n16499), .B(n16225), .ZN(
        n16226) );
  AOI21_X1 U19481 ( .B1(n19654), .B2(n19946), .A(n16226), .ZN(n16227) );
  OAI211_X1 U19482 ( .C1(n16229), .C2(n17292), .A(n16228), .B(n16227), .ZN(
        P2_U2998) );
  AND2_X1 U19483 ( .A1(n16232), .A2(n16231), .ZN(n16233) );
  XNOR2_X1 U19484 ( .A(n16230), .B(n16233), .ZN(n16515) );
  NAND2_X1 U19485 ( .A1(n9622), .A2(n14555), .ZN(n16506) );
  NAND3_X1 U19486 ( .A1(n16506), .A2(n16335), .A3(n16224), .ZN(n16237) );
  NOR2_X1 U19487 ( .A1(n19701), .A2(n20531), .ZN(n16507) );
  AOI21_X1 U19488 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16507), .ZN(n16234) );
  OAI21_X1 U19489 ( .B1(n19939), .B2(n19663), .A(n16234), .ZN(n16235) );
  AOI21_X1 U19490 ( .B1(n19664), .B2(n19946), .A(n16235), .ZN(n16236) );
  OAI211_X1 U19491 ( .C1(n16515), .C2(n17292), .A(n16237), .B(n16236), .ZN(
        P2_U2999) );
  INV_X1 U19492 ( .A(n16527), .ZN(n16517) );
  OAI21_X1 U19493 ( .B1(n16253), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n9622), .ZN(n16525) );
  NAND2_X1 U19494 ( .A1(n16239), .A2(n16238), .ZN(n16240) );
  XNOR2_X1 U19495 ( .A(n16241), .B(n16240), .ZN(n16522) );
  NOR2_X1 U19496 ( .A1(n19701), .A2(n20529), .ZN(n16518) );
  NOR2_X1 U19497 ( .A1(n19939), .A2(n16242), .ZN(n16243) );
  AOI211_X1 U19498 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17289), .A(
        n16518), .B(n16243), .ZN(n16244) );
  OAI21_X1 U19499 ( .B1(n16245), .B2(n19928), .A(n16244), .ZN(n16246) );
  AOI21_X1 U19500 ( .B1(n16522), .B2(n19936), .A(n16246), .ZN(n16247) );
  OAI21_X1 U19501 ( .B1(n16525), .B2(n19941), .A(n16247), .ZN(P2_U3000) );
  NAND2_X1 U19502 ( .A1(n16248), .A2(n16263), .ZN(n16252) );
  NAND2_X1 U19503 ( .A1(n16250), .A2(n16249), .ZN(n16251) );
  XNOR2_X1 U19504 ( .A(n16252), .B(n16251), .ZN(n16537) );
  NAND2_X1 U19505 ( .A1(n19917), .A2(n16255), .ZN(n16256) );
  NAND2_X1 U19506 ( .A1(n16341), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n16530) );
  OAI211_X1 U19507 ( .C1(n16257), .C2(n19950), .A(n16256), .B(n16530), .ZN(
        n16258) );
  AOI21_X1 U19508 ( .B1(n16259), .B2(n19946), .A(n16258), .ZN(n16260) );
  OAI211_X1 U19509 ( .C1(n17292), .C2(n16537), .A(n16261), .B(n16260), .ZN(
        P2_U3001) );
  INV_X1 U19510 ( .A(n16263), .ZN(n16265) );
  NOR2_X1 U19511 ( .A1(n16265), .A2(n16264), .ZN(n16266) );
  XNOR2_X1 U19512 ( .A(n16262), .B(n16266), .ZN(n16548) );
  NAND2_X1 U19513 ( .A1(n16268), .A2(n16526), .ZN(n16538) );
  NAND3_X1 U19514 ( .A1(n16539), .A2(n16335), .A3(n16538), .ZN(n16272) );
  NOR2_X1 U19515 ( .A1(n19701), .A2(n20526), .ZN(n16540) );
  AOI21_X1 U19516 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16540), .ZN(n16269) );
  OAI21_X1 U19517 ( .B1(n19690), .B2(n19939), .A(n16269), .ZN(n16270) );
  AOI21_X1 U19518 ( .B1(n19697), .B2(n19946), .A(n16270), .ZN(n16271) );
  OAI211_X1 U19519 ( .C1(n16548), .C2(n17292), .A(n16272), .B(n16271), .ZN(
        P2_U3002) );
  NAND2_X1 U19520 ( .A1(n16274), .A2(n16273), .ZN(n16283) );
  XNOR2_X1 U19521 ( .A(n16277), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16343) );
  NAND2_X1 U19522 ( .A1(n16305), .A2(n16303), .ZN(n16292) );
  INV_X1 U19523 ( .A(n16291), .ZN(n16281) );
  OAI21_X1 U19524 ( .B1(n16292), .B2(n16281), .A(n16280), .ZN(n16282) );
  XOR2_X1 U19525 ( .A(n16283), .B(n16282), .Z(n16561) );
  AOI21_X1 U19526 ( .B1(n16551), .B2(n16284), .A(n16285), .ZN(n16559) );
  NOR2_X1 U19527 ( .A1(n19701), .A2(n19703), .ZN(n16554) );
  NOR2_X1 U19528 ( .A1(n19939), .A2(n19715), .ZN(n16286) );
  AOI211_X1 U19529 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17289), .A(
        n16554), .B(n16286), .ZN(n16287) );
  OAI21_X1 U19530 ( .B1(n16553), .B2(n19928), .A(n16287), .ZN(n16288) );
  AOI21_X1 U19531 ( .B1(n16559), .B2(n16335), .A(n16288), .ZN(n16289) );
  OAI21_X1 U19532 ( .B1(n16561), .B2(n17292), .A(n16289), .ZN(P2_U3003) );
  NAND2_X1 U19533 ( .A1(n16291), .A2(n16290), .ZN(n16294) );
  NAND2_X1 U19534 ( .A1(n16292), .A2(n16302), .ZN(n16293) );
  XOR2_X1 U19535 ( .A(n16294), .B(n16293), .Z(n16575) );
  AOI21_X1 U19536 ( .B1(n13663), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16295) );
  NOR2_X1 U19537 ( .A1(n13581), .A2(n16295), .ZN(n16573) );
  OR2_X1 U19538 ( .A1(n19701), .A2(n20523), .ZN(n16565) );
  OAI21_X1 U19539 ( .B1(n19950), .B2(n16296), .A(n16565), .ZN(n16297) );
  AOI21_X1 U19540 ( .B1(n19917), .B2(n16298), .A(n16297), .ZN(n16299) );
  OAI21_X1 U19541 ( .B1(n16566), .B2(n19928), .A(n16299), .ZN(n16300) );
  AOI21_X1 U19542 ( .B1(n16573), .B2(n16335), .A(n16300), .ZN(n16301) );
  OAI21_X1 U19543 ( .B1(n16575), .B2(n17292), .A(n16301), .ZN(P2_U3004) );
  XNOR2_X1 U19544 ( .A(n13663), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16588) );
  NAND2_X1 U19545 ( .A1(n16303), .A2(n16302), .ZN(n16304) );
  XNOR2_X1 U19546 ( .A(n16305), .B(n16304), .ZN(n16586) );
  NOR2_X1 U19547 ( .A1(n19701), .A2(n16306), .ZN(n16579) );
  NOR2_X1 U19548 ( .A1(n19939), .A2(n16307), .ZN(n16308) );
  AOI211_X1 U19549 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17289), .A(
        n16579), .B(n16308), .ZN(n16309) );
  OAI21_X1 U19550 ( .B1(n16310), .B2(n19928), .A(n16309), .ZN(n16311) );
  AOI21_X1 U19551 ( .B1(n16586), .B2(n19936), .A(n16311), .ZN(n16312) );
  OAI21_X1 U19552 ( .B1(n16588), .B2(n19941), .A(n16312), .ZN(P2_U3005) );
  NAND2_X1 U19553 ( .A1(n16315), .A2(n16314), .ZN(n16333) );
  NOR2_X1 U19554 ( .A1(n16334), .A2(n16333), .ZN(n16332) );
  XNOR2_X1 U19555 ( .A(n16315), .B(n16593), .ZN(n16316) );
  XNOR2_X1 U19556 ( .A(n16317), .B(n16316), .ZN(n16601) );
  NAND2_X1 U19557 ( .A1(n16319), .A2(n16318), .ZN(n16322) );
  NAND2_X1 U19558 ( .A1(n16320), .A2(n16330), .ZN(n16321) );
  XOR2_X1 U19559 ( .A(n16322), .B(n16321), .Z(n16599) );
  NAND2_X1 U19560 ( .A1(n16341), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16592) );
  OAI21_X1 U19561 ( .B1(n19950), .B2(n19721), .A(n16592), .ZN(n16323) );
  AOI21_X1 U19562 ( .B1(n19917), .B2(n19719), .A(n16323), .ZN(n16324) );
  OAI21_X1 U19563 ( .B1(n19726), .B2(n19928), .A(n16324), .ZN(n16325) );
  AOI21_X1 U19564 ( .B1(n16599), .B2(n19936), .A(n16325), .ZN(n16326) );
  OAI21_X1 U19565 ( .B1(n16601), .B2(n19941), .A(n16326), .ZN(P2_U3006) );
  AOI21_X1 U19566 ( .B1(n16330), .B2(n16328), .A(n16327), .ZN(n16329) );
  AOI21_X1 U19567 ( .B1(n16331), .B2(n16330), .A(n16329), .ZN(n16615) );
  INV_X1 U19568 ( .A(n16332), .ZN(n16604) );
  NAND2_X1 U19569 ( .A1(n16334), .A2(n16333), .ZN(n16602) );
  NAND3_X1 U19570 ( .A1(n16604), .A2(n16335), .A3(n16602), .ZN(n16339) );
  INV_X1 U19571 ( .A(n19740), .ZN(n16608) );
  NOR2_X1 U19572 ( .A1(n19701), .A2(n20518), .ZN(n16607) );
  AOI21_X1 U19573 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16607), .ZN(n16336) );
  OAI21_X1 U19574 ( .B1(n19733), .B2(n19939), .A(n16336), .ZN(n16337) );
  AOI21_X1 U19575 ( .B1(n16608), .B2(n19946), .A(n16337), .ZN(n16338) );
  OAI211_X1 U19576 ( .C1(n16615), .C2(n17292), .A(n16339), .B(n16338), .ZN(
        P2_U3007) );
  NAND2_X1 U19577 ( .A1(n19917), .A2(n19747), .ZN(n16342) );
  NAND2_X1 U19578 ( .A1(n16341), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n16616) );
  OAI211_X1 U19579 ( .C1(n19748), .C2(n19950), .A(n16342), .B(n16616), .ZN(
        n16345) );
  XNOR2_X1 U19580 ( .A(n16276), .B(n16343), .ZN(n16620) );
  NOR2_X1 U19581 ( .A1(n16620), .A2(n17292), .ZN(n16344) );
  AOI211_X1 U19582 ( .C1(n19946), .C2(n19755), .A(n16345), .B(n16344), .ZN(
        n16346) );
  OAI21_X1 U19583 ( .B1(n19941), .B2(n16626), .A(n16346), .ZN(P2_U3008) );
  XNOR2_X1 U19584 ( .A(n16348), .B(n16347), .ZN(n17301) );
  NAND2_X1 U19585 ( .A1(n16350), .A2(n16349), .ZN(n16352) );
  INV_X1 U19586 ( .A(n16352), .ZN(n16351) );
  NAND2_X1 U19587 ( .A1(n16351), .A2(n17306), .ZN(n19924) );
  NAND2_X1 U19588 ( .A1(n16352), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19922) );
  NAND2_X1 U19589 ( .A1(n19924), .A2(n19922), .ZN(n16353) );
  XNOR2_X1 U19590 ( .A(n16353), .B(n19920), .ZN(n17303) );
  NAND2_X1 U19591 ( .A1(n17303), .A2(n19936), .ZN(n16359) );
  NOR2_X1 U19592 ( .A1(n19939), .A2(n16354), .ZN(n16357) );
  OR2_X1 U19593 ( .A1(n19701), .A2(n20513), .ZN(n17298) );
  OAI21_X1 U19594 ( .B1(n19950), .B2(n16355), .A(n17298), .ZN(n16356) );
  AOI211_X1 U19595 ( .C1(n15822), .C2(n19946), .A(n16357), .B(n16356), .ZN(
        n16358) );
  OAI211_X1 U19596 ( .C1(n17301), .C2(n19941), .A(n16359), .B(n16358), .ZN(
        P2_U3011) );
  NOR2_X1 U19597 ( .A1(n16360), .A2(n19959), .ZN(n16368) );
  NOR2_X1 U19598 ( .A1(n16385), .A2(n16362), .ZN(n16361) );
  NOR2_X1 U19599 ( .A1(n16388), .A2(n16361), .ZN(n16375) );
  INV_X1 U19600 ( .A(n16385), .ZN(n16363) );
  NAND3_X1 U19601 ( .A1(n16363), .A2(n16362), .A3(n16366), .ZN(n16364) );
  OAI211_X1 U19602 ( .C1(n16375), .C2(n16366), .A(n16365), .B(n16364), .ZN(
        n16367) );
  NAND2_X1 U19603 ( .A1(n16370), .A2(n16603), .ZN(n16371) );
  NOR2_X1 U19604 ( .A1(n16374), .A2(n19959), .ZN(n16381) );
  OAI21_X1 U19605 ( .B1(n16385), .B2(n16377), .A(n16376), .ZN(n16379) );
  OAI21_X1 U19606 ( .B1(n19967), .B2(n16384), .A(n16383), .ZN(P2_U3018) );
  NOR2_X1 U19607 ( .A1(n16385), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16386) );
  AOI211_X1 U19608 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n16388), .A(
        n16387), .B(n16386), .ZN(n16391) );
  NAND2_X1 U19609 ( .A1(n16389), .A2(n16645), .ZN(n16390) );
  OAI211_X1 U19610 ( .C1(n16392), .C2(n16639), .A(n16391), .B(n16390), .ZN(
        n16393) );
  AOI21_X1 U19611 ( .B1(n19962), .B2(n16394), .A(n16393), .ZN(n16395) );
  OAI21_X1 U19612 ( .B1(n19967), .B2(n16396), .A(n16395), .ZN(P2_U3019) );
  AOI21_X1 U19613 ( .B1(n16400), .B2(n16399), .A(n16398), .ZN(n16404) );
  AND2_X1 U19614 ( .A1(n16401), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16402) );
  AND2_X1 U19615 ( .A1(n16420), .A2(n16402), .ZN(n16410) );
  OAI21_X1 U19616 ( .B1(n16412), .B2(n16410), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16403) );
  OAI211_X1 U19617 ( .C1(n16405), .C2(n16639), .A(n16404), .B(n16403), .ZN(
        n16406) );
  AOI211_X1 U19618 ( .C1(n16412), .C2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n16411), .B(n16410), .ZN(n16413) );
  OAI21_X1 U19619 ( .B1(n16414), .B2(n16639), .A(n16413), .ZN(n16415) );
  AOI21_X1 U19620 ( .B1(n16420), .B2(n16419), .A(n16418), .ZN(n16423) );
  NAND2_X1 U19621 ( .A1(n16421), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16422) );
  OAI211_X1 U19622 ( .C1(n16424), .C2(n16639), .A(n16423), .B(n16422), .ZN(
        n16425) );
  AOI21_X1 U19623 ( .B1(n16645), .B2(n16426), .A(n16425), .ZN(n16429) );
  NAND2_X1 U19624 ( .A1(n16427), .A2(n16603), .ZN(n16428) );
  OAI211_X1 U19625 ( .C1(n16430), .C2(n16648), .A(n16429), .B(n16428), .ZN(
        P2_U3022) );
  NAND2_X1 U19626 ( .A1(n16431), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16444) );
  OAI21_X1 U19627 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16432), .ZN(n16434) );
  OAI21_X1 U19628 ( .B1(n16444), .B2(n16434), .A(n16433), .ZN(n16435) );
  AOI21_X1 U19629 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16447), .A(
        n16435), .ZN(n16436) );
  OAI21_X1 U19630 ( .B1(n16437), .B2(n16639), .A(n16436), .ZN(n16438) );
  AOI21_X1 U19631 ( .B1(n16645), .B2(n16439), .A(n16438), .ZN(n16442) );
  NAND3_X1 U19632 ( .A1(n16440), .A2(n16175), .A3(n19962), .ZN(n16441) );
  OAI211_X1 U19633 ( .C1(n16443), .C2(n19967), .A(n16442), .B(n16441), .ZN(
        P2_U3023) );
  NOR2_X1 U19634 ( .A1(n16444), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16445) );
  AOI211_X1 U19635 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n16447), .A(
        n16446), .B(n16445), .ZN(n16448) );
  OAI21_X1 U19636 ( .B1(n16449), .B2(n16639), .A(n16448), .ZN(n16450) );
  AOI21_X1 U19637 ( .B1(n16645), .B2(n16451), .A(n16450), .ZN(n16455) );
  NAND3_X1 U19638 ( .A1(n16453), .A2(n16603), .A3(n16452), .ZN(n16454) );
  OAI211_X1 U19639 ( .C1(n16456), .C2(n16648), .A(n16455), .B(n16454), .ZN(
        P2_U3024) );
  AOI21_X1 U19640 ( .B1(n16458), .B2(n16480), .A(n16545), .ZN(n16475) );
  OR3_X1 U19641 ( .A1(n16543), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n16458), .ZN(n16470) );
  AOI21_X1 U19642 ( .B1(n16475), .B2(n16470), .A(n16457), .ZN(n16465) );
  NOR4_X1 U19643 ( .A1(n16543), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n16458), .A4(n16474), .ZN(n16459) );
  AOI211_X1 U19644 ( .C1(n16461), .C2(n19952), .A(n16460), .B(n16459), .ZN(
        n16462) );
  OAI21_X1 U19645 ( .B1(n19959), .B2(n16463), .A(n16462), .ZN(n16464) );
  INV_X1 U19646 ( .A(n16467), .ZN(n16477) );
  INV_X1 U19647 ( .A(n16468), .ZN(n16469) );
  NAND2_X1 U19648 ( .A1(n16470), .A2(n16469), .ZN(n16472) );
  NOR2_X1 U19649 ( .A1(n19619), .A2(n19959), .ZN(n16471) );
  AOI211_X1 U19650 ( .C1(n19621), .C2(n19952), .A(n16472), .B(n16471), .ZN(
        n16473) );
  OAI21_X1 U19651 ( .B1(n16475), .B2(n16474), .A(n16473), .ZN(n16476) );
  AOI21_X1 U19652 ( .B1(n16477), .B2(n16603), .A(n16476), .ZN(n16478) );
  OAI21_X1 U19653 ( .B1(n16479), .B2(n16648), .A(n16478), .ZN(P2_U3027) );
  NAND2_X1 U19654 ( .A1(n16480), .A2(n16484), .ZN(n16482) );
  AOI21_X1 U19655 ( .B1(n16509), .B2(n16482), .A(n16481), .ZN(n16490) );
  INV_X1 U19656 ( .A(n16483), .ZN(n19637) );
  NOR3_X1 U19657 ( .A1(n16485), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n16484), .ZN(n16486) );
  AOI211_X1 U19658 ( .C1(n19637), .C2(n19952), .A(n16487), .B(n16486), .ZN(
        n16488) );
  OAI21_X1 U19659 ( .B1(n19959), .B2(n19635), .A(n16488), .ZN(n16489) );
  AOI211_X1 U19660 ( .C1(n16491), .C2(n16603), .A(n16490), .B(n16489), .ZN(
        n16492) );
  AOI22_X1 U19661 ( .A1(n16494), .A2(n16603), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16512), .ZN(n16505) );
  NAND2_X1 U19662 ( .A1(n16495), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16504) );
  AOI21_X1 U19663 ( .B1(n16497), .B2(n16496), .A(n14563), .ZN(n19803) );
  NAND2_X1 U19664 ( .A1(n19803), .A2(n16645), .ZN(n16498) );
  OAI211_X1 U19665 ( .C1(n16500), .C2(n16639), .A(n16499), .B(n16498), .ZN(
        n16501) );
  AOI21_X1 U19666 ( .B1(n16502), .B2(n19962), .A(n16501), .ZN(n16503) );
  OAI211_X1 U19667 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16505), .A(
        n16504), .B(n16503), .ZN(P2_U3030) );
  NAND3_X1 U19668 ( .A1(n16506), .A2(n16603), .A3(n16224), .ZN(n16514) );
  AOI21_X1 U19669 ( .B1(n19664), .B2(n19952), .A(n16507), .ZN(n16508) );
  OAI21_X1 U19670 ( .B1(n19959), .B2(n19665), .A(n16508), .ZN(n16511) );
  NOR2_X1 U19671 ( .A1(n16509), .A2(n14555), .ZN(n16510) );
  AOI211_X1 U19672 ( .C1(n16512), .C2(n14555), .A(n16511), .B(n16510), .ZN(
        n16513) );
  OAI211_X1 U19673 ( .C1(n16515), .C2(n16648), .A(n16514), .B(n16513), .ZN(
        P2_U3031) );
  INV_X1 U19674 ( .A(n16545), .ZN(n16516) );
  OAI21_X1 U19675 ( .B1(n16527), .B2(n16543), .A(n16516), .ZN(n16534) );
  NOR3_X1 U19676 ( .A1(n16543), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n16517), .ZN(n16521) );
  AOI21_X1 U19677 ( .B1(n19682), .B2(n19952), .A(n16518), .ZN(n16519) );
  OAI21_X1 U19678 ( .B1(n19959), .B2(n19680), .A(n16519), .ZN(n16520) );
  AOI211_X1 U19679 ( .C1(n16534), .C2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16521), .B(n16520), .ZN(n16524) );
  NAND2_X1 U19680 ( .A1(n16522), .A2(n19962), .ZN(n16523) );
  OAI211_X1 U19681 ( .C1(n16525), .C2(n19967), .A(n16524), .B(n16523), .ZN(
        P2_U3032) );
  NOR3_X1 U19682 ( .A1(n16543), .A2(n16527), .A3(n16526), .ZN(n16533) );
  NAND2_X1 U19683 ( .A1(n16528), .A2(n16645), .ZN(n16529) );
  OAI211_X1 U19684 ( .C1(n16531), .C2(n16639), .A(n16530), .B(n16529), .ZN(
        n16532) );
  AOI211_X1 U19685 ( .C1(n16534), .C2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n16533), .B(n16532), .ZN(n16535) );
  OAI211_X1 U19686 ( .C1(n16537), .C2(n16648), .A(n16536), .B(n16535), .ZN(
        P2_U3033) );
  NAND3_X1 U19687 ( .A1(n16539), .A2(n16603), .A3(n16538), .ZN(n16547) );
  AOI21_X1 U19688 ( .B1(n19697), .B2(n19952), .A(n16540), .ZN(n16542) );
  NAND2_X1 U19689 ( .A1(n19696), .A2(n16645), .ZN(n16541) );
  OAI211_X1 U19690 ( .C1(n16543), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16542), .B(n16541), .ZN(n16544) );
  AOI21_X1 U19691 ( .B1(n16545), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n16544), .ZN(n16546) );
  OAI211_X1 U19692 ( .C1(n16548), .C2(n16648), .A(n16547), .B(n16546), .ZN(
        P2_U3034) );
  NAND2_X1 U19693 ( .A1(n16562), .A2(n16549), .ZN(n16550) );
  NAND3_X1 U19694 ( .A1(n16578), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n16563), .ZN(n16569) );
  AOI21_X1 U19695 ( .B1(n16550), .B2(n16569), .A(n16551), .ZN(n16558) );
  NAND3_X1 U19696 ( .A1(n16578), .A2(n16552), .A3(n16551), .ZN(n16556) );
  INV_X1 U19697 ( .A(n16553), .ZN(n19710) );
  AOI21_X1 U19698 ( .B1(n19710), .B2(n19952), .A(n16554), .ZN(n16555) );
  OAI211_X1 U19699 ( .C1(n19959), .C2(n19707), .A(n16556), .B(n16555), .ZN(
        n16557) );
  AOI211_X1 U19700 ( .C1(n16559), .C2(n16603), .A(n16558), .B(n16557), .ZN(
        n16560) );
  OAI21_X1 U19701 ( .B1(n16561), .B2(n16648), .A(n16560), .ZN(P2_U3035) );
  INV_X1 U19702 ( .A(n16562), .ZN(n16564) );
  NOR3_X1 U19703 ( .A1(n16564), .A2(n16637), .A3(n16563), .ZN(n16572) );
  OAI21_X1 U19704 ( .B1(n16566), .B2(n16639), .A(n16565), .ZN(n16567) );
  INV_X1 U19705 ( .A(n16567), .ZN(n16568) );
  OAI211_X1 U19706 ( .C1(n19959), .C2(n16570), .A(n16569), .B(n16568), .ZN(
        n16571) );
  AOI211_X1 U19707 ( .C1(n16573), .C2(n16603), .A(n16572), .B(n16571), .ZN(
        n16574) );
  OAI21_X1 U19708 ( .B1(n16575), .B2(n16648), .A(n16574), .ZN(P2_U3036) );
  NOR2_X1 U19709 ( .A1(n16576), .A2(n16577), .ZN(n16585) );
  NAND2_X1 U19710 ( .A1(n16578), .A2(n16577), .ZN(n16582) );
  AOI21_X1 U19711 ( .B1(n16580), .B2(n19952), .A(n16579), .ZN(n16581) );
  OAI211_X1 U19712 ( .C1(n16583), .C2(n19959), .A(n16582), .B(n16581), .ZN(
        n16584) );
  AOI211_X1 U19713 ( .C1(n16586), .C2(n19962), .A(n16585), .B(n16584), .ZN(
        n16587) );
  OAI21_X1 U19714 ( .B1(n16588), .B2(n19967), .A(n16587), .ZN(P2_U3037) );
  INV_X1 U19715 ( .A(n16589), .ZN(n16623) );
  NAND2_X1 U19716 ( .A1(n16623), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16605) );
  AOI211_X1 U19717 ( .C1(n16593), .C2(n16611), .A(n16590), .B(n16605), .ZN(
        n16598) );
  OR2_X1 U19718 ( .A1(n16637), .A2(n16591), .ZN(n16617) );
  OAI21_X1 U19719 ( .B1(n16617), .B2(n16593), .A(n16592), .ZN(n16594) );
  AOI21_X1 U19720 ( .B1(n16595), .B2(n19952), .A(n16594), .ZN(n16596) );
  OAI21_X1 U19721 ( .B1(n19959), .B2(n19725), .A(n16596), .ZN(n16597) );
  AOI211_X1 U19722 ( .C1(n16599), .C2(n19962), .A(n16598), .B(n16597), .ZN(
        n16600) );
  OAI21_X1 U19723 ( .B1(n16601), .B2(n19967), .A(n16600), .ZN(P2_U3038) );
  NAND3_X1 U19724 ( .A1(n16604), .A2(n16603), .A3(n16602), .ZN(n16614) );
  INV_X1 U19725 ( .A(n16605), .ZN(n16612) );
  NOR2_X1 U19726 ( .A1(n16611), .A2(n16617), .ZN(n16606) );
  AOI211_X1 U19727 ( .C1(n16608), .C2(n19952), .A(n16607), .B(n16606), .ZN(
        n16609) );
  OAI21_X1 U19728 ( .B1(n19959), .B2(n19739), .A(n16609), .ZN(n16610) );
  AOI21_X1 U19729 ( .B1(n16612), .B2(n16611), .A(n16610), .ZN(n16613) );
  OAI211_X1 U19730 ( .C1(n16615), .C2(n16648), .A(n16614), .B(n16613), .ZN(
        P2_U3039) );
  OAI21_X1 U19731 ( .B1(n16617), .B2(n16624), .A(n16616), .ZN(n16618) );
  AOI21_X1 U19732 ( .B1(n19755), .B2(n19952), .A(n16618), .ZN(n16619) );
  OAI21_X1 U19733 ( .B1(n19959), .B2(n19752), .A(n16619), .ZN(n16622) );
  NOR2_X1 U19734 ( .A1(n16620), .A2(n16648), .ZN(n16621) );
  AOI211_X1 U19735 ( .C1(n16624), .C2(n16623), .A(n16622), .B(n16621), .ZN(
        n16625) );
  OAI21_X1 U19736 ( .B1(n19967), .B2(n16626), .A(n16625), .ZN(P2_U3040) );
  AND2_X1 U19737 ( .A1(n16628), .A2(n16627), .ZN(n16630) );
  XNOR2_X1 U19738 ( .A(n16630), .B(n16629), .ZN(n17293) );
  INV_X1 U19739 ( .A(n16635), .ZN(n16631) );
  NOR2_X1 U19740 ( .A1(n16632), .A2(n16631), .ZN(n17291) );
  AOI21_X1 U19741 ( .B1(n16635), .B2(n16634), .A(n16633), .ZN(n17290) );
  OR3_X1 U19742 ( .A1(n17291), .A2(n17290), .A3(n19967), .ZN(n16647) );
  INV_X1 U19743 ( .A(n16636), .ZN(n17307) );
  NOR2_X1 U19744 ( .A1(n16637), .A2(n17307), .ZN(n19957) );
  NAND2_X1 U19745 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n19957), .ZN(
        n16638) );
  OR2_X1 U19746 ( .A1(n19701), .A2(n19759), .ZN(n17287) );
  OAI211_X1 U19747 ( .C1(n19769), .C2(n16639), .A(n16638), .B(n17287), .ZN(
        n16643) );
  OAI211_X1 U19748 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n19955), .B(n16640), .ZN(n16641) );
  INV_X1 U19749 ( .A(n16641), .ZN(n16642) );
  AOI211_X1 U19750 ( .C1(n16645), .C2(n16644), .A(n16643), .B(n16642), .ZN(
        n16646) );
  OAI211_X1 U19751 ( .C1(n17293), .C2(n16648), .A(n16647), .B(n16646), .ZN(
        P2_U3041) );
  INV_X1 U19752 ( .A(n16649), .ZN(n16689) );
  NAND2_X1 U19753 ( .A1(n16650), .A2(n13118), .ZN(n16659) );
  MUX2_X1 U19754 ( .A(n16659), .B(n16694), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16651) );
  AOI21_X1 U19755 ( .B1(n16652), .B2(n16689), .A(n16651), .ZN(n16806) );
  MUX2_X1 U19756 ( .A(n16653), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .S(
        n19764), .Z(n16685) );
  OAI222_X1 U19757 ( .A1(n16836), .A2(n16654), .B1(n16705), .B2(n16806), .C1(
        n13787), .C2(n16685), .ZN(n16655) );
  MUX2_X1 U19758 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n16655), .S(
        n16707), .Z(P2_U3601) );
  NAND2_X1 U19759 ( .A1(n16694), .A2(n16656), .ZN(n16663) );
  INV_X1 U19760 ( .A(n16657), .ZN(n16658) );
  NAND2_X1 U19761 ( .A1(n16659), .A2(n16658), .ZN(n16662) );
  AOI21_X1 U19762 ( .B1(n16663), .B2(n16662), .A(n16661), .ZN(n16664) );
  AOI21_X1 U19763 ( .B1(n16665), .B2(n16689), .A(n16664), .ZN(n16807) );
  INV_X1 U19764 ( .A(n16807), .ZN(n16669) );
  NAND2_X1 U19765 ( .A1(n19764), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16666) );
  NAND2_X1 U19766 ( .A1(n16667), .A2(n16666), .ZN(n16684) );
  NOR2_X1 U19767 ( .A1(n16684), .A2(n13787), .ZN(n16668) );
  AOI22_X1 U19768 ( .A1(n16669), .A2(n20579), .B1(n16685), .B2(n16668), .ZN(
        n16670) );
  OAI21_X1 U19769 ( .B1(n19968), .B2(n16836), .A(n16670), .ZN(n16671) );
  MUX2_X1 U19770 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n16671), .S(
        n16707), .Z(P2_U3600) );
  NOR2_X1 U19771 ( .A1(n16661), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16690) );
  NAND2_X1 U19772 ( .A1(n16673), .A2(n16672), .ZN(n16675) );
  NAND2_X1 U19773 ( .A1(n16675), .A2(n16674), .ZN(n16697) );
  INV_X1 U19774 ( .A(n16676), .ZN(n16801) );
  OR2_X1 U19775 ( .A1(n16798), .A2(n16801), .ZN(n16691) );
  OAI21_X1 U19776 ( .B1(n16692), .B2(n16690), .A(n16691), .ZN(n16680) );
  INV_X1 U19777 ( .A(n16693), .ZN(n16677) );
  NAND2_X1 U19778 ( .A1(n16694), .A2(n16677), .ZN(n16699) );
  NOR2_X1 U19779 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16678) );
  OR2_X1 U19780 ( .A1(n16699), .A2(n16678), .ZN(n16679) );
  OAI211_X1 U19781 ( .C1(n16690), .C2(n16697), .A(n16680), .B(n16679), .ZN(
        n16681) );
  AOI21_X1 U19782 ( .B1(n19945), .B2(n16689), .A(n16681), .ZN(n16796) );
  INV_X1 U19783 ( .A(n16836), .ZN(n16682) );
  NAND2_X1 U19784 ( .A1(n16683), .A2(n16682), .ZN(n16687) );
  NAND3_X1 U19785 ( .A1(n16685), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n16684), 
        .ZN(n16686) );
  OAI211_X1 U19786 ( .C1(n16796), .C2(n16705), .A(n16687), .B(n16686), .ZN(
        n16688) );
  MUX2_X1 U19787 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n16688), .S(
        n16707), .Z(P2_U3599) );
  NAND2_X1 U19788 ( .A1(n15822), .A2(n16689), .ZN(n16704) );
  INV_X1 U19789 ( .A(n16690), .ZN(n16698) );
  NAND2_X1 U19790 ( .A1(n16691), .A2(n16698), .ZN(n16696) );
  AOI21_X1 U19791 ( .B1(n16694), .B2(n16693), .A(n16692), .ZN(n16695) );
  NAND2_X1 U19792 ( .A1(n16696), .A2(n16695), .ZN(n16701) );
  NAND3_X1 U19793 ( .A1(n16699), .A2(n16698), .A3(n16697), .ZN(n16700) );
  MUX2_X1 U19794 ( .A(n16701), .B(n16700), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n16702) );
  INV_X1 U19795 ( .A(n16702), .ZN(n16703) );
  NAND2_X1 U19796 ( .A1(n16704), .A2(n16703), .ZN(n16795) );
  INV_X1 U19797 ( .A(n16795), .ZN(n16706) );
  OAI22_X1 U19798 ( .A1(n20582), .A2(n16836), .B1(n16706), .B2(n16705), .ZN(
        n16708) );
  MUX2_X1 U19799 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16708), .S(
        n16707), .Z(P2_U3596) );
  AND3_X1 U19800 ( .A1(n16748), .A2(n20586), .A3(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16716) );
  INV_X1 U19801 ( .A(n20156), .ZN(n16711) );
  OAI21_X1 U19802 ( .B1(n16717), .B2(n20392), .A(n20581), .ZN(n16710) );
  NAND2_X1 U19803 ( .A1(n20582), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20576) );
  OAI21_X1 U19804 ( .B1(n20576), .B2(n16765), .A(n20382), .ZN(n16719) );
  NOR2_X1 U19805 ( .A1(n16719), .A2(n16716), .ZN(n16709) );
  INV_X1 U19806 ( .A(n20162), .ZN(n16712) );
  NAND2_X1 U19807 ( .A1(n16712), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n16724) );
  INV_X1 U19808 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18997) );
  OAI22_X2 U19809 ( .A1(n17344), .A2(n20007), .B1(n18997), .B2(n20005), .ZN(
        n20435) );
  NOR2_X2 U19810 ( .A1(n20004), .A2(n16815), .ZN(n20433) );
  AOI22_X1 U19811 ( .A1(n20435), .A2(n10453), .B1(n20156), .B2(n20433), .ZN(
        n16723) );
  INV_X1 U19812 ( .A(n16716), .ZN(n20114) );
  OAI21_X1 U19813 ( .B1(n16717), .B2(n20156), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16718) );
  NAND2_X1 U19814 ( .A1(n20397), .A2(n19797), .ZN(n20401) );
  NAND2_X1 U19815 ( .A1(n20158), .A2(n20434), .ZN(n16722) );
  INV_X1 U19816 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n17333) );
  OAI22_X2 U19817 ( .A1(n17333), .A2(n20007), .B1(n16026), .B2(n20005), .ZN(
        n20436) );
  NAND2_X1 U19818 ( .A1(n20436), .A2(n20157), .ZN(n16721) );
  NAND4_X1 U19819 ( .A1(n16724), .A2(n16723), .A3(n16722), .A4(n16721), .ZN(
        P2_U3088) );
  OAI21_X1 U19820 ( .B1(n10453), .B2(n20202), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16727) );
  NAND2_X1 U19821 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16725) );
  NOR2_X1 U19822 ( .A1(n16725), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20181) );
  AND2_X1 U19823 ( .A1(n20181), .A2(n20604), .ZN(n20173) );
  NOR2_X1 U19824 ( .A1(n20156), .A2(n20173), .ZN(n16730) );
  AOI211_X1 U19825 ( .C1(n16728), .C2(n20581), .A(n20382), .B(n20173), .ZN(
        n16726) );
  INV_X1 U19826 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19827 ( .A1(n10453), .A2(n20436), .B1(n20202), .B2(n20435), .ZN(
        n16732) );
  OAI21_X1 U19828 ( .B1(n16728), .B2(n20173), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16729) );
  AOI22_X1 U19829 ( .A1(n20174), .A2(n20434), .B1(n20173), .B2(n20433), .ZN(
        n16731) );
  OAI211_X1 U19830 ( .C1(n20177), .C2(n16733), .A(n16732), .B(n16731), .ZN(
        P2_U3096) );
  INV_X1 U19831 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16738) );
  INV_X1 U19832 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19021) );
  OAI22_X2 U19833 ( .A1(n16039), .A2(n20007), .B1(n19021), .B2(n20005), .ZN(
        n20422) );
  INV_X1 U19834 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n17326) );
  OAI22_X2 U19835 ( .A1(n17326), .A2(n20007), .B1(n14609), .B2(n20005), .ZN(
        n20421) );
  AOI22_X1 U19836 ( .A1(n20202), .A2(n20422), .B1(n10453), .B2(n20421), .ZN(
        n16737) );
  NAND2_X1 U19837 ( .A1(n20397), .A2(n16734), .ZN(n20425) );
  NOR2_X2 U19838 ( .A1(n20004), .A2(n16735), .ZN(n20420) );
  AOI22_X1 U19839 ( .A1(n20174), .A2(n20376), .B1(n20173), .B2(n20420), .ZN(
        n16736) );
  OAI211_X1 U19840 ( .C1(n20177), .C2(n16738), .A(n16737), .B(n16736), .ZN(
        P2_U3102) );
  INV_X1 U19841 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16743) );
  INV_X1 U19842 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n17335) );
  OAI22_X2 U19843 ( .A1(n17335), .A2(n20007), .B1(n16031), .B2(n20005), .ZN(
        n20474) );
  INV_X1 U19844 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17404) );
  OAI22_X2 U19845 ( .A1(n17324), .A2(n20007), .B1(n17404), .B2(n20005), .ZN(
        n20472) );
  AOI22_X1 U19846 ( .A1(n20202), .A2(n20474), .B1(n10453), .B2(n20472), .ZN(
        n16742) );
  NAND2_X1 U19847 ( .A1(n20397), .A2(n16739), .ZN(n20431) );
  NOR2_X2 U19848 ( .A1(n20004), .A2(n16740), .ZN(n20468) );
  AOI22_X1 U19849 ( .A1(n20174), .A2(n20470), .B1(n20173), .B2(n20468), .ZN(
        n16741) );
  OAI211_X1 U19850 ( .C1(n20177), .C2(n16743), .A(n16742), .B(n16741), .ZN(
        P2_U3103) );
  OAI21_X1 U19851 ( .B1(n20358), .B2(n20378), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n16754) );
  NOR2_X1 U19852 ( .A1(n16747), .A2(n20272), .ZN(n20117) );
  NAND2_X1 U19853 ( .A1(n20117), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16753) );
  AND2_X1 U19854 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16776) );
  AND2_X1 U19855 ( .A1(n16776), .A2(n16748), .ZN(n16766) );
  NAND2_X1 U19856 ( .A1(n16766), .A2(n20604), .ZN(n16749) );
  INV_X1 U19857 ( .A(n16749), .ZN(n20356) );
  AND2_X1 U19858 ( .A1(n16749), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16750) );
  NAND2_X1 U19859 ( .A1(n16751), .A2(n16750), .ZN(n16755) );
  OAI211_X1 U19860 ( .C1(n20356), .C2(n20581), .A(n16755), .B(n20397), .ZN(
        n16752) );
  INV_X1 U19861 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16760) );
  AOI22_X1 U19862 ( .A1(n20378), .A2(n20422), .B1(n20358), .B2(n20421), .ZN(
        n16759) );
  NAND3_X1 U19863 ( .A1(n20117), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n20581), .ZN(n16757) );
  INV_X1 U19864 ( .A(n16755), .ZN(n16756) );
  AOI22_X1 U19865 ( .A1(n20357), .A2(n20376), .B1(n20420), .B2(n20356), .ZN(
        n16758) );
  OAI211_X1 U19866 ( .C1(n20362), .C2(n16760), .A(n16759), .B(n16758), .ZN(
        P2_U3150) );
  INV_X1 U19867 ( .A(n16765), .ZN(n16761) );
  AOI21_X1 U19868 ( .B1(n20306), .B2(n16761), .A(n16766), .ZN(n16764) );
  AOI211_X1 U19869 ( .C1(n16767), .C2(n20581), .A(n20382), .B(n20387), .ZN(
        n16763) );
  NOR3_X2 U19870 ( .A1(n16764), .A2(n16763), .A3(n20183), .ZN(n20381) );
  INV_X1 U19871 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16772) );
  AOI22_X1 U19872 ( .A1(n20378), .A2(n20436), .B1(n20427), .B2(n20435), .ZN(
        n16771) );
  INV_X1 U19873 ( .A(n16766), .ZN(n16769) );
  OAI21_X1 U19874 ( .B1(n16767), .B2(n20387), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16768) );
  AOI22_X1 U19875 ( .A1(n20377), .A2(n20434), .B1(n20433), .B2(n20387), .ZN(
        n16770) );
  OAI211_X1 U19876 ( .C1(n20381), .C2(n16772), .A(n16771), .B(n16770), .ZN(
        P2_U3152) );
  INV_X1 U19877 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16775) );
  AOI22_X1 U19878 ( .A1(n20427), .A2(n20474), .B1(n20378), .B2(n20472), .ZN(
        n16774) );
  AOI22_X1 U19879 ( .A1(n20377), .A2(n20470), .B1(n20468), .B2(n20387), .ZN(
        n16773) );
  OAI211_X1 U19880 ( .C1(n20381), .C2(n16775), .A(n16774), .B(n16773), .ZN(
        P2_U3159) );
  INV_X1 U19881 ( .A(n20574), .ZN(n20577) );
  AND2_X1 U19882 ( .A1(n16776), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20389) );
  AOI21_X1 U19883 ( .B1(n20306), .B2(n20577), .A(n20389), .ZN(n16780) );
  INV_X1 U19884 ( .A(n19978), .ZN(n20469) );
  AND2_X1 U19885 ( .A1(n19978), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16777) );
  NAND2_X1 U19886 ( .A1(n16778), .A2(n16777), .ZN(n16781) );
  OAI211_X1 U19887 ( .C1(n20469), .C2(n20581), .A(n16781), .B(n20397), .ZN(
        n16779) );
  INV_X1 U19888 ( .A(n16781), .ZN(n16783) );
  AOI21_X1 U19889 ( .B1(n20389), .B2(n20581), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n16782) );
  NAND2_X1 U19890 ( .A1(n20397), .A2(n16784), .ZN(n20419) );
  NOR2_X2 U19891 ( .A1(n20004), .A2(n9575), .ZN(n20414) );
  INV_X1 U19892 ( .A(n20414), .ZN(n16786) );
  INV_X1 U19893 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n17328) );
  OAI22_X2 U19894 ( .A1(n17328), .A2(n20007), .B1(n12390), .B2(n20005), .ZN(
        n20415) );
  INV_X1 U19895 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n17338) );
  OAI22_X2 U19896 ( .A1(n17338), .A2(n20007), .B1(n16046), .B2(n20005), .ZN(
        n20416) );
  AOI22_X1 U19897 ( .A1(n20473), .A2(n20415), .B1(n20475), .B2(n20416), .ZN(
        n16785) );
  OAI21_X1 U19898 ( .B1(n16786), .B2(n19978), .A(n16785), .ZN(n16787) );
  AOI21_X1 U19899 ( .B1(n20471), .B2(n20373), .A(n16787), .ZN(n16788) );
  OAI21_X1 U19900 ( .B1(n20479), .B2(n16789), .A(n16788), .ZN(P2_U3173) );
  INV_X1 U19901 ( .A(n20420), .ZN(n16791) );
  AOI22_X1 U19902 ( .A1(n20475), .A2(n20422), .B1(n20473), .B2(n20421), .ZN(
        n16790) );
  OAI21_X1 U19903 ( .B1(n16791), .B2(n19978), .A(n16790), .ZN(n16792) );
  AOI21_X1 U19904 ( .B1(n20471), .B2(n20376), .A(n16792), .ZN(n16793) );
  OAI21_X1 U19905 ( .B1(n20479), .B2(n16794), .A(n16793), .ZN(P2_U3174) );
  MUX2_X1 U19906 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16795), .S(
        n16825), .Z(n16828) );
  MUX2_X1 U19907 ( .A(n16797), .B(n16796), .S(n16825), .Z(n16804) );
  INV_X1 U19908 ( .A(n16804), .ZN(n16827) );
  INV_X1 U19909 ( .A(n16798), .ZN(n16802) );
  NOR2_X1 U19910 ( .A1(P2_MORE_REG_SCAN_IN), .A2(P2_FLUSH_REG_SCAN_IN), .ZN(
        n16821) );
  INV_X1 U19911 ( .A(n16803), .ZN(n16818) );
  NOR2_X1 U19912 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16804), .ZN(
        n16813) );
  INV_X1 U19913 ( .A(n16828), .ZN(n16811) );
  OAI21_X1 U19914 ( .B1(n16813), .B2(n20594), .A(n16825), .ZN(n16805) );
  AOI21_X1 U19915 ( .B1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16807), .A(
        n16805), .ZN(n16809) );
  OAI211_X1 U19916 ( .C1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n16807), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n16806), .ZN(n16808) );
  OAI211_X1 U19917 ( .C1(n16828), .C2(n20586), .A(n16809), .B(n16808), .ZN(
        n16810) );
  OAI21_X1 U19918 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16811), .A(
        n16810), .ZN(n16812) );
  AOI21_X1 U19919 ( .B1(n16813), .B2(n20594), .A(n16812), .ZN(n16814) );
  OAI22_X1 U19920 ( .A1(n16816), .A2(n16815), .B1(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16814), .ZN(n16817) );
  AOI21_X1 U19921 ( .B1(n16819), .B2(n16818), .A(n16817), .ZN(n16820) );
  OAI21_X1 U19922 ( .B1(n16822), .B2(n16821), .A(n16820), .ZN(n16823) );
  NOR2_X1 U19923 ( .A1(n20607), .A2(n16823), .ZN(n16824) );
  OAI21_X1 U19924 ( .B1(n16825), .B2(n12127), .A(n16824), .ZN(n16826) );
  AOI21_X1 U19925 ( .B1(n16828), .B2(n16827), .A(n16826), .ZN(n16845) );
  AOI21_X1 U19926 ( .B1(n16845), .B2(n13787), .A(n9587), .ZN(n16833) );
  NOR2_X1 U19927 ( .A1(n16830), .A2(n20392), .ZN(n16831) );
  OAI21_X1 U19928 ( .B1(n13788), .B2(n16832), .A(n16831), .ZN(n16834) );
  OAI22_X1 U19929 ( .A1(n16836), .A2(n16835), .B1(n20480), .B2(n16834), .ZN(
        n16838) );
  MUX2_X1 U19930 ( .A(n20487), .B(n16838), .S(n9587), .Z(n16844) );
  INV_X1 U19931 ( .A(n16839), .ZN(n16841) );
  AOI211_X1 U19932 ( .C1(n20615), .C2(n16842), .A(n16841), .B(n16840), .ZN(
        n16843) );
  OAI211_X1 U19933 ( .C1(n16845), .C2(n20481), .A(n16844), .B(n16843), .ZN(
        P2_U3176) );
  INV_X1 U19934 ( .A(n16846), .ZN(n16847) );
  OAI21_X1 U19935 ( .B1(n20487), .B2(n20581), .A(n16847), .ZN(P2_U3593) );
  AND2_X1 U19936 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16851) );
  NAND2_X1 U19937 ( .A1(n18438), .A2(n17135), .ZN(n16848) );
  INV_X1 U19938 ( .A(n16850), .ZN(n16849) );
  AOI22_X1 U19939 ( .A1(n18450), .A2(n16851), .B1(n16849), .B2(n18565), .ZN(
        n17178) );
  OAI21_X1 U19940 ( .B1(n17178), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16855), .ZN(n16854) );
  OAI21_X1 U19941 ( .B1(n16873), .B2(n18565), .A(n16854), .ZN(n16861) );
  OAI211_X1 U19942 ( .C1(n16855), .C2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18565), .B(n16873), .ZN(n16857) );
  NAND3_X1 U19943 ( .A1(n16855), .A2(n18659), .A3(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16856) );
  NAND2_X1 U19944 ( .A1(n16857), .A2(n16856), .ZN(n16858) );
  NOR2_X1 U19945 ( .A1(n16873), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16940) );
  INV_X1 U19946 ( .A(n16940), .ZN(n16872) );
  NAND2_X1 U19947 ( .A1(n16858), .A2(n16872), .ZN(n16860) );
  AOI21_X1 U19948 ( .B1(n16861), .B2(n16860), .A(n16859), .ZN(n16959) );
  NAND2_X1 U19949 ( .A1(n17177), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16951) );
  NOR2_X1 U19950 ( .A1(n18843), .A2(n16951), .ZN(n16862) );
  XOR2_X1 U19951 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n16862), .Z(
        n16957) );
  NAND2_X1 U19952 ( .A1(n16863), .A2(n18432), .ZN(n17311) );
  INV_X1 U19953 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17457) );
  XOR2_X1 U19954 ( .A(n17457), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16866) );
  INV_X1 U19955 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19536) );
  OR2_X1 U19956 ( .A1(n18981), .A2(n19536), .ZN(n16947) );
  INV_X1 U19957 ( .A(n16947), .ZN(n16864) );
  AOI21_X1 U19958 ( .B1(n18529), .B2(n14217), .A(n16864), .ZN(n16865) );
  OAI21_X1 U19959 ( .B1(n17311), .B2(n16866), .A(n16865), .ZN(n16870) );
  NOR2_X1 U19960 ( .A1(n16868), .A2(n16867), .ZN(n17310) );
  NOR2_X1 U19961 ( .A1(n17310), .A2(n17457), .ZN(n16869) );
  AOI211_X1 U19962 ( .C1(n16957), .C2(n18647), .A(n16870), .B(n16869), .ZN(
        n16875) );
  NAND3_X1 U19963 ( .A1(n17315), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16873), .ZN(n16871) );
  OAI211_X1 U19964 ( .C1(n17315), .C2(n16873), .A(n16872), .B(n16871), .ZN(
        n16953) );
  NAND2_X1 U19965 ( .A1(n16953), .A2(n18645), .ZN(n16874) );
  INV_X1 U19966 ( .A(n16876), .ZN(n16877) );
  AOI21_X1 U19967 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n16878), .A(
        n16877), .ZN(n16989) );
  OR2_X1 U19968 ( .A1(n18904), .A2(n18727), .ZN(n16880) );
  NAND2_X1 U19969 ( .A1(n18645), .A2(n18901), .ZN(n16879) );
  NAND2_X2 U19970 ( .A1(n16880), .A2(n16879), .ZN(n18654) );
  NAND2_X2 U19971 ( .A1(n18810), .A2(n18654), .ZN(n18579) );
  NOR4_X1 U19972 ( .A1(n18478), .A2(n18737), .A3(n18743), .A4(n18579), .ZN(
        n16889) );
  OAI22_X1 U19973 ( .A1(n16979), .A2(n17314), .B1(n16978), .B2(n18727), .ZN(
        n18455) );
  NOR2_X1 U19974 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18495), .ZN(
        n18430) );
  NOR2_X1 U19975 ( .A1(n18529), .A2(n18430), .ZN(n16887) );
  INV_X1 U19976 ( .A(n16896), .ZN(n18459) );
  NOR2_X1 U19977 ( .A1(n16927), .A2(n18459), .ZN(n17444) );
  INV_X1 U19978 ( .A(n17444), .ZN(n16895) );
  NOR2_X1 U19979 ( .A1(n18465), .A2(n16895), .ZN(n16882) );
  NAND2_X1 U19980 ( .A1(n16881), .A2(n17444), .ZN(n17440) );
  OAI21_X1 U19981 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16882), .A(
        n17440), .ZN(n17441) );
  NAND2_X1 U19982 ( .A1(n18954), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n16985) );
  NOR3_X1 U19983 ( .A1(n19180), .A2(n18459), .A3(n18465), .ZN(n16885) );
  INV_X1 U19984 ( .A(n16882), .ZN(n17442) );
  NAND2_X1 U19985 ( .A1(n16883), .A2(n17442), .ZN(n16884) );
  OAI211_X1 U19986 ( .C1(n18431), .C2(n16928), .A(n18708), .B(n16884), .ZN(
        n18429) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n16885), .A(
        n18429), .ZN(n16886) );
  OAI211_X1 U19988 ( .C1(n16887), .C2(n17441), .A(n16985), .B(n16886), .ZN(
        n16888) );
  AOI221_X1 U19989 ( .B1(n16889), .B2(n10054), .C1(n18455), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n16888), .ZN(n16890) );
  OAI21_X1 U19990 ( .B1(n16989), .B2(n18653), .A(n16890), .ZN(P3_U2804) );
  INV_X1 U19991 ( .A(n16891), .ZN(n16892) );
  AOI21_X1 U19992 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16893), .A(
        n16892), .ZN(n17004) );
  NOR2_X1 U19993 ( .A1(n18844), .A2(n16894), .ZN(n18467) );
  NOR2_X1 U19994 ( .A1(n18843), .A2(n16894), .ZN(n16992) );
  OAI22_X1 U19995 ( .A1(n18467), .A2(n17314), .B1(n16992), .B2(n18727), .ZN(
        n18486) );
  NOR2_X1 U19996 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n16894), .ZN(
        n17001) );
  AOI22_X1 U19997 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18486), .B1(
        n18559), .B2(n17001), .ZN(n16900) );
  INV_X1 U19998 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n18460) );
  NOR2_X1 U19999 ( .A1(n18460), .A2(n16895), .ZN(n17443) );
  AOI21_X1 U20000 ( .B1(n18460), .B2(n16895), .A(n17443), .ZN(n17531) );
  NAND2_X1 U20001 ( .A1(n16896), .A2(n18432), .ZN(n16897) );
  NOR2_X1 U20002 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18495), .ZN(
        n18481) );
  NOR2_X1 U20003 ( .A1(n16927), .A2(n10441), .ZN(n17447) );
  NAND2_X1 U20004 ( .A1(n19351), .A2(n18459), .ZN(n18484) );
  OAI211_X1 U20005 ( .C1(n17447), .C2(n18608), .A(n18708), .B(n18484), .ZN(
        n18479) );
  NOR2_X1 U20006 ( .A1(n18481), .A2(n18479), .ZN(n18463) );
  NAND2_X1 U20007 ( .A1(n18954), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17002) );
  OAI221_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16897), .C1(
        n18460), .C2(n18463), .A(n17002), .ZN(n16898) );
  AOI21_X1 U20009 ( .B1(n18529), .B2(n17531), .A(n16898), .ZN(n16899) );
  OAI211_X1 U20010 ( .C1(n17004), .C2(n18653), .A(n16900), .B(n16899), .ZN(
        P3_U2806) );
  OAI21_X1 U20011 ( .B1(n16901), .B2(n16928), .A(n18708), .ZN(n16915) );
  NAND2_X1 U20012 ( .A1(n16901), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16903) );
  AOI211_X1 U20013 ( .C1(n17721), .C2(n16903), .A(n18637), .B(n19180), .ZN(
        n16905) );
  INV_X1 U20014 ( .A(n18495), .ZN(n16902) );
  OR2_X2 U20015 ( .A1(n18529), .A2(n16902), .ZN(n18714) );
  NOR2_X1 U20016 ( .A1(n16927), .A2(n16903), .ZN(n16912) );
  NAND2_X1 U20017 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16912), .ZN(
        n17646) );
  OAI21_X1 U20018 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16912), .A(
        n17646), .ZN(n17714) );
  OAI22_X1 U20019 ( .A1(n18720), .A2(n17714), .B1(n18981), .B2(n14261), .ZN(
        n16904) );
  AOI211_X1 U20020 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n16915), .A(
        n16905), .B(n16904), .ZN(n16909) );
  AOI22_X1 U20021 ( .A1(n18645), .A2(n16907), .B1(n16906), .B2(n18647), .ZN(
        n16908) );
  OAI211_X1 U20022 ( .C1(n18653), .C2(n16910), .A(n16909), .B(n16908), .ZN(
        P3_U2822) );
  NOR2_X1 U20023 ( .A1(n16927), .A2(n16911), .ZN(n17747) );
  NAND2_X1 U20024 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17747), .ZN(
        n17737) );
  AOI21_X1 U20025 ( .B1(n17713), .B2(n17737), .A(n16912), .ZN(n17730) );
  AOI22_X1 U20026 ( .A1(n18714), .A2(n17730), .B1(n16923), .B2(n16913), .ZN(
        n16917) );
  NOR3_X1 U20027 ( .A1(n19180), .A2(n16911), .A3(n18685), .ZN(n18636) );
  AOI221_X1 U20028 ( .B1(n18636), .B2(n17713), .C1(n16915), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n16914), .ZN(n16916) );
  OAI211_X1 U20029 ( .C1(n18727), .C2(n16918), .A(n16917), .B(n16916), .ZN(
        P3_U2823) );
  OR2_X1 U20030 ( .A1(n16920), .A2(n16919), .ZN(n16921) );
  AND2_X1 U20031 ( .A1(n16922), .A2(n16921), .ZN(n18950) );
  INV_X1 U20032 ( .A(n16923), .ZN(n18717) );
  OAI21_X1 U20033 ( .B1(n16926), .B2(n16925), .A(n16924), .ZN(n18957) );
  OAI22_X1 U20034 ( .A1(n18727), .A2(n18957), .B1(n18981), .B2(n19485), .ZN(
        n16930) );
  NAND2_X1 U20035 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18701), .ZN(
        n17748) );
  OAI21_X1 U20036 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17774), .A(
        n17748), .ZN(n17769) );
  INV_X1 U20037 ( .A(n16928), .ZN(n18606) );
  INV_X1 U20038 ( .A(n18708), .ZN(n18722) );
  OAI22_X1 U20039 ( .A1(n18720), .A2(n17769), .B1(n17761), .B2(n18712), .ZN(
        n16929) );
  AOI211_X1 U20040 ( .C1(n19351), .C2(n17767), .A(n16930), .B(n16929), .ZN(
        n16931) );
  OAI21_X1 U20041 ( .B1(n18950), .B2(n18717), .A(n16931), .ZN(P3_U2826) );
  OAI21_X1 U20042 ( .B1(n16936), .B2(n16933), .A(n16932), .ZN(n18970) );
  INV_X1 U20043 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19554) );
  OAI22_X1 U20044 ( .A1(n18717), .A2(n18970), .B1(n19554), .B2(n18981), .ZN(
        n16938) );
  AOI21_X1 U20045 ( .B1(n16936), .B2(n16935), .A(n16934), .ZN(n18972) );
  NOR2_X1 U20046 ( .A1(n18727), .A2(n18972), .ZN(n16937) );
  AOI211_X1 U20047 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18674), .A(
        n16938), .B(n16937), .ZN(n16939) );
  OAI21_X1 U20048 ( .B1(n18720), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n16939), .ZN(P3_U2829) );
  AOI21_X1 U20049 ( .B1(n17179), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n16940), .ZN(n16949) );
  AND2_X1 U20050 ( .A1(n18836), .A2(n18958), .ZN(n18977) );
  INV_X1 U20051 ( .A(n18977), .ZN(n18949) );
  INV_X1 U20052 ( .A(n18437), .ZN(n16942) );
  NAND4_X1 U20053 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n16944), .A4(n16941), .ZN(
        n18880) );
  NOR2_X1 U20054 ( .A1(n10159), .A2(n18880), .ZN(n16995) );
  AOI21_X1 U20055 ( .B1(n16942), .B2(n16995), .A(n18762), .ZN(n16982) );
  NAND3_X1 U20056 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n16944), .A3(
        n16943), .ZN(n18928) );
  NOR2_X1 U20057 ( .A1(n13334), .A2(n18928), .ZN(n18856) );
  NAND2_X1 U20058 ( .A1(n18810), .A2(n18856), .ZN(n18759) );
  NOR2_X1 U20059 ( .A1(n18437), .A2(n18759), .ZN(n16945) );
  OAI22_X1 U20060 ( .A1(n18926), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n18817), .B2(n16945), .ZN(n16946) );
  NOR4_X1 U20061 ( .A1(n18976), .A2(n16976), .A3(n16982), .A4(n16946), .ZN(
        n16965) );
  NOR2_X1 U20062 ( .A1(n16965), .A2(n18954), .ZN(n17131) );
  NAND2_X1 U20063 ( .A1(n17131), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16948) );
  OAI211_X1 U20064 ( .C1(n16949), .C2(n18949), .A(n16948), .B(n16947), .ZN(
        n16956) );
  INV_X1 U20065 ( .A(n18759), .ZN(n18756) );
  AOI22_X1 U20066 ( .A1(n19400), .A2(n16995), .B1(n16950), .B2(n18756), .ZN(
        n18738) );
  NOR3_X1 U20067 ( .A1(n18738), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16951), .ZN(n16952) );
  AOI21_X1 U20068 ( .B1(n16953), .B2(n18878), .A(n16952), .ZN(n16954) );
  NOR2_X1 U20069 ( .A1(n16954), .A2(n18888), .ZN(n16955) );
  AOI211_X1 U20070 ( .C1(n16957), .C2(n18870), .A(n16956), .B(n16955), .ZN(
        n16958) );
  OAI21_X1 U20071 ( .B1(n16959), .B2(n18913), .A(n16958), .ZN(P3_U2831) );
  NAND2_X1 U20072 ( .A1(n16960), .A2(n18446), .ZN(n18440) );
  XNOR2_X1 U20073 ( .A(n18565), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n18439) );
  INV_X1 U20074 ( .A(n16961), .ZN(n19406) );
  NOR4_X1 U20075 ( .A1(n18441), .A2(n18450), .A3(n18302), .A4(n19406), .ZN(
        n16967) );
  AOI22_X1 U20076 ( .A1(n19399), .A2(n16963), .B1(n18878), .B2(n16962), .ZN(
        n16964) );
  OAI211_X1 U20077 ( .C1(n18882), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16965), .B(n16964), .ZN(n16966) );
  OAI211_X1 U20078 ( .C1(n16967), .C2(n16966), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18981), .ZN(n16974) );
  NOR2_X1 U20079 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n13355), .ZN(
        n18443) );
  NAND2_X1 U20080 ( .A1(n18878), .A2(n18901), .ZN(n16969) );
  INV_X1 U20081 ( .A(n18904), .ZN(n18646) );
  NAND2_X1 U20082 ( .A1(n19399), .A2(n18646), .ZN(n16968) );
  OAI21_X1 U20083 ( .B1(n18808), .B2(n10159), .A(n18738), .ZN(n18771) );
  NAND2_X1 U20084 ( .A1(n18958), .A2(n18771), .ZN(n17185) );
  NOR2_X1 U20085 ( .A1(n18437), .A2(n17185), .ZN(n18730) );
  INV_X1 U20086 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19531) );
  NOR2_X1 U20087 ( .A1(n18981), .A2(n19531), .ZN(n18435) );
  NOR3_X1 U20088 ( .A1(n18446), .A2(n18439), .A3(n18913), .ZN(n16970) );
  AOI211_X1 U20089 ( .C1(n18443), .C2(n18730), .A(n18435), .B(n16970), .ZN(
        n16973) );
  INV_X1 U20090 ( .A(n18971), .ZN(n16971) );
  NAND3_X1 U20091 ( .A1(n18450), .A2(n16971), .A3(n18438), .ZN(n16972) );
  NAND3_X1 U20092 ( .A1(n16974), .A2(n16973), .A3(n16972), .ZN(P3_U2834) );
  OR2_X1 U20093 ( .A1(n18737), .A2(n18743), .ZN(n16975) );
  INV_X1 U20094 ( .A(n18478), .ZN(n16990) );
  NAND2_X1 U20095 ( .A1(n16990), .A2(n18771), .ZN(n18751) );
  NOR2_X1 U20096 ( .A1(n16975), .A2(n18751), .ZN(n16984) );
  NOR2_X1 U20097 ( .A1(n16976), .A2(n18759), .ZN(n18811) );
  AOI21_X1 U20098 ( .B1(n18741), .B2(n18811), .A(n18817), .ZN(n18736) );
  OAI22_X1 U20099 ( .A1(n18927), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18926), .B2(n16977), .ZN(n16981) );
  OAI22_X1 U20100 ( .A1(n16979), .A2(n18902), .B1(n16978), .B2(n16991), .ZN(
        n16980) );
  INV_X1 U20101 ( .A(n18728), .ZN(n16983) );
  MUX2_X1 U20102 ( .A(n16984), .B(n16983), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n16987) );
  OAI21_X1 U20103 ( .B1(n10054), .B2(n18969), .A(n16985), .ZN(n16986) );
  AOI21_X1 U20104 ( .B1(n16987), .B2(n18958), .A(n16986), .ZN(n16988) );
  OAI21_X1 U20105 ( .B1(n16989), .B2(n18913), .A(n16988), .ZN(P3_U2836) );
  INV_X1 U20106 ( .A(n17185), .ZN(n18779) );
  AOI21_X1 U20107 ( .B1(n16990), .B2(n18811), .A(n18817), .ZN(n16994) );
  OAI22_X1 U20108 ( .A1(n18467), .A2(n18902), .B1(n16992), .B2(n16991), .ZN(
        n16993) );
  NOR3_X1 U20109 ( .A1(n18976), .A2(n16994), .A3(n16993), .ZN(n16998) );
  NAND2_X1 U20110 ( .A1(n18813), .A2(n16995), .ZN(n18816) );
  NOR2_X1 U20111 ( .A1(n18818), .A2(n18816), .ZN(n18763) );
  AOI21_X1 U20112 ( .B1(n16996), .B2(n18763), .A(n18762), .ZN(n18735) );
  NOR2_X1 U20113 ( .A1(n18735), .A2(n18750), .ZN(n16997) );
  AOI21_X1 U20114 ( .B1(n16998), .B2(n16997), .A(n18954), .ZN(n18753) );
  AOI21_X1 U20115 ( .B1(n16999), .B2(n16998), .A(n9886), .ZN(n17000) );
  AOI22_X1 U20116 ( .A1(n18779), .A2(n17001), .B1(n18753), .B2(n17000), .ZN(
        n17003) );
  OAI211_X1 U20117 ( .C1(n17004), .C2(n18913), .A(n17003), .B(n17002), .ZN(
        P3_U2838) );
  NAND3_X1 U20118 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n18168) );
  NOR2_X1 U20119 ( .A1(n17787), .A2(n18168), .ZN(n18159) );
  NOR2_X2 U20120 ( .A1(n18155), .A2(n17754), .ZN(n18158) );
  INV_X1 U20121 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17633) );
  INV_X1 U20122 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17973) );
  NAND2_X1 U20123 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17941), .ZN(n17927) );
  NAND3_X1 U20124 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .ZN(n17823) );
  NAND2_X1 U20125 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .ZN(n17822) );
  INV_X1 U20126 ( .A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20127 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18081), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17009) );
  NAND2_X1 U20128 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n17008) );
  OAI211_X1 U20129 ( .C1(n17010), .C2(n10442), .A(n17009), .B(n17008), .ZN(
        n17011) );
  INV_X1 U20130 ( .A(n17011), .ZN(n17014) );
  AOI22_X1 U20131 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20132 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17012) );
  NAND3_X1 U20133 ( .A1(n17014), .A2(n17013), .A3(n17012), .ZN(n17020) );
  AOI22_X1 U20134 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20135 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20136 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20137 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17015) );
  NAND4_X1 U20138 ( .A1(n17018), .A2(n17017), .A3(n17016), .A4(n17015), .ZN(
        n17019) );
  OR2_X1 U20139 ( .A1(n17020), .A2(n17019), .ZN(n17867) );
  INV_X1 U20140 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20141 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17022) );
  NAND2_X1 U20142 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n17021) );
  OAI211_X1 U20143 ( .C1(n17023), .C2(n18086), .A(n17022), .B(n17021), .ZN(
        n17024) );
  INV_X1 U20144 ( .A(n17024), .ZN(n17027) );
  AOI22_X1 U20145 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20146 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17025) );
  NAND3_X1 U20147 ( .A1(n17027), .A2(n17026), .A3(n17025), .ZN(n17033) );
  AOI22_X1 U20148 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20149 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20150 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20151 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U20152 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17032) );
  NOR2_X1 U20153 ( .A1(n17033), .A2(n17032), .ZN(n17878) );
  INV_X1 U20154 ( .A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n18137) );
  OAI22_X1 U20155 ( .A1(n10448), .A2(n17993), .B1(n17045), .B2(n18137), .ZN(
        n17034) );
  AOI21_X1 U20156 ( .B1(n13168), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17034), .ZN(n17038) );
  AOI22_X1 U20157 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20158 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17036) );
  NAND2_X1 U20159 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n17035) );
  NAND4_X1 U20160 ( .A1(n17038), .A2(n17037), .A3(n17036), .A4(n17035), .ZN(
        n17044) );
  AOI22_X1 U20161 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17897), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20162 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20163 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20164 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17039) );
  NAND4_X1 U20165 ( .A1(n17042), .A2(n17041), .A3(n17040), .A4(n17039), .ZN(
        n17043) );
  NOR2_X1 U20166 ( .A1(n17044), .A2(n17043), .ZN(n17888) );
  INV_X1 U20167 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n18016) );
  OAI22_X1 U20168 ( .A1(n17087), .A2(n18016), .B1(n17045), .B2(n18014), .ZN(
        n17046) );
  AOI21_X1 U20169 ( .B1(n18091), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n17046), .ZN(n17050) );
  AOI22_X1 U20170 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20171 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17048) );
  NAND2_X1 U20172 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n17047) );
  NAND4_X1 U20173 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17056) );
  AOI22_X1 U20174 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9573), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17054) );
  AOI22_X1 U20175 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20176 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20177 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17051) );
  NAND4_X1 U20178 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17055) );
  NOR2_X1 U20179 ( .A1(n17056), .A2(n17055), .ZN(n17887) );
  NOR2_X1 U20180 ( .A1(n17888), .A2(n17887), .ZN(n17883) );
  AOI22_X1 U20181 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20182 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17060) );
  AOI22_X1 U20183 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17059) );
  AOI22_X1 U20184 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17058) );
  NAND4_X1 U20185 ( .A1(n17061), .A2(n17060), .A3(n17059), .A4(n17058), .ZN(
        n17071) );
  INV_X1 U20186 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U20187 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17063) );
  NAND2_X1 U20188 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n17062) );
  OAI211_X1 U20189 ( .C1(n18172), .C2(n18135), .A(n17063), .B(n17062), .ZN(
        n17070) );
  INV_X1 U20190 ( .A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17065) );
  INV_X1 U20191 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17064) );
  OAI22_X1 U20192 ( .A1(n18067), .A2(n17065), .B1(n18138), .B2(n17064), .ZN(
        n17069) );
  INV_X1 U20193 ( .A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17067) );
  INV_X1 U20194 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17066) );
  OAI22_X1 U20195 ( .A1(n17112), .A2(n17067), .B1(n18141), .B2(n17066), .ZN(
        n17068) );
  OR4_X1 U20196 ( .A1(n17071), .A2(n17070), .A3(n17069), .A4(n17068), .ZN(
        n17882) );
  NAND2_X1 U20197 ( .A1(n17883), .A2(n17882), .ZN(n17881) );
  NOR2_X1 U20198 ( .A1(n17878), .A2(n17881), .ZN(n17875) );
  AOI22_X1 U20199 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17075) );
  AOI22_X1 U20200 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20201 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20202 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17072) );
  NAND4_X1 U20203 ( .A1(n17075), .A2(n17074), .A3(n17073), .A4(n17072), .ZN(
        n17086) );
  INV_X1 U20204 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20205 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17077) );
  NAND2_X1 U20206 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n17076) );
  OAI211_X1 U20207 ( .C1(n17078), .C2(n18086), .A(n17077), .B(n17076), .ZN(
        n17085) );
  INV_X1 U20208 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17080) );
  INV_X1 U20209 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17079) );
  OAI22_X1 U20210 ( .A1(n18067), .A2(n17080), .B1(n18138), .B2(n17079), .ZN(
        n17084) );
  OAI22_X1 U20211 ( .A1(n17112), .A2(n17082), .B1(n18141), .B2(n17081), .ZN(
        n17083) );
  NAND2_X1 U20212 ( .A1(n17875), .A2(n17874), .ZN(n17873) );
  INV_X1 U20213 ( .A(n17873), .ZN(n17868) );
  NAND2_X1 U20214 ( .A1(n17867), .A2(n17868), .ZN(n17866) );
  INV_X1 U20215 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17920) );
  OAI22_X1 U20216 ( .A1(n10448), .A2(n17917), .B1(n17087), .B2(n17920), .ZN(
        n17088) );
  AOI21_X1 U20217 ( .B1(n18080), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n17088), .ZN(n17093) );
  AOI22_X1 U20218 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20219 ( .A1(n17089), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17091) );
  NAND2_X1 U20220 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n17090) );
  NAND4_X1 U20221 ( .A1(n17093), .A2(n17092), .A3(n17091), .A4(n17090), .ZN(
        n17099) );
  AOI22_X1 U20222 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20223 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20224 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20225 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17094) );
  NAND4_X1 U20226 ( .A1(n17097), .A2(n17096), .A3(n17095), .A4(n17094), .ZN(
        n17098) );
  NOR2_X1 U20227 ( .A1(n17099), .A2(n17098), .ZN(n17861) );
  XNOR2_X1 U20228 ( .A(n17866), .B(n17861), .ZN(n18201) );
  NAND3_X1 U20229 ( .A1(n9632), .A2(P3_EBX_REG_28__SCAN_IN), .A3(n18163), .ZN(
        n17100) );
  OAI221_X1 U20230 ( .B1(n9632), .B2(P3_EBX_REG_28__SCAN_IN), .C1(n18171), 
        .C2(n18201), .A(n17100), .ZN(P3_U2675) );
  NAND2_X1 U20231 ( .A1(n18163), .A2(n17117), .ZN(n18063) );
  AOI22_X1 U20232 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20233 ( .A1(n13178), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20234 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13200), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20235 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17101) );
  NAND4_X1 U20236 ( .A1(n17104), .A2(n17103), .A3(n17102), .A4(n17101), .ZN(
        n17116) );
  AOI22_X1 U20237 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18081), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17106) );
  NAND2_X1 U20238 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n17105) );
  OAI211_X1 U20239 ( .C1(n18156), .C2(n18086), .A(n17106), .B(n17105), .ZN(
        n17115) );
  INV_X1 U20240 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17108) );
  OAI22_X1 U20241 ( .A1(n18067), .A2(n17108), .B1(n18138), .B2(n17107), .ZN(
        n17114) );
  OAI22_X1 U20242 ( .A1(n17112), .A2(n17111), .B1(n18141), .B2(n17110), .ZN(
        n17113) );
  OR4_X1 U20243 ( .A1(n17116), .A2(n17115), .A3(n17114), .A4(n17113), .ZN(
        n18275) );
  NOR2_X1 U20244 ( .A1(n19024), .A2(n17117), .ZN(n18048) );
  AOI22_X1 U20245 ( .A1(n18177), .A2(n18275), .B1(n18048), .B2(n17653), .ZN(
        n17118) );
  OAI21_X1 U20246 ( .B1(n17653), .B2(n18063), .A(n17118), .ZN(P3_U2690) );
  NOR2_X1 U20247 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19552), .ZN(
        n19031) );
  NOR2_X1 U20248 ( .A1(n17119), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n17126) );
  AND2_X1 U20249 ( .A1(n10442), .A2(n17126), .ZN(n18982) );
  AOI21_X1 U20250 ( .B1(n18982), .B2(n17424), .A(n19551), .ZN(n17120) );
  NOR2_X1 U20251 ( .A1(n19323), .A2(n17120), .ZN(n18986) );
  NOR2_X1 U20252 ( .A1(n19031), .A2(n18986), .ZN(n17122) );
  INV_X1 U20253 ( .A(n19271), .ZN(n19320) );
  INV_X1 U20254 ( .A(n18986), .ZN(n18990) );
  OAI22_X1 U20255 ( .A1(n19567), .A2(n18606), .B1(n13509), .B2(n19552), .ZN(
        n17125) );
  NAND3_X1 U20256 ( .A1(n13491), .A2(n18990), .A3(n17125), .ZN(n17121) );
  OAI221_X1 U20257 ( .B1(n13491), .B2(n17122), .C1(n13491), .C2(n19320), .A(
        n17121), .ZN(P3_U2864) );
  NAND2_X1 U20258 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19158) );
  NOR2_X1 U20259 ( .A1(n19567), .A2(n18606), .ZN(n17124) );
  INV_X1 U20260 ( .A(n17122), .ZN(n17123) );
  AOI221_X1 U20261 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n19158), .C1(n17124), 
        .C2(n19158), .A(n17123), .ZN(n18989) );
  OAI221_X1 U20262 ( .B1(n19271), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n19271), .C2(n17125), .A(n18990), .ZN(n18987) );
  AOI22_X1 U20263 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18989), .B1(
        n18987), .B2(n19430), .ZN(P3_U2865) );
  NOR2_X1 U20264 ( .A1(n17127), .A2(n17126), .ZN(n19439) );
  NAND3_X1 U20265 ( .A1(n17129), .A2(n19584), .A3(n19439), .ZN(n17128) );
  OAI21_X1 U20266 ( .B1(n17129), .B2(n19410), .A(n17128), .ZN(P3_U3284) );
  NOR3_X1 U20267 ( .A1(n17315), .A2(n17130), .A3(n18971), .ZN(n17132) );
  AOI211_X1 U20268 ( .C1(n18870), .C2(n17133), .A(n17132), .B(n17131), .ZN(
        n17182) );
  OAI221_X1 U20269 ( .B1(n18949), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n18949), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17182), .ZN(
        n17134) );
  AOI22_X1 U20270 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17134), .B1(
        n18954), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n17138) );
  NAND3_X1 U20271 ( .A1(n17136), .A2(n18730), .A3(n17135), .ZN(n17137) );
  OAI211_X1 U20272 ( .C1(n17139), .C2(n18913), .A(n17138), .B(n17137), .ZN(
        P3_U2833) );
  AOI21_X1 U20273 ( .B1(n17140), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n21264), .ZN(n17141) );
  AND2_X1 U20274 ( .A1(n17142), .A2(n17141), .ZN(n17146) );
  NAND2_X1 U20275 ( .A1(n17144), .A2(n17143), .ZN(n17145) );
  OAI21_X1 U20276 ( .B1(n17146), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n17145), .ZN(n17148) );
  NAND2_X1 U20277 ( .A1(n17146), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n17147) );
  AND2_X1 U20278 ( .A1(n17148), .A2(n17147), .ZN(n17150) );
  INV_X1 U20279 ( .A(n17150), .ZN(n17152) );
  OAI21_X1 U20280 ( .B1(n17150), .B2(n21143), .A(n17149), .ZN(n17151) );
  OAI21_X1 U20281 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n17152), .A(
        n17151), .ZN(n17153) );
  AOI222_X1 U20282 ( .A1(n21184), .A2(n17154), .B1(n21184), .B2(n17153), .C1(
        n17154), .C2(n17153), .ZN(n17164) );
  INV_X1 U20283 ( .A(n17155), .ZN(n17160) );
  AOI21_X1 U20284 ( .B1(n21646), .B2(n17157), .A(n17156), .ZN(n17159) );
  NOR4_X1 U20285 ( .A1(n17161), .A2(n17160), .A3(n17159), .A4(n17158), .ZN(
        n17162) );
  OAI211_X1 U20286 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n17164), .A(
        n17163), .B(n17162), .ZN(n17169) );
  NOR3_X1 U20287 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n11005), .A3(n21419), 
        .ZN(n17167) );
  OAI22_X1 U20288 ( .A1(n17170), .A2(n17167), .B1(n17166), .B2(n17165), .ZN(
        n17279) );
  AOI221_X1 U20289 ( .B1(n10276), .B2(n21403), .C1(n17169), .C2(n21403), .A(
        n17279), .ZN(n17171) );
  NOR2_X1 U20290 ( .A1(n17171), .A2(n10276), .ZN(n17286) );
  OAI21_X1 U20291 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21419), .A(n17286), 
        .ZN(n17284) );
  AOI211_X1 U20292 ( .C1(n17170), .C2(n17169), .A(n17168), .B(n17284), .ZN(
        n17176) );
  AOI21_X1 U20293 ( .B1(n17173), .B2(n17172), .A(n17171), .ZN(n17174) );
  INV_X1 U20294 ( .A(n17174), .ZN(n17175) );
  AOI22_X1 U20295 ( .A1(n17176), .A2(n17281), .B1(n10276), .B2(n17175), .ZN(
        P1_U3161) );
  INV_X1 U20296 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n17180) );
  NAND2_X1 U20297 ( .A1(n17177), .A2(n17180), .ZN(n17320) );
  XNOR2_X1 U20298 ( .A(n17178), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n17317) );
  NAND2_X1 U20299 ( .A1(n18977), .A2(n17179), .ZN(n17181) );
  AOI21_X1 U20300 ( .B1(n17182), .B2(n17181), .A(n17180), .ZN(n17183) );
  AOI21_X1 U20301 ( .B1(n17317), .B2(n18936), .A(n17183), .ZN(n17184) );
  NAND2_X1 U20302 ( .A1(n18954), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n17309) );
  OAI211_X1 U20303 ( .C1(n17185), .C2(n17320), .A(n17184), .B(n17309), .ZN(
        P3_U2832) );
  INV_X1 U20304 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21421) );
  NOR2_X1 U20305 ( .A1(n21415), .A2(n21421), .ZN(n21417) );
  INV_X1 U20306 ( .A(n21417), .ZN(n17188) );
  INV_X1 U20307 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20621) );
  NOR2_X1 U20308 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20621), .ZN(n21418) );
  NOR2_X1 U20309 ( .A1(n20621), .A2(n21419), .ZN(n21414) );
  AOI211_X1 U20310 ( .C1(HOLD), .C2(n21418), .A(n17186), .B(n21414), .ZN(
        n17187) );
  OAI221_X1 U20311 ( .B1(n17188), .B2(HOLD), .C1(n17188), .C2(
        P1_STATE_REG_2__SCAN_IN), .A(n17187), .ZN(P1_U3195) );
  AND2_X1 U20312 ( .A1(n20737), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U20313 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U20314 ( .A1(n17189), .A2(n20602), .ZN(P2_U3047) );
  INV_X1 U20315 ( .A(n17190), .ZN(n17199) );
  OAI21_X1 U20316 ( .B1(n20646), .B2(n17191), .A(n20688), .ZN(n17192) );
  AOI21_X1 U20317 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(n20685), .A(n17192), .ZN(
        n17193) );
  OAI21_X1 U20318 ( .B1(n17212), .B2(n21447), .A(n17193), .ZN(n17194) );
  AOI21_X1 U20319 ( .B1(n17195), .B2(n20705), .A(n17194), .ZN(n17196) );
  OAI21_X1 U20320 ( .B1(n20691), .B2(n17197), .A(n17196), .ZN(n17198) );
  AOI21_X1 U20321 ( .B1(n17199), .B2(n13732), .A(n17198), .ZN(n17200) );
  OAI21_X1 U20322 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n17201), .A(n17200), 
        .ZN(P1_U2825) );
  AOI21_X1 U20323 ( .B1(n17202), .B2(n20652), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n17211) );
  AOI21_X1 U20324 ( .B1(n20698), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20662), .ZN(n17203) );
  OAI21_X1 U20325 ( .B1(n17214), .B2(n17204), .A(n17203), .ZN(n17205) );
  AOI21_X1 U20326 ( .B1(n17206), .B2(n20705), .A(n17205), .ZN(n17210) );
  INV_X1 U20327 ( .A(n17207), .ZN(n17208) );
  AOI22_X1 U20328 ( .A1(n17228), .A2(n13732), .B1(n17208), .B2(n20709), .ZN(
        n17209) );
  OAI211_X1 U20329 ( .C1(n17212), .C2(n17211), .A(n17210), .B(n17209), .ZN(
        P1_U2826) );
  OAI21_X1 U20330 ( .B1(n20646), .B2(n11138), .A(n20688), .ZN(n17217) );
  OAI22_X1 U20331 ( .A1(n17215), .A2(n17214), .B1(n20650), .B2(n17213), .ZN(
        n17216) );
  AOI211_X1 U20332 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n17218), .A(n17217), 
        .B(n17216), .ZN(n17222) );
  AOI22_X1 U20333 ( .A1(n17220), .A2(n13732), .B1(n17219), .B2(n15336), .ZN(
        n17221) );
  OAI211_X1 U20334 ( .C1(n17223), .C2(n20691), .A(n17222), .B(n17221), .ZN(
        P1_U2829) );
  INV_X1 U20335 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21625) );
  INV_X1 U20336 ( .A(n17224), .ZN(n20756) );
  INV_X1 U20337 ( .A(n17225), .ZN(n17226) );
  AOI22_X1 U20338 ( .A1(n17228), .A2(n17227), .B1(n20756), .B2(n17226), .ZN(
        n17229) );
  OAI21_X1 U20339 ( .B1(n21625), .B2(n17230), .A(n17229), .ZN(P1_U2890) );
  AOI22_X1 U20340 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20786), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n17236) );
  NAND2_X1 U20341 ( .A1(n17232), .A2(n17231), .ZN(n17233) );
  XNOR2_X1 U20342 ( .A(n17234), .B(n17233), .ZN(n17261) );
  AOI22_X1 U20343 ( .A1(n17261), .A2(n20780), .B1(n20779), .B2(n20668), .ZN(
        n17235) );
  OAI211_X1 U20344 ( .C1(n20784), .C2(n20666), .A(n17236), .B(n17235), .ZN(
        P1_U2992) );
  AOI22_X1 U20345 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20786), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n17243) );
  XNOR2_X1 U20346 ( .A(n17238), .B(n17237), .ZN(n17239) );
  XNOR2_X1 U20347 ( .A(n17240), .B(n17239), .ZN(n17267) );
  AOI22_X1 U20348 ( .A1(n17241), .A2(n20779), .B1(n17267), .B2(n20780), .ZN(
        n17242) );
  OAI211_X1 U20349 ( .C1(n20784), .C2(n20683), .A(n17243), .B(n17242), .ZN(
        P1_U2993) );
  AOI22_X1 U20350 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20786), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n17249) );
  OAI22_X1 U20351 ( .A1(n17246), .A2(n20631), .B1(n17245), .B2(n17244), .ZN(
        n17247) );
  INV_X1 U20352 ( .A(n17247), .ZN(n17248) );
  OAI211_X1 U20353 ( .C1(n20784), .C2(n17250), .A(n17249), .B(n17248), .ZN(
        P1_U2994) );
  NAND2_X1 U20354 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17266), .ZN(
        n17264) );
  AOI22_X1 U20355 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17251), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n11592), .ZN(n17259) );
  INV_X1 U20356 ( .A(n17252), .ZN(n17254) );
  AOI21_X1 U20357 ( .B1(n17254), .B2(n20801), .A(n17253), .ZN(n17258) );
  OAI21_X1 U20358 ( .B1(n17255), .B2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17270), .ZN(n17260) );
  AOI22_X1 U20359 ( .A1(n17256), .A2(n20795), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17260), .ZN(n17257) );
  OAI211_X1 U20360 ( .C1(n17264), .C2(n17259), .A(n17258), .B(n17257), .ZN(
        P1_U3023) );
  AOI22_X1 U20361 ( .A1(n20801), .A2(n20663), .B1(n20786), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n17263) );
  AOI22_X1 U20362 ( .A1(n17261), .A2(n20795), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17260), .ZN(n17262) );
  OAI211_X1 U20363 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n17264), .A(
        n17263), .B(n17262), .ZN(P1_U3024) );
  INV_X1 U20364 ( .A(n17265), .ZN(n20674) );
  AOI22_X1 U20365 ( .A1(n20801), .A2(n20674), .B1(n20786), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20366 ( .A1(n17267), .A2(n20795), .B1(n17237), .B2(n17266), .ZN(
        n17268) );
  OAI211_X1 U20367 ( .C1(n17270), .C2(n17237), .A(n17269), .B(n17268), .ZN(
        P1_U3025) );
  OR4_X1 U20368 ( .A1(n17273), .A2(n20690), .A3(n17272), .A4(n17271), .ZN(
        n17274) );
  OAI21_X1 U20369 ( .B1(n17276), .B2(n17275), .A(n17274), .ZN(P1_U3468) );
  NAND4_X1 U20370 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n11005), .A4(n21419), .ZN(n17277) );
  NAND2_X1 U20371 ( .A1(n17278), .A2(n17277), .ZN(n21404) );
  OAI21_X1 U20372 ( .B1(n21404), .B2(n17280), .A(n17279), .ZN(n17282) );
  NAND2_X1 U20373 ( .A1(n17282), .A2(n17281), .ZN(n17283) );
  AOI21_X1 U20374 ( .B1(n21403), .B2(n17284), .A(n17283), .ZN(P1_U3162) );
  OAI21_X1 U20375 ( .B1(n17286), .B2(n21222), .A(n17285), .ZN(P1_U3466) );
  INV_X1 U20376 ( .A(n17287), .ZN(n17288) );
  AOI21_X1 U20377 ( .B1(n17289), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n17288), .ZN(n17297) );
  NOR3_X1 U20378 ( .A1(n17291), .A2(n17290), .A3(n19941), .ZN(n17295) );
  OAI22_X1 U20379 ( .A1(n17293), .A2(n17292), .B1(n19928), .B2(n19769), .ZN(
        n17294) );
  NOR2_X1 U20380 ( .A1(n17295), .A2(n17294), .ZN(n17296) );
  OAI211_X1 U20381 ( .C1(n19939), .C2(n19766), .A(n17297), .B(n17296), .ZN(
        P2_U3009) );
  OAI21_X1 U20382 ( .B1(n19959), .B2(n20580), .A(n17298), .ZN(n17299) );
  AOI21_X1 U20383 ( .B1(n15822), .B2(n19952), .A(n17299), .ZN(n17300) );
  OAI21_X1 U20384 ( .B1(n17301), .B2(n19967), .A(n17300), .ZN(n17302) );
  AOI21_X1 U20385 ( .B1(n17303), .B2(n19962), .A(n17302), .ZN(n17304) );
  OAI221_X1 U20386 ( .B1(n17307), .B2(n17306), .C1(n17307), .C2(n17305), .A(
        n17304), .ZN(P2_U3043) );
  XOR2_X1 U20387 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n17308), .Z(
        n17460) );
  INV_X1 U20388 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n17461) );
  OAI221_X1 U20389 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17311), .C1(
        n17461), .C2(n17310), .A(n17309), .ZN(n17312) );
  AOI21_X1 U20390 ( .B1(n18529), .B2(n17460), .A(n17312), .ZN(n17319) );
  OAI21_X1 U20391 ( .B1(n17315), .B2(n17314), .A(n17313), .ZN(n17316) );
  AOI22_X1 U20392 ( .A1(n17317), .A2(n18681), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17316), .ZN(n17318) );
  OAI211_X1 U20393 ( .C1(n17320), .C2(n18579), .A(n17319), .B(n17318), .ZN(
        P3_U2800) );
  NOR3_X1 U20394 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n17322) );
  NOR4_X1 U20395 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n17321) );
  INV_X2 U20396 ( .A(n17405), .ZN(U215) );
  NAND4_X1 U20397 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n17322), .A3(n17321), .A4(
        U215), .ZN(U213) );
  INV_X1 U20398 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19838) );
  INV_X2 U20399 ( .A(U214), .ZN(n17369) );
  INV_X1 U20400 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n17407) );
  OAI222_X1 U20401 ( .A1(U212), .A2(n19838), .B1(n17371), .B2(n17324), .C1(
        U214), .C2(n17407), .ZN(U216) );
  INV_X1 U20402 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19843) );
  INV_X1 U20403 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n17325) );
  OAI222_X1 U20404 ( .A1(U212), .A2(n19843), .B1(n17371), .B2(n17326), .C1(
        U214), .C2(n17325), .ZN(U217) );
  AOI22_X1 U20405 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n17366), .ZN(n17327) );
  OAI21_X1 U20406 ( .B1(n17328), .B2(n17371), .A(n17327), .ZN(U218) );
  INV_X1 U20407 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U20408 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n17366), .ZN(n17329) );
  OAI21_X1 U20409 ( .B1(n20002), .B2(n17371), .A(n17329), .ZN(U219) );
  INV_X1 U20410 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19996) );
  AOI22_X1 U20411 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n17366), .ZN(n17330) );
  OAI21_X1 U20412 ( .B1(n19996), .B2(n17371), .A(n17330), .ZN(U220) );
  INV_X1 U20413 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n21644) );
  INV_X1 U20414 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n17331) );
  OAI222_X1 U20415 ( .A1(U212), .A2(n21644), .B1(n17371), .B2(n19991), .C1(
        U214), .C2(n17331), .ZN(U221) );
  INV_X1 U20416 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U20417 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n17366), .ZN(n17332) );
  OAI21_X1 U20418 ( .B1(n19984), .B2(n17371), .A(n17332), .ZN(U222) );
  INV_X1 U20419 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n17398) );
  INV_X1 U20420 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n21552) );
  OAI222_X1 U20421 ( .A1(U212), .A2(n17398), .B1(n17371), .B2(n17333), .C1(
        U214), .C2(n21552), .ZN(U223) );
  AOI22_X1 U20422 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n17366), .ZN(n17334) );
  OAI21_X1 U20423 ( .B1(n17335), .B2(n17371), .A(n17334), .ZN(U224) );
  AOI22_X1 U20424 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n17366), .ZN(n17336) );
  OAI21_X1 U20425 ( .B1(n16039), .B2(n17371), .A(n17336), .ZN(U225) );
  AOI22_X1 U20426 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n17366), .ZN(n17337) );
  OAI21_X1 U20427 ( .B1(n17338), .B2(n17371), .A(n17337), .ZN(U226) );
  AOI22_X1 U20428 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n17366), .ZN(n17339) );
  OAI21_X1 U20429 ( .B1(n16053), .B2(n17371), .A(n17339), .ZN(U227) );
  INV_X1 U20430 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n19998) );
  AOI22_X1 U20431 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n17366), .ZN(n17340) );
  OAI21_X1 U20432 ( .B1(n19998), .B2(n17371), .A(n17340), .ZN(U228) );
  INV_X1 U20433 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n21551) );
  AOI22_X1 U20434 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n17366), .ZN(n17341) );
  OAI21_X1 U20435 ( .B1(n21551), .B2(n17371), .A(n17341), .ZN(U229) );
  INV_X1 U20436 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19986) );
  AOI22_X1 U20437 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n17366), .ZN(n17342) );
  OAI21_X1 U20438 ( .B1(n19986), .B2(n17371), .A(n17342), .ZN(U230) );
  AOI22_X1 U20439 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n17366), .ZN(n17343) );
  OAI21_X1 U20440 ( .B1(n17344), .B2(n17371), .A(n17343), .ZN(U231) );
  AOI22_X1 U20441 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n17366), .ZN(n17345) );
  OAI21_X1 U20442 ( .B1(n14181), .B2(n17371), .A(n17345), .ZN(U232) );
  AOI22_X1 U20443 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n17366), .ZN(n17346) );
  OAI21_X1 U20444 ( .B1(n15109), .B2(n17371), .A(n17346), .ZN(U233) );
  AOI22_X1 U20445 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n17366), .ZN(n17347) );
  OAI21_X1 U20446 ( .B1(n14712), .B2(n17371), .A(n17347), .ZN(U234) );
  AOI22_X1 U20447 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n17366), .ZN(n17348) );
  OAI21_X1 U20448 ( .B1(n15115), .B2(n17371), .A(n17348), .ZN(U235) );
  INV_X1 U20449 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n17350) );
  AOI22_X1 U20450 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n17366), .ZN(n17349) );
  OAI21_X1 U20451 ( .B1(n17350), .B2(n17371), .A(n17349), .ZN(U236) );
  AOI22_X1 U20452 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n17366), .ZN(n17351) );
  OAI21_X1 U20453 ( .B1(n21596), .B2(n17371), .A(n17351), .ZN(U237) );
  AOI22_X1 U20454 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n17366), .ZN(n17352) );
  OAI21_X1 U20455 ( .B1(n15136), .B2(n17371), .A(n17352), .ZN(U238) );
  INV_X1 U20456 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20457 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n17366), .ZN(n17353) );
  OAI21_X1 U20458 ( .B1(n17354), .B2(n17371), .A(n17353), .ZN(U239) );
  INV_X1 U20459 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n21583) );
  AOI22_X1 U20460 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n17366), .ZN(n17355) );
  OAI21_X1 U20461 ( .B1(n21583), .B2(n17371), .A(n17355), .ZN(U240) );
  INV_X1 U20462 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20463 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n17366), .ZN(n17356) );
  OAI21_X1 U20464 ( .B1(n17357), .B2(n17371), .A(n17356), .ZN(U241) );
  INV_X1 U20465 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20466 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n17366), .ZN(n17358) );
  OAI21_X1 U20467 ( .B1(n17359), .B2(n17371), .A(n17358), .ZN(U242) );
  INV_X1 U20468 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n17361) );
  AOI22_X1 U20469 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n17366), .ZN(n17360) );
  OAI21_X1 U20470 ( .B1(n17361), .B2(n17371), .A(n17360), .ZN(U243) );
  INV_X1 U20471 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20472 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n17366), .ZN(n17362) );
  OAI21_X1 U20473 ( .B1(n17363), .B2(n17371), .A(n17362), .ZN(U244) );
  INV_X1 U20474 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20475 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n17366), .ZN(n17364) );
  OAI21_X1 U20476 ( .B1(n17365), .B2(n17371), .A(n17364), .ZN(U245) );
  INV_X1 U20477 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20478 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n17366), .ZN(n17367) );
  OAI21_X1 U20479 ( .B1(n17368), .B2(n17371), .A(n17367), .ZN(U246) );
  INV_X1 U20480 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U20481 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n17369), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n17366), .ZN(n17370) );
  OAI21_X1 U20482 ( .B1(n17372), .B2(n17371), .A(n17370), .ZN(U247) );
  INV_X1 U20483 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n17373) );
  INV_X1 U20484 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18993) );
  AOI22_X1 U20485 ( .A1(n17405), .A2(n17373), .B1(n18993), .B2(U215), .ZN(U251) );
  OAI22_X1 U20486 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17405), .ZN(n17374) );
  INV_X1 U20487 ( .A(n17374), .ZN(U252) );
  INV_X1 U20488 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U20489 ( .A1(n17405), .A2(n17375), .B1(n19005), .B2(U215), .ZN(U253) );
  INV_X1 U20490 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n17376) );
  AOI22_X1 U20491 ( .A1(n17393), .A2(n17376), .B1(n19009), .B2(U215), .ZN(U254) );
  INV_X1 U20492 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20493 ( .A1(n17405), .A2(n17377), .B1(n19013), .B2(U215), .ZN(U255) );
  OAI22_X1 U20494 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n17405), .ZN(n17378) );
  INV_X1 U20495 ( .A(n17378), .ZN(U256) );
  INV_X1 U20496 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n17379) );
  AOI22_X1 U20497 ( .A1(n17393), .A2(n17379), .B1(n19020), .B2(U215), .ZN(U257) );
  INV_X1 U20498 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20499 ( .A1(n17393), .A2(n17380), .B1(n13836), .B2(U215), .ZN(U258) );
  OAI22_X1 U20500 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n17405), .ZN(n17381) );
  INV_X1 U20501 ( .A(n17381), .ZN(U259) );
  INV_X1 U20502 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U20503 ( .A1(n17393), .A2(n17382), .B1(n13820), .B2(U215), .ZN(U260) );
  INV_X1 U20504 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20505 ( .A1(n17393), .A2(n17383), .B1(n21539), .B2(U215), .ZN(U261) );
  INV_X1 U20506 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20507 ( .A1(n17393), .A2(n17384), .B1(n13842), .B2(U215), .ZN(U262) );
  INV_X1 U20508 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20509 ( .A1(n17393), .A2(n17385), .B1(n13823), .B2(U215), .ZN(U263) );
  OAI22_X1 U20510 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n17405), .ZN(n17386) );
  INV_X1 U20511 ( .A(n17386), .ZN(U264) );
  OAI22_X1 U20512 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n17405), .ZN(n17387) );
  INV_X1 U20513 ( .A(n17387), .ZN(U265) );
  INV_X1 U20514 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n17388) );
  INV_X1 U20515 ( .A(BUF2_REG_15__SCAN_IN), .ZN(n21571) );
  AOI22_X1 U20516 ( .A1(n17393), .A2(n17388), .B1(n21571), .B2(U215), .ZN(U266) );
  INV_X1 U20517 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20518 ( .A1(n17405), .A2(n17389), .B1(n18997), .B2(U215), .ZN(U267) );
  INV_X1 U20519 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20520 ( .A1(n17393), .A2(n17390), .B1(n16076), .B2(U215), .ZN(U268) );
  INV_X1 U20521 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n17391) );
  AOI22_X1 U20522 ( .A1(n17405), .A2(n17391), .B1(n16070), .B2(U215), .ZN(U269) );
  INV_X1 U20523 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n17392) );
  AOI22_X1 U20524 ( .A1(n17393), .A2(n17392), .B1(n16061), .B2(U215), .ZN(U270) );
  INV_X1 U20525 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n17394) );
  INV_X1 U20526 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n20006) );
  AOI22_X1 U20527 ( .A1(n17405), .A2(n17394), .B1(n20006), .B2(U215), .ZN(U271) );
  INV_X1 U20528 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20529 ( .A1(n17405), .A2(n17395), .B1(n16046), .B2(U215), .ZN(U272) );
  INV_X1 U20530 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20531 ( .A1(n17405), .A2(n17396), .B1(n19021), .B2(U215), .ZN(U273) );
  INV_X1 U20532 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20533 ( .A1(n17405), .A2(n17397), .B1(n16031), .B2(U215), .ZN(U274) );
  AOI22_X1 U20534 ( .A1(n17405), .A2(n17398), .B1(n16026), .B2(U215), .ZN(U275) );
  INV_X1 U20535 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20536 ( .A1(n17405), .A2(n17399), .B1(n16018), .B2(U215), .ZN(U276) );
  INV_X1 U20537 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n19990) );
  AOI22_X1 U20538 ( .A1(n17405), .A2(n21644), .B1(n19990), .B2(U215), .ZN(U277) );
  INV_X1 U20539 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20540 ( .A1(n17405), .A2(n17400), .B1(n14536), .B2(U215), .ZN(U278) );
  INV_X1 U20541 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20542 ( .A1(n17405), .A2(n17401), .B1(n16005), .B2(U215), .ZN(U279) );
  INV_X1 U20543 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U20544 ( .A1(n17405), .A2(n17402), .B1(n12390), .B2(U215), .ZN(U280) );
  AOI22_X1 U20545 ( .A1(n17405), .A2(n19843), .B1(n14609), .B2(U215), .ZN(U281) );
  AOI22_X1 U20546 ( .A1(n17405), .A2(n19838), .B1(n17404), .B2(U215), .ZN(U282) );
  INV_X1 U20547 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17406) );
  AOI222_X1 U20548 ( .A1(n17407), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19838), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17406), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n17408) );
  INV_X2 U20549 ( .A(n17410), .ZN(n17409) );
  INV_X1 U20550 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19496) );
  INV_X1 U20551 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20524) );
  AOI22_X1 U20552 ( .A1(n17409), .A2(n19496), .B1(n20524), .B2(n17410), .ZN(
        U347) );
  INV_X1 U20553 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19494) );
  INV_X1 U20554 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20522) );
  AOI22_X1 U20555 ( .A1(n17408), .A2(n19494), .B1(n20522), .B2(n17410), .ZN(
        U348) );
  INV_X1 U20556 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19492) );
  INV_X1 U20557 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20521) );
  AOI22_X1 U20558 ( .A1(n17409), .A2(n19492), .B1(n20521), .B2(n17410), .ZN(
        U349) );
  INV_X1 U20559 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19491) );
  INV_X1 U20560 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20519) );
  AOI22_X1 U20561 ( .A1(n17409), .A2(n19491), .B1(n20519), .B2(n17410), .ZN(
        U350) );
  INV_X1 U20562 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19489) );
  INV_X1 U20563 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20517) );
  AOI22_X1 U20564 ( .A1(n17409), .A2(n19489), .B1(n20517), .B2(n17410), .ZN(
        U351) );
  INV_X1 U20565 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19487) );
  INV_X1 U20566 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20515) );
  AOI22_X1 U20567 ( .A1(n17409), .A2(n19487), .B1(n20515), .B2(n17410), .ZN(
        U352) );
  INV_X1 U20568 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19486) );
  INV_X1 U20569 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20514) );
  AOI22_X1 U20570 ( .A1(n17409), .A2(n19486), .B1(n20514), .B2(n17410), .ZN(
        U353) );
  INV_X1 U20571 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19484) );
  AOI22_X1 U20572 ( .A1(n17409), .A2(n19484), .B1(n20512), .B2(n17410), .ZN(
        U354) );
  INV_X1 U20573 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n21582) );
  INV_X1 U20574 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20560) );
  AOI22_X1 U20575 ( .A1(n17409), .A2(n21582), .B1(n20560), .B2(n17410), .ZN(
        U355) );
  INV_X1 U20576 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19533) );
  INV_X1 U20577 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20557) );
  AOI22_X1 U20578 ( .A1(n17409), .A2(n19533), .B1(n20557), .B2(n17410), .ZN(
        U356) );
  INV_X1 U20579 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19530) );
  INV_X1 U20580 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20555) );
  AOI22_X1 U20581 ( .A1(n17409), .A2(n19530), .B1(n20555), .B2(n17410), .ZN(
        U357) );
  INV_X1 U20582 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19529) );
  INV_X1 U20583 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20553) );
  AOI22_X1 U20584 ( .A1(n17409), .A2(n19529), .B1(n20553), .B2(n17410), .ZN(
        U358) );
  INV_X1 U20585 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19527) );
  INV_X1 U20586 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20552) );
  AOI22_X1 U20587 ( .A1(n17409), .A2(n19527), .B1(n20552), .B2(n17410), .ZN(
        U359) );
  INV_X1 U20588 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19525) );
  INV_X1 U20589 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20551) );
  AOI22_X1 U20590 ( .A1(n17409), .A2(n19525), .B1(n20551), .B2(n17410), .ZN(
        U360) );
  INV_X1 U20591 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19523) );
  INV_X1 U20592 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20549) );
  AOI22_X1 U20593 ( .A1(n17409), .A2(n19523), .B1(n20549), .B2(n17410), .ZN(
        U361) );
  INV_X1 U20594 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19520) );
  INV_X1 U20595 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20547) );
  AOI22_X1 U20596 ( .A1(n17409), .A2(n19520), .B1(n20547), .B2(n17410), .ZN(
        U362) );
  INV_X1 U20597 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19519) );
  INV_X1 U20598 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20545) );
  AOI22_X1 U20599 ( .A1(n17409), .A2(n19519), .B1(n20545), .B2(n17410), .ZN(
        U363) );
  INV_X1 U20600 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19517) );
  INV_X1 U20601 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20543) );
  AOI22_X1 U20602 ( .A1(n17409), .A2(n19517), .B1(n20543), .B2(n17410), .ZN(
        U364) );
  INV_X1 U20603 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19482) );
  INV_X1 U20604 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20510) );
  AOI22_X1 U20605 ( .A1(n17409), .A2(n19482), .B1(n20510), .B2(n17410), .ZN(
        U365) );
  INV_X1 U20606 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19516) );
  INV_X1 U20607 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20541) );
  AOI22_X1 U20608 ( .A1(n17409), .A2(n19516), .B1(n20541), .B2(n17410), .ZN(
        U366) );
  INV_X1 U20609 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19513) );
  INV_X1 U20610 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20539) );
  AOI22_X1 U20611 ( .A1(n17409), .A2(n19513), .B1(n20539), .B2(n17410), .ZN(
        U367) );
  INV_X1 U20612 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19512) );
  INV_X1 U20613 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20537) );
  AOI22_X1 U20614 ( .A1(n17409), .A2(n19512), .B1(n20537), .B2(n17410), .ZN(
        U368) );
  INV_X1 U20615 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19509) );
  INV_X1 U20616 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20536) );
  AOI22_X1 U20617 ( .A1(n17409), .A2(n19509), .B1(n20536), .B2(n17410), .ZN(
        U369) );
  INV_X1 U20618 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19508) );
  INV_X1 U20619 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20534) );
  AOI22_X1 U20620 ( .A1(n17409), .A2(n19508), .B1(n20534), .B2(n17410), .ZN(
        U370) );
  INV_X1 U20621 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19506) );
  INV_X1 U20622 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20532) );
  AOI22_X1 U20623 ( .A1(n17408), .A2(n19506), .B1(n20532), .B2(n17410), .ZN(
        U371) );
  INV_X1 U20624 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19503) );
  INV_X1 U20625 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20530) );
  AOI22_X1 U20626 ( .A1(n17409), .A2(n19503), .B1(n20530), .B2(n17410), .ZN(
        U372) );
  INV_X1 U20627 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19502) );
  INV_X1 U20628 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20528) );
  AOI22_X1 U20629 ( .A1(n17409), .A2(n19502), .B1(n20528), .B2(n17410), .ZN(
        U373) );
  INV_X1 U20630 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19500) );
  INV_X1 U20631 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20527) );
  AOI22_X1 U20632 ( .A1(n17409), .A2(n19500), .B1(n20527), .B2(n17410), .ZN(
        U374) );
  INV_X1 U20633 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19498) );
  INV_X1 U20634 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20525) );
  AOI22_X1 U20635 ( .A1(n17408), .A2(n19498), .B1(n20525), .B2(n17410), .ZN(
        U375) );
  INV_X1 U20636 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19481) );
  INV_X1 U20637 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20508) );
  AOI22_X1 U20638 ( .A1(n17408), .A2(n19481), .B1(n20508), .B2(n17410), .ZN(
        U376) );
  INV_X1 U20639 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n17412) );
  NAND2_X1 U20640 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19480), .ZN(n19468) );
  NOR2_X1 U20641 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(P3_STATE_REG_1__SCAN_IN), 
        .ZN(n19465) );
  INV_X1 U20642 ( .A(n19465), .ZN(n17411) );
  OAI21_X1 U20643 ( .B1(n19468), .B2(n19479), .A(n17411), .ZN(n19550) );
  OAI21_X1 U20644 ( .B1(n19479), .B2(n17412), .A(n19547), .ZN(P3_U2633) );
  NOR2_X1 U20645 ( .A1(n18379), .A2(n17413), .ZN(n17414) );
  OAI21_X1 U20646 ( .B1(n17414), .B2(n18380), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17415) );
  OAI21_X1 U20647 ( .B1(n17417), .B2(n17416), .A(n17415), .ZN(P3_U2634) );
  AOI21_X1 U20648 ( .B1(n19479), .B2(n19480), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n17418) );
  AOI22_X1 U20649 ( .A1(n19583), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n17418), 
        .B2(n19581), .ZN(P3_U2635) );
  OAI21_X1 U20650 ( .B1(n19463), .B2(BS16), .A(n19550), .ZN(n19548) );
  OAI21_X1 U20651 ( .B1(n19550), .B2(n19571), .A(n19548), .ZN(P3_U2636) );
  INV_X1 U20652 ( .A(n19404), .ZN(n17419) );
  AOI211_X1 U20653 ( .C1(n17422), .C2(n17421), .A(n17420), .B(n17419), .ZN(
        n19407) );
  NOR2_X1 U20654 ( .A1(n19407), .A2(n19449), .ZN(n19563) );
  OAI21_X1 U20655 ( .B1(n19563), .B2(n17424), .A(n17423), .ZN(P3_U2637) );
  NOR4_X1 U20656 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n17428) );
  NOR4_X1 U20657 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n17427) );
  NOR4_X1 U20658 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n17426) );
  NOR4_X1 U20659 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n17425) );
  NAND4_X1 U20660 ( .A1(n17428), .A2(n17427), .A3(n17426), .A4(n17425), .ZN(
        n17434) );
  NOR4_X1 U20661 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n17432) );
  AOI211_X1 U20662 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_26__SCAN_IN), .B(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n17431) );
  NOR4_X1 U20663 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A3(P3_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n17430) );
  NOR4_X1 U20664 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20665 ( .A1(n17432), .A2(n17431), .A3(n17430), .A4(n17429), .ZN(
        n17433) );
  NOR2_X1 U20666 ( .A1(n17434), .A2(n17433), .ZN(n19561) );
  INV_X1 U20667 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19543) );
  NOR3_X1 U20668 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n17436) );
  OAI21_X1 U20669 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n17436), .A(n19561), .ZN(
        n17435) );
  OAI21_X1 U20670 ( .B1(n19561), .B2(n19543), .A(n17435), .ZN(P3_U2638) );
  INV_X1 U20671 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19549) );
  AOI21_X1 U20672 ( .B1(n19554), .B2(n19549), .A(n17436), .ZN(n17437) );
  INV_X1 U20673 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19540) );
  INV_X1 U20674 ( .A(n19561), .ZN(n19556) );
  AOI22_X1 U20675 ( .A1(n19561), .A2(n17437), .B1(n19540), .B2(n19556), .ZN(
        P3_U2639) );
  INV_X1 U20676 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19537) );
  INV_X1 U20677 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19528) );
  INV_X1 U20678 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19526) );
  INV_X1 U20679 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19522) );
  NAND2_X1 U20680 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n17549), .ZN(n17554) );
  NOR2_X1 U20681 ( .A1(n21548), .A2(n17554), .ZN(n17536) );
  NAND2_X1 U20682 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n17536), .ZN(n17514) );
  NOR2_X1 U20683 ( .A1(n19522), .A2(n17514), .ZN(n17520) );
  NAND2_X1 U20684 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n17520), .ZN(n17513) );
  NOR2_X1 U20685 ( .A1(n19526), .A2(n17513), .ZN(n17452) );
  NAND2_X1 U20686 ( .A1(n17807), .A2(n17452), .ZN(n17496) );
  NOR3_X1 U20687 ( .A1(n19531), .A2(n19528), .A3(n17496), .ZN(n17477) );
  NAND2_X1 U20688 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n17477), .ZN(n17454) );
  NOR3_X1 U20689 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19537), .A3(n17454), 
        .ZN(n17438) );
  AOI21_X1 U20690 ( .B1(n17764), .B2(P3_EBX_REG_31__SCAN_IN), .A(n17438), .ZN(
        n17456) );
  INV_X1 U20691 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17891) );
  NAND2_X1 U20692 ( .A1(n17568), .A2(n17891), .ZN(n17567) );
  NOR2_X2 U20693 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17567), .ZN(n17550) );
  INV_X1 U20694 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U20695 ( .A1(n17550), .A2(n17544), .ZN(n17543) );
  INV_X1 U20696 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17872) );
  NAND2_X1 U20697 ( .A1(n17527), .A2(n17872), .ZN(n17519) );
  INV_X1 U20698 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n17825) );
  NAND2_X1 U20699 ( .A1(n17503), .A2(n17825), .ZN(n17499) );
  NOR2_X1 U20700 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17499), .ZN(n17484) );
  INV_X1 U20701 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17480) );
  NAND2_X1 U20702 ( .A1(n17484), .A2(n17480), .ZN(n17458) );
  NOR2_X1 U20703 ( .A1(n17811), .A2(n17458), .ZN(n17466) );
  INV_X1 U20704 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U20705 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n9726), .A(
        n17439), .ZN(n18445) );
  INV_X1 U20706 ( .A(n18445), .ZN(n17487) );
  AOI21_X1 U20707 ( .B1(n10228), .B2(n17440), .A(n9726), .ZN(n18452) );
  INV_X1 U20708 ( .A(n17441), .ZN(n17506) );
  OAI21_X1 U20709 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17443), .A(
        n17442), .ZN(n18461) );
  INV_X1 U20710 ( .A(n18461), .ZN(n17517) );
  INV_X1 U20711 ( .A(n17447), .ZN(n17445) );
  AOI21_X1 U20712 ( .B1(n17540), .B2(n17445), .A(n17444), .ZN(n18480) );
  XOR2_X1 U20713 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n17448), .Z(
        n18504) );
  INV_X1 U20714 ( .A(n18504), .ZN(n17563) );
  INV_X1 U20715 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18507) );
  INV_X1 U20716 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17555) );
  AOI221_X1 U20717 ( .B1(n18507), .B2(n17555), .C1(n17448), .C2(n17555), .A(
        n17447), .ZN(n18496) );
  NOR2_X1 U20718 ( .A1(n17538), .A2(n17775), .ZN(n17530) );
  INV_X1 U20719 ( .A(n17530), .ZN(n17450) );
  INV_X1 U20720 ( .A(n17531), .ZN(n17449) );
  NAND2_X1 U20721 ( .A1(n17450), .A2(n17449), .ZN(n17528) );
  NOR2_X1 U20722 ( .A1(n17504), .A2(n17775), .ZN(n17495) );
  INV_X1 U20723 ( .A(n17473), .ZN(n17451) );
  INV_X1 U20724 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19532) );
  NAND2_X1 U20725 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .ZN(n17453) );
  OR2_X1 U20726 ( .A1(n17712), .A2(n17452), .ZN(n17512) );
  NAND2_X1 U20727 ( .A1(n17816), .A2(n17512), .ZN(n17509) );
  AOI221_X1 U20728 ( .B1(n19532), .B2(n17807), .C1(n17453), .C2(n17807), .A(
        n17509), .ZN(n17483) );
  AOI21_X1 U20729 ( .B1(n17483), .B2(n10428), .A(n19536), .ZN(n17455) );
  NAND2_X1 U20730 ( .A1(n17786), .A2(n17458), .ZN(n17478) );
  XNOR2_X1 U20731 ( .A(n17460), .B(n17459), .ZN(n17464) );
  OAI22_X1 U20732 ( .A1(n17483), .A2(n19537), .B1(n17461), .B2(n17791), .ZN(
        n17462) );
  INV_X1 U20733 ( .A(n17462), .ZN(n17463) );
  INV_X1 U20734 ( .A(n17465), .ZN(n17468) );
  OAI21_X1 U20735 ( .B1(n17764), .B2(n17466), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n17467) );
  OAI211_X1 U20736 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n17478), .A(n17468), .B(
        n17467), .ZN(P3_U2641) );
  INV_X1 U20737 ( .A(n17469), .ZN(n17472) );
  INV_X1 U20738 ( .A(n17470), .ZN(n17471) );
  AOI211_X1 U20739 ( .C1(n17473), .C2(n17472), .A(n17471), .B(n19459), .ZN(
        n17476) );
  OAI22_X1 U20740 ( .A1(n17474), .A2(n17791), .B1(n17812), .B2(n17480), .ZN(
        n17475) );
  AOI211_X1 U20741 ( .C1(n17477), .C2(n19532), .A(n17476), .B(n17475), .ZN(
        n17482) );
  INV_X1 U20742 ( .A(n17478), .ZN(n17479) );
  OAI21_X1 U20743 ( .B1(n17484), .B2(n17480), .A(n17479), .ZN(n17481) );
  OAI211_X1 U20744 ( .C1(n17483), .C2(n19532), .A(n17482), .B(n17481), .ZN(
        P3_U2642) );
  NAND2_X1 U20745 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n19531), .ZN(n17493) );
  AOI22_X1 U20746 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n17492) );
  INV_X1 U20747 ( .A(n17509), .ZN(n17502) );
  OAI21_X1 U20748 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n17496), .A(n17502), 
        .ZN(n17490) );
  AOI211_X1 U20749 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n17499), .A(n17484), .B(
        n17811), .ZN(n17489) );
  AOI211_X1 U20750 ( .C1(n17487), .C2(n17486), .A(n17485), .B(n19459), .ZN(
        n17488) );
  AOI211_X1 U20751 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n17490), .A(n17489), 
        .B(n17488), .ZN(n17491) );
  OAI211_X1 U20752 ( .C1(n17496), .C2(n17493), .A(n17492), .B(n17491), .ZN(
        P3_U2643) );
  AOI211_X1 U20753 ( .C1(n18452), .C2(n17495), .A(n17494), .B(n19459), .ZN(
        n17498) );
  OAI22_X1 U20754 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n17496), .B1(n17825), 
        .B2(n17812), .ZN(n17497) );
  AOI211_X1 U20755 ( .C1(n17805), .C2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n17498), .B(n17497), .ZN(n17501) );
  OAI211_X1 U20756 ( .C1(n17503), .C2(n17825), .A(n17786), .B(n17499), .ZN(
        n17500) );
  OAI211_X1 U20757 ( .C1(n17502), .C2(n19528), .A(n17501), .B(n17500), .ZN(
        P3_U2644) );
  AOI22_X1 U20758 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n17511) );
  AOI211_X1 U20759 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n17519), .A(n17503), .B(
        n17811), .ZN(n17508) );
  AOI211_X1 U20760 ( .C1(n17506), .C2(n17505), .A(n17504), .B(n19459), .ZN(
        n17507) );
  AOI211_X1 U20761 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n17509), .A(n17508), 
        .B(n17507), .ZN(n17510) );
  OAI211_X1 U20762 ( .C1(n17513), .C2(n17512), .A(n17511), .B(n17510), .ZN(
        P3_U2645) );
  AOI22_X1 U20763 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_25__SCAN_IN), .ZN(n17524) );
  INV_X1 U20764 ( .A(n17514), .ZN(n17526) );
  OAI21_X1 U20765 ( .B1(n17526), .B2(n17712), .A(n17816), .ZN(n17537) );
  NOR2_X1 U20766 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17712), .ZN(n17525) );
  AOI211_X1 U20767 ( .C1(n17517), .C2(n17516), .A(n17515), .B(n19459), .ZN(
        n17518) );
  AOI221_X1 U20768 ( .B1(n17537), .B2(P3_REIP_REG_25__SCAN_IN), .C1(n17525), 
        .C2(P3_REIP_REG_25__SCAN_IN), .A(n17518), .ZN(n17523) );
  OAI211_X1 U20769 ( .C1(n17527), .C2(n17872), .A(n17786), .B(n17519), .ZN(
        n17522) );
  INV_X1 U20770 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19524) );
  NAND3_X1 U20771 ( .A1(n17807), .A2(n17520), .A3(n19524), .ZN(n17521) );
  NAND4_X1 U20772 ( .A1(n17524), .A2(n17523), .A3(n17522), .A4(n17521), .ZN(
        P3_U2646) );
  AOI22_X1 U20773 ( .A1(n17764), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n17526), 
        .B2(n17525), .ZN(n17535) );
  AOI211_X1 U20774 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n17543), .A(n17527), .B(
        n17811), .ZN(n17533) );
  INV_X1 U20775 ( .A(n17528), .ZN(n17529) );
  AOI211_X1 U20776 ( .C1(n17531), .C2(n17530), .A(n17529), .B(n19459), .ZN(
        n17532) );
  AOI211_X1 U20777 ( .C1(n17537), .C2(P3_REIP_REG_24__SCAN_IN), .A(n17533), 
        .B(n17532), .ZN(n17534) );
  OAI211_X1 U20778 ( .C1(n18460), .C2(n17791), .A(n17535), .B(n17534), .ZN(
        P3_U2647) );
  AOI21_X1 U20779 ( .B1(n17807), .B2(n17536), .A(P3_REIP_REG_23__SCAN_IN), 
        .ZN(n17548) );
  INV_X1 U20780 ( .A(n17537), .ZN(n17547) );
  AOI211_X1 U20781 ( .C1(n18480), .C2(n17539), .A(n17538), .B(n19459), .ZN(
        n17542) );
  OAI22_X1 U20782 ( .A1(n17540), .A2(n17791), .B1(n17812), .B2(n17544), .ZN(
        n17541) );
  NOR2_X1 U20783 ( .A1(n17542), .A2(n17541), .ZN(n17546) );
  OAI211_X1 U20784 ( .C1(n17550), .C2(n17544), .A(n17786), .B(n17543), .ZN(
        n17545) );
  OAI211_X1 U20785 ( .C1(n17548), .C2(n17547), .A(n17546), .B(n17545), .ZN(
        P3_U2648) );
  INV_X1 U20786 ( .A(n17566), .ZN(n17561) );
  INV_X1 U20787 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19518) );
  NAND3_X1 U20788 ( .A1(n17807), .A2(n17549), .A3(n19518), .ZN(n17570) );
  AOI211_X1 U20789 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n17567), .A(n17550), .B(
        n17811), .ZN(n17559) );
  INV_X1 U20790 ( .A(n17551), .ZN(n17552) );
  AOI211_X1 U20791 ( .C1(n18496), .C2(n17553), .A(n17552), .B(n19459), .ZN(
        n17558) );
  NOR3_X1 U20792 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17712), .A3(n17554), 
        .ZN(n17557) );
  INV_X1 U20793 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n17886) );
  OAI22_X1 U20794 ( .A1(n17555), .A2(n17791), .B1(n17812), .B2(n17886), .ZN(
        n17556) );
  NOR4_X1 U20795 ( .A1(n17559), .A2(n17558), .A3(n17557), .A4(n17556), .ZN(
        n17560) );
  OAI221_X1 U20796 ( .B1(n21548), .B2(n17561), .C1(n21548), .C2(n17570), .A(
        n17560), .ZN(P3_U2649) );
  AOI211_X1 U20797 ( .C1(n17563), .C2(n9730), .A(n17562), .B(n19459), .ZN(
        n17565) );
  OAI22_X1 U20798 ( .A1(n18507), .A2(n17791), .B1(n17812), .B2(n17891), .ZN(
        n17564) );
  AOI211_X1 U20799 ( .C1(n17566), .C2(P3_REIP_REG_21__SCAN_IN), .A(n17565), 
        .B(n17564), .ZN(n17571) );
  OAI211_X1 U20800 ( .C1(n17568), .C2(n17891), .A(n17786), .B(n17567), .ZN(
        n17569) );
  NAND3_X1 U20801 ( .A1(n17571), .A2(n17570), .A3(n17569), .ZN(P3_U2650) );
  AOI22_X1 U20802 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n17584) );
  OAI21_X1 U20803 ( .B1(n17572), .B2(n17712), .A(n17816), .ZN(n17603) );
  INV_X1 U20804 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19514) );
  INV_X1 U20805 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19511) );
  AOI211_X1 U20806 ( .C1(n19514), .C2(n19511), .A(n17573), .B(n17594), .ZN(
        n17579) );
  INV_X1 U20807 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17575) );
  NAND2_X1 U20808 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17574), .ZN(
        n17595) );
  NOR2_X1 U20809 ( .A1(n10231), .A2(n17595), .ZN(n18527) );
  NAND2_X1 U20810 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n18527), .ZN(
        n17585) );
  AOI21_X1 U20811 ( .B1(n17575), .B2(n17585), .A(n18493), .ZN(n18528) );
  INV_X1 U20812 ( .A(n17597), .ZN(n17614) );
  OAI21_X1 U20813 ( .B1(n17585), .B2(n17614), .A(n14217), .ZN(n17587) );
  INV_X1 U20814 ( .A(n17587), .ZN(n17577) );
  OAI21_X1 U20815 ( .B1(n18528), .B2(n17577), .A(n17784), .ZN(n17576) );
  AOI21_X1 U20816 ( .B1(n18528), .B2(n17577), .A(n17576), .ZN(n17578) );
  AOI211_X1 U20817 ( .C1(n17603), .C2(P3_REIP_REG_19__SCAN_IN), .A(n17579), 
        .B(n17578), .ZN(n17583) );
  OAI211_X1 U20818 ( .C1(n17588), .C2(n17581), .A(n17786), .B(n17580), .ZN(
        n17582) );
  NAND4_X1 U20819 ( .A1(n17584), .A2(n17583), .A3(n18981), .A4(n17582), .ZN(
        P3_U2652) );
  INV_X1 U20820 ( .A(n17603), .ZN(n17593) );
  OAI21_X1 U20821 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18527), .A(
        n17585), .ZN(n18542) );
  NAND2_X1 U20822 ( .A1(n17784), .A2(n17775), .ZN(n17802) );
  INV_X1 U20823 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n18545) );
  OAI221_X1 U20824 ( .B1(n18542), .B2(n17597), .C1(n18542), .C2(n18545), .A(
        n17784), .ZN(n17586) );
  AOI22_X1 U20825 ( .A1(n17587), .A2(n18542), .B1(n17802), .B2(n17586), .ZN(
        n17591) );
  AOI211_X1 U20826 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17604), .A(n17588), .B(
        n17811), .ZN(n17590) );
  OAI22_X1 U20827 ( .A1(n18545), .A2(n17791), .B1(n17812), .B2(n17973), .ZN(
        n17589) );
  NOR4_X1 U20828 ( .A1(n18954), .A2(n17591), .A3(n17590), .A4(n17589), .ZN(
        n17592) );
  OAI221_X1 U20829 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17594), .C1(n19511), 
        .C2(n17593), .A(n17592), .ZN(P3_U2653) );
  AOI21_X1 U20830 ( .B1(n10231), .B2(n17595), .A(n18527), .ZN(n18557) );
  INV_X1 U20831 ( .A(n17618), .ZN(n17596) );
  OAI21_X1 U20832 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17596), .A(
        n17595), .ZN(n18575) );
  AOI21_X1 U20833 ( .B1(n17597), .B2(n18575), .A(n17775), .ZN(n17599) );
  OAI21_X1 U20834 ( .B1(n18557), .B2(n17599), .A(n17784), .ZN(n17598) );
  AOI21_X1 U20835 ( .B1(n18557), .B2(n17599), .A(n17598), .ZN(n17602) );
  NAND4_X1 U20836 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17625), .A4(n19510), .ZN(n17600) );
  OAI211_X1 U20837 ( .C1(n17812), .C2(n17605), .A(n18981), .B(n17600), .ZN(
        n17601) );
  AOI211_X1 U20838 ( .C1(n17603), .C2(P3_REIP_REG_17__SCAN_IN), .A(n17602), 
        .B(n17601), .ZN(n17607) );
  OAI211_X1 U20839 ( .C1(n17609), .C2(n17605), .A(n17786), .B(n17604), .ZN(
        n17606) );
  OAI211_X1 U20840 ( .C1(n17791), .C2(n10231), .A(n17607), .B(n17606), .ZN(
        P3_U2654) );
  AOI21_X1 U20841 ( .B1(n17807), .B2(n17608), .A(n17796), .ZN(n17642) );
  AOI211_X1 U20842 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17626), .A(n17609), .B(
        n17811), .ZN(n17613) );
  NAND2_X1 U20843 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n17610) );
  OAI211_X1 U20844 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n17625), .B(n17610), .ZN(n17611) );
  OAI211_X1 U20845 ( .C1(n17812), .C2(n18006), .A(n18981), .B(n17611), .ZN(
        n17612) );
  AOI211_X1 U20846 ( .C1(n17805), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n17613), .B(n17612), .ZN(n17617) );
  NAND2_X1 U20847 ( .A1(n14217), .A2(n17614), .ZN(n17619) );
  NAND2_X1 U20848 ( .A1(n18575), .A2(n17619), .ZN(n17615) );
  OAI211_X1 U20849 ( .C1(n18575), .C2(n17619), .A(n17784), .B(n17615), .ZN(
        n17616) );
  OAI211_X1 U20850 ( .C1(n17642), .C2(n19507), .A(n17617), .B(n17616), .ZN(
        P3_U2655) );
  AOI22_X1 U20851 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_15__SCAN_IN), .ZN(n17630) );
  OAI21_X1 U20852 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n18570), .A(
        n17618), .ZN(n18580) );
  INV_X1 U20853 ( .A(n18580), .ZN(n17620) );
  NOR3_X1 U20854 ( .A1(n17620), .A2(n19459), .A3(n17619), .ZN(n17624) );
  NOR2_X1 U20855 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19459), .ZN(
        n17621) );
  INV_X1 U20856 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n18583) );
  INV_X1 U20857 ( .A(n17802), .ZN(n17671) );
  AOI21_X1 U20858 ( .B1(n17621), .B2(n18583), .A(n17671), .ZN(n17622) );
  OAI22_X1 U20859 ( .A1(n17622), .A2(n18580), .B1(n19505), .B2(n17642), .ZN(
        n17623) );
  AOI211_X1 U20860 ( .C1(n17625), .C2(n19505), .A(n17624), .B(n17623), .ZN(
        n17629) );
  OAI211_X1 U20861 ( .C1(n17632), .C2(n17627), .A(n17786), .B(n17626), .ZN(
        n17628) );
  NAND4_X1 U20862 ( .A1(n17630), .A2(n17629), .A3(n18981), .A4(n17628), .ZN(
        P3_U2656) );
  NOR2_X1 U20863 ( .A1(n17712), .A2(n17631), .ZN(n17656) );
  AOI21_X1 U20864 ( .B1(P3_REIP_REG_13__SCAN_IN), .B2(n17656), .A(
        P3_REIP_REG_14__SCAN_IN), .ZN(n17643) );
  AOI211_X1 U20865 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17650), .A(n17632), .B(
        n17811), .ZN(n17640) );
  OAI22_X1 U20866 ( .A1(n17634), .A2(n17791), .B1(n17812), .B2(n17633), .ZN(
        n17639) );
  AOI21_X1 U20867 ( .B1(n17634), .B2(n17647), .A(n18570), .ZN(n18600) );
  NAND2_X1 U20868 ( .A1(n17635), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17798) );
  INV_X1 U20869 ( .A(n17798), .ZN(n17799) );
  NAND2_X1 U20870 ( .A1(n16901), .A2(n17799), .ZN(n17739) );
  OAI21_X1 U20871 ( .B1(n17636), .B2(n17739), .A(n14217), .ZN(n17681) );
  OAI21_X1 U20872 ( .B1(n10222), .B2(n17775), .A(n17681), .ZN(n17657) );
  OAI21_X1 U20873 ( .B1(n18600), .B2(n17657), .A(n17784), .ZN(n17637) );
  AOI21_X1 U20874 ( .B1(n18600), .B2(n17657), .A(n17637), .ZN(n17638) );
  NOR4_X1 U20875 ( .A1(n18954), .A2(n17640), .A3(n17639), .A4(n17638), .ZN(
        n17641) );
  OAI21_X1 U20876 ( .B1(n17643), .B2(n17642), .A(n17641), .ZN(P3_U2657) );
  INV_X1 U20877 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19499) );
  INV_X1 U20878 ( .A(n17644), .ZN(n17645) );
  NOR2_X1 U20879 ( .A1(n17796), .A2(n17690), .ZN(n17689) );
  NOR2_X1 U20880 ( .A1(n17807), .A2(n17796), .ZN(n17813) );
  AOI21_X1 U20881 ( .B1(n17645), .B2(n17689), .A(n17813), .ZN(n17673) );
  AOI21_X1 U20882 ( .B1(n17807), .B2(n19499), .A(n17673), .ZN(n17660) );
  INV_X1 U20883 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18625) );
  INV_X1 U20884 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18658) );
  INV_X1 U20885 ( .A(n17646), .ZN(n17698) );
  NAND2_X1 U20886 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17698), .ZN(
        n17697) );
  NOR2_X1 U20887 ( .A1(n18658), .A2(n17697), .ZN(n17683) );
  NAND2_X1 U20888 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17683), .ZN(
        n17670) );
  NOR2_X1 U20889 ( .A1(n18625), .A2(n17670), .ZN(n17648) );
  INV_X1 U20890 ( .A(n17648), .ZN(n17665) );
  OAI21_X1 U20891 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17648), .A(
        n17647), .ZN(n18613) );
  AOI211_X1 U20892 ( .C1(n17665), .C2(n17802), .A(n17649), .B(n18613), .ZN(
        n17655) );
  AOI21_X1 U20893 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17805), .A(
        n18954), .ZN(n17652) );
  OAI211_X1 U20894 ( .C1(n17661), .C2(n17653), .A(n17786), .B(n17650), .ZN(
        n17651) );
  OAI211_X1 U20895 ( .C1(n17653), .C2(n17812), .A(n17652), .B(n17651), .ZN(
        n17654) );
  AOI211_X1 U20896 ( .C1(n17656), .C2(n19501), .A(n17655), .B(n17654), .ZN(
        n17659) );
  NAND3_X1 U20897 ( .A1(n17784), .A2(n18613), .A3(n17657), .ZN(n17658) );
  OAI211_X1 U20898 ( .C1(n17660), .C2(n19501), .A(n17659), .B(n17658), .ZN(
        P3_U2658) );
  AOI22_X1 U20899 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17805), .B1(
        n17764), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n17669) );
  NOR2_X1 U20900 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17712), .ZN(n17663) );
  AOI211_X1 U20901 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17674), .A(n17661), .B(
        n17811), .ZN(n17662) );
  AOI211_X1 U20902 ( .C1(n17664), .C2(n17663), .A(n18954), .B(n17662), .ZN(
        n17668) );
  INV_X1 U20903 ( .A(n17670), .ZN(n18609) );
  OAI21_X1 U20904 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18609), .A(
        n17665), .ZN(n18621) );
  XOR2_X1 U20905 ( .A(n18621), .B(n17681), .Z(n17666) );
  AOI22_X1 U20906 ( .A1(n17784), .A2(n17666), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n17673), .ZN(n17667) );
  NAND3_X1 U20907 ( .A1(n17669), .A2(n17668), .A3(n17667), .ZN(P3_U2659) );
  OAI21_X1 U20908 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17683), .A(
        n17670), .ZN(n18639) );
  OR2_X1 U20909 ( .A1(n17683), .A2(n17671), .ZN(n17672) );
  AOI22_X1 U20910 ( .A1(n17784), .A2(n18639), .B1(n17740), .B2(n17672), .ZN(
        n17682) );
  INV_X1 U20911 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17678) );
  INV_X1 U20912 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19493) );
  NOR3_X1 U20913 ( .A1(n17712), .A2(n17690), .A3(n19493), .ZN(n17688) );
  OAI221_X1 U20914 ( .B1(P3_REIP_REG_11__SCAN_IN), .B2(P3_REIP_REG_10__SCAN_IN), .C1(P3_REIP_REG_11__SCAN_IN), .C2(n17688), .A(n17673), .ZN(n17677) );
  OAI211_X1 U20915 ( .C1(n17684), .C2(n17675), .A(n17786), .B(n17674), .ZN(
        n17676) );
  OAI211_X1 U20916 ( .C1(n17791), .C2(n17678), .A(n17677), .B(n17676), .ZN(
        n17679) );
  AOI211_X1 U20917 ( .C1(n17764), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18954), .B(
        n17679), .ZN(n17680) );
  OAI221_X1 U20918 ( .B1(n17682), .B2(n18639), .C1(n17682), .C2(n17681), .A(
        n17680), .ZN(P3_U2660) );
  AOI21_X1 U20919 ( .B1(n18658), .B2(n17697), .A(n17683), .ZN(n18666) );
  OAI21_X1 U20920 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17697), .A(
        n14217), .ZN(n17701) );
  XOR2_X1 U20921 ( .A(n18666), .B(n17701), .Z(n17695) );
  AOI211_X1 U20922 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17685), .A(n17684), .B(
        n17811), .ZN(n17687) );
  OAI21_X1 U20923 ( .B1(n18658), .B2(n17791), .A(n18981), .ZN(n17686) );
  AOI211_X1 U20924 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17764), .A(n17687), .B(
        n17686), .ZN(n17694) );
  INV_X1 U20925 ( .A(n17688), .ZN(n17692) );
  NOR2_X1 U20926 ( .A1(n17813), .A2(n17689), .ZN(n17696) );
  NOR3_X1 U20927 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17690), .A3(n17712), .ZN(
        n17704) );
  NOR2_X1 U20928 ( .A1(n17696), .A2(n17704), .ZN(n17691) );
  MUX2_X1 U20929 ( .A(n17692), .B(n17691), .S(P3_REIP_REG_10__SCAN_IN), .Z(
        n17693) );
  OAI211_X1 U20930 ( .C1(n19459), .C2(n17695), .A(n17694), .B(n17693), .ZN(
        P3_U2661) );
  INV_X1 U20931 ( .A(n17696), .ZN(n17716) );
  OAI21_X1 U20932 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17698), .A(
        n17697), .ZN(n18678) );
  NOR2_X1 U20933 ( .A1(n17713), .A2(n17739), .ZN(n17699) );
  OAI221_X1 U20934 ( .B1(n18678), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n18678), .C2(n17699), .A(n17784), .ZN(n17700) );
  AOI22_X1 U20935 ( .A1(n18678), .A2(n17701), .B1(n17802), .B2(n17700), .ZN(
        n17702) );
  AOI211_X1 U20936 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17805), .A(
        n18954), .B(n17702), .ZN(n17709) );
  INV_X1 U20937 ( .A(n17710), .ZN(n17703) );
  OAI21_X1 U20938 ( .B1(n17811), .B2(n17703), .A(n17812), .ZN(n17707) );
  NOR2_X1 U20939 ( .A1(n17710), .A2(n17811), .ZN(n17706) );
  AOI221_X1 U20940 ( .B1(n17707), .B2(P3_EBX_REG_9__SCAN_IN), .C1(n17706), 
        .C2(n17705), .A(n17704), .ZN(n17708) );
  OAI211_X1 U20941 ( .C1(n19493), .C2(n17716), .A(n17709), .B(n17708), .ZN(
        P3_U2662) );
  AOI211_X1 U20942 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17731), .A(n17710), .B(
        n17811), .ZN(n17719) );
  NOR2_X1 U20943 ( .A1(n19490), .A2(n14303), .ZN(n17724) );
  INV_X1 U20944 ( .A(n17711), .ZN(n17723) );
  NOR2_X1 U20945 ( .A1(n17712), .A2(n17723), .ZN(n17744) );
  AOI21_X1 U20946 ( .B1(n17724), .B2(n17744), .A(P3_REIP_REG_8__SCAN_IN), .ZN(
        n17717) );
  OAI21_X1 U20947 ( .B1(n17713), .B2(n17739), .A(n14217), .ZN(n17722) );
  XNOR2_X1 U20948 ( .A(n17714), .B(n17722), .ZN(n17715) );
  OAI22_X1 U20949 ( .A1(n17717), .A2(n17716), .B1(n19459), .B2(n17715), .ZN(
        n17718) );
  AOI211_X1 U20950 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17764), .A(n17719), .B(
        n17718), .ZN(n17720) );
  OAI211_X1 U20951 ( .C1(n17721), .C2(n17791), .A(n17720), .B(n18981), .ZN(
        P3_U2663) );
  OAI221_X1 U20952 ( .B1(n19459), .B2(n17730), .C1(n19459), .C2(n17739), .A(
        n17802), .ZN(n17729) );
  INV_X1 U20953 ( .A(n17722), .ZN(n17728) );
  AOI21_X1 U20954 ( .B1(n17807), .B2(n17723), .A(n17796), .ZN(n17750) );
  AOI21_X1 U20955 ( .B1(n19490), .B2(n14303), .A(n17724), .ZN(n17725) );
  AOI22_X1 U20956 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17805), .B1(
        n17744), .B2(n17725), .ZN(n17726) );
  OAI211_X1 U20957 ( .C1(n17750), .C2(n19490), .A(n17726), .B(n18981), .ZN(
        n17727) );
  AOI221_X1 U20958 ( .B1(n17730), .B2(n17729), .C1(n17728), .C2(n17729), .A(
        n17727), .ZN(n17733) );
  OAI211_X1 U20959 ( .C1(n17735), .C2(n17734), .A(n17786), .B(n17731), .ZN(
        n17732) );
  OAI211_X1 U20960 ( .C1(n17734), .C2(n17812), .A(n17733), .B(n17732), .ZN(
        P3_U2664) );
  AOI211_X1 U20961 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17753), .A(n17735), .B(
        n17811), .ZN(n17736) );
  AOI211_X1 U20962 ( .C1(n17764), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18954), .B(
        n17736), .ZN(n17746) );
  OAI21_X1 U20963 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17747), .A(
        n17737), .ZN(n18689) );
  INV_X1 U20964 ( .A(n17738), .ZN(n17797) );
  AND3_X1 U20965 ( .A1(n18689), .A2(n17739), .A3(n17797), .ZN(n17743) );
  OAI21_X1 U20966 ( .B1(n17747), .B2(n17775), .A(n17740), .ZN(n17741) );
  OAI22_X1 U20967 ( .A1(n17750), .A2(n14303), .B1(n18689), .B2(n17741), .ZN(
        n17742) );
  AOI211_X1 U20968 ( .C1(n17744), .C2(n14303), .A(n17743), .B(n17742), .ZN(
        n17745) );
  OAI211_X1 U20969 ( .C1(n18685), .C2(n17791), .A(n17746), .B(n17745), .ZN(
        P3_U2665) );
  INV_X1 U20970 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17757) );
  INV_X1 U20971 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19483) );
  NAND3_X1 U20972 ( .A1(n17807), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n17778) );
  NOR2_X1 U20973 ( .A1(n19483), .A2(n17778), .ZN(n17770) );
  AOI21_X1 U20974 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n17770), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17751) );
  AOI21_X1 U20975 ( .B1(n17757), .B2(n17748), .A(n17747), .ZN(n18699) );
  OAI21_X1 U20976 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17748), .A(
        n14217), .ZN(n17765) );
  XOR2_X1 U20977 ( .A(n18699), .B(n17765), .Z(n17749) );
  OAI22_X1 U20978 ( .A1(n17751), .A2(n17750), .B1(n19459), .B2(n17749), .ZN(
        n17752) );
  AOI211_X1 U20979 ( .C1(n17764), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18954), .B(
        n17752), .ZN(n17756) );
  OAI211_X1 U20980 ( .C1(n17759), .C2(n17754), .A(n17786), .B(n17753), .ZN(
        n17755) );
  OAI211_X1 U20981 ( .C1(n17791), .C2(n17757), .A(n17756), .B(n17755), .ZN(
        P3_U2666) );
  AOI21_X1 U20982 ( .B1(n17807), .B2(n17758), .A(n17796), .ZN(n17777) );
  AOI211_X1 U20983 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17785), .A(n17759), .B(
        n17811), .ZN(n17763) );
  OAI21_X1 U20984 ( .B1(n18112), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n19588), .ZN(n17760) );
  OAI211_X1 U20985 ( .C1(n17791), .C2(n17761), .A(n18981), .B(n17760), .ZN(
        n17762) );
  AOI211_X1 U20986 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17764), .A(n17763), .B(
        n17762), .ZN(n17773) );
  INV_X1 U20987 ( .A(n17765), .ZN(n17766) );
  AOI22_X1 U20988 ( .A1(n17799), .A2(n17767), .B1(n17766), .B2(n17769), .ZN(
        n17768) );
  OAI21_X1 U20989 ( .B1(n14217), .B2(n17769), .A(n17768), .ZN(n17771) );
  AOI22_X1 U20990 ( .A1(n17784), .A2(n17771), .B1(n17770), .B2(n19485), .ZN(
        n17772) );
  OAI211_X1 U20991 ( .C1(n19485), .C2(n17777), .A(n17773), .B(n17772), .ZN(
        P3_U2667) );
  INV_X1 U20992 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17790) );
  NAND2_X1 U20993 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17794) );
  AOI21_X1 U20994 ( .B1(n17790), .B2(n17794), .A(n17774), .ZN(n18715) );
  AOI21_X1 U20995 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17799), .A(
        n17775), .ZN(n17776) );
  XOR2_X1 U20996 ( .A(n18715), .B(n17776), .Z(n17783) );
  AOI21_X1 U20997 ( .B1(n19483), .B2(n17778), .A(n17777), .ZN(n17782) );
  INV_X1 U20998 ( .A(n17779), .ZN(n17780) );
  OAI22_X1 U20999 ( .A1(n17820), .A2(n17780), .B1(n17787), .B2(n17812), .ZN(
        n17781) );
  AOI211_X1 U21000 ( .C1(n17784), .C2(n17783), .A(n17782), .B(n17781), .ZN(
        n17789) );
  OAI211_X1 U21001 ( .C1(n17792), .C2(n17787), .A(n17786), .B(n17785), .ZN(
        n17788) );
  OAI211_X1 U21002 ( .C1(n17791), .C2(n17790), .A(n17789), .B(n17788), .ZN(
        P3_U2668) );
  INV_X1 U21003 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17810) );
  AOI211_X1 U21004 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17793), .A(n17792), .B(
        n17811), .ZN(n17804) );
  OAI21_X1 U21005 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17794), .ZN(n18719) );
  AOI22_X1 U21006 ( .A1(n17796), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n19588), 
        .B2(n17795), .ZN(n17801) );
  INV_X1 U21007 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18723) );
  OAI221_X1 U21008 ( .B1(n17799), .B2(n18719), .C1(n17798), .C2(n18723), .A(
        n17797), .ZN(n17800) );
  OAI211_X1 U21009 ( .C1(n17802), .C2(n18719), .A(n17801), .B(n17800), .ZN(
        n17803) );
  AOI211_X1 U21010 ( .C1(n17805), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n17804), .B(n17803), .ZN(n17809) );
  NAND2_X1 U21011 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17806) );
  OAI211_X1 U21012 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n17807), .B(n17806), .ZN(n17808) );
  OAI211_X1 U21013 ( .C1(n17810), .C2(n17812), .A(n17809), .B(n17808), .ZN(
        P3_U2669) );
  NAND2_X1 U21014 ( .A1(n17812), .A2(n17811), .ZN(n17815) );
  INV_X1 U21015 ( .A(n17813), .ZN(n17814) );
  AOI22_X1 U21016 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17815), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n17814), .ZN(n17819) );
  NAND3_X1 U21017 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17817), .A3(
        n17816), .ZN(n17818) );
  OAI211_X1 U21018 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n17820), .A(
        n17819), .B(n17818), .ZN(P3_U2671) );
  NOR2_X1 U21019 ( .A1(n17821), .A2(n17955), .ZN(n17910) );
  INV_X1 U21020 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n17824) );
  NOR4_X1 U21021 ( .A1(n17825), .A2(n17824), .A3(n17823), .A4(n17822), .ZN(
        n17826) );
  NAND4_X1 U21022 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_28__SCAN_IN), 
        .A3(n17910), .A4(n17826), .ZN(n17829) );
  NAND2_X1 U21023 ( .A1(n18163), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17828) );
  NAND2_X1 U21024 ( .A1(n17860), .A2(n18120), .ZN(n17827) );
  OAI22_X1 U21025 ( .A1(n17860), .A2(n17828), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17827), .ZN(P3_U2672) );
  NAND2_X1 U21026 ( .A1(n17830), .A2(n17829), .ZN(n17831) );
  NAND2_X1 U21027 ( .A1(n17831), .A2(n18171), .ZN(n17859) );
  AOI22_X1 U21028 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17835) );
  AOI22_X1 U21029 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18056), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17833) );
  AOI22_X1 U21031 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17832) );
  NAND4_X1 U21032 ( .A1(n17835), .A2(n17834), .A3(n17833), .A4(n17832), .ZN(
        n17843) );
  AOI22_X1 U21033 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n9573), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17837) );
  NAND2_X1 U21034 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n17836) );
  OAI211_X1 U21035 ( .C1(n18151), .C2(n18135), .A(n17837), .B(n17836), .ZN(
        n17842) );
  INV_X1 U21036 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17839) );
  INV_X1 U21037 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17838) );
  OAI22_X1 U21038 ( .A1(n18067), .A2(n17839), .B1(n18138), .B2(n17838), .ZN(
        n17841) );
  OAI22_X1 U21039 ( .A1(n17112), .A2(n18016), .B1(n18141), .B2(n18014), .ZN(
        n17840) );
  OR4_X1 U21040 ( .A1(n17843), .A2(n17842), .A3(n17841), .A4(n17840), .ZN(
        n17858) );
  INV_X1 U21041 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17894) );
  AOI22_X1 U21042 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17845) );
  NAND2_X1 U21043 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n17844) );
  OAI211_X1 U21044 ( .C1(n17894), .C2(n18067), .A(n17845), .B(n17844), .ZN(
        n17850) );
  INV_X1 U21045 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n18036) );
  OAI22_X1 U21046 ( .A1(n9620), .A2(n17846), .B1(n18141), .B2(n18036), .ZN(
        n17849) );
  INV_X1 U21047 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18034) );
  INV_X1 U21048 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17847) );
  OAI22_X1 U21049 ( .A1(n9626), .A2(n18034), .B1(n18035), .B2(n17847), .ZN(
        n17848) );
  OR3_X1 U21050 ( .A1(n17850), .A2(n17849), .A3(n17848), .ZN(n17856) );
  AOI22_X1 U21051 ( .A1(n18091), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17854) );
  AOI22_X1 U21052 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U21053 ( .A1(n13178), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17852) );
  AOI22_X1 U21054 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17851) );
  NAND4_X1 U21055 ( .A1(n17854), .A2(n17853), .A3(n17852), .A4(n17851), .ZN(
        n17855) );
  NOR2_X1 U21056 ( .A1(n17856), .A2(n17855), .ZN(n17863) );
  NOR3_X1 U21057 ( .A1(n17863), .A2(n17861), .A3(n17866), .ZN(n17857) );
  XNOR2_X1 U21058 ( .A(n17858), .B(n17857), .ZN(n18193) );
  OAI22_X1 U21059 ( .A1(n17860), .A2(n17859), .B1(n18193), .B2(n18171), .ZN(
        P3_U2673) );
  INV_X1 U21060 ( .A(n9632), .ZN(n17870) );
  NAND2_X1 U21061 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17870), .ZN(n17865) );
  NOR2_X1 U21062 ( .A1(n17861), .A2(n17866), .ZN(n17862) );
  XOR2_X1 U21063 ( .A(n17863), .B(n17862), .Z(n18197) );
  NAND3_X1 U21064 ( .A1(n17865), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n18171), 
        .ZN(n17864) );
  OAI221_X1 U21065 ( .B1(n17865), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n18171), 
        .C2(n18197), .A(n17864), .ZN(P3_U2674) );
  AOI21_X1 U21066 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n18163), .A(n17877), .ZN(
        n17869) );
  OAI21_X1 U21067 ( .B1(n17868), .B2(n17867), .A(n17866), .ZN(n18205) );
  OAI22_X1 U21068 ( .A1(n17870), .A2(n17869), .B1(n18171), .B2(n18205), .ZN(
        P3_U2676) );
  INV_X1 U21069 ( .A(n17885), .ZN(n17871) );
  NOR2_X1 U21070 ( .A1(n17872), .A2(n17871), .ZN(n17880) );
  AOI21_X1 U21071 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n18163), .A(n17880), .ZN(
        n17876) );
  OAI21_X1 U21072 ( .B1(n17875), .B2(n17874), .A(n17873), .ZN(n18210) );
  OAI22_X1 U21073 ( .A1(n17877), .A2(n17876), .B1(n18171), .B2(n18210), .ZN(
        P3_U2677) );
  AOI21_X1 U21074 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n18163), .A(n17885), .ZN(
        n17879) );
  XNOR2_X1 U21075 ( .A(n17878), .B(n17881), .ZN(n18215) );
  OAI22_X1 U21076 ( .A1(n17880), .A2(n17879), .B1(n18171), .B2(n18215), .ZN(
        P3_U2678) );
  AOI21_X1 U21077 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n18163), .A(n17890), .ZN(
        n17884) );
  OAI21_X1 U21078 ( .B1(n17883), .B2(n17882), .A(n17881), .ZN(n18220) );
  OAI22_X1 U21079 ( .A1(n17885), .A2(n17884), .B1(n18171), .B2(n18220), .ZN(
        P3_U2679) );
  NOR3_X1 U21080 ( .A1(n17886), .A2(n17891), .A3(n17927), .ZN(n17909) );
  AOI21_X1 U21081 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n18163), .A(n17909), .ZN(
        n17889) );
  XNOR2_X1 U21082 ( .A(n17888), .B(n17887), .ZN(n18224) );
  OAI22_X1 U21083 ( .A1(n17890), .A2(n17889), .B1(n18171), .B2(n18224), .ZN(
        P3_U2680) );
  NOR2_X1 U21084 ( .A1(n17891), .A2(n17927), .ZN(n17892) );
  AOI21_X1 U21085 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n18163), .A(n17892), .ZN(
        n17908) );
  NOR2_X1 U21086 ( .A1(n18135), .A2(n17893), .ZN(n17896) );
  OAI22_X1 U21087 ( .A1(n9620), .A2(n17894), .B1(n18138), .B2(n18034), .ZN(
        n17895) );
  AOI211_X1 U21088 ( .C1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .C2(n18112), .A(
        n17896), .B(n17895), .ZN(n17901) );
  AOI22_X1 U21089 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17900) );
  NAND2_X1 U21090 ( .A1(n17897), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n17899) );
  INV_X1 U21091 ( .A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n18031) );
  OR2_X1 U21092 ( .A1(n18086), .A2(n18031), .ZN(n17898) );
  NAND4_X1 U21093 ( .A1(n17901), .A2(n17900), .A3(n17899), .A4(n17898), .ZN(
        n17907) );
  AOI22_X1 U21094 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17905) );
  AOI22_X1 U21095 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n18056), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17904) );
  AOI22_X1 U21096 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17903) );
  AOI22_X1 U21097 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17902) );
  NAND4_X1 U21098 ( .A1(n17905), .A2(n17904), .A3(n17903), .A4(n17902), .ZN(
        n17906) );
  NOR2_X1 U21099 ( .A1(n17907), .A2(n17906), .ZN(n18226) );
  OAI22_X1 U21100 ( .A1(n17909), .A2(n17908), .B1(n18226), .B2(n18163), .ZN(
        P3_U2681) );
  NOR2_X1 U21101 ( .A1(n18177), .A2(n17910), .ZN(n17940) );
  AOI22_X1 U21102 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17914) );
  AOI22_X1 U21103 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17913) );
  AOI22_X1 U21104 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17912) );
  AOI22_X1 U21105 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17911) );
  NAND4_X1 U21106 ( .A1(n17914), .A2(n17913), .A3(n17912), .A4(n17911), .ZN(
        n17925) );
  AOI22_X1 U21107 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17916) );
  NAND2_X1 U21108 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n17915) );
  OAI211_X1 U21109 ( .C1(n17917), .C2(n18135), .A(n17916), .B(n17915), .ZN(
        n17924) );
  INV_X1 U21110 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17918) );
  OAI22_X1 U21111 ( .A1(n18067), .A2(n17919), .B1(n18138), .B2(n17918), .ZN(
        n17923) );
  INV_X1 U21112 ( .A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17921) );
  OAI22_X1 U21113 ( .A1(n17112), .A2(n17921), .B1(n18141), .B2(n17920), .ZN(
        n17922) );
  OR4_X1 U21114 ( .A1(n17925), .A2(n17924), .A3(n17923), .A4(n17922), .ZN(
        n18231) );
  AOI22_X1 U21115 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17940), .B1(n18177), 
        .B2(n18231), .ZN(n17926) );
  OAI21_X1 U21116 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17927), .A(n17926), .ZN(
        P3_U2682) );
  INV_X1 U21117 ( .A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17929) );
  AOI22_X1 U21118 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17928) );
  OAI21_X1 U21119 ( .B1(n18067), .B2(n17929), .A(n17928), .ZN(n17930) );
  AOI21_X1 U21120 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n17930), .ZN(n17933) );
  AOI22_X1 U21121 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17932) );
  AOI22_X1 U21122 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17931) );
  NAND3_X1 U21123 ( .A1(n17933), .A2(n17932), .A3(n17931), .ZN(n17939) );
  AOI22_X1 U21124 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17937) );
  AOI22_X1 U21125 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17936) );
  AOI22_X1 U21126 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17935) );
  AOI22_X1 U21127 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17934) );
  NAND4_X1 U21128 ( .A1(n17937), .A2(n17936), .A3(n17935), .A4(n17934), .ZN(
        n17938) );
  NOR2_X1 U21129 ( .A1(n17939), .A2(n17938), .ZN(n18237) );
  OAI21_X1 U21130 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17941), .A(n17940), .ZN(
        n17942) );
  OAI21_X1 U21131 ( .B1(n18237), .B2(n18163), .A(n17942), .ZN(P3_U2683) );
  INV_X1 U21132 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17944) );
  AOI22_X1 U21133 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17943) );
  OAI21_X1 U21134 ( .B1(n17112), .B2(n17944), .A(n17943), .ZN(n17945) );
  AOI21_X1 U21135 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n17945), .ZN(n17948) );
  AOI22_X1 U21136 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17947) );
  AOI22_X1 U21137 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17946) );
  NAND3_X1 U21138 ( .A1(n17948), .A2(n17947), .A3(n17946), .ZN(n17954) );
  AOI22_X1 U21139 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17952) );
  AOI22_X1 U21140 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U21141 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17950) );
  AOI22_X1 U21142 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17949) );
  NAND4_X1 U21143 ( .A1(n17952), .A2(n17951), .A3(n17950), .A4(n17949), .ZN(
        n17953) );
  NOR2_X1 U21144 ( .A1(n17954), .A2(n17953), .ZN(n18245) );
  OAI21_X1 U21145 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17972), .A(n17955), .ZN(
        n17956) );
  AOI22_X1 U21146 ( .A1(n18177), .A2(n18245), .B1(n17956), .B2(n18163), .ZN(
        P3_U2684) );
  NOR3_X1 U21147 ( .A1(n19024), .A2(n18006), .A3(n18026), .ZN(n17989) );
  NAND2_X1 U21148 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17989), .ZN(n17988) );
  AOI22_X1 U21149 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17960) );
  AOI22_X1 U21150 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17959) );
  AOI22_X1 U21151 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17958) );
  AOI22_X1 U21152 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17957) );
  NAND4_X1 U21153 ( .A1(n17960), .A2(n17959), .A3(n17958), .A4(n17957), .ZN(
        n17971) );
  AOI22_X1 U21154 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17962) );
  NAND2_X1 U21155 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n17961) );
  OAI211_X1 U21156 ( .C1(n17963), .C2(n18135), .A(n17962), .B(n17961), .ZN(
        n17970) );
  INV_X1 U21157 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17965) );
  INV_X1 U21158 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17964) );
  OAI22_X1 U21159 ( .A1(n18067), .A2(n17965), .B1(n18138), .B2(n17964), .ZN(
        n17969) );
  INV_X1 U21160 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17967) );
  INV_X1 U21161 ( .A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17966) );
  OAI22_X1 U21162 ( .A1(n17112), .A2(n17967), .B1(n18141), .B2(n17966), .ZN(
        n17968) );
  OR4_X1 U21163 ( .A1(n17971), .A2(n17970), .A3(n17969), .A4(n17968), .ZN(
        n18246) );
  OAI21_X1 U21164 ( .B1(n17973), .B2(n17972), .A(n18171), .ZN(n17974) );
  OAI21_X1 U21165 ( .B1(n18163), .B2(n18246), .A(n17974), .ZN(n17975) );
  OAI21_X1 U21166 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17988), .A(n17975), .ZN(
        P3_U2685) );
  INV_X1 U21167 ( .A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17977) );
  AOI22_X1 U21168 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17976) );
  OAI21_X1 U21169 ( .B1(n18067), .B2(n17977), .A(n17976), .ZN(n17978) );
  AOI21_X1 U21170 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n17978), .ZN(n17981) );
  AOI22_X1 U21171 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17980) );
  AOI22_X1 U21172 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17979) );
  NAND3_X1 U21173 ( .A1(n17981), .A2(n17980), .A3(n17979), .ZN(n17987) );
  AOI22_X1 U21174 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17985) );
  AOI22_X1 U21175 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17984) );
  AOI22_X1 U21176 ( .A1(n18092), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U21177 ( .A1(n18091), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17982) );
  NAND4_X1 U21178 ( .A1(n17985), .A2(n17984), .A3(n17983), .A4(n17982), .ZN(
        n17986) );
  NOR2_X1 U21179 ( .A1(n17987), .A2(n17986), .ZN(n18256) );
  OAI211_X1 U21180 ( .C1(n17989), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18163), .B(
        n17988), .ZN(n17990) );
  OAI21_X1 U21181 ( .B1(n18256), .B2(n18163), .A(n17990), .ZN(P3_U2686) );
  INV_X1 U21182 ( .A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n21618) );
  AOI22_X1 U21183 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17992) );
  NAND2_X1 U21184 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n17991) );
  OAI211_X1 U21185 ( .C1(n21618), .C2(n18086), .A(n17992), .B(n17991), .ZN(
        n17999) );
  INV_X1 U21186 ( .A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17994) );
  OAI22_X1 U21187 ( .A1(n9620), .A2(n17994), .B1(n18135), .B2(n17993), .ZN(
        n17998) );
  INV_X1 U21188 ( .A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n18142) );
  INV_X1 U21189 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17995) );
  OAI22_X1 U21190 ( .A1(n17996), .A2(n18142), .B1(n18030), .B2(n17995), .ZN(
        n17997) );
  OR3_X1 U21191 ( .A1(n17999), .A2(n17998), .A3(n17997), .ZN(n18005) );
  AOI22_X1 U21192 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18003) );
  AOI22_X1 U21193 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18002) );
  AOI22_X1 U21194 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n18001) );
  AOI22_X1 U21195 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18000) );
  NAND4_X1 U21196 ( .A1(n18003), .A2(n18002), .A3(n18001), .A4(n18000), .ZN(
        n18004) );
  NOR2_X1 U21197 ( .A1(n18005), .A2(n18004), .ZN(n18263) );
  NAND2_X1 U21198 ( .A1(n18120), .A2(n18180), .ZN(n18174) );
  OAI22_X1 U21199 ( .A1(n18177), .A2(n9570), .B1(P3_EBX_REG_15__SCAN_IN), .B2(
        n18174), .ZN(n18008) );
  NOR2_X1 U21200 ( .A1(n19024), .A2(n18026), .ZN(n18007) );
  AOI22_X1 U21201 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n18008), .B1(n18007), 
        .B2(n18006), .ZN(n18009) );
  OAI21_X1 U21202 ( .B1(n18263), .B2(n18163), .A(n18009), .ZN(P3_U2687) );
  INV_X1 U21203 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n18012) );
  AOI22_X1 U21204 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n18011) );
  NAND2_X1 U21205 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n18010) );
  OAI211_X1 U21206 ( .C1(n18135), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        n18019) );
  INV_X1 U21207 ( .A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n18013) );
  OAI22_X1 U21208 ( .A1(n9626), .A2(n18014), .B1(n18138), .B2(n18013), .ZN(
        n18018) );
  INV_X1 U21209 ( .A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n18015) );
  OAI22_X1 U21210 ( .A1(n18141), .A2(n18016), .B1(n18030), .B2(n18015), .ZN(
        n18017) );
  OR3_X1 U21211 ( .A1(n18019), .A2(n18018), .A3(n18017), .ZN(n18025) );
  AOI22_X1 U21212 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n18023) );
  AOI22_X1 U21213 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18080), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n18022) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9573), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n18021) );
  AOI22_X1 U21215 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18020) );
  NAND4_X1 U21216 ( .A1(n18023), .A2(n18022), .A3(n18021), .A4(n18020), .ZN(
        n18024) );
  NOR2_X1 U21217 ( .A1(n18025), .A2(n18024), .ZN(n18269) );
  OAI21_X1 U21218 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n9570), .A(n18026), .ZN(
        n18027) );
  AOI22_X1 U21219 ( .A1(n18177), .A2(n18269), .B1(n18027), .B2(n18163), .ZN(
        P3_U2688) );
  AOI22_X1 U21220 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n18029) );
  NAND2_X1 U21221 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n18028) );
  OAI211_X1 U21222 ( .C1(n18031), .C2(n18030), .A(n18029), .B(n18028), .ZN(
        n18039) );
  INV_X1 U21223 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n18033) );
  INV_X1 U21224 ( .A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n18032) );
  OAI22_X1 U21225 ( .A1(n9620), .A2(n18033), .B1(n18141), .B2(n18032), .ZN(
        n18038) );
  OAI22_X1 U21226 ( .A1(n9626), .A2(n18036), .B1(n18035), .B2(n18034), .ZN(
        n18037) );
  OR3_X1 U21227 ( .A1(n18039), .A2(n18038), .A3(n18037), .ZN(n18045) );
  AOI22_X1 U21228 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n18043) );
  AOI22_X1 U21229 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n18111), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n18042) );
  AOI22_X1 U21230 ( .A1(n18123), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n18041) );
  AOI22_X1 U21231 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n18040) );
  NAND4_X1 U21232 ( .A1(n18043), .A2(n18042), .A3(n18041), .A4(n18040), .ZN(
        n18044) );
  NOR2_X1 U21233 ( .A1(n18045), .A2(n18044), .ZN(n18271) );
  NOR2_X1 U21234 ( .A1(n18177), .A2(n9570), .ZN(n18047) );
  OAI221_X1 U21235 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n18048), .C1(
        P3_EBX_REG_14__SCAN_IN), .C2(P3_EBX_REG_13__SCAN_IN), .A(n18047), .ZN(
        n18049) );
  OAI21_X1 U21236 ( .B1(n18271), .B2(n18163), .A(n18049), .ZN(P3_U2689) );
  NOR2_X1 U21237 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n18079), .ZN(n18064) );
  AOI22_X1 U21238 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n18050) );
  OAI21_X1 U21239 ( .B1(n18135), .B2(n18051), .A(n18050), .ZN(n18052) );
  AOI21_X1 U21240 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A(
        n18052), .ZN(n18055) );
  AOI22_X1 U21241 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n18054) );
  AOI22_X1 U21242 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n18053) );
  NAND3_X1 U21243 ( .A1(n18055), .A2(n18054), .A3(n18053), .ZN(n18062) );
  AOI22_X1 U21244 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n18060) );
  AOI22_X1 U21245 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18059) );
  AOI22_X1 U21246 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n18058) );
  AOI22_X1 U21247 ( .A1(n18091), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n18057) );
  NAND4_X1 U21248 ( .A1(n18060), .A2(n18059), .A3(n18058), .A4(n18057), .ZN(
        n18061) );
  NOR2_X1 U21249 ( .A1(n18062), .A2(n18061), .ZN(n18279) );
  OAI22_X1 U21250 ( .A1(n18064), .A2(n18063), .B1(n18279), .B2(n18171), .ZN(
        P3_U2691) );
  INV_X1 U21251 ( .A(n18099), .ZN(n18065) );
  OAI21_X1 U21252 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n18065), .A(n18171), .ZN(
        n18078) );
  INV_X1 U21253 ( .A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n21609) );
  AOI22_X1 U21254 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n18066) );
  OAI21_X1 U21255 ( .B1(n18067), .B2(n21609), .A(n18066), .ZN(n18068) );
  AOI21_X1 U21256 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A(
        n18068), .ZN(n18071) );
  AOI22_X1 U21257 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9580), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18070) );
  AOI22_X1 U21258 ( .A1(n13168), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n18069) );
  NAND3_X1 U21259 ( .A1(n18071), .A2(n18070), .A3(n18069), .ZN(n18077) );
  AOI22_X1 U21260 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n18075) );
  AOI22_X1 U21261 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n18074) );
  AOI22_X1 U21262 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n18073) );
  AOI22_X1 U21263 ( .A1(n18122), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n18072) );
  NAND4_X1 U21264 ( .A1(n18075), .A2(n18074), .A3(n18073), .A4(n18072), .ZN(
        n18076) );
  NOR2_X1 U21265 ( .A1(n18077), .A2(n18076), .ZN(n18282) );
  OAI22_X1 U21266 ( .A1(n18079), .A2(n18078), .B1(n18282), .B2(n18171), .ZN(
        P3_U2692) );
  AOI22_X1 U21267 ( .A1(n18080), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n18090) );
  NAND2_X1 U21268 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n18084) );
  NAND2_X1 U21269 ( .A1(n18081), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n18083) );
  NAND2_X1 U21270 ( .A1(n13412), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n18082) );
  AND3_X1 U21271 ( .A1(n18084), .A2(n18083), .A3(n18082), .ZN(n18089) );
  AOI22_X1 U21272 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n18088) );
  INV_X1 U21273 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18085) );
  OR2_X1 U21274 ( .A1(n18086), .A2(n18085), .ZN(n18087) );
  NAND4_X1 U21275 ( .A1(n18090), .A2(n18089), .A3(n18088), .A4(n18087), .ZN(
        n18098) );
  AOI22_X1 U21276 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n18091), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n18096) );
  AOI22_X1 U21277 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n18095) );
  AOI22_X1 U21278 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n18092), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18094) );
  AOI22_X1 U21279 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n18093) );
  NAND4_X1 U21280 ( .A1(n18096), .A2(n18095), .A3(n18094), .A4(n18093), .ZN(
        n18097) );
  OR2_X1 U21281 ( .A1(n18098), .A2(n18097), .ZN(n18286) );
  INV_X1 U21282 ( .A(n18286), .ZN(n18101) );
  OAI21_X1 U21283 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n9595), .A(n18099), .ZN(
        n18100) );
  AOI22_X1 U21284 ( .A1(n18177), .A2(n18101), .B1(n18100), .B2(n18163), .ZN(
        P3_U2693) );
  OAI21_X1 U21285 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n9735), .A(n18171), .ZN(
        n18119) );
  AOI22_X1 U21286 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n18103) );
  OAI21_X1 U21287 ( .B1(n10442), .B2(n18104), .A(n18103), .ZN(n18105) );
  AOI21_X1 U21288 ( .B1(n18132), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A(
        n18105), .ZN(n18110) );
  AOI22_X1 U21289 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18109) );
  AOI22_X1 U21290 ( .A1(n18107), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n18106), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n18108) );
  NAND3_X1 U21291 ( .A1(n18110), .A2(n18109), .A3(n18108), .ZN(n18118) );
  AOI22_X1 U21292 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n18116) );
  AOI22_X1 U21293 ( .A1(n18111), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13168), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n18115) );
  AOI22_X1 U21294 ( .A1(n18056), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n18112), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n18114) );
  AOI22_X1 U21295 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13412), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n18113) );
  NAND4_X1 U21296 ( .A1(n18116), .A2(n18115), .A3(n18114), .A4(n18113), .ZN(
        n18117) );
  NOR2_X1 U21297 ( .A1(n18118), .A2(n18117), .ZN(n18291) );
  OAI22_X1 U21298 ( .A1(n9595), .A2(n18119), .B1(n18291), .B2(n18171), .ZN(
        P3_U2694) );
  NAND2_X1 U21299 ( .A1(n18120), .A2(n18121), .ZN(n18148) );
  NOR2_X1 U21300 ( .A1(n18177), .A2(n18121), .ZN(n18149) );
  AOI22_X1 U21301 ( .A1(n18106), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n18122), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n18130) );
  AOI22_X1 U21302 ( .A1(n18102), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n18123), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n18129) );
  AOI22_X1 U21303 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n18124), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18128) );
  AOI22_X1 U21304 ( .A1(n9580), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n18125), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n18127) );
  NAND4_X1 U21305 ( .A1(n18130), .A2(n18129), .A3(n18128), .A4(n18127), .ZN(
        n18146) );
  AOI22_X1 U21306 ( .A1(n9573), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n18131), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n18134) );
  NAND2_X1 U21307 ( .A1(n18132), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n18133) );
  OAI211_X1 U21308 ( .C1(n18136), .C2(n18135), .A(n18134), .B(n18133), .ZN(
        n18145) );
  INV_X1 U21309 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n18139) );
  OAI22_X1 U21310 ( .A1(n18067), .A2(n18139), .B1(n18138), .B2(n18137), .ZN(
        n18144) );
  INV_X1 U21311 ( .A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n18140) );
  OAI22_X1 U21312 ( .A1(n17112), .A2(n18142), .B1(n18141), .B2(n18140), .ZN(
        n18143) );
  OR4_X1 U21313 ( .A1(n18146), .A2(n18145), .A3(n18144), .A4(n18143), .ZN(
        n18294) );
  AOI22_X1 U21314 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18149), .B1(n18177), .B2(
        n18294), .ZN(n18147) );
  OAI21_X1 U21315 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n18148), .A(n18147), .ZN(
        P3_U2695) );
  OAI21_X1 U21316 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n9979), .A(n18149), .ZN(
        n18150) );
  OAI21_X1 U21317 ( .B1(n18171), .B2(n18151), .A(n18150), .ZN(P3_U2696) );
  INV_X1 U21318 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18154) );
  OAI21_X1 U21319 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n18158), .A(n18152), .ZN(
        n18153) );
  AOI22_X1 U21320 ( .A1(n18177), .A2(n18154), .B1(n18153), .B2(n18163), .ZN(
        P3_U2697) );
  INV_X1 U21321 ( .A(n18155), .ZN(n18162) );
  OAI21_X1 U21322 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n18162), .A(n18171), .ZN(
        n18157) );
  OAI22_X1 U21323 ( .A1(n18158), .A2(n18157), .B1(n18156), .B2(n18171), .ZN(
        P3_U2698) );
  INV_X1 U21324 ( .A(n18174), .ZN(n18176) );
  AOI22_X1 U21325 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n18163), .B1(n18159), .B2(
        n18176), .ZN(n18161) );
  INV_X1 U21326 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18160) );
  OAI22_X1 U21327 ( .A1(n18162), .A2(n18161), .B1(n18160), .B2(n18171), .ZN(
        P3_U2699) );
  OR2_X1 U21328 ( .A1(n18168), .A2(n18174), .ZN(n18166) );
  INV_X1 U21329 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18165) );
  NAND3_X1 U21330 ( .A1(n18166), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n18163), .ZN(
        n18164) );
  OAI221_X1 U21331 ( .B1(n18166), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n18171), 
        .C2(n18165), .A(n18164), .ZN(P3_U2700) );
  NOR2_X1 U21332 ( .A1(n18179), .A2(n18173), .ZN(n18167) );
  AOI21_X1 U21333 ( .B1(n18180), .B2(n18167), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n18170) );
  OAI21_X1 U21334 ( .B1(n18168), .B2(n18174), .A(n18171), .ZN(n18169) );
  OAI22_X1 U21335 ( .A1(n18170), .A2(n18169), .B1(n18085), .B2(n18171), .ZN(
        P3_U2701) );
  OAI222_X1 U21336 ( .A1(n18175), .A2(n18174), .B1(n18173), .B2(n18180), .C1(
        n18172), .C2(n18171), .ZN(P3_U2702) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18177), .B1(
        n18176), .B2(n18179), .ZN(n18178) );
  OAI21_X1 U21338 ( .B1(n18180), .B2(n18179), .A(n18178), .ZN(P3_U2703) );
  INV_X1 U21339 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18327) );
  INV_X1 U21340 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n18331) );
  INV_X1 U21341 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18362) );
  INV_X1 U21342 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18368) );
  INV_X1 U21343 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n18370) );
  NOR4_X1 U21344 ( .A1(n18362), .A2(n18368), .A3(n18370), .A4(n18372), .ZN(
        n18181) );
  NAND4_X1 U21345 ( .A1(n18182), .A2(P3_EAX_REG_6__SCAN_IN), .A3(
        P3_EAX_REG_5__SCAN_IN), .A4(n18181), .ZN(n18301) );
  NAND2_X1 U21346 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n18296), .ZN(n18295) );
  NAND3_X1 U21347 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .ZN(n18270) );
  NOR2_X1 U21348 ( .A1(n18295), .A2(n18270), .ZN(n18184) );
  INV_X1 U21349 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n18428) );
  INV_X1 U21350 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n18388) );
  INV_X1 U21351 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n18341) );
  NOR2_X1 U21352 ( .A1(n18388), .A2(n18341), .ZN(n18185) );
  NAND4_X1 U21353 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n18185), .ZN(n18225) );
  INV_X1 U21354 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n18338) );
  NAND2_X1 U21355 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n18217), .ZN(n18216) );
  NAND2_X1 U21356 ( .A1(n18190), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n18189) );
  OAI22_X1 U21357 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n18300), .B1(n18312), 
        .B2(n18190), .ZN(n18187) );
  AOI22_X1 U21358 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18257), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n18187), .ZN(n18188) );
  OAI21_X1 U21359 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n18189), .A(n18188), .ZN(
        P3_U2704) );
  AOI22_X1 U21360 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n18257), .ZN(n18192) );
  OAI211_X1 U21361 ( .C1(n18190), .C2(P3_EAX_REG_30__SCAN_IN), .A(n18316), .B(
        n18189), .ZN(n18191) );
  OAI211_X1 U21362 ( .C1(n18193), .C2(n18318), .A(n18192), .B(n18191), .ZN(
        P3_U2705) );
  AOI22_X1 U21363 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n18257), .ZN(n18196) );
  OAI211_X1 U21364 ( .C1(n9623), .C2(P3_EAX_REG_29__SCAN_IN), .A(n18316), .B(
        n18194), .ZN(n18195) );
  OAI211_X1 U21365 ( .C1(n18318), .C2(n18197), .A(n18196), .B(n18195), .ZN(
        P3_U2706) );
  AOI22_X1 U21366 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n18257), .ZN(n18200) );
  AOI211_X1 U21367 ( .C1(n18327), .C2(n18202), .A(n9623), .B(n18312), .ZN(
        n18198) );
  INV_X1 U21368 ( .A(n18198), .ZN(n18199) );
  OAI211_X1 U21369 ( .C1(n18318), .C2(n18201), .A(n18200), .B(n18199), .ZN(
        P3_U2707) );
  AOI22_X1 U21370 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n18257), .ZN(n18204) );
  OAI211_X1 U21371 ( .C1(n18206), .C2(P3_EAX_REG_27__SCAN_IN), .A(n18316), .B(
        n18202), .ZN(n18203) );
  OAI211_X1 U21372 ( .C1(n18318), .C2(n18205), .A(n18204), .B(n18203), .ZN(
        P3_U2708) );
  AOI22_X1 U21373 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n18257), .ZN(n18209) );
  AOI211_X1 U21374 ( .C1(n18331), .C2(n18211), .A(n18206), .B(n18312), .ZN(
        n18207) );
  INV_X1 U21375 ( .A(n18207), .ZN(n18208) );
  OAI211_X1 U21376 ( .C1(n18318), .C2(n18210), .A(n18209), .B(n18208), .ZN(
        P3_U2709) );
  AOI22_X1 U21377 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n18257), .ZN(n18214) );
  OAI211_X1 U21378 ( .C1(n18212), .C2(P3_EAX_REG_25__SCAN_IN), .A(n18316), .B(
        n18211), .ZN(n18213) );
  OAI211_X1 U21379 ( .C1(n18215), .C2(n18318), .A(n18214), .B(n18213), .ZN(
        P3_U2710) );
  AOI22_X1 U21380 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n18257), .ZN(n18219) );
  OAI211_X1 U21381 ( .C1(n18217), .C2(P3_EAX_REG_24__SCAN_IN), .A(n18316), .B(
        n18216), .ZN(n18218) );
  OAI211_X1 U21382 ( .C1(n18220), .C2(n18318), .A(n18219), .B(n18218), .ZN(
        P3_U2711) );
  AOI22_X1 U21383 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n18257), .ZN(n18223) );
  OAI211_X1 U21384 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n9638), .A(n18316), .B(
        n18221), .ZN(n18222) );
  OAI211_X1 U21385 ( .C1(n18224), .C2(n18318), .A(n18223), .B(n18222), .ZN(
        P3_U2712) );
  INV_X1 U21386 ( .A(n18258), .ZN(n18250) );
  NOR3_X1 U21387 ( .A1(n19024), .A2(n18259), .A3(n18225), .ZN(n18229) );
  INV_X1 U21388 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n18343) );
  INV_X1 U21389 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n18383) );
  NAND2_X1 U21390 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n18251), .ZN(n18247) );
  NOR2_X1 U21391 ( .A1(n18343), .A2(n18247), .ZN(n18241) );
  NAND2_X1 U21392 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n18241), .ZN(n18235) );
  NAND2_X1 U21393 ( .A1(n18316), .A2(n18235), .ZN(n18232) );
  OAI21_X1 U21394 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n18300), .A(n18232), .ZN(
        n18228) );
  INV_X1 U21395 ( .A(n18257), .ZN(n18236) );
  OAI22_X1 U21396 ( .A1(n18226), .A2(n18318), .B1(n19021), .B2(n18236), .ZN(
        n18227) );
  AOI221_X1 U21397 ( .B1(n18229), .B2(n18338), .C1(n18228), .C2(
        P3_EAX_REG_22__SCAN_IN), .A(n18227), .ZN(n18230) );
  OAI21_X1 U21398 ( .B1(n19020), .B2(n18250), .A(n18230), .ZN(P3_U2713) );
  AOI22_X1 U21399 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18257), .B1(n18309), .B2(
        n18231), .ZN(n18234) );
  INV_X1 U21400 ( .A(n18232), .ZN(n18239) );
  AOI22_X1 U21401 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18258), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n18239), .ZN(n18233) );
  OAI211_X1 U21402 ( .C1(P3_EAX_REG_21__SCAN_IN), .C2(n18235), .A(n18234), .B(
        n18233), .ZN(P3_U2714) );
  OAI22_X1 U21403 ( .A1(n18237), .A2(n18318), .B1(n20006), .B2(n18236), .ZN(
        n18238) );
  AOI221_X1 U21404 ( .B1(n18239), .B2(P3_EAX_REG_20__SCAN_IN), .C1(n18241), 
        .C2(n18341), .A(n18238), .ZN(n18240) );
  OAI21_X1 U21405 ( .B1(n19013), .B2(n18250), .A(n18240), .ZN(P3_U2715) );
  AOI22_X1 U21406 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18257), .ZN(n18244) );
  AOI211_X1 U21407 ( .C1(n18343), .C2(n18247), .A(n18241), .B(n18312), .ZN(
        n18242) );
  INV_X1 U21408 ( .A(n18242), .ZN(n18243) );
  OAI211_X1 U21409 ( .C1(n18245), .C2(n18318), .A(n18244), .B(n18243), .ZN(
        P3_U2716) );
  AOI22_X1 U21410 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18257), .B1(n18309), .B2(
        n18246), .ZN(n18249) );
  OAI211_X1 U21411 ( .C1(n18251), .C2(P3_EAX_REG_18__SCAN_IN), .A(n18316), .B(
        n18247), .ZN(n18248) );
  OAI211_X1 U21412 ( .C1(n18250), .C2(n19005), .A(n18249), .B(n18248), .ZN(
        P3_U2717) );
  AOI22_X1 U21413 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18257), .ZN(n18255) );
  INV_X1 U21414 ( .A(n18259), .ZN(n18253) );
  INV_X1 U21415 ( .A(n18251), .ZN(n18252) );
  OAI211_X1 U21416 ( .C1(n18253), .C2(P3_EAX_REG_17__SCAN_IN), .A(n18316), .B(
        n18252), .ZN(n18254) );
  OAI211_X1 U21417 ( .C1(n18256), .C2(n18318), .A(n18255), .B(n18254), .ZN(
        P3_U2718) );
  AOI22_X1 U21418 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n18258), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n18257), .ZN(n18262) );
  OAI211_X1 U21419 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n18260), .A(n18316), .B(
        n18259), .ZN(n18261) );
  OAI211_X1 U21420 ( .C1(n18263), .C2(n18318), .A(n18262), .B(n18261), .ZN(
        P3_U2719) );
  NOR2_X1 U21421 ( .A1(n19024), .A2(n18264), .ZN(n18266) );
  NAND2_X1 U21422 ( .A1(n18316), .A2(n18264), .ZN(n18274) );
  INV_X1 U21423 ( .A(n18274), .ZN(n18265) );
  MUX2_X1 U21424 ( .A(n18266), .B(n18265), .S(P3_EAX_REG_15__SCAN_IN), .Z(
        n18267) );
  AOI21_X1 U21425 ( .B1(BUF2_REG_15__SCAN_IN), .B2(n18310), .A(n18267), .ZN(
        n18268) );
  OAI21_X1 U21426 ( .B1(n18269), .B2(n18318), .A(n18268), .ZN(P3_U2720) );
  NOR2_X1 U21427 ( .A1(n19024), .A2(n18295), .ZN(n18290) );
  INV_X1 U21428 ( .A(n18290), .ZN(n18285) );
  NOR2_X1 U21429 ( .A1(n18270), .A2(n18285), .ZN(n18284) );
  NAND2_X1 U21430 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n18281), .ZN(n18276) );
  INV_X1 U21431 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n18423) );
  INV_X1 U21432 ( .A(n18271), .ZN(n18272) );
  AOI22_X1 U21433 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18310), .B1(n18309), .B2(
        n18272), .ZN(n18273) );
  OAI221_X1 U21434 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n18276), .C1(n18423), 
        .C2(n18274), .A(n18273), .ZN(P3_U2721) );
  AOI22_X1 U21435 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18310), .B1(n18309), .B2(
        n18275), .ZN(n18278) );
  OAI211_X1 U21436 ( .C1(n18281), .C2(P3_EAX_REG_13__SCAN_IN), .A(n18316), .B(
        n18276), .ZN(n18277) );
  NAND2_X1 U21437 ( .A1(n18278), .A2(n18277), .ZN(P3_U2722) );
  AOI21_X1 U21438 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n18316), .A(n18284), .ZN(
        n18280) );
  OAI222_X1 U21439 ( .A1(n18321), .A2(n13823), .B1(n18281), .B2(n18280), .C1(
        n18318), .C2(n18279), .ZN(P3_U2723) );
  INV_X1 U21440 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18357) );
  INV_X1 U21441 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n18359) );
  NOR3_X1 U21442 ( .A1(n18357), .A2(n18359), .A3(n18285), .ZN(n18289) );
  AOI21_X1 U21443 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n18316), .A(n18289), .ZN(
        n18283) );
  OAI222_X1 U21444 ( .A1(n18321), .A2(n13842), .B1(n18284), .B2(n18283), .C1(
        n18318), .C2(n18282), .ZN(P3_U2724) );
  NOR2_X1 U21445 ( .A1(n18359), .A2(n18285), .ZN(n18293) );
  OAI21_X1 U21446 ( .B1(P3_EAX_REG_10__SCAN_IN), .B2(n18293), .A(n18316), .ZN(
        n18288) );
  AOI22_X1 U21447 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n18310), .B1(n18309), .B2(
        n18286), .ZN(n18287) );
  OAI21_X1 U21448 ( .B1(n18289), .B2(n18288), .A(n18287), .ZN(P3_U2725) );
  AOI21_X1 U21449 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n18316), .A(n18290), .ZN(
        n18292) );
  OAI222_X1 U21450 ( .A1(n18321), .A2(n13820), .B1(n18293), .B2(n18292), .C1(
        n18318), .C2(n18291), .ZN(P3_U2726) );
  AOI22_X1 U21451 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18310), .B1(n18309), .B2(
        n18294), .ZN(n18298) );
  OAI211_X1 U21452 ( .C1(P3_EAX_REG_8__SCAN_IN), .C2(n18296), .A(n18316), .B(
        n18295), .ZN(n18297) );
  NAND2_X1 U21453 ( .A1(n18298), .A2(n18297), .ZN(P3_U2727) );
  NAND2_X1 U21454 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n18299) );
  NAND2_X1 U21455 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n18315), .ZN(n18314) );
  NOR2_X1 U21456 ( .A1(n18299), .A2(n18314), .ZN(n18307) );
  AOI21_X1 U21457 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n18316), .A(n18307), .ZN(
        n18304) );
  NOR2_X1 U21458 ( .A1(n18301), .A2(n18300), .ZN(n18303) );
  OAI222_X1 U21459 ( .A1(n18321), .A2(n13836), .B1(n18304), .B2(n18303), .C1(
        n18318), .C2(n18302), .ZN(P3_U2728) );
  INV_X1 U21460 ( .A(n18314), .ZN(n18320) );
  AOI22_X1 U21461 ( .A1(n18320), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n18316), .ZN(n18306) );
  OAI222_X1 U21462 ( .A1(n19020), .A2(n18321), .B1(n18307), .B2(n18306), .C1(
        n18318), .C2(n18305), .ZN(P3_U2729) );
  NAND2_X1 U21463 ( .A1(n18314), .A2(P3_EAX_REG_5__SCAN_IN), .ZN(n18313) );
  AOI22_X1 U21464 ( .A1(n18310), .A2(BUF2_REG_5__SCAN_IN), .B1(n18309), .B2(
        n18308), .ZN(n18311) );
  OAI221_X1 U21465 ( .B1(n18314), .B2(P3_EAX_REG_5__SCAN_IN), .C1(n18313), 
        .C2(n18312), .A(n18311), .ZN(P3_U2730) );
  AOI21_X1 U21466 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n18316), .A(n18315), .ZN(
        n18319) );
  OAI222_X1 U21467 ( .A1(n19013), .A2(n18321), .B1(n18320), .B2(n18319), .C1(
        n18318), .C2(n18317), .ZN(P3_U2731) );
  NOR2_X2 U21468 ( .A1(n19451), .A2(n18608), .ZN(n19565) );
  NOR2_X4 U21469 ( .A1(n19565), .A2(n18323), .ZN(n18363) );
  AND2_X1 U21470 ( .A1(n18363), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U21471 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n18400) );
  AOI22_X1 U21472 ( .A1(n19565), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18324) );
  OAI21_X1 U21473 ( .B1(n18400), .B2(n18348), .A(n18324), .ZN(P3_U2737) );
  INV_X1 U21474 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n18398) );
  AOI22_X1 U21475 ( .A1(n19565), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18325) );
  OAI21_X1 U21476 ( .B1(n18398), .B2(n18348), .A(n18325), .ZN(P3_U2738) );
  AOI22_X1 U21477 ( .A1(n19565), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18326) );
  OAI21_X1 U21478 ( .B1(n18327), .B2(n18348), .A(n18326), .ZN(P3_U2739) );
  INV_X1 U21479 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n18329) );
  AOI22_X1 U21480 ( .A1(n19565), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18328) );
  OAI21_X1 U21481 ( .B1(n18329), .B2(n18348), .A(n18328), .ZN(P3_U2740) );
  AOI22_X1 U21482 ( .A1(n19565), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18330) );
  OAI21_X1 U21483 ( .B1(n18331), .B2(n18348), .A(n18330), .ZN(P3_U2741) );
  INV_X1 U21484 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n18333) );
  AOI22_X1 U21485 ( .A1(n19565), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18332) );
  OAI21_X1 U21486 ( .B1(n18333), .B2(n18348), .A(n18332), .ZN(P3_U2742) );
  INV_X1 U21487 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n18392) );
  AOI22_X1 U21488 ( .A1(n19565), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18334) );
  OAI21_X1 U21489 ( .B1(n18392), .B2(n18348), .A(n18334), .ZN(P3_U2743) );
  INV_X1 U21490 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18336) );
  AOI22_X1 U21491 ( .A1(n19565), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18335) );
  OAI21_X1 U21492 ( .B1(n18336), .B2(n18348), .A(n18335), .ZN(P3_U2744) );
  AOI22_X1 U21493 ( .A1(n18374), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18337) );
  OAI21_X1 U21494 ( .B1(n18338), .B2(n18348), .A(n18337), .ZN(P3_U2745) );
  AOI22_X1 U21495 ( .A1(n18374), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18339) );
  OAI21_X1 U21496 ( .B1(n18388), .B2(n18348), .A(n18339), .ZN(P3_U2746) );
  AOI22_X1 U21497 ( .A1(n18374), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18340) );
  OAI21_X1 U21498 ( .B1(n18341), .B2(n18348), .A(n18340), .ZN(P3_U2747) );
  AOI22_X1 U21499 ( .A1(n18374), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18342) );
  OAI21_X1 U21500 ( .B1(n18343), .B2(n18348), .A(n18342), .ZN(P3_U2748) );
  INV_X1 U21501 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n18345) );
  AOI22_X1 U21502 ( .A1(n18374), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18344) );
  OAI21_X1 U21503 ( .B1(n18345), .B2(n18348), .A(n18344), .ZN(P3_U2749) );
  AOI22_X1 U21504 ( .A1(n18374), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18346) );
  OAI21_X1 U21505 ( .B1(n18383), .B2(n18348), .A(n18346), .ZN(P3_U2750) );
  AOI22_X1 U21506 ( .A1(n18374), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18347) );
  OAI21_X1 U21507 ( .B1(n9967), .B2(n18348), .A(n18347), .ZN(P3_U2751) );
  AOI22_X1 U21508 ( .A1(n18374), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18349) );
  OAI21_X1 U21509 ( .B1(n18428), .B2(n18376), .A(n18349), .ZN(P3_U2752) );
  AOI22_X1 U21510 ( .A1(n18374), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18350) );
  OAI21_X1 U21511 ( .B1(n18423), .B2(n18376), .A(n18350), .ZN(P3_U2753) );
  INV_X1 U21512 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18421) );
  AOI22_X1 U21513 ( .A1(n18374), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18351) );
  OAI21_X1 U21514 ( .B1(n18421), .B2(n18376), .A(n18351), .ZN(P3_U2754) );
  INV_X1 U21515 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n18353) );
  AOI22_X1 U21516 ( .A1(n18374), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18352) );
  OAI21_X1 U21517 ( .B1(n18353), .B2(n18376), .A(n18352), .ZN(P3_U2755) );
  INV_X1 U21518 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n18355) );
  AOI22_X1 U21519 ( .A1(n18374), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18354) );
  OAI21_X1 U21520 ( .B1(n18355), .B2(n18376), .A(n18354), .ZN(P3_U2756) );
  AOI22_X1 U21521 ( .A1(n18374), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18356) );
  OAI21_X1 U21522 ( .B1(n18357), .B2(n18376), .A(n18356), .ZN(P3_U2757) );
  AOI22_X1 U21523 ( .A1(n18374), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18358) );
  OAI21_X1 U21524 ( .B1(n18359), .B2(n18376), .A(n18358), .ZN(P3_U2758) );
  INV_X1 U21525 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n18412) );
  AOI22_X1 U21526 ( .A1(n18374), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18360) );
  OAI21_X1 U21527 ( .B1(n18412), .B2(n18376), .A(n18360), .ZN(P3_U2759) );
  AOI22_X1 U21528 ( .A1(n18374), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18361) );
  OAI21_X1 U21529 ( .B1(n18362), .B2(n18376), .A(n18361), .ZN(P3_U2760) );
  INV_X1 U21530 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n18365) );
  AOI22_X1 U21531 ( .A1(n18374), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18364) );
  OAI21_X1 U21532 ( .B1(n18365), .B2(n18376), .A(n18364), .ZN(P3_U2761) );
  INV_X1 U21533 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n18408) );
  AOI22_X1 U21534 ( .A1(n18374), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18366) );
  OAI21_X1 U21535 ( .B1(n18408), .B2(n18376), .A(n18366), .ZN(P3_U2762) );
  AOI22_X1 U21536 ( .A1(n18374), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18367) );
  OAI21_X1 U21537 ( .B1(n18368), .B2(n18376), .A(n18367), .ZN(P3_U2763) );
  AOI22_X1 U21538 ( .A1(n18374), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18369) );
  OAI21_X1 U21539 ( .B1(n18370), .B2(n18376), .A(n18369), .ZN(P3_U2764) );
  AOI22_X1 U21540 ( .A1(n18374), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18371) );
  OAI21_X1 U21541 ( .B1(n18372), .B2(n18376), .A(n18371), .ZN(P3_U2765) );
  AOI22_X1 U21542 ( .A1(n18374), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18373) );
  OAI21_X1 U21543 ( .B1(n18403), .B2(n18376), .A(n18373), .ZN(P3_U2766) );
  AOI22_X1 U21544 ( .A1(n18374), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18363), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18375) );
  OAI21_X1 U21545 ( .B1(n18377), .B2(n18376), .A(n18375), .ZN(P3_U2767) );
  AOI22_X1 U21546 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n18424), .ZN(n18381) );
  OAI21_X1 U21547 ( .B1(n18993), .B2(n18419), .A(n18381), .ZN(P3_U2768) );
  INV_X1 U21548 ( .A(n9566), .ZN(n18427) );
  AOI22_X1 U21549 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18425), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n18424), .ZN(n18382) );
  OAI21_X1 U21550 ( .B1(n18383), .B2(n18427), .A(n18382), .ZN(P3_U2769) );
  AOI22_X1 U21551 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n18424), .ZN(n18384) );
  OAI21_X1 U21552 ( .B1(n19005), .B2(n18419), .A(n18384), .ZN(P3_U2770) );
  AOI22_X1 U21553 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n18424), .ZN(n18385) );
  OAI21_X1 U21554 ( .B1(n19009), .B2(n18419), .A(n18385), .ZN(P3_U2771) );
  AOI22_X1 U21555 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n18424), .ZN(n18386) );
  OAI21_X1 U21556 ( .B1(n19013), .B2(n18419), .A(n18386), .ZN(P3_U2772) );
  AOI22_X1 U21557 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18425), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n18424), .ZN(n18387) );
  OAI21_X1 U21558 ( .B1(n18388), .B2(n18427), .A(n18387), .ZN(P3_U2773) );
  AOI22_X1 U21559 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n18424), .ZN(n18389) );
  OAI21_X1 U21560 ( .B1(n19020), .B2(n18419), .A(n18389), .ZN(P3_U2774) );
  AOI22_X1 U21561 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n18424), .ZN(n18390) );
  OAI21_X1 U21562 ( .B1(n13836), .B2(n18419), .A(n18390), .ZN(P3_U2775) );
  AOI22_X1 U21563 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18425), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n18424), .ZN(n18391) );
  OAI21_X1 U21564 ( .B1(n18392), .B2(n18427), .A(n18391), .ZN(P3_U2776) );
  AOI22_X1 U21565 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n18424), .ZN(n18393) );
  OAI21_X1 U21566 ( .B1(n13820), .B2(n18419), .A(n18393), .ZN(P3_U2777) );
  AOI22_X1 U21567 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n18424), .ZN(n18394) );
  OAI21_X1 U21568 ( .B1(n21539), .B2(n18419), .A(n18394), .ZN(P3_U2778) );
  AOI22_X1 U21569 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n18424), .ZN(n18395) );
  OAI21_X1 U21570 ( .B1(n13842), .B2(n18419), .A(n18395), .ZN(P3_U2779) );
  AOI22_X1 U21571 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n9566), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n18424), .ZN(n18396) );
  OAI21_X1 U21572 ( .B1(n13823), .B2(n18419), .A(n18396), .ZN(P3_U2780) );
  AOI22_X1 U21573 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18425), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n18417), .ZN(n18397) );
  OAI21_X1 U21574 ( .B1(n18398), .B2(n18427), .A(n18397), .ZN(P3_U2781) );
  AOI22_X1 U21575 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18425), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n18417), .ZN(n18399) );
  OAI21_X1 U21576 ( .B1(n18400), .B2(n18427), .A(n18399), .ZN(P3_U2782) );
  AOI22_X1 U21577 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n18424), .ZN(n18401) );
  OAI21_X1 U21578 ( .B1(n18993), .B2(n18419), .A(n18401), .ZN(P3_U2783) );
  AOI22_X1 U21579 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n18417), .ZN(n18402) );
  OAI21_X1 U21580 ( .B1(n18403), .B2(n18427), .A(n18402), .ZN(P3_U2784) );
  AOI22_X1 U21581 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n18424), .ZN(n18404) );
  OAI21_X1 U21582 ( .B1(n19005), .B2(n18419), .A(n18404), .ZN(P3_U2785) );
  AOI22_X1 U21583 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n18417), .ZN(n18405) );
  OAI21_X1 U21584 ( .B1(n19009), .B2(n18419), .A(n18405), .ZN(P3_U2786) );
  AOI22_X1 U21585 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n18424), .ZN(n18406) );
  OAI21_X1 U21586 ( .B1(n19013), .B2(n18419), .A(n18406), .ZN(P3_U2787) );
  AOI22_X1 U21587 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n18417), .ZN(n18407) );
  OAI21_X1 U21588 ( .B1(n18408), .B2(n18427), .A(n18407), .ZN(P3_U2788) );
  AOI22_X1 U21589 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n18424), .ZN(n18409) );
  OAI21_X1 U21590 ( .B1(n19020), .B2(n18419), .A(n18409), .ZN(P3_U2789) );
  AOI22_X1 U21591 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n18424), .ZN(n18410) );
  OAI21_X1 U21592 ( .B1(n13836), .B2(n18419), .A(n18410), .ZN(P3_U2790) );
  AOI22_X1 U21593 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n18424), .ZN(n18411) );
  OAI21_X1 U21594 ( .B1(n18412), .B2(n18427), .A(n18411), .ZN(P3_U2791) );
  AOI22_X1 U21595 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n18417), .ZN(n18414) );
  OAI21_X1 U21596 ( .B1(n13820), .B2(n18419), .A(n18414), .ZN(P3_U2792) );
  AOI22_X1 U21597 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n18417), .ZN(n18415) );
  OAI21_X1 U21598 ( .B1(n21539), .B2(n18419), .A(n18415), .ZN(P3_U2793) );
  AOI22_X1 U21599 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n18417), .ZN(n18416) );
  OAI21_X1 U21600 ( .B1(n13842), .B2(n18419), .A(n18416), .ZN(P3_U2794) );
  AOI22_X1 U21601 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n9566), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n18417), .ZN(n18418) );
  OAI21_X1 U21602 ( .B1(n13823), .B2(n18419), .A(n18418), .ZN(P3_U2795) );
  AOI22_X1 U21603 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n18424), .ZN(n18420) );
  OAI21_X1 U21604 ( .B1(n18421), .B2(n18427), .A(n18420), .ZN(P3_U2796) );
  AOI22_X1 U21605 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n18424), .ZN(n18422) );
  OAI21_X1 U21606 ( .B1(n18423), .B2(n18427), .A(n18422), .ZN(P3_U2797) );
  AOI22_X1 U21607 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n18425), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n18424), .ZN(n18426) );
  OAI21_X1 U21608 ( .B1(n18428), .B2(n18427), .A(n18426), .ZN(P3_U2798) );
  NOR2_X1 U21609 ( .A1(n18430), .A2(n18429), .ZN(n18457) );
  NAND3_X1 U21610 ( .A1(n18431), .A2(n18432), .A3(n10228), .ZN(n18453) );
  NAND2_X1 U21611 ( .A1(n18457), .A2(n18453), .ZN(n18436) );
  NOR3_X1 U21612 ( .A1(n18610), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        n18433), .ZN(n18434) );
  AOI211_X1 U21613 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n18436), .A(
        n18435), .B(n18434), .ZN(n18444) );
  NOR2_X1 U21614 ( .A1(n18437), .A2(n18579), .ZN(n18456) );
  NOR2_X1 U21615 ( .A1(n18645), .A2(n18647), .ZN(n18520) );
  OAI21_X1 U21616 ( .B1(n18440), .B2(n18439), .A(n18681), .ZN(n18442) );
  INV_X1 U21617 ( .A(n18446), .ZN(n18449) );
  NOR2_X1 U21618 ( .A1(n18447), .A2(n18449), .ZN(n18448) );
  MUX2_X1 U21619 ( .A(n18449), .B(n18448), .S(n18565), .Z(n18451) );
  AOI22_X1 U21620 ( .A1(n18954), .A2(P3_REIP_REG_27__SCAN_IN), .B1(n18529), 
        .B2(n18452), .ZN(n18454) );
  XNOR2_X1 U21621 ( .A(n18743), .B(n18458), .ZN(n18749) );
  INV_X1 U21622 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n18462) );
  AOI211_X1 U21623 ( .C1(n18460), .C2(n18462), .A(n18610), .B(n18459), .ZN(
        n18466) );
  NOR2_X1 U21624 ( .A1(n18981), .A2(n19524), .ZN(n18734) );
  OAI22_X1 U21625 ( .A1(n18463), .A2(n18462), .B1(n18622), .B2(n18461), .ZN(
        n18464) );
  AOI211_X1 U21626 ( .C1(n18466), .C2(n18465), .A(n18734), .B(n18464), .ZN(
        n18473) );
  NAND2_X1 U21627 ( .A1(n18467), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18468) );
  XNOR2_X1 U21628 ( .A(n18468), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18739) );
  NAND2_X1 U21629 ( .A1(n18470), .A2(n18469), .ZN(n18471) );
  XNOR2_X1 U21630 ( .A(n18471), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n18745) );
  AOI22_X1 U21631 ( .A1(n18645), .A2(n18739), .B1(n18681), .B2(n18745), .ZN(
        n18472) );
  OAI211_X1 U21632 ( .C1(n18727), .C2(n18749), .A(n18473), .B(n18472), .ZN(
        P3_U2805) );
  INV_X1 U21633 ( .A(n18489), .ZN(n18475) );
  NAND2_X1 U21634 ( .A1(n18565), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18474) );
  OAI211_X1 U21635 ( .C1(n18476), .C2(n18475), .A(n18522), .B(n18474), .ZN(
        n18477) );
  XNOR2_X1 U21636 ( .A(n18477), .B(n18750), .ZN(n18755) );
  NOR2_X1 U21637 ( .A1(n18478), .A2(n18579), .ZN(n18487) );
  AOI22_X1 U21638 ( .A1(n18954), .A2(P3_REIP_REG_23__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18479), .ZN(n18483) );
  OAI21_X1 U21639 ( .B1(n18529), .B2(n18481), .A(n18480), .ZN(n18482) );
  OAI211_X1 U21640 ( .C1(n18484), .C2(n10441), .A(n18483), .B(n18482), .ZN(
        n18485) );
  AOI221_X1 U21641 ( .B1(n18487), .B2(n18750), .C1(n18486), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n18485), .ZN(n18488) );
  OAI21_X1 U21642 ( .B1(n18653), .B2(n18755), .A(n18488), .ZN(P3_U2807) );
  INV_X1 U21643 ( .A(n18772), .ZN(n18490) );
  OAI21_X1 U21644 ( .B1(n18510), .B2(n18490), .A(n18489), .ZN(n18491) );
  NAND2_X1 U21645 ( .A1(n18522), .A2(n18491), .ZN(n18492) );
  XNOR2_X1 U21646 ( .A(n18492), .B(n18765), .ZN(n18778) );
  AOI22_X1 U21647 ( .A1(n18645), .A2(n18844), .B1(n18647), .B2(n18843), .ZN(
        n18578) );
  OAI21_X1 U21648 ( .B1(n18772), .B2(n18520), .A(n18578), .ZN(n18513) );
  OAI21_X1 U21649 ( .B1(n18493), .B2(n18608), .A(n18708), .ZN(n18494) );
  AOI21_X1 U21650 ( .B1(n18606), .B2(n18497), .A(n18494), .ZN(n18516) );
  OAI21_X1 U21651 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n18495), .A(
        n18516), .ZN(n18506) );
  AOI22_X1 U21652 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18506), .B1(
        n18529), .B2(n18496), .ZN(n18500) );
  NOR2_X1 U21653 ( .A1(n18610), .A2(n18497), .ZN(n18508) );
  OAI211_X1 U21654 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n18508), .B(n18498), .ZN(n18499) );
  OAI211_X1 U21655 ( .C1(n21548), .C2(n18981), .A(n18500), .B(n18499), .ZN(
        n18501) );
  AOI21_X1 U21656 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18513), .A(
        n18501), .ZN(n18503) );
  NAND3_X1 U21657 ( .A1(n18772), .A2(n18559), .A3(n18765), .ZN(n18502) );
  OAI211_X1 U21658 ( .C1(n18653), .C2(n18778), .A(n18503), .B(n18502), .ZN(
        P3_U2808) );
  NAND2_X1 U21659 ( .A1(n18784), .A2(n18770), .ZN(n18788) );
  INV_X1 U21660 ( .A(n18757), .ZN(n18780) );
  NAND2_X1 U21661 ( .A1(n18780), .A2(n18559), .ZN(n18534) );
  OAI22_X1 U21662 ( .A1(n18981), .A2(n19518), .B1(n18622), .B2(n18504), .ZN(
        n18505) );
  AOI221_X1 U21663 ( .B1(n18508), .B2(n18507), .C1(n18506), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n18505), .ZN(n18515) );
  INV_X1 U21664 ( .A(n18548), .ZN(n18531) );
  OR4_X1 U21665 ( .A1(n18510), .A2(n18818), .A3(n18565), .A4(n18509), .ZN(
        n18532) );
  INV_X1 U21666 ( .A(n18532), .ZN(n18523) );
  AOI22_X1 U21667 ( .A1(n18531), .A2(n18511), .B1(n18784), .B2(n18523), .ZN(
        n18512) );
  XNOR2_X1 U21668 ( .A(n18512), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18781) );
  AOI22_X1 U21669 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18513), .B1(
        n18681), .B2(n18781), .ZN(n18514) );
  OAI211_X1 U21670 ( .C1(n18788), .C2(n18534), .A(n18515), .B(n18514), .ZN(
        P3_U2809) );
  NAND2_X1 U21671 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21624), .ZN(
        n18798) );
  AOI221_X1 U21672 ( .B1(n9624), .B2(n18517), .C1(n19180), .C2(n18517), .A(
        n18516), .ZN(n18518) );
  INV_X1 U21673 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19515) );
  NOR2_X1 U21674 ( .A1(n18981), .A2(n19515), .ZN(n18789) );
  AOI211_X1 U21675 ( .C1(n18519), .C2(n18714), .A(n18518), .B(n18789), .ZN(
        n18526) );
  NOR2_X1 U21676 ( .A1(n18757), .A2(n18800), .ZN(n18758) );
  OAI21_X1 U21677 ( .B1(n18520), .B2(n18758), .A(n18578), .ZN(n18536) );
  INV_X1 U21678 ( .A(n18530), .ZN(n18547) );
  NAND2_X1 U21679 ( .A1(n18547), .A2(n18800), .ZN(n18521) );
  OAI211_X1 U21680 ( .C1(n18800), .C2(n18523), .A(n18522), .B(n18521), .ZN(
        n18524) );
  XNOR2_X1 U21681 ( .A(n18524), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18790) );
  AOI22_X1 U21682 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n18536), .B1(
        n18681), .B2(n18790), .ZN(n18525) );
  OAI211_X1 U21683 ( .C1(n18534), .C2(n18798), .A(n18526), .B(n18525), .ZN(
        P3_U2810) );
  AOI21_X1 U21684 ( .B1(n18606), .B2(n18537), .A(n18722), .ZN(n18560) );
  OAI21_X1 U21685 ( .B1(n18527), .B2(n18608), .A(n18560), .ZN(n18544) );
  AOI22_X1 U21686 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18544), .B1(
        n18529), .B2(n18528), .ZN(n18541) );
  NAND2_X1 U21687 ( .A1(n18531), .A2(n18530), .ZN(n18551) );
  NAND2_X1 U21688 ( .A1(n18551), .A2(n18532), .ZN(n18533) );
  XOR2_X1 U21689 ( .A(n18800), .B(n18533), .Z(n18805) );
  OAI22_X1 U21690 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18534), .B1(
        n18805), .B2(n18653), .ZN(n18535) );
  AOI21_X1 U21691 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n18536), .A(
        n18535), .ZN(n18540) );
  NAND2_X1 U21692 ( .A1(n18954), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18803) );
  NOR2_X1 U21693 ( .A1(n18610), .A2(n18537), .ZN(n18546) );
  OAI211_X1 U21694 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n18546), .B(n18538), .ZN(n18539) );
  NAND4_X1 U21695 ( .A1(n18541), .A2(n18540), .A3(n18803), .A4(n18539), .ZN(
        P3_U2811) );
  NAND2_X1 U21696 ( .A1(n18813), .A2(n18818), .ZN(n18824) );
  OAI22_X1 U21697 ( .A1(n18981), .A2(n19511), .B1(n18622), .B2(n18542), .ZN(
        n18543) );
  AOI221_X1 U21698 ( .B1(n18546), .B2(n18545), .C1(n18544), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n18543), .ZN(n18554) );
  OAI21_X1 U21699 ( .B1(n18813), .B2(n18579), .A(n18578), .ZN(n18558) );
  NAND2_X1 U21700 ( .A1(n18659), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18550) );
  NAND2_X1 U21701 ( .A1(n18547), .A2(n18550), .ZN(n18549) );
  MUX2_X1 U21702 ( .A(n18550), .B(n18549), .S(n18548), .Z(n18552) );
  NAND2_X1 U21703 ( .A1(n18552), .A2(n18551), .ZN(n18819) );
  AOI22_X1 U21704 ( .A1(n18558), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n18681), .B2(n18819), .ZN(n18553) );
  OAI211_X1 U21705 ( .C1(n18579), .C2(n18824), .A(n18554), .B(n18553), .ZN(
        P3_U2812) );
  XNOR2_X1 U21706 ( .A(n18555), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18829) );
  INV_X1 U21707 ( .A(n18829), .ZN(n18556) );
  AOI22_X1 U21708 ( .A1(n18714), .A2(n18557), .B1(n18681), .B2(n18556), .ZN(
        n18564) );
  OAI221_X1 U21709 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n18559), .A(n18558), .ZN(
        n18563) );
  NAND2_X1 U21710 ( .A1(n18954), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18831) );
  INV_X1 U21711 ( .A(n18560), .ZN(n18561) );
  OAI221_X1 U21712 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n19351), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n17574), .A(n18561), .ZN(
        n18562) );
  NAND4_X1 U21713 ( .A1(n18564), .A2(n18563), .A3(n18831), .A4(n18562), .ZN(
        P3_U2813) );
  NAND2_X1 U21714 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18807) );
  NOR2_X1 U21715 ( .A1(n18565), .A2(n18807), .ZN(n18566) );
  NAND2_X1 U21716 ( .A1(n18567), .A2(n18566), .ZN(n18671) );
  OAI21_X1 U21717 ( .B1(n10159), .B2(n18671), .A(n18568), .ZN(n18569) );
  XOR2_X1 U21718 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n18569), .Z(
        n18838) );
  AOI21_X1 U21719 ( .B1(n18606), .B2(n18571), .A(n18722), .ZN(n18598) );
  OAI21_X1 U21720 ( .B1(n18570), .B2(n18608), .A(n18598), .ZN(n18582) );
  AOI22_X1 U21721 ( .A1(n18954), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18582), .ZN(n18574) );
  NOR2_X1 U21722 ( .A1(n18610), .A2(n18571), .ZN(n18584) );
  OAI211_X1 U21723 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n18584), .B(n18572), .ZN(n18573) );
  OAI211_X1 U21724 ( .C1(n18622), .C2(n18575), .A(n18574), .B(n18573), .ZN(
        n18576) );
  AOI21_X1 U21725 ( .B1(n18681), .B2(n18838), .A(n18576), .ZN(n18577) );
  OAI221_X1 U21726 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18579), 
        .C1(n10157), .C2(n18578), .A(n18577), .ZN(P3_U2814) );
  NOR3_X1 U21727 ( .A1(n18904), .A2(n18861), .A3(n18868), .ZN(n18602) );
  NOR2_X1 U21728 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18602), .ZN(
        n18851) );
  NAND2_X1 U21729 ( .A1(n18647), .A2(n18843), .ZN(n18592) );
  NAND2_X1 U21730 ( .A1(n18954), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18853) );
  OAI21_X1 U21731 ( .B1(n18622), .B2(n18580), .A(n18853), .ZN(n18581) );
  AOI221_X1 U21732 ( .B1(n18584), .B2(n18583), .C1(n18582), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n18581), .ZN(n18591) );
  NAND2_X1 U21733 ( .A1(n18594), .A2(n18868), .ZN(n18586) );
  INV_X1 U21734 ( .A(n18908), .ZN(n18655) );
  OR2_X1 U21735 ( .A1(n18671), .A2(n18655), .ZN(n18661) );
  AND2_X1 U21736 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n13336), .ZN(
        n18593) );
  AOI21_X1 U21737 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18615), .A(
        n18593), .ZN(n18585) );
  NAND2_X1 U21738 ( .A1(n18586), .A2(n18585), .ZN(n18587) );
  XNOR2_X1 U21739 ( .A(n18587), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18842) );
  AND2_X1 U21740 ( .A1(n18844), .A2(n18645), .ZN(n18589) );
  OR2_X1 U21741 ( .A1(n18845), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18588) );
  AOI22_X1 U21742 ( .A1(n18681), .A2(n18842), .B1(n18589), .B2(n18588), .ZN(
        n18590) );
  OAI211_X1 U21743 ( .C1(n18851), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2815) );
  AOI21_X1 U21744 ( .B1(n18594), .B2(n18615), .A(n18593), .ZN(n18595) );
  XNOR2_X1 U21745 ( .A(n18595), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n18874) );
  AOI21_X1 U21746 ( .B1(n18596), .B2(n19351), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18597) );
  OAI22_X1 U21747 ( .A1(n18598), .A2(n18597), .B1(n18981), .B2(n19504), .ZN(
        n18599) );
  AOI21_X1 U21748 ( .B1(n18600), .B2(n18714), .A(n18599), .ZN(n18605) );
  AOI21_X1 U21749 ( .B1(n18868), .B2(n18601), .A(n18845), .ZN(n18864) );
  NAND2_X1 U21750 ( .A1(n18858), .A2(n18646), .ZN(n18603) );
  AOI21_X1 U21751 ( .B1(n18868), .B2(n18603), .A(n18602), .ZN(n18869) );
  AOI22_X1 U21752 ( .A1(n18645), .A2(n18864), .B1(n18647), .B2(n18869), .ZN(
        n18604) );
  OAI211_X1 U21753 ( .C1(n18653), .C2(n18874), .A(n18605), .B(n18604), .ZN(
        P3_U2816) );
  NAND2_X1 U21754 ( .A1(n18901), .A2(n18617), .ZN(n18877) );
  NAND2_X1 U21755 ( .A1(n18617), .A2(n18646), .ZN(n18879) );
  AOI22_X1 U21756 ( .A1(n18645), .A2(n18877), .B1(n18647), .B2(n18879), .ZN(
        n18627) );
  AOI21_X1 U21757 ( .B1(n18606), .B2(n18638), .A(n18722), .ZN(n18607) );
  OAI21_X1 U21758 ( .B1(n18609), .B2(n18608), .A(n18607), .ZN(n18624) );
  NOR2_X1 U21759 ( .A1(n18610), .A2(n18638), .ZN(n18626) );
  OAI211_X1 U21760 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18626), .B(n18611), .ZN(n18612) );
  NAND2_X1 U21761 ( .A1(n18954), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18886) );
  OAI211_X1 U21762 ( .C1(n18622), .C2(n18613), .A(n18612), .B(n18886), .ZN(
        n18614) );
  AOI21_X1 U21763 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18624), .A(
        n18614), .ZN(n18619) );
  OAI21_X1 U21764 ( .B1(n9690), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18615), .ZN(n18616) );
  XNOR2_X1 U21765 ( .A(n18616), .B(n13336), .ZN(n18876) );
  INV_X1 U21766 ( .A(n18617), .ZN(n18860) );
  NOR2_X1 U21767 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18860), .ZN(
        n18875) );
  AOI22_X1 U21768 ( .A1(n18681), .A2(n18876), .B1(n18875), .B2(n18654), .ZN(
        n18618) );
  OAI211_X1 U21769 ( .C1(n18627), .C2(n13336), .A(n18619), .B(n18618), .ZN(
        P3_U2817) );
  NAND2_X1 U21770 ( .A1(n9690), .A2(n18634), .ZN(n18620) );
  XNOR2_X1 U21771 ( .A(n18620), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18898) );
  NAND2_X1 U21772 ( .A1(n18954), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18896) );
  OAI21_X1 U21773 ( .B1(n18622), .B2(n18621), .A(n18896), .ZN(n18623) );
  AOI221_X1 U21774 ( .B1(n18626), .B2(n18625), .C1(n18624), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18623), .ZN(n18631) );
  INV_X1 U21775 ( .A(n18627), .ZN(n18629) );
  NOR2_X1 U21776 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18889), .ZN(
        n18628) );
  AOI22_X1 U21777 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18629), .B1(
        n18628), .B2(n18654), .ZN(n18630) );
  OAI211_X1 U21778 ( .C1(n18898), .C2(n18653), .A(n18631), .B(n18630), .ZN(
        P3_U2818) );
  NAND2_X1 U21779 ( .A1(n18661), .A2(n10057), .ZN(n18633) );
  MUX2_X1 U21780 ( .A(n10057), .B(n18633), .S(n18632), .Z(n18635) );
  NAND2_X1 U21781 ( .A1(n18635), .A2(n18634), .ZN(n18914) );
  NOR2_X1 U21782 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18655), .ZN(
        n18899) );
  INV_X1 U21783 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19497) );
  NOR2_X1 U21784 ( .A1(n18981), .A2(n19497), .ZN(n18643) );
  INV_X1 U21785 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18676) );
  NAND2_X1 U21786 ( .A1(n18637), .A2(n18636), .ZN(n18677) );
  NOR2_X1 U21787 ( .A1(n18676), .A2(n18677), .ZN(n18675) );
  AOI22_X1 U21788 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18675), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18674), .ZN(n18641) );
  NOR2_X1 U21789 ( .A1(n19180), .A2(n18638), .ZN(n18640) );
  OAI22_X1 U21790 ( .A1(n18641), .A2(n18640), .B1(n18720), .B2(n18639), .ZN(
        n18642) );
  AOI211_X1 U21791 ( .C1(n18899), .C2(n18654), .A(n18643), .B(n18642), .ZN(
        n18652) );
  INV_X1 U21792 ( .A(n18654), .ZN(n18684) );
  NOR2_X1 U21793 ( .A1(n18908), .A2(n18684), .ZN(n18650) );
  INV_X1 U21794 ( .A(n18901), .ZN(n18644) );
  NAND2_X1 U21795 ( .A1(n18645), .A2(n18644), .ZN(n18649) );
  NAND2_X1 U21796 ( .A1(n18647), .A2(n18904), .ZN(n18648) );
  AND2_X1 U21797 ( .A1(n18649), .A2(n18648), .ZN(n18683) );
  INV_X1 U21798 ( .A(n18683), .ZN(n18656) );
  OAI21_X1 U21799 ( .B1(n18650), .B2(n18656), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18651) );
  OAI211_X1 U21800 ( .C1(n18914), .C2(n18653), .A(n18652), .B(n18651), .ZN(
        P3_U2819) );
  AOI22_X1 U21801 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18656), .B1(
        n18655), .B2(n18654), .ZN(n18669) );
  NOR2_X1 U21802 ( .A1(n18675), .A2(n18658), .ZN(n18657) );
  INV_X1 U21803 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19495) );
  NOR2_X1 U21804 ( .A1(n18981), .A2(n19495), .ZN(n18922) );
  AOI221_X1 U21805 ( .B1(n18675), .B2(n18658), .C1(n18657), .C2(n18674), .A(
        n18922), .ZN(n18668) );
  NOR4_X1 U21806 ( .A1(n18660), .A2(n18659), .A3(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A4(n18919), .ZN(n18665) );
  INV_X1 U21807 ( .A(n18661), .ZN(n18664) );
  OAI21_X1 U21808 ( .B1(n18671), .B2(n18931), .A(n18919), .ZN(n18662) );
  AOI21_X1 U21809 ( .B1(n13335), .B2(n18931), .A(n18662), .ZN(n18663) );
  NOR3_X1 U21810 ( .A1(n18665), .A2(n18664), .A3(n18663), .ZN(n18923) );
  AOI22_X1 U21811 ( .A1(n18681), .A2(n18923), .B1(n18666), .B2(n18714), .ZN(
        n18667) );
  OAI211_X1 U21812 ( .C1(n18670), .C2(n18669), .A(n18668), .B(n18667), .ZN(
        P3_U2820) );
  NAND2_X1 U21813 ( .A1(n18672), .A2(n18671), .ZN(n18673) );
  XNOR2_X1 U21814 ( .A(n18673), .B(n18931), .ZN(n18935) );
  INV_X1 U21815 ( .A(n18674), .ZN(n18687) );
  AOI211_X1 U21816 ( .C1(n18677), .C2(n18676), .A(n18687), .B(n18675), .ZN(
        n18680) );
  NAND2_X1 U21817 ( .A1(n18954), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18937) );
  OAI21_X1 U21818 ( .B1(n18720), .B2(n18678), .A(n18937), .ZN(n18679) );
  AOI211_X1 U21819 ( .C1(n18681), .C2(n18935), .A(n18680), .B(n18679), .ZN(
        n18682) );
  OAI221_X1 U21820 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18684), .C1(
        n18931), .C2(n18683), .A(n18682), .ZN(P3_U2821) );
  NOR2_X1 U21821 ( .A1(n19180), .A2(n16911), .ZN(n18686) );
  AOI22_X1 U21822 ( .A1(n18954), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18686), 
        .B2(n18685), .ZN(n18692) );
  NOR2_X1 U21823 ( .A1(n18687), .A2(n18686), .ZN(n18700) );
  OAI22_X1 U21824 ( .A1(n18720), .A2(n18689), .B1(n18717), .B2(n18688), .ZN(
        n18690) );
  AOI21_X1 U21825 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18700), .A(
        n18690), .ZN(n18691) );
  OAI211_X1 U21826 ( .C1(n18693), .C2(n18727), .A(n18692), .B(n18691), .ZN(
        P3_U2824) );
  OAI21_X1 U21827 ( .B1(n18696), .B2(n18695), .A(n18694), .ZN(n18948) );
  XNOR2_X1 U21828 ( .A(n18697), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18941) );
  OAI22_X1 U21829 ( .A1(n18717), .A2(n18941), .B1(n19488), .B2(n18981), .ZN(
        n18698) );
  AOI21_X1 U21830 ( .B1(n18699), .B2(n18714), .A(n18698), .ZN(n18703) );
  OAI221_X1 U21831 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18701), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18708), .A(n18700), .ZN(n18702) );
  OAI211_X1 U21832 ( .C1(n18727), .C2(n18948), .A(n18703), .B(n18702), .ZN(
        P3_U2825) );
  OR2_X1 U21833 ( .A1(n18705), .A2(n18704), .ZN(n18707) );
  NAND2_X1 U21834 ( .A1(n18707), .A2(n18706), .ZN(n18963) );
  AOI21_X1 U21835 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18708), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18711) );
  XNOR2_X1 U21836 ( .A(n18710), .B(n18709), .ZN(n18962) );
  OAI22_X1 U21837 ( .A1(n18712), .A2(n18711), .B1(n18717), .B2(n18962), .ZN(
        n18713) );
  AOI21_X1 U21838 ( .B1(n18715), .B2(n18714), .A(n18713), .ZN(n18716) );
  NAND2_X1 U21839 ( .A1(n18954), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18966) );
  OAI211_X1 U21840 ( .C1(n18727), .C2(n18963), .A(n18716), .B(n18966), .ZN(
        P3_U2827) );
  OAI22_X1 U21841 ( .A1(n18720), .A2(n18719), .B1(n18718), .B2(n18717), .ZN(
        n18721) );
  AOI221_X1 U21842 ( .B1(n19351), .B2(n18723), .C1(n18722), .C2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n18721), .ZN(n18725) );
  OAI211_X1 U21843 ( .C1(n18727), .C2(n18726), .A(n18725), .B(n18724), .ZN(
        P3_U2828) );
  AOI22_X1 U21844 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18976), .B1(
        n18954), .B2(P3_REIP_REG_27__SCAN_IN), .ZN(n18732) );
  OAI211_X1 U21845 ( .C1(n18927), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18728), .ZN(n18729) );
  OAI211_X1 U21846 ( .C1(n18730), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18958), .B(n18729), .ZN(n18731) );
  OAI211_X1 U21847 ( .C1(n18733), .C2(n18913), .A(n18732), .B(n18731), .ZN(
        P3_U2835) );
  AOI21_X1 U21848 ( .B1(n18976), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18734), .ZN(n18748) );
  AOI211_X1 U21849 ( .C1(n19400), .C2(n18737), .A(n18736), .B(n18735), .ZN(
        n18744) );
  NOR2_X1 U21850 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18738), .ZN(
        n18740) );
  AOI22_X1 U21851 ( .A1(n18741), .A2(n18740), .B1(n18878), .B2(n18739), .ZN(
        n18742) );
  OAI21_X1 U21852 ( .B1(n18744), .B2(n18743), .A(n18742), .ZN(n18746) );
  AOI22_X1 U21853 ( .A1(n18958), .A2(n18746), .B1(n18936), .B2(n18745), .ZN(
        n18747) );
  OAI211_X1 U21854 ( .C1(n18973), .C2(n18749), .A(n18748), .B(n18747), .ZN(
        P3_U2837) );
  OAI21_X1 U21855 ( .B1(n18976), .B2(n18751), .A(n18750), .ZN(n18752) );
  AOI22_X1 U21856 ( .A1(n18954), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n18753), 
        .B2(n18752), .ZN(n18754) );
  OAI21_X1 U21857 ( .B1(n18913), .B2(n18755), .A(n18754), .ZN(P3_U2839) );
  NOR2_X1 U21858 ( .A1(n18981), .A2(n21548), .ZN(n18776) );
  AOI22_X1 U21859 ( .A1(n19399), .A2(n18843), .B1(n18878), .B2(n18844), .ZN(
        n18782) );
  INV_X1 U21860 ( .A(n18817), .ZN(n18769) );
  NAND2_X1 U21861 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18756), .ZN(
        n18833) );
  OAI21_X1 U21862 ( .B1(n18757), .B2(n18833), .A(n18905), .ZN(n18761) );
  INV_X1 U21863 ( .A(n18758), .ZN(n18793) );
  OAI21_X1 U21864 ( .B1(n18759), .B2(n18793), .A(n18978), .ZN(n18760) );
  OAI211_X1 U21865 ( .C1(n18763), .C2(n18762), .A(n18761), .B(n18760), .ZN(
        n18791) );
  NOR2_X1 U21866 ( .A1(n19399), .A2(n18878), .ZN(n18907) );
  OAI22_X1 U21867 ( .A1(n18927), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18772), .B2(n18907), .ZN(n18764) );
  NOR2_X1 U21868 ( .A1(n18791), .A2(n18764), .ZN(n18783) );
  AOI21_X1 U21869 ( .B1(n19400), .B2(n18766), .A(n18765), .ZN(n18767) );
  OAI211_X1 U21870 ( .C1(n18926), .C2(n18784), .A(n18783), .B(n18767), .ZN(
        n18768) );
  AOI21_X1 U21871 ( .B1(n18770), .B2(n18769), .A(n18768), .ZN(n18774) );
  AOI21_X1 U21872 ( .B1(n18772), .B2(n18771), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18773) );
  AOI211_X1 U21873 ( .C1(n18782), .C2(n18774), .A(n18773), .B(n18888), .ZN(
        n18775) );
  AOI211_X1 U21874 ( .C1(n18976), .C2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n18776), .B(n18775), .ZN(n18777) );
  OAI21_X1 U21875 ( .B1(n18913), .B2(n18778), .A(n18777), .ZN(P3_U2840) );
  NAND2_X1 U21876 ( .A1(n18780), .A2(n18779), .ZN(n18799) );
  AOI22_X1 U21877 ( .A1(n18954), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18936), 
        .B2(n18781), .ZN(n18787) );
  NAND2_X1 U21878 ( .A1(n18958), .A2(n18782), .ZN(n18837) );
  OAI21_X1 U21879 ( .B1(n18784), .B2(n18857), .A(n18783), .ZN(n18785) );
  OAI211_X1 U21880 ( .C1(n18837), .C2(n18785), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18981), .ZN(n18786) );
  OAI211_X1 U21881 ( .C1(n18799), .C2(n18788), .A(n18787), .B(n18786), .ZN(
        P3_U2841) );
  AOI21_X1 U21882 ( .B1(n18790), .B2(n18936), .A(n18789), .ZN(n18797) );
  INV_X1 U21883 ( .A(n18907), .ZN(n18792) );
  AOI211_X1 U21884 ( .C1(n18793), .C2(n18792), .A(n18837), .B(n18791), .ZN(
        n18794) );
  NOR2_X1 U21885 ( .A1(n18954), .A2(n18794), .ZN(n18802) );
  NOR3_X1 U21886 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18857), .A3(
        n21628), .ZN(n18795) );
  OAI21_X1 U21887 ( .B1(n18802), .B2(n18795), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18796) );
  OAI211_X1 U21888 ( .C1(n18798), .C2(n18799), .A(n18797), .B(n18796), .ZN(
        P3_U2842) );
  INV_X1 U21889 ( .A(n18799), .ZN(n18801) );
  AOI22_X1 U21890 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18802), .B1(
        n18801), .B2(n18800), .ZN(n18804) );
  OAI211_X1 U21891 ( .C1(n18805), .C2(n18913), .A(n18804), .B(n18803), .ZN(
        P3_U2843) );
  NAND2_X1 U21892 ( .A1(n18810), .A2(n18915), .ZN(n18841) );
  AOI21_X1 U21893 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18811), .A(
        n18817), .ZN(n18815) );
  INV_X1 U21894 ( .A(n18837), .ZN(n18812) );
  OAI21_X1 U21895 ( .B1(n18813), .B2(n18907), .A(n18812), .ZN(n18814) );
  AOI211_X1 U21896 ( .C1(n19400), .C2(n18816), .A(n18815), .B(n18814), .ZN(
        n18826) );
  OAI21_X1 U21897 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18817), .A(
        n18826), .ZN(n18821) );
  NOR2_X1 U21898 ( .A1(n18954), .A2(n18818), .ZN(n18820) );
  AOI22_X1 U21899 ( .A1(n18821), .A2(n18820), .B1(n18936), .B2(n18819), .ZN(
        n18823) );
  NAND2_X1 U21900 ( .A1(n18954), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n18822) );
  OAI211_X1 U21901 ( .C1(n18824), .C2(n18841), .A(n18823), .B(n18822), .ZN(
        P3_U2844) );
  NAND2_X1 U21902 ( .A1(n18981), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n18825) );
  OR2_X1 U21903 ( .A1(n18826), .A2(n18825), .ZN(n18828) );
  OR3_X1 U21904 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n10157), .A3(
        n18841), .ZN(n18827) );
  OAI211_X1 U21905 ( .C1(n18829), .C2(n18913), .A(n18828), .B(n18827), .ZN(
        n18830) );
  INV_X1 U21906 ( .A(n18830), .ZN(n18832) );
  NAND2_X1 U21907 ( .A1(n18832), .A2(n18831), .ZN(P3_U2845) );
  NOR2_X1 U21908 ( .A1(n18927), .A2(n18856), .ZN(n18917) );
  AOI21_X1 U21909 ( .B1(n19400), .B2(n18880), .A(n18917), .ZN(n18867) );
  OAI21_X1 U21910 ( .B1(n18834), .B2(n18905), .A(n18833), .ZN(n18835) );
  OAI211_X1 U21911 ( .C1(n18882), .C2(n18847), .A(n18867), .B(n18835), .ZN(
        n18846) );
  OAI221_X1 U21912 ( .B1(n18837), .B2(n18836), .C1(n18837), .C2(n18846), .A(
        n18981), .ZN(n18840) );
  AOI22_X1 U21913 ( .A1(n18954), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18936), 
        .B2(n18838), .ZN(n18839) );
  OAI221_X1 U21914 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18841), 
        .C1(n10157), .C2(n18840), .A(n18839), .ZN(P3_U2846) );
  INV_X1 U21915 ( .A(n18842), .ZN(n18855) );
  NAND2_X1 U21916 ( .A1(n19399), .A2(n18843), .ZN(n18850) );
  OAI211_X1 U21917 ( .C1(n18845), .C2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n18878), .B(n18844), .ZN(n18849) );
  OAI221_X1 U21918 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18847), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18863), .A(n18846), .ZN(
        n18848) );
  OAI211_X1 U21919 ( .C1(n18851), .C2(n18850), .A(n18849), .B(n18848), .ZN(
        n18852) );
  AOI22_X1 U21920 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18976), .B1(
        n18958), .B2(n18852), .ZN(n18854) );
  OAI211_X1 U21921 ( .C1(n18913), .C2(n18855), .A(n18854), .B(n18853), .ZN(
        P3_U2847) );
  AOI22_X1 U21922 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18976), .B1(
        n18954), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18873) );
  NAND2_X1 U21923 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18856), .ZN(
        n18929) );
  NOR2_X1 U21924 ( .A1(n18860), .A2(n18929), .ZN(n18893) );
  NOR2_X1 U21925 ( .A1(n18926), .A2(n18893), .ZN(n18884) );
  OAI22_X1 U21926 ( .A1(n18927), .A2(n18858), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n18857), .ZN(n18859) );
  AOI211_X1 U21927 ( .C1(n19400), .C2(n18860), .A(n18884), .B(n18859), .ZN(
        n18866) );
  NOR2_X1 U21928 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18861), .ZN(
        n18862) );
  AOI22_X1 U21929 ( .A1(n18878), .A2(n18864), .B1(n18863), .B2(n18862), .ZN(
        n18865) );
  OAI221_X1 U21930 ( .B1(n18868), .B2(n18867), .C1(n18868), .C2(n18866), .A(
        n18865), .ZN(n18871) );
  AOI22_X1 U21931 ( .A1(n18958), .A2(n18871), .B1(n18870), .B2(n18869), .ZN(
        n18872) );
  OAI211_X1 U21932 ( .C1(n18913), .C2(n18874), .A(n18873), .B(n18872), .ZN(
        P3_U2848) );
  AOI22_X1 U21933 ( .A1(n18936), .A2(n18876), .B1(n18915), .B2(n18875), .ZN(
        n18887) );
  AOI22_X1 U21934 ( .A1(n19399), .A2(n18879), .B1(n18878), .B2(n18877), .ZN(
        n18881) );
  NAND2_X1 U21935 ( .A1(n19400), .A2(n18880), .ZN(n18900) );
  INV_X1 U21936 ( .A(n18882), .ZN(n18918) );
  OAI21_X1 U21937 ( .B1(n18917), .B2(n18889), .A(n18918), .ZN(n18909) );
  AND3_X1 U21938 ( .A1(n18881), .A2(n18900), .A3(n18909), .ZN(n18892) );
  OAI211_X1 U21939 ( .C1(n18882), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18958), .B(n18892), .ZN(n18883) );
  OAI211_X1 U21940 ( .C1(n18884), .C2(n18883), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18981), .ZN(n18885) );
  NAND3_X1 U21941 ( .A1(n18887), .A2(n18886), .A3(n18885), .ZN(P3_U2849) );
  AOI221_X1 U21942 ( .B1(n18891), .B2(n18890), .C1(n18889), .C2(n18890), .A(
        n18888), .ZN(n18895) );
  OAI211_X1 U21943 ( .C1(n18893), .C2(n18926), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18892), .ZN(n18894) );
  AOI22_X1 U21944 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18976), .B1(
        n18895), .B2(n18894), .ZN(n18897) );
  OAI211_X1 U21945 ( .C1(n18898), .C2(n18913), .A(n18897), .B(n18896), .ZN(
        P3_U2850) );
  AOI22_X1 U21946 ( .A1(n18954), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18915), 
        .B2(n18899), .ZN(n18912) );
  OAI211_X1 U21947 ( .C1(n18902), .C2(n18901), .A(n18958), .B(n18900), .ZN(
        n18903) );
  AOI21_X1 U21948 ( .B1(n19399), .B2(n18904), .A(n18903), .ZN(n18933) );
  OAI21_X1 U21949 ( .B1(n18931), .B2(n18929), .A(n18905), .ZN(n18906) );
  OAI211_X1 U21950 ( .C1(n18908), .C2(n18907), .A(n18933), .B(n18906), .ZN(
        n18916) );
  OAI21_X1 U21951 ( .B1(n18926), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18909), .ZN(n18910) );
  OAI211_X1 U21952 ( .C1(n18916), .C2(n18910), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18981), .ZN(n18911) );
  OAI211_X1 U21953 ( .C1(n18914), .C2(n18913), .A(n18912), .B(n18911), .ZN(
        P3_U2851) );
  INV_X1 U21954 ( .A(n18915), .ZN(n18939) );
  NAND2_X1 U21955 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18919), .ZN(
        n18925) );
  AOI211_X1 U21956 ( .C1(n18918), .C2(n18931), .A(n18917), .B(n18916), .ZN(
        n18920) );
  NOR3_X1 U21957 ( .A1(n18954), .A2(n18920), .A3(n18919), .ZN(n18921) );
  AOI211_X1 U21958 ( .C1(n18923), .C2(n18936), .A(n18922), .B(n18921), .ZN(
        n18924) );
  OAI21_X1 U21959 ( .B1(n18939), .B2(n18925), .A(n18924), .ZN(P3_U2852) );
  OAI21_X1 U21960 ( .B1(n18927), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n18926), .ZN(n18930) );
  AOI22_X1 U21961 ( .A1(n18930), .A2(n18929), .B1(n18978), .B2(n18928), .ZN(
        n18932) );
  AOI211_X1 U21962 ( .C1(n18933), .C2(n18932), .A(n18954), .B(n18931), .ZN(
        n18934) );
  AOI21_X1 U21963 ( .B1(n18936), .B2(n18935), .A(n18934), .ZN(n18938) );
  OAI211_X1 U21964 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18939), .A(
        n18938), .B(n18937), .ZN(P3_U2853) );
  NAND3_X1 U21965 ( .A1(n18940), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18958), .ZN(n18951) );
  NOR2_X1 U21966 ( .A1(n18951), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18945) );
  OAI22_X1 U21967 ( .A1(n18943), .A2(n18942), .B1(n18941), .B2(n18971), .ZN(
        n18944) );
  AOI21_X1 U21968 ( .B1(n18945), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18944), .ZN(n18947) );
  NAND2_X1 U21969 ( .A1(n18954), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18946) );
  OAI211_X1 U21970 ( .C1(n18948), .C2(n18973), .A(n18947), .B(n18946), .ZN(
        P3_U2857) );
  AOI21_X1 U21971 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18961), .A(
        n18949), .ZN(n18953) );
  OAI22_X1 U21972 ( .A1(n18951), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n18950), .B2(n18971), .ZN(n18952) );
  AOI221_X1 U21973 ( .B1(n18976), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n18953), .C2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18952), .ZN(
        n18956) );
  NAND2_X1 U21974 ( .A1(n18954), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18955) );
  OAI211_X1 U21975 ( .C1(n18973), .C2(n18957), .A(n18956), .B(n18955), .ZN(
        P3_U2858) );
  NAND2_X1 U21976 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18958), .ZN(
        n18959) );
  AOI22_X1 U21977 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18959), .ZN(n18965) );
  OAI22_X1 U21978 ( .A1(n18973), .A2(n18963), .B1(n18971), .B2(n18962), .ZN(
        n18964) );
  NOR2_X1 U21979 ( .A1(n18965), .A2(n18964), .ZN(n18967) );
  OAI211_X1 U21980 ( .C1(n18969), .C2(n18968), .A(n18967), .B(n18966), .ZN(
        P3_U2859) );
  OAI22_X1 U21981 ( .A1(n18973), .A2(n18972), .B1(n18971), .B2(n18970), .ZN(
        n18974) );
  AOI221_X1 U21982 ( .B1(n18976), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18975), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n18974), .ZN(
        n18980) );
  OAI211_X1 U21983 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18978), .A(
        n18977), .B(n9830), .ZN(n18979) );
  OAI211_X1 U21984 ( .C1(n19554), .C2(n18981), .A(n18980), .B(n18979), .ZN(
        P3_U2861) );
  OAI211_X1 U21985 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18982), .A(
        P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .ZN(n19443)
         );
  INV_X1 U21986 ( .A(n19031), .ZN(n18985) );
  OAI21_X1 U21987 ( .B1(n18986), .B2(n18983), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18984) );
  OAI221_X1 U21988 ( .B1(n18986), .B2(n19443), .C1(n18986), .C2(n18985), .A(
        n18984), .ZN(P3_U2863) );
  INV_X1 U21989 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19432) );
  NOR2_X1 U21990 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19432), .ZN(
        n19270) );
  NOR2_X1 U21991 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19430), .ZN(
        n19131) );
  NOR2_X1 U21992 ( .A1(n19270), .A2(n19131), .ZN(n18988) );
  OAI22_X1 U21993 ( .A1(n18989), .A2(n19432), .B1(n18988), .B2(n18987), .ZN(
        P3_U2866) );
  NOR2_X1 U21994 ( .A1(n19433), .A2(n18990), .ZN(P3_U2867) );
  NAND2_X1 U21995 ( .A1(n13491), .A2(n13509), .ZN(n19425) );
  NAND2_X1 U21996 ( .A1(n19430), .A2(n19432), .ZN(n19067) );
  NOR2_X2 U21997 ( .A1(n19425), .A2(n19067), .ZN(n21666) );
  INV_X1 U21998 ( .A(n21666), .ZN(n19030) );
  NOR3_X2 U21999 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18991), .A3(n19552), 
        .ZN(n19025) );
  NAND2_X1 U22000 ( .A1(n19025), .A2(n18992), .ZN(n19355) );
  NOR2_X2 U22001 ( .A1(n19179), .A2(n18993), .ZN(n19347) );
  NAND2_X1 U22002 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19419) );
  NAND2_X1 U22003 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18994) );
  NOR2_X2 U22004 ( .A1(n19419), .A2(n18994), .ZN(n19345) );
  NOR2_X1 U22005 ( .A1(n21666), .A2(n19345), .ZN(n19051) );
  NOR2_X1 U22006 ( .A1(n19318), .A2(n19051), .ZN(n19026) );
  INV_X1 U22007 ( .A(n18994), .ZN(n18998) );
  NAND2_X1 U22008 ( .A1(n18998), .A2(n13491), .ZN(n19296) );
  NOR2_X2 U22009 ( .A1(n13509), .A2(n19296), .ZN(n19395) );
  NOR2_X2 U22010 ( .A1(n16026), .A2(n19180), .ZN(n19346) );
  AOI22_X1 U22011 ( .A1(n19347), .A2(n19026), .B1(n19395), .B2(n19346), .ZN(
        n19000) );
  AOI21_X1 U22012 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n19051), .ZN(n18996) );
  NOR2_X1 U22013 ( .A1(n13491), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19269) );
  NOR2_X1 U22014 ( .A1(n13509), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19268) );
  OAI21_X1 U22015 ( .B1(n19269), .B2(n19268), .A(n18998), .ZN(n19319) );
  INV_X1 U22016 ( .A(n19319), .ZN(n18995) );
  AOI22_X1 U22017 ( .A1(n19323), .A2(n18996), .B1(n19351), .B2(n18995), .ZN(
        n19027) );
  NOR2_X2 U22018 ( .A1(n19180), .A2(n18997), .ZN(n19352) );
  NAND2_X1 U22019 ( .A1(n18998), .A2(n19269), .ZN(n19344) );
  AOI22_X1 U22020 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19027), .B1(
        n19352), .B2(n19324), .ZN(n18999) );
  OAI211_X1 U22021 ( .C1(n19030), .C2(n19355), .A(n19000), .B(n18999), .ZN(
        P3_U2868) );
  NAND2_X1 U22022 ( .A1(n19025), .A2(n19001), .ZN(n19361) );
  AND2_X1 U22023 ( .A1(n19323), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19356) );
  NOR2_X2 U22024 ( .A1(n16018), .A2(n19180), .ZN(n19358) );
  AOI22_X1 U22025 ( .A1(n19026), .A2(n19356), .B1(n19395), .B2(n19358), .ZN(
        n19003) );
  NOR2_X2 U22026 ( .A1(n19180), .A2(n16076), .ZN(n19357) );
  AOI22_X1 U22027 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19027), .B1(
        n19324), .B2(n19357), .ZN(n19002) );
  OAI211_X1 U22028 ( .C1(n19030), .C2(n19361), .A(n19003), .B(n19002), .ZN(
        P3_U2869) );
  NAND2_X1 U22029 ( .A1(n19025), .A2(n19004), .ZN(n19367) );
  NOR2_X2 U22030 ( .A1(n19180), .A2(n16070), .ZN(n19364) );
  NOR2_X2 U22031 ( .A1(n19179), .A2(n19005), .ZN(n19362) );
  AOI22_X1 U22032 ( .A1(n19324), .A2(n19364), .B1(n19026), .B2(n19362), .ZN(
        n19007) );
  NOR2_X2 U22033 ( .A1(n19990), .A2(n19180), .ZN(n19363) );
  AOI22_X1 U22034 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19027), .B1(
        n19395), .B2(n19363), .ZN(n19006) );
  OAI211_X1 U22035 ( .C1(n19030), .C2(n19367), .A(n19007), .B(n19006), .ZN(
        P3_U2870) );
  NAND2_X1 U22036 ( .A1(n19025), .A2(n19008), .ZN(n19373) );
  NOR2_X2 U22037 ( .A1(n19179), .A2(n19009), .ZN(n19368) );
  NOR2_X2 U22038 ( .A1(n14536), .A2(n19180), .ZN(n19370) );
  AOI22_X1 U22039 ( .A1(n19026), .A2(n19368), .B1(n19395), .B2(n19370), .ZN(
        n19011) );
  NOR2_X2 U22040 ( .A1(n19180), .A2(n16061), .ZN(n19369) );
  AOI22_X1 U22041 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19027), .B1(
        n19324), .B2(n19369), .ZN(n19010) );
  OAI211_X1 U22042 ( .C1(n19030), .C2(n19373), .A(n19011), .B(n19010), .ZN(
        P3_U2871) );
  NAND2_X1 U22043 ( .A1(n19025), .A2(n19012), .ZN(n19379) );
  NOR2_X2 U22044 ( .A1(n19179), .A2(n19013), .ZN(n19374) );
  NOR2_X2 U22045 ( .A1(n16005), .A2(n19180), .ZN(n19376) );
  AOI22_X1 U22046 ( .A1(n19026), .A2(n19374), .B1(n19395), .B2(n19376), .ZN(
        n19015) );
  NOR2_X2 U22047 ( .A1(n19180), .A2(n20006), .ZN(n19375) );
  AOI22_X1 U22048 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19027), .B1(
        n19324), .B2(n19375), .ZN(n19014) );
  OAI211_X1 U22049 ( .C1(n19030), .C2(n19379), .A(n19015), .B(n19014), .ZN(
        P3_U2872) );
  NAND2_X1 U22050 ( .A1(n19025), .A2(n19016), .ZN(n19385) );
  AND2_X1 U22051 ( .A1(n19323), .A2(BUF2_REG_5__SCAN_IN), .ZN(n19380) );
  NOR2_X2 U22052 ( .A1(n12390), .A2(n19180), .ZN(n19382) );
  AOI22_X1 U22053 ( .A1(n19026), .A2(n19380), .B1(n19395), .B2(n19382), .ZN(
        n19018) );
  NOR2_X2 U22054 ( .A1(n19180), .A2(n16046), .ZN(n19381) );
  AOI22_X1 U22055 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19027), .B1(
        n19324), .B2(n19381), .ZN(n19017) );
  OAI211_X1 U22056 ( .C1(n19030), .C2(n19385), .A(n19018), .B(n19017), .ZN(
        P3_U2873) );
  NAND2_X1 U22057 ( .A1(n19025), .A2(n19019), .ZN(n19391) );
  NOR2_X2 U22058 ( .A1(n19179), .A2(n19020), .ZN(n19386) );
  NOR2_X2 U22059 ( .A1(n14609), .A2(n19180), .ZN(n19388) );
  AOI22_X1 U22060 ( .A1(n19026), .A2(n19386), .B1(n19395), .B2(n19388), .ZN(
        n19023) );
  NOR2_X2 U22061 ( .A1(n19180), .A2(n19021), .ZN(n19387) );
  AOI22_X1 U22062 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19027), .B1(
        n19324), .B2(n19387), .ZN(n19022) );
  OAI211_X1 U22063 ( .C1(n19030), .C2(n19391), .A(n19023), .B(n19022), .ZN(
        P3_U2874) );
  NAND2_X1 U22064 ( .A1(n19025), .A2(n19024), .ZN(n21668) );
  NAND2_X1 U22065 ( .A1(n19351), .A2(BUF2_REG_31__SCAN_IN), .ZN(n21670) );
  INV_X1 U22066 ( .A(n21670), .ZN(n19394) );
  NOR2_X2 U22067 ( .A1(n13836), .A2(n19179), .ZN(n21663) );
  AOI22_X1 U22068 ( .A1(n19394), .A2(n19395), .B1(n21663), .B2(n19026), .ZN(
        n19029) );
  NOR2_X2 U22069 ( .A1(n16031), .A2(n19180), .ZN(n21665) );
  AOI22_X1 U22070 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19027), .B1(
        n21665), .B2(n19324), .ZN(n19028) );
  OAI211_X1 U22071 ( .C1(n19030), .C2(n21668), .A(n19029), .B(n19028), .ZN(
        P3_U2875) );
  INV_X1 U22072 ( .A(n19067), .ZN(n19068) );
  NAND2_X1 U22073 ( .A1(n19068), .A2(n19268), .ZN(n19050) );
  NAND2_X1 U22074 ( .A1(n13491), .A2(n19454), .ZN(n19203) );
  NOR2_X1 U22075 ( .A1(n19067), .A2(n19203), .ZN(n19046) );
  AOI22_X1 U22076 ( .A1(n19345), .A2(n19352), .B1(n19347), .B2(n19046), .ZN(
        n19033) );
  NOR2_X1 U22077 ( .A1(n19432), .A2(n19158), .ZN(n19349) );
  NOR2_X1 U22078 ( .A1(n19179), .A2(n19031), .ZN(n19348) );
  AND2_X1 U22079 ( .A1(n13491), .A2(n19348), .ZN(n19110) );
  AOI22_X1 U22080 ( .A1(n19351), .A2(n19349), .B1(n19068), .B2(n19110), .ZN(
        n19047) );
  AOI22_X1 U22081 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19047), .B1(
        n19324), .B2(n19346), .ZN(n19032) );
  OAI211_X1 U22082 ( .C1(n19050), .C2(n19355), .A(n19033), .B(n19032), .ZN(
        P3_U2876) );
  AOI22_X1 U22083 ( .A1(n19324), .A2(n19358), .B1(n19356), .B2(n19046), .ZN(
        n19035) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19047), .B1(
        n19345), .B2(n19357), .ZN(n19034) );
  OAI211_X1 U22085 ( .C1(n19050), .C2(n19361), .A(n19035), .B(n19034), .ZN(
        P3_U2877) );
  AOI22_X1 U22086 ( .A1(n19345), .A2(n19364), .B1(n19362), .B2(n19046), .ZN(
        n19037) );
  AOI22_X1 U22087 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19047), .B1(
        n19324), .B2(n19363), .ZN(n19036) );
  OAI211_X1 U22088 ( .C1(n19050), .C2(n19367), .A(n19037), .B(n19036), .ZN(
        P3_U2878) );
  AOI22_X1 U22089 ( .A1(n19345), .A2(n19369), .B1(n19368), .B2(n19046), .ZN(
        n19039) );
  AOI22_X1 U22090 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19047), .B1(
        n19324), .B2(n19370), .ZN(n19038) );
  OAI211_X1 U22091 ( .C1(n19050), .C2(n19373), .A(n19039), .B(n19038), .ZN(
        P3_U2879) );
  AOI22_X1 U22092 ( .A1(n19324), .A2(n19376), .B1(n19374), .B2(n19046), .ZN(
        n19041) );
  AOI22_X1 U22093 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19047), .B1(
        n19345), .B2(n19375), .ZN(n19040) );
  OAI211_X1 U22094 ( .C1(n19050), .C2(n19379), .A(n19041), .B(n19040), .ZN(
        P3_U2880) );
  AOI22_X1 U22095 ( .A1(n19345), .A2(n19381), .B1(n19380), .B2(n19046), .ZN(
        n19043) );
  AOI22_X1 U22096 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19047), .B1(
        n19324), .B2(n19382), .ZN(n19042) );
  OAI211_X1 U22097 ( .C1(n19050), .C2(n19385), .A(n19043), .B(n19042), .ZN(
        P3_U2881) );
  AOI22_X1 U22098 ( .A1(n19345), .A2(n19387), .B1(n19386), .B2(n19046), .ZN(
        n19045) );
  AOI22_X1 U22099 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19047), .B1(
        n19324), .B2(n19388), .ZN(n19044) );
  OAI211_X1 U22100 ( .C1(n19050), .C2(n19391), .A(n19045), .B(n19044), .ZN(
        P3_U2882) );
  AOI22_X1 U22101 ( .A1(n19394), .A2(n19324), .B1(n21663), .B2(n19046), .ZN(
        n19049) );
  AOI22_X1 U22102 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19047), .B1(
        n19345), .B2(n21665), .ZN(n19048) );
  OAI211_X1 U22103 ( .C1(n19050), .C2(n21668), .A(n19049), .B(n19048), .ZN(
        P3_U2883) );
  NAND2_X1 U22104 ( .A1(n19068), .A2(n19269), .ZN(n21669) );
  NOR2_X1 U22105 ( .A1(n19127), .A2(n19104), .ZN(n19087) );
  NOR2_X1 U22106 ( .A1(n19318), .A2(n19087), .ZN(n21664) );
  AOI22_X1 U22107 ( .A1(n19345), .A2(n19346), .B1(n21664), .B2(n19347), .ZN(
        n19054) );
  OAI21_X1 U22108 ( .B1(n19051), .B2(n19320), .A(n19087), .ZN(n19052) );
  OAI211_X1 U22109 ( .C1(n19127), .C2(n19552), .A(n19323), .B(n19052), .ZN(
        n21674) );
  AOI22_X1 U22110 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n21674), .B1(
        n21666), .B2(n19352), .ZN(n19053) );
  OAI211_X1 U22111 ( .C1(n21669), .C2(n19355), .A(n19054), .B(n19053), .ZN(
        P3_U2884) );
  AOI22_X1 U22112 ( .A1(n19345), .A2(n19358), .B1(n21664), .B2(n19356), .ZN(
        n19056) );
  AOI22_X1 U22113 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n21674), .B1(
        n21666), .B2(n19357), .ZN(n19055) );
  OAI211_X1 U22114 ( .C1(n21669), .C2(n19361), .A(n19056), .B(n19055), .ZN(
        P3_U2885) );
  AOI22_X1 U22115 ( .A1(n21666), .A2(n19364), .B1(n21664), .B2(n19362), .ZN(
        n19058) );
  AOI22_X1 U22116 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n21674), .B1(
        n19345), .B2(n19363), .ZN(n19057) );
  OAI211_X1 U22117 ( .C1(n21669), .C2(n19367), .A(n19058), .B(n19057), .ZN(
        P3_U2886) );
  AOI22_X1 U22118 ( .A1(n21666), .A2(n19369), .B1(n21664), .B2(n19368), .ZN(
        n19060) );
  AOI22_X1 U22119 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n21674), .B1(
        n19345), .B2(n19370), .ZN(n19059) );
  OAI211_X1 U22120 ( .C1(n21669), .C2(n19373), .A(n19060), .B(n19059), .ZN(
        P3_U2887) );
  AOI22_X1 U22121 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n21674), .B1(
        n21664), .B2(n19374), .ZN(n19062) );
  AOI22_X1 U22122 ( .A1(n21666), .A2(n19375), .B1(n19345), .B2(n19376), .ZN(
        n19061) );
  OAI211_X1 U22123 ( .C1(n21669), .C2(n19379), .A(n19062), .B(n19061), .ZN(
        P3_U2888) );
  AOI22_X1 U22124 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n21674), .B1(
        n21664), .B2(n19380), .ZN(n19064) );
  AOI22_X1 U22125 ( .A1(n21666), .A2(n19381), .B1(n19345), .B2(n19382), .ZN(
        n19063) );
  OAI211_X1 U22126 ( .C1(n21669), .C2(n19385), .A(n19064), .B(n19063), .ZN(
        P3_U2889) );
  AOI22_X1 U22127 ( .A1(n19345), .A2(n19388), .B1(n21664), .B2(n19386), .ZN(
        n19066) );
  AOI22_X1 U22128 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n21674), .B1(
        n21666), .B2(n19387), .ZN(n19065) );
  OAI211_X1 U22129 ( .C1(n21669), .C2(n19391), .A(n19066), .B(n19065), .ZN(
        P3_U2890) );
  NOR2_X1 U22130 ( .A1(n13491), .A2(n19067), .ZN(n19111) );
  NAND2_X1 U22131 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19111), .ZN(
        n19109) );
  AND2_X1 U22132 ( .A1(n19454), .A2(n19111), .ZN(n19083) );
  AOI22_X1 U22133 ( .A1(n21666), .A2(n19346), .B1(n19347), .B2(n19083), .ZN(
        n19070) );
  NAND2_X1 U22134 ( .A1(n13491), .A2(n19320), .ZN(n19156) );
  NAND3_X1 U22135 ( .A1(n19068), .A2(n19348), .A3(n19156), .ZN(n19084) );
  AOI22_X1 U22136 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19084), .B1(
        n19104), .B2(n19352), .ZN(n19069) );
  OAI211_X1 U22137 ( .C1(n19355), .C2(n19109), .A(n19070), .B(n19069), .ZN(
        P3_U2892) );
  AOI22_X1 U22138 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19084), .B1(
        n19356), .B2(n19083), .ZN(n19072) );
  AOI22_X1 U22139 ( .A1(n21666), .A2(n19358), .B1(n19104), .B2(n19357), .ZN(
        n19071) );
  OAI211_X1 U22140 ( .C1(n19361), .C2(n19109), .A(n19072), .B(n19071), .ZN(
        P3_U2893) );
  AOI22_X1 U22141 ( .A1(n21666), .A2(n19363), .B1(n19362), .B2(n19083), .ZN(
        n19074) );
  AOI22_X1 U22142 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19084), .B1(
        n19104), .B2(n19364), .ZN(n19073) );
  OAI211_X1 U22143 ( .C1(n19367), .C2(n19109), .A(n19074), .B(n19073), .ZN(
        P3_U2894) );
  AOI22_X1 U22144 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19084), .B1(
        n19368), .B2(n19083), .ZN(n19076) );
  AOI22_X1 U22145 ( .A1(n21666), .A2(n19370), .B1(n19104), .B2(n19369), .ZN(
        n19075) );
  OAI211_X1 U22146 ( .C1(n19373), .C2(n19109), .A(n19076), .B(n19075), .ZN(
        P3_U2895) );
  AOI22_X1 U22147 ( .A1(n19104), .A2(n19375), .B1(n19374), .B2(n19083), .ZN(
        n19078) );
  AOI22_X1 U22148 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19084), .B1(
        n21666), .B2(n19376), .ZN(n19077) );
  OAI211_X1 U22149 ( .C1(n19379), .C2(n19109), .A(n19078), .B(n19077), .ZN(
        P3_U2896) );
  AOI22_X1 U22150 ( .A1(n19104), .A2(n19381), .B1(n19380), .B2(n19083), .ZN(
        n19080) );
  AOI22_X1 U22151 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19084), .B1(
        n21666), .B2(n19382), .ZN(n19079) );
  OAI211_X1 U22152 ( .C1(n19385), .C2(n19109), .A(n19080), .B(n19079), .ZN(
        P3_U2897) );
  AOI22_X1 U22153 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19084), .B1(
        n19386), .B2(n19083), .ZN(n19082) );
  AOI22_X1 U22154 ( .A1(n21666), .A2(n19388), .B1(n19104), .B2(n19387), .ZN(
        n19081) );
  OAI211_X1 U22155 ( .C1(n19391), .C2(n19109), .A(n19082), .B(n19081), .ZN(
        P3_U2898) );
  AOI22_X1 U22156 ( .A1(n21666), .A2(n19394), .B1(n21663), .B2(n19083), .ZN(
        n19086) );
  AOI22_X1 U22157 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19084), .B1(
        n19104), .B2(n21665), .ZN(n19085) );
  OAI211_X1 U22158 ( .C1(n21668), .C2(n19109), .A(n19086), .B(n19085), .ZN(
        P3_U2899) );
  INV_X1 U22159 ( .A(n19131), .ZN(n19155) );
  NOR2_X2 U22160 ( .A1(n19425), .A2(n19155), .ZN(n19175) );
  AOI21_X1 U22161 ( .B1(n19109), .B2(n19108), .A(n19318), .ZN(n19103) );
  AOI22_X1 U22162 ( .A1(n19127), .A2(n19352), .B1(n19347), .B2(n19103), .ZN(
        n19090) );
  AOI221_X1 U22163 ( .B1(n19087), .B2(n19109), .C1(n19320), .C2(n19109), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n19088) );
  OAI21_X1 U22164 ( .B1(n19175), .B2(n19088), .A(n19323), .ZN(n19105) );
  AOI22_X1 U22165 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19346), .ZN(n19089) );
  OAI211_X1 U22166 ( .C1(n19355), .C2(n19108), .A(n19090), .B(n19089), .ZN(
        P3_U2900) );
  AOI22_X1 U22167 ( .A1(n19127), .A2(n19357), .B1(n19356), .B2(n19103), .ZN(
        n19092) );
  AOI22_X1 U22168 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19358), .ZN(n19091) );
  OAI211_X1 U22169 ( .C1(n19361), .C2(n19108), .A(n19092), .B(n19091), .ZN(
        P3_U2901) );
  AOI22_X1 U22170 ( .A1(n19127), .A2(n19364), .B1(n19362), .B2(n19103), .ZN(
        n19094) );
  AOI22_X1 U22171 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19363), .ZN(n19093) );
  OAI211_X1 U22172 ( .C1(n19367), .C2(n19108), .A(n19094), .B(n19093), .ZN(
        P3_U2902) );
  AOI22_X1 U22173 ( .A1(n19127), .A2(n19369), .B1(n19368), .B2(n19103), .ZN(
        n19096) );
  AOI22_X1 U22174 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19370), .ZN(n19095) );
  OAI211_X1 U22175 ( .C1(n19373), .C2(n19108), .A(n19096), .B(n19095), .ZN(
        P3_U2903) );
  AOI22_X1 U22176 ( .A1(n19104), .A2(n19376), .B1(n19374), .B2(n19103), .ZN(
        n19098) );
  AOI22_X1 U22177 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19105), .B1(
        n19127), .B2(n19375), .ZN(n19097) );
  OAI211_X1 U22178 ( .C1(n19379), .C2(n19108), .A(n19098), .B(n19097), .ZN(
        P3_U2904) );
  AOI22_X1 U22179 ( .A1(n19104), .A2(n19382), .B1(n19380), .B2(n19103), .ZN(
        n19100) );
  AOI22_X1 U22180 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19105), .B1(
        n19127), .B2(n19381), .ZN(n19099) );
  OAI211_X1 U22181 ( .C1(n19385), .C2(n19108), .A(n19100), .B(n19099), .ZN(
        P3_U2905) );
  AOI22_X1 U22182 ( .A1(n19104), .A2(n19388), .B1(n19386), .B2(n19103), .ZN(
        n19102) );
  AOI22_X1 U22183 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19105), .B1(
        n19127), .B2(n19387), .ZN(n19101) );
  OAI211_X1 U22184 ( .C1(n19391), .C2(n19108), .A(n19102), .B(n19101), .ZN(
        P3_U2906) );
  AOI22_X1 U22185 ( .A1(n19127), .A2(n21665), .B1(n21663), .B2(n19103), .ZN(
        n19107) );
  AOI22_X1 U22186 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19105), .B1(
        n19104), .B2(n19394), .ZN(n19106) );
  OAI211_X1 U22187 ( .C1(n21668), .C2(n19108), .A(n19107), .B(n19106), .ZN(
        P3_U2907) );
  NAND2_X1 U22188 ( .A1(n19268), .A2(n19131), .ZN(n19132) );
  NOR2_X1 U22189 ( .A1(n19155), .A2(n19203), .ZN(n19126) );
  AOI22_X1 U22190 ( .A1(n19352), .A2(n19150), .B1(n19347), .B2(n19126), .ZN(
        n19113) );
  AOI22_X1 U22191 ( .A1(n19351), .A2(n19111), .B1(n19131), .B2(n19110), .ZN(
        n19128) );
  AOI22_X1 U22192 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19128), .B1(
        n19127), .B2(n19346), .ZN(n19112) );
  OAI211_X1 U22193 ( .C1(n19355), .C2(n19132), .A(n19113), .B(n19112), .ZN(
        P3_U2908) );
  AOI22_X1 U22194 ( .A1(n19127), .A2(n19358), .B1(n19356), .B2(n19126), .ZN(
        n19115) );
  AOI22_X1 U22195 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19128), .B1(
        n19357), .B2(n19150), .ZN(n19114) );
  OAI211_X1 U22196 ( .C1(n19361), .C2(n19132), .A(n19115), .B(n19114), .ZN(
        P3_U2909) );
  AOI22_X1 U22197 ( .A1(n19127), .A2(n19363), .B1(n19362), .B2(n19126), .ZN(
        n19117) );
  AOI22_X1 U22198 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19128), .B1(
        n19364), .B2(n19150), .ZN(n19116) );
  OAI211_X1 U22199 ( .C1(n19367), .C2(n19132), .A(n19117), .B(n19116), .ZN(
        P3_U2910) );
  AOI22_X1 U22200 ( .A1(n19127), .A2(n19370), .B1(n19368), .B2(n19126), .ZN(
        n19119) );
  AOI22_X1 U22201 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19128), .B1(
        n19369), .B2(n19150), .ZN(n19118) );
  OAI211_X1 U22202 ( .C1(n19373), .C2(n19132), .A(n19119), .B(n19118), .ZN(
        P3_U2911) );
  AOI22_X1 U22203 ( .A1(n19375), .A2(n19150), .B1(n19374), .B2(n19126), .ZN(
        n19121) );
  AOI22_X1 U22204 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19128), .B1(
        n19127), .B2(n19376), .ZN(n19120) );
  OAI211_X1 U22205 ( .C1(n19379), .C2(n19132), .A(n19121), .B(n19120), .ZN(
        P3_U2912) );
  AOI22_X1 U22206 ( .A1(n19127), .A2(n19382), .B1(n19380), .B2(n19126), .ZN(
        n19123) );
  AOI22_X1 U22207 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19128), .B1(
        n19381), .B2(n19150), .ZN(n19122) );
  OAI211_X1 U22208 ( .C1(n19385), .C2(n19132), .A(n19123), .B(n19122), .ZN(
        P3_U2913) );
  AOI22_X1 U22209 ( .A1(n19387), .A2(n19150), .B1(n19386), .B2(n19126), .ZN(
        n19125) );
  AOI22_X1 U22210 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19128), .B1(
        n19127), .B2(n19388), .ZN(n19124) );
  OAI211_X1 U22211 ( .C1(n19391), .C2(n19132), .A(n19125), .B(n19124), .ZN(
        P3_U2914) );
  AOI22_X1 U22212 ( .A1(n19127), .A2(n19394), .B1(n21663), .B2(n19126), .ZN(
        n19130) );
  AOI22_X1 U22213 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19128), .B1(
        n21665), .B2(n19150), .ZN(n19129) );
  OAI211_X1 U22214 ( .C1(n21668), .C2(n19132), .A(n19130), .B(n19129), .ZN(
        P3_U2915) );
  NAND2_X1 U22215 ( .A1(n19269), .A2(n19131), .ZN(n19154) );
  NOR2_X1 U22216 ( .A1(n19198), .A2(n19220), .ZN(n19181) );
  NOR2_X1 U22217 ( .A1(n19318), .A2(n19181), .ZN(n19149) );
  AOI22_X1 U22218 ( .A1(n19352), .A2(n19175), .B1(n19347), .B2(n19149), .ZN(
        n19136) );
  NOR2_X1 U22219 ( .A1(n19150), .A2(n19175), .ZN(n19133) );
  OAI21_X1 U22220 ( .B1(n19133), .B2(n19320), .A(n19181), .ZN(n19134) );
  OAI211_X1 U22221 ( .C1(n19220), .C2(n19552), .A(n19323), .B(n19134), .ZN(
        n19151) );
  AOI22_X1 U22222 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19151), .B1(
        n19346), .B2(n19150), .ZN(n19135) );
  OAI211_X1 U22223 ( .C1(n19355), .C2(n19154), .A(n19136), .B(n19135), .ZN(
        P3_U2916) );
  AOI22_X1 U22224 ( .A1(n19357), .A2(n19175), .B1(n19356), .B2(n19149), .ZN(
        n19138) );
  AOI22_X1 U22225 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19151), .B1(
        n19358), .B2(n19150), .ZN(n19137) );
  OAI211_X1 U22226 ( .C1(n19361), .C2(n19154), .A(n19138), .B(n19137), .ZN(
        P3_U2917) );
  AOI22_X1 U22227 ( .A1(n19363), .A2(n19150), .B1(n19362), .B2(n19149), .ZN(
        n19140) );
  AOI22_X1 U22228 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19151), .B1(
        n19364), .B2(n19175), .ZN(n19139) );
  OAI211_X1 U22229 ( .C1(n19367), .C2(n19154), .A(n19140), .B(n19139), .ZN(
        P3_U2918) );
  AOI22_X1 U22230 ( .A1(n19369), .A2(n19175), .B1(n19368), .B2(n19149), .ZN(
        n19142) );
  AOI22_X1 U22231 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19151), .B1(
        n19370), .B2(n19150), .ZN(n19141) );
  OAI211_X1 U22232 ( .C1(n19373), .C2(n19154), .A(n19142), .B(n19141), .ZN(
        P3_U2919) );
  AOI22_X1 U22233 ( .A1(n19376), .A2(n19150), .B1(n19374), .B2(n19149), .ZN(
        n19144) );
  AOI22_X1 U22234 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19151), .B1(
        n19375), .B2(n19175), .ZN(n19143) );
  OAI211_X1 U22235 ( .C1(n19379), .C2(n19154), .A(n19144), .B(n19143), .ZN(
        P3_U2920) );
  AOI22_X1 U22236 ( .A1(n19381), .A2(n19175), .B1(n19380), .B2(n19149), .ZN(
        n19146) );
  AOI22_X1 U22237 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19151), .B1(
        n19382), .B2(n19150), .ZN(n19145) );
  OAI211_X1 U22238 ( .C1(n19385), .C2(n19154), .A(n19146), .B(n19145), .ZN(
        P3_U2921) );
  AOI22_X1 U22239 ( .A1(n19388), .A2(n19150), .B1(n19386), .B2(n19149), .ZN(
        n19148) );
  AOI22_X1 U22240 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19151), .B1(
        n19387), .B2(n19175), .ZN(n19147) );
  OAI211_X1 U22241 ( .C1(n19391), .C2(n19154), .A(n19148), .B(n19147), .ZN(
        P3_U2922) );
  AOI22_X1 U22242 ( .A1(n21665), .A2(n19175), .B1(n21663), .B2(n19149), .ZN(
        n19153) );
  AOI22_X1 U22243 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19151), .B1(
        n19394), .B2(n19150), .ZN(n19152) );
  OAI211_X1 U22244 ( .C1(n21668), .C2(n19154), .A(n19153), .B(n19152), .ZN(
        P3_U2923) );
  NOR2_X1 U22245 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19158), .ZN(
        n19204) );
  NAND2_X1 U22246 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19204), .ZN(
        n19178) );
  AOI211_X1 U22247 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n19419), .A(n19179), 
        .B(n19155), .ZN(n19157) );
  NAND2_X1 U22248 ( .A1(n19157), .A2(n19156), .ZN(n19174) );
  AOI22_X1 U22249 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19174), .B1(
        n19347), .B2(n19173), .ZN(n19160) );
  AOI22_X1 U22250 ( .A1(n19352), .A2(n19198), .B1(n19346), .B2(n19175), .ZN(
        n19159) );
  OAI211_X1 U22251 ( .C1(n19355), .C2(n19178), .A(n19160), .B(n19159), .ZN(
        P3_U2924) );
  AOI22_X1 U22252 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19174), .B1(
        n19356), .B2(n19173), .ZN(n19162) );
  AOI22_X1 U22253 ( .A1(n19357), .A2(n19198), .B1(n19358), .B2(n19175), .ZN(
        n19161) );
  OAI211_X1 U22254 ( .C1(n19361), .C2(n19178), .A(n19162), .B(n19161), .ZN(
        P3_U2925) );
  AOI22_X1 U22255 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19174), .B1(
        n19362), .B2(n19173), .ZN(n19164) );
  AOI22_X1 U22256 ( .A1(n19363), .A2(n19175), .B1(n19364), .B2(n19198), .ZN(
        n19163) );
  OAI211_X1 U22257 ( .C1(n19367), .C2(n19178), .A(n19164), .B(n19163), .ZN(
        P3_U2926) );
  AOI22_X1 U22258 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19174), .B1(
        n19368), .B2(n19173), .ZN(n19166) );
  AOI22_X1 U22259 ( .A1(n19369), .A2(n19198), .B1(n19370), .B2(n19175), .ZN(
        n19165) );
  OAI211_X1 U22260 ( .C1(n19373), .C2(n19178), .A(n19166), .B(n19165), .ZN(
        P3_U2927) );
  AOI22_X1 U22261 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19174), .B1(
        n19374), .B2(n19173), .ZN(n19168) );
  AOI22_X1 U22262 ( .A1(n19375), .A2(n19198), .B1(n19376), .B2(n19175), .ZN(
        n19167) );
  OAI211_X1 U22263 ( .C1(n19379), .C2(n19178), .A(n19168), .B(n19167), .ZN(
        P3_U2928) );
  AOI22_X1 U22264 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19174), .B1(
        n19380), .B2(n19173), .ZN(n19170) );
  AOI22_X1 U22265 ( .A1(n19381), .A2(n19198), .B1(n19382), .B2(n19175), .ZN(
        n19169) );
  OAI211_X1 U22266 ( .C1(n19385), .C2(n19178), .A(n19170), .B(n19169), .ZN(
        P3_U2929) );
  AOI22_X1 U22267 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19174), .B1(
        n19386), .B2(n19173), .ZN(n19172) );
  AOI22_X1 U22268 ( .A1(n19387), .A2(n19198), .B1(n19388), .B2(n19175), .ZN(
        n19171) );
  OAI211_X1 U22269 ( .C1(n19391), .C2(n19178), .A(n19172), .B(n19171), .ZN(
        P3_U2930) );
  AOI22_X1 U22270 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19174), .B1(
        n21663), .B2(n19173), .ZN(n19177) );
  AOI22_X1 U22271 ( .A1(n19394), .A2(n19175), .B1(n21665), .B2(n19198), .ZN(
        n19176) );
  OAI211_X1 U22272 ( .C1(n21668), .C2(n19178), .A(n19177), .B(n19176), .ZN(
        P3_U2931) );
  NOR2_X2 U22273 ( .A1(n19425), .A2(n19246), .ZN(n19264) );
  INV_X1 U22274 ( .A(n19264), .ZN(n19202) );
  NOR2_X1 U22275 ( .A1(n19241), .A2(n19264), .ZN(n19224) );
  NOR2_X1 U22276 ( .A1(n19318), .A2(n19224), .ZN(n19197) );
  AOI22_X1 U22277 ( .A1(n19352), .A2(n19220), .B1(n19347), .B2(n19197), .ZN(
        n19184) );
  OAI22_X1 U22278 ( .A1(n19181), .A2(n19180), .B1(n19224), .B2(n19179), .ZN(
        n19182) );
  OAI21_X1 U22279 ( .B1(n19264), .B2(n19552), .A(n19182), .ZN(n19199) );
  AOI22_X1 U22280 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19199), .B1(
        n19346), .B2(n19198), .ZN(n19183) );
  OAI211_X1 U22281 ( .C1(n19355), .C2(n19202), .A(n19184), .B(n19183), .ZN(
        P3_U2932) );
  AOI22_X1 U22282 ( .A1(n19357), .A2(n19220), .B1(n19356), .B2(n19197), .ZN(
        n19186) );
  AOI22_X1 U22283 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19199), .B1(
        n19358), .B2(n19198), .ZN(n19185) );
  OAI211_X1 U22284 ( .C1(n19361), .C2(n19202), .A(n19186), .B(n19185), .ZN(
        P3_U2933) );
  AOI22_X1 U22285 ( .A1(n19362), .A2(n19197), .B1(n19364), .B2(n19220), .ZN(
        n19188) );
  AOI22_X1 U22286 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19199), .B1(
        n19363), .B2(n19198), .ZN(n19187) );
  OAI211_X1 U22287 ( .C1(n19367), .C2(n19202), .A(n19188), .B(n19187), .ZN(
        P3_U2934) );
  AOI22_X1 U22288 ( .A1(n19369), .A2(n19220), .B1(n19368), .B2(n19197), .ZN(
        n19190) );
  AOI22_X1 U22289 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19199), .B1(
        n19370), .B2(n19198), .ZN(n19189) );
  OAI211_X1 U22290 ( .C1(n19373), .C2(n19202), .A(n19190), .B(n19189), .ZN(
        P3_U2935) );
  AOI22_X1 U22291 ( .A1(n19376), .A2(n19198), .B1(n19374), .B2(n19197), .ZN(
        n19192) );
  AOI22_X1 U22292 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19199), .B1(
        n19375), .B2(n19220), .ZN(n19191) );
  OAI211_X1 U22293 ( .C1(n19379), .C2(n19202), .A(n19192), .B(n19191), .ZN(
        P3_U2936) );
  AOI22_X1 U22294 ( .A1(n19382), .A2(n19198), .B1(n19380), .B2(n19197), .ZN(
        n19194) );
  AOI22_X1 U22295 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19199), .B1(
        n19381), .B2(n19220), .ZN(n19193) );
  OAI211_X1 U22296 ( .C1(n19385), .C2(n19202), .A(n19194), .B(n19193), .ZN(
        P3_U2937) );
  AOI22_X1 U22297 ( .A1(n19387), .A2(n19220), .B1(n19386), .B2(n19197), .ZN(
        n19196) );
  AOI22_X1 U22298 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19199), .B1(
        n19388), .B2(n19198), .ZN(n19195) );
  OAI211_X1 U22299 ( .C1(n19391), .C2(n19202), .A(n19196), .B(n19195), .ZN(
        P3_U2938) );
  AOI22_X1 U22300 ( .A1(n21665), .A2(n19220), .B1(n21663), .B2(n19197), .ZN(
        n19201) );
  AOI22_X1 U22301 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19199), .B1(
        n19394), .B2(n19198), .ZN(n19200) );
  OAI211_X1 U22302 ( .C1(n21668), .C2(n19202), .A(n19201), .B(n19200), .ZN(
        P3_U2939) );
  NAND2_X1 U22303 ( .A1(n19268), .A2(n19270), .ZN(n19247) );
  NOR2_X1 U22304 ( .A1(n19246), .A2(n19203), .ZN(n19219) );
  AOI22_X1 U22305 ( .A1(n19352), .A2(n19241), .B1(n19347), .B2(n19219), .ZN(
        n19206) );
  NOR2_X1 U22306 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19246), .ZN(
        n19248) );
  AOI22_X1 U22307 ( .A1(n19351), .A2(n19204), .B1(n19348), .B2(n19248), .ZN(
        n19221) );
  AOI22_X1 U22308 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19221), .B1(
        n19346), .B2(n19220), .ZN(n19205) );
  OAI211_X1 U22309 ( .C1(n19355), .C2(n19247), .A(n19206), .B(n19205), .ZN(
        P3_U2940) );
  AOI22_X1 U22310 ( .A1(n19356), .A2(n19219), .B1(n19358), .B2(n19220), .ZN(
        n19208) );
  AOI22_X1 U22311 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19221), .B1(
        n19357), .B2(n19241), .ZN(n19207) );
  OAI211_X1 U22312 ( .C1(n19361), .C2(n19247), .A(n19208), .B(n19207), .ZN(
        P3_U2941) );
  AOI22_X1 U22313 ( .A1(n19363), .A2(n19220), .B1(n19362), .B2(n19219), .ZN(
        n19210) );
  AOI22_X1 U22314 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19221), .B1(
        n19364), .B2(n19241), .ZN(n19209) );
  OAI211_X1 U22315 ( .C1(n19367), .C2(n19247), .A(n19210), .B(n19209), .ZN(
        P3_U2942) );
  AOI22_X1 U22316 ( .A1(n19370), .A2(n19220), .B1(n19368), .B2(n19219), .ZN(
        n19212) );
  AOI22_X1 U22317 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19221), .B1(
        n19369), .B2(n19241), .ZN(n19211) );
  OAI211_X1 U22318 ( .C1(n19373), .C2(n19247), .A(n19212), .B(n19211), .ZN(
        P3_U2943) );
  AOI22_X1 U22319 ( .A1(n19376), .A2(n19220), .B1(n19374), .B2(n19219), .ZN(
        n19214) );
  AOI22_X1 U22320 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19221), .B1(
        n19375), .B2(n19241), .ZN(n19213) );
  OAI211_X1 U22321 ( .C1(n19379), .C2(n19247), .A(n19214), .B(n19213), .ZN(
        P3_U2944) );
  AOI22_X1 U22322 ( .A1(n19382), .A2(n19220), .B1(n19380), .B2(n19219), .ZN(
        n19216) );
  AOI22_X1 U22323 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19221), .B1(
        n19381), .B2(n19241), .ZN(n19215) );
  OAI211_X1 U22324 ( .C1(n19385), .C2(n19247), .A(n19216), .B(n19215), .ZN(
        P3_U2945) );
  AOI22_X1 U22325 ( .A1(n19387), .A2(n19241), .B1(n19386), .B2(n19219), .ZN(
        n19218) );
  AOI22_X1 U22326 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19221), .B1(
        n19388), .B2(n19220), .ZN(n19217) );
  OAI211_X1 U22327 ( .C1(n19391), .C2(n19247), .A(n19218), .B(n19217), .ZN(
        P3_U2946) );
  AOI22_X1 U22328 ( .A1(n19394), .A2(n19220), .B1(n21663), .B2(n19219), .ZN(
        n19223) );
  AOI22_X1 U22329 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19221), .B1(
        n21665), .B2(n19241), .ZN(n19222) );
  OAI211_X1 U22330 ( .C1(n21668), .C2(n19247), .A(n19223), .B(n19222), .ZN(
        P3_U2947) );
  NAND2_X1 U22331 ( .A1(n19269), .A2(n19270), .ZN(n19245) );
  AOI21_X1 U22332 ( .B1(n19247), .B2(n19245), .A(n19318), .ZN(n19240) );
  AOI22_X1 U22333 ( .A1(n19347), .A2(n19240), .B1(n19346), .B2(n19241), .ZN(
        n19227) );
  INV_X1 U22334 ( .A(n19245), .ZN(n19313) );
  OAI211_X1 U22335 ( .C1(n19224), .C2(n19320), .A(n19247), .B(n19245), .ZN(
        n19225) );
  OAI211_X1 U22336 ( .C1(n19313), .C2(n19552), .A(n19323), .B(n19225), .ZN(
        n19242) );
  AOI22_X1 U22337 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19242), .B1(
        n19352), .B2(n19264), .ZN(n19226) );
  OAI211_X1 U22338 ( .C1(n19355), .C2(n19245), .A(n19227), .B(n19226), .ZN(
        P3_U2948) );
  AOI22_X1 U22339 ( .A1(n19357), .A2(n19264), .B1(n19356), .B2(n19240), .ZN(
        n19229) );
  AOI22_X1 U22340 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19242), .B1(
        n19358), .B2(n19241), .ZN(n19228) );
  OAI211_X1 U22341 ( .C1(n19361), .C2(n19245), .A(n19229), .B(n19228), .ZN(
        P3_U2949) );
  AOI22_X1 U22342 ( .A1(n19362), .A2(n19240), .B1(n19364), .B2(n19264), .ZN(
        n19231) );
  AOI22_X1 U22343 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19242), .B1(
        n19363), .B2(n19241), .ZN(n19230) );
  OAI211_X1 U22344 ( .C1(n19367), .C2(n19245), .A(n19231), .B(n19230), .ZN(
        P3_U2950) );
  AOI22_X1 U22345 ( .A1(n19370), .A2(n19241), .B1(n19368), .B2(n19240), .ZN(
        n19233) );
  AOI22_X1 U22346 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19242), .B1(
        n19369), .B2(n19264), .ZN(n19232) );
  OAI211_X1 U22347 ( .C1(n19373), .C2(n19245), .A(n19233), .B(n19232), .ZN(
        P3_U2951) );
  AOI22_X1 U22348 ( .A1(n19376), .A2(n19241), .B1(n19374), .B2(n19240), .ZN(
        n19235) );
  AOI22_X1 U22349 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19242), .B1(
        n19375), .B2(n19264), .ZN(n19234) );
  OAI211_X1 U22350 ( .C1(n19379), .C2(n19245), .A(n19235), .B(n19234), .ZN(
        P3_U2952) );
  AOI22_X1 U22351 ( .A1(n19382), .A2(n19241), .B1(n19380), .B2(n19240), .ZN(
        n19237) );
  AOI22_X1 U22352 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19242), .B1(
        n19381), .B2(n19264), .ZN(n19236) );
  OAI211_X1 U22353 ( .C1(n19385), .C2(n19245), .A(n19237), .B(n19236), .ZN(
        P3_U2953) );
  AOI22_X1 U22354 ( .A1(n19388), .A2(n19241), .B1(n19386), .B2(n19240), .ZN(
        n19239) );
  AOI22_X1 U22355 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19242), .B1(
        n19387), .B2(n19264), .ZN(n19238) );
  OAI211_X1 U22356 ( .C1(n19391), .C2(n19245), .A(n19239), .B(n19238), .ZN(
        P3_U2954) );
  AOI22_X1 U22357 ( .A1(n19394), .A2(n19241), .B1(n21663), .B2(n19240), .ZN(
        n19244) );
  AOI22_X1 U22358 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19242), .B1(
        n21665), .B2(n19264), .ZN(n19243) );
  OAI211_X1 U22359 ( .C1(n21668), .C2(n19245), .A(n19244), .B(n19243), .ZN(
        P3_U2955) );
  NOR2_X1 U22360 ( .A1(n13491), .A2(n19246), .ZN(n19297) );
  NAND2_X1 U22361 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19297), .ZN(
        n19272) );
  INV_X1 U22362 ( .A(n19247), .ZN(n19292) );
  AND2_X1 U22363 ( .A1(n19454), .A2(n19297), .ZN(n19263) );
  AOI22_X1 U22364 ( .A1(n19352), .A2(n19292), .B1(n19347), .B2(n19263), .ZN(
        n19250) );
  AOI22_X1 U22365 ( .A1(n19351), .A2(n19248), .B1(n19348), .B2(n19297), .ZN(
        n19265) );
  AOI22_X1 U22366 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19265), .B1(
        n19346), .B2(n19264), .ZN(n19249) );
  OAI211_X1 U22367 ( .C1(n19355), .C2(n19272), .A(n19250), .B(n19249), .ZN(
        P3_U2956) );
  AOI22_X1 U22368 ( .A1(n19356), .A2(n19263), .B1(n19358), .B2(n19264), .ZN(
        n19252) );
  AOI22_X1 U22369 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19265), .B1(
        n19357), .B2(n19292), .ZN(n19251) );
  OAI211_X1 U22370 ( .C1(n19361), .C2(n19272), .A(n19252), .B(n19251), .ZN(
        P3_U2957) );
  AOI22_X1 U22371 ( .A1(n19362), .A2(n19263), .B1(n19364), .B2(n19292), .ZN(
        n19254) );
  AOI22_X1 U22372 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19265), .B1(
        n19363), .B2(n19264), .ZN(n19253) );
  OAI211_X1 U22373 ( .C1(n19367), .C2(n19272), .A(n19254), .B(n19253), .ZN(
        P3_U2958) );
  AOI22_X1 U22374 ( .A1(n19370), .A2(n19264), .B1(n19368), .B2(n19263), .ZN(
        n19256) );
  AOI22_X1 U22375 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19265), .B1(
        n19369), .B2(n19292), .ZN(n19255) );
  OAI211_X1 U22376 ( .C1(n19373), .C2(n19272), .A(n19256), .B(n19255), .ZN(
        P3_U2959) );
  AOI22_X1 U22377 ( .A1(n19376), .A2(n19264), .B1(n19374), .B2(n19263), .ZN(
        n19258) );
  AOI22_X1 U22378 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19265), .B1(
        n19375), .B2(n19292), .ZN(n19257) );
  OAI211_X1 U22379 ( .C1(n19379), .C2(n19272), .A(n19258), .B(n19257), .ZN(
        P3_U2960) );
  AOI22_X1 U22380 ( .A1(n19382), .A2(n19264), .B1(n19380), .B2(n19263), .ZN(
        n19260) );
  AOI22_X1 U22381 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19265), .B1(
        n19381), .B2(n19292), .ZN(n19259) );
  OAI211_X1 U22382 ( .C1(n19385), .C2(n19272), .A(n19260), .B(n19259), .ZN(
        P3_U2961) );
  AOI22_X1 U22383 ( .A1(n19388), .A2(n19264), .B1(n19386), .B2(n19263), .ZN(
        n19262) );
  AOI22_X1 U22384 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19265), .B1(
        n19387), .B2(n19292), .ZN(n19261) );
  OAI211_X1 U22385 ( .C1(n19391), .C2(n19272), .A(n19262), .B(n19261), .ZN(
        P3_U2962) );
  AOI22_X1 U22386 ( .A1(n19394), .A2(n19264), .B1(n21663), .B2(n19263), .ZN(
        n19267) );
  AOI22_X1 U22387 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19265), .B1(
        n21665), .B2(n19292), .ZN(n19266) );
  OAI211_X1 U22388 ( .C1(n21668), .C2(n19272), .A(n19267), .B(n19266), .ZN(
        P3_U2963) );
  INV_X1 U22389 ( .A(n19296), .ZN(n19350) );
  NAND2_X1 U22390 ( .A1(n19350), .A2(n13509), .ZN(n19295) );
  INV_X1 U22391 ( .A(n19295), .ZN(n19393) );
  NOR2_X1 U22392 ( .A1(n19269), .A2(n19268), .ZN(n19274) );
  NAND2_X1 U22393 ( .A1(n19271), .A2(n19270), .ZN(n19273) );
  NOR2_X1 U22394 ( .A1(n19340), .A2(n19393), .ZN(n19321) );
  OAI21_X1 U22395 ( .B1(n19274), .B2(n19273), .A(n19321), .ZN(n19275) );
  OAI211_X1 U22396 ( .C1(n19393), .C2(n19552), .A(n19323), .B(n19275), .ZN(
        n19291) );
  NOR2_X1 U22397 ( .A1(n19318), .A2(n19321), .ZN(n19290) );
  AOI22_X1 U22398 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19291), .B1(
        n19347), .B2(n19290), .ZN(n19277) );
  AOI22_X1 U22399 ( .A1(n19352), .A2(n19313), .B1(n19346), .B2(n19292), .ZN(
        n19276) );
  OAI211_X1 U22400 ( .C1(n19355), .C2(n19295), .A(n19277), .B(n19276), .ZN(
        P3_U2964) );
  AOI22_X1 U22401 ( .A1(n19356), .A2(n19290), .B1(n19358), .B2(n19292), .ZN(
        n19279) );
  AOI22_X1 U22402 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19291), .B1(
        n19357), .B2(n19313), .ZN(n19278) );
  OAI211_X1 U22403 ( .C1(n19361), .C2(n19295), .A(n19279), .B(n19278), .ZN(
        P3_U2965) );
  AOI22_X1 U22404 ( .A1(n19363), .A2(n19292), .B1(n19362), .B2(n19290), .ZN(
        n19281) );
  AOI22_X1 U22405 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19291), .B1(
        n19364), .B2(n19313), .ZN(n19280) );
  OAI211_X1 U22406 ( .C1(n19367), .C2(n19295), .A(n19281), .B(n19280), .ZN(
        P3_U2966) );
  AOI22_X1 U22407 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19291), .B1(
        n19368), .B2(n19290), .ZN(n19283) );
  AOI22_X1 U22408 ( .A1(n19369), .A2(n19313), .B1(n19370), .B2(n19292), .ZN(
        n19282) );
  OAI211_X1 U22409 ( .C1(n19373), .C2(n19295), .A(n19283), .B(n19282), .ZN(
        P3_U2967) );
  AOI22_X1 U22410 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19291), .B1(
        n19374), .B2(n19290), .ZN(n19285) );
  AOI22_X1 U22411 ( .A1(n19375), .A2(n19313), .B1(n19376), .B2(n19292), .ZN(
        n19284) );
  OAI211_X1 U22412 ( .C1(n19379), .C2(n19295), .A(n19285), .B(n19284), .ZN(
        P3_U2968) );
  AOI22_X1 U22413 ( .A1(n19382), .A2(n19292), .B1(n19380), .B2(n19290), .ZN(
        n19287) );
  AOI22_X1 U22414 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19291), .B1(
        n19381), .B2(n19313), .ZN(n19286) );
  OAI211_X1 U22415 ( .C1(n19385), .C2(n19295), .A(n19287), .B(n19286), .ZN(
        P3_U2969) );
  AOI22_X1 U22416 ( .A1(n19387), .A2(n19313), .B1(n19386), .B2(n19290), .ZN(
        n19289) );
  AOI22_X1 U22417 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19291), .B1(
        n19388), .B2(n19292), .ZN(n19288) );
  OAI211_X1 U22418 ( .C1(n19391), .C2(n19295), .A(n19289), .B(n19288), .ZN(
        P3_U2970) );
  AOI22_X1 U22419 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19291), .B1(
        n21663), .B2(n19290), .ZN(n19294) );
  AOI22_X1 U22420 ( .A1(n19394), .A2(n19292), .B1(n21665), .B2(n19313), .ZN(
        n19293) );
  OAI211_X1 U22421 ( .C1(n21668), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P3_U2971) );
  NOR2_X1 U22422 ( .A1(n19318), .A2(n19296), .ZN(n19312) );
  AOI22_X1 U22423 ( .A1(n19352), .A2(n19340), .B1(n19347), .B2(n19312), .ZN(
        n19299) );
  AOI22_X1 U22424 ( .A1(n19351), .A2(n19297), .B1(n19350), .B2(n19348), .ZN(
        n19314) );
  AOI22_X1 U22425 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19314), .B1(
        n19346), .B2(n19313), .ZN(n19298) );
  OAI211_X1 U22426 ( .C1(n19355), .C2(n19317), .A(n19299), .B(n19298), .ZN(
        P3_U2972) );
  AOI22_X1 U22427 ( .A1(n19357), .A2(n19340), .B1(n19356), .B2(n19312), .ZN(
        n19301) );
  AOI22_X1 U22428 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19314), .B1(
        n19358), .B2(n19313), .ZN(n19300) );
  OAI211_X1 U22429 ( .C1(n19317), .C2(n19361), .A(n19301), .B(n19300), .ZN(
        P3_U2973) );
  AOI22_X1 U22430 ( .A1(n19362), .A2(n19312), .B1(n19364), .B2(n19340), .ZN(
        n19303) );
  AOI22_X1 U22431 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19314), .B1(
        n19363), .B2(n19313), .ZN(n19302) );
  OAI211_X1 U22432 ( .C1(n19317), .C2(n19367), .A(n19303), .B(n19302), .ZN(
        P3_U2974) );
  AOI22_X1 U22433 ( .A1(n19369), .A2(n19340), .B1(n19368), .B2(n19312), .ZN(
        n19305) );
  AOI22_X1 U22434 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19314), .B1(
        n19370), .B2(n19313), .ZN(n19304) );
  OAI211_X1 U22435 ( .C1(n19317), .C2(n19373), .A(n19305), .B(n19304), .ZN(
        P3_U2975) );
  AOI22_X1 U22436 ( .A1(n19375), .A2(n19340), .B1(n19374), .B2(n19312), .ZN(
        n19307) );
  AOI22_X1 U22437 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19314), .B1(
        n19376), .B2(n19313), .ZN(n19306) );
  OAI211_X1 U22438 ( .C1(n19317), .C2(n19379), .A(n19307), .B(n19306), .ZN(
        P3_U2976) );
  AOI22_X1 U22439 ( .A1(n19382), .A2(n19313), .B1(n19380), .B2(n19312), .ZN(
        n19309) );
  AOI22_X1 U22440 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19314), .B1(
        n19381), .B2(n19340), .ZN(n19308) );
  OAI211_X1 U22441 ( .C1(n19317), .C2(n19385), .A(n19309), .B(n19308), .ZN(
        P3_U2977) );
  AOI22_X1 U22442 ( .A1(n19387), .A2(n19340), .B1(n19386), .B2(n19312), .ZN(
        n19311) );
  AOI22_X1 U22443 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19314), .B1(
        n19388), .B2(n19313), .ZN(n19310) );
  OAI211_X1 U22444 ( .C1(n19317), .C2(n19391), .A(n19311), .B(n19310), .ZN(
        P3_U2978) );
  AOI22_X1 U22445 ( .A1(n19394), .A2(n19313), .B1(n21663), .B2(n19312), .ZN(
        n19316) );
  AOI22_X1 U22446 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19314), .B1(
        n21665), .B2(n19340), .ZN(n19315) );
  OAI211_X1 U22447 ( .C1(n21668), .C2(n19317), .A(n19316), .B(n19315), .ZN(
        P3_U2979) );
  NOR2_X1 U22448 ( .A1(n19318), .A2(n19319), .ZN(n19339) );
  AOI22_X1 U22449 ( .A1(n19347), .A2(n19339), .B1(n19346), .B2(n19340), .ZN(
        n19326) );
  OAI21_X1 U22450 ( .B1(n19321), .B2(n19320), .A(n19319), .ZN(n19322) );
  OAI211_X1 U22451 ( .C1(n19324), .C2(n19552), .A(n19323), .B(n19322), .ZN(
        n19341) );
  AOI22_X1 U22452 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19341), .B1(
        n19352), .B2(n19393), .ZN(n19325) );
  OAI211_X1 U22453 ( .C1(n19344), .C2(n19355), .A(n19326), .B(n19325), .ZN(
        P3_U2980) );
  AOI22_X1 U22454 ( .A1(n19357), .A2(n19393), .B1(n19356), .B2(n19339), .ZN(
        n19328) );
  AOI22_X1 U22455 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19341), .B1(
        n19358), .B2(n19340), .ZN(n19327) );
  OAI211_X1 U22456 ( .C1(n19344), .C2(n19361), .A(n19328), .B(n19327), .ZN(
        P3_U2981) );
  AOI22_X1 U22457 ( .A1(n19363), .A2(n19340), .B1(n19362), .B2(n19339), .ZN(
        n19330) );
  AOI22_X1 U22458 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19341), .B1(
        n19364), .B2(n19393), .ZN(n19329) );
  OAI211_X1 U22459 ( .C1(n19344), .C2(n19367), .A(n19330), .B(n19329), .ZN(
        P3_U2982) );
  AOI22_X1 U22460 ( .A1(n19370), .A2(n19340), .B1(n19368), .B2(n19339), .ZN(
        n19332) );
  AOI22_X1 U22461 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19341), .B1(
        n19369), .B2(n19393), .ZN(n19331) );
  OAI211_X1 U22462 ( .C1(n19344), .C2(n19373), .A(n19332), .B(n19331), .ZN(
        P3_U2983) );
  AOI22_X1 U22463 ( .A1(n19376), .A2(n19340), .B1(n19374), .B2(n19339), .ZN(
        n19334) );
  AOI22_X1 U22464 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19341), .B1(
        n19375), .B2(n19393), .ZN(n19333) );
  OAI211_X1 U22465 ( .C1(n19344), .C2(n19379), .A(n19334), .B(n19333), .ZN(
        P3_U2984) );
  AOI22_X1 U22466 ( .A1(n19381), .A2(n19393), .B1(n19380), .B2(n19339), .ZN(
        n19336) );
  AOI22_X1 U22467 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19341), .B1(
        n19382), .B2(n19340), .ZN(n19335) );
  OAI211_X1 U22468 ( .C1(n19344), .C2(n19385), .A(n19336), .B(n19335), .ZN(
        P3_U2985) );
  AOI22_X1 U22469 ( .A1(n19388), .A2(n19340), .B1(n19386), .B2(n19339), .ZN(
        n19338) );
  AOI22_X1 U22470 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19341), .B1(
        n19387), .B2(n19393), .ZN(n19337) );
  OAI211_X1 U22471 ( .C1(n19344), .C2(n19391), .A(n19338), .B(n19337), .ZN(
        P3_U2986) );
  AOI22_X1 U22472 ( .A1(n19394), .A2(n19340), .B1(n21663), .B2(n19339), .ZN(
        n19343) );
  AOI22_X1 U22473 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19341), .B1(
        n21665), .B2(n19393), .ZN(n19342) );
  OAI211_X1 U22474 ( .C1(n21668), .C2(n19344), .A(n19343), .B(n19342), .ZN(
        P3_U2987) );
  INV_X1 U22475 ( .A(n19345), .ZN(n21671) );
  AND2_X1 U22476 ( .A1(n19454), .A2(n19349), .ZN(n19392) );
  AOI22_X1 U22477 ( .A1(n19347), .A2(n19392), .B1(n19346), .B2(n19393), .ZN(
        n19354) );
  AOI22_X1 U22478 ( .A1(n19351), .A2(n19350), .B1(n19349), .B2(n19348), .ZN(
        n19396) );
  AOI22_X1 U22479 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19396), .B1(
        n19352), .B2(n19395), .ZN(n19353) );
  OAI211_X1 U22480 ( .C1(n21671), .C2(n19355), .A(n19354), .B(n19353), .ZN(
        P3_U2988) );
  AOI22_X1 U22481 ( .A1(n19395), .A2(n19357), .B1(n19356), .B2(n19392), .ZN(
        n19360) );
  AOI22_X1 U22482 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19396), .B1(
        n19358), .B2(n19393), .ZN(n19359) );
  OAI211_X1 U22483 ( .C1(n21671), .C2(n19361), .A(n19360), .B(n19359), .ZN(
        P3_U2989) );
  AOI22_X1 U22484 ( .A1(n19363), .A2(n19393), .B1(n19362), .B2(n19392), .ZN(
        n19366) );
  AOI22_X1 U22485 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19396), .B1(
        n19395), .B2(n19364), .ZN(n19365) );
  OAI211_X1 U22486 ( .C1(n21671), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P3_U2990) );
  AOI22_X1 U22487 ( .A1(n19395), .A2(n19369), .B1(n19368), .B2(n19392), .ZN(
        n19372) );
  AOI22_X1 U22488 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19396), .B1(
        n19370), .B2(n19393), .ZN(n19371) );
  OAI211_X1 U22489 ( .C1(n21671), .C2(n19373), .A(n19372), .B(n19371), .ZN(
        P3_U2991) );
  AOI22_X1 U22490 ( .A1(n19395), .A2(n19375), .B1(n19374), .B2(n19392), .ZN(
        n19378) );
  AOI22_X1 U22491 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19396), .B1(
        n19376), .B2(n19393), .ZN(n19377) );
  OAI211_X1 U22492 ( .C1(n21671), .C2(n19379), .A(n19378), .B(n19377), .ZN(
        P3_U2992) );
  AOI22_X1 U22493 ( .A1(n19395), .A2(n19381), .B1(n19380), .B2(n19392), .ZN(
        n19384) );
  AOI22_X1 U22494 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19396), .B1(
        n19382), .B2(n19393), .ZN(n19383) );
  OAI211_X1 U22495 ( .C1(n21671), .C2(n19385), .A(n19384), .B(n19383), .ZN(
        P3_U2993) );
  AOI22_X1 U22496 ( .A1(n19395), .A2(n19387), .B1(n19386), .B2(n19392), .ZN(
        n19390) );
  AOI22_X1 U22497 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19396), .B1(
        n19388), .B2(n19393), .ZN(n19389) );
  OAI211_X1 U22498 ( .C1(n21671), .C2(n19391), .A(n19390), .B(n19389), .ZN(
        P3_U2994) );
  AOI22_X1 U22499 ( .A1(n19394), .A2(n19393), .B1(n21663), .B2(n19392), .ZN(
        n19398) );
  AOI22_X1 U22500 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19396), .B1(
        n21665), .B2(n19395), .ZN(n19397) );
  OAI211_X1 U22501 ( .C1(n21671), .C2(n21668), .A(n19398), .B(n19397), .ZN(
        P3_U2995) );
  NOR2_X1 U22502 ( .A1(n19400), .A2(n19399), .ZN(n19402) );
  OAI222_X1 U22503 ( .A1(n19406), .A2(n19405), .B1(n19404), .B2(n19403), .C1(
        n19402), .C2(n19401), .ZN(n19564) );
  OAI21_X1 U22504 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n19407), .ZN(n19408) );
  OAI211_X1 U22505 ( .C1(n19410), .C2(n19418), .A(n19409), .B(n19408), .ZN(
        n19438) );
  INV_X1 U22506 ( .A(n19411), .ZN(n19413) );
  AOI21_X1 U22507 ( .B1(n19418), .B2(n19413), .A(n19412), .ZN(n19415) );
  OAI22_X1 U22508 ( .A1(n19415), .A2(n19414), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19418), .ZN(n19436) );
  NOR2_X1 U22509 ( .A1(n19418), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n19416) );
  AOI21_X1 U22510 ( .B1(n19418), .B2(n19417), .A(n19416), .ZN(n19431) );
  INV_X1 U22511 ( .A(n19419), .ZN(n19420) );
  NAND2_X1 U22512 ( .A1(n19421), .A2(n19420), .ZN(n19423) );
  INV_X1 U22513 ( .A(n19421), .ZN(n19422) );
  AOI22_X1 U22514 ( .A1(n19424), .A2(n19423), .B1(n19422), .B2(n13491), .ZN(
        n19428) );
  NAND2_X1 U22515 ( .A1(n19431), .A2(n19430), .ZN(n19426) );
  OAI211_X1 U22516 ( .C1(n19428), .C2(n19427), .A(n19426), .B(n19425), .ZN(
        n19429) );
  OAI211_X1 U22517 ( .C1(n19430), .C2(n19431), .A(n19429), .B(n19433), .ZN(
        n19435) );
  AOI21_X1 U22518 ( .B1(n19433), .B2(n19432), .A(n19431), .ZN(n19434) );
  AOI222_X1 U22519 ( .A1(n19436), .A2(n19435), .B1(n19436), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19435), .C2(n19434), .ZN(
        n19437) );
  NOR4_X1 U22520 ( .A1(n19439), .A2(n19564), .A3(n19438), .A4(n19437), .ZN(
        n19450) );
  INV_X1 U22521 ( .A(n19440), .ZN(n19448) );
  OAI211_X1 U22522 ( .C1(n19442), .C2(n19441), .A(n19568), .B(n19450), .ZN(
        n19455) );
  AND2_X1 U22523 ( .A1(n19455), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19553) );
  OAI211_X1 U22524 ( .C1(P3_STATE2_REG_2__SCAN_IN), .C2(n19572), .A(n19553), 
        .B(n19443), .ZN(n19446) );
  NOR2_X1 U22525 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19577) );
  AOI22_X1 U22526 ( .A1(n19444), .A2(n19577), .B1(n19467), .B2(n19565), .ZN(
        n19445) );
  NAND2_X1 U22527 ( .A1(n19446), .A2(n19445), .ZN(n19447) );
  OAI211_X1 U22528 ( .C1(n19450), .C2(n19449), .A(n19448), .B(n19447), .ZN(
        P3_U2996) );
  NAND2_X1 U22529 ( .A1(n19467), .A2(n19565), .ZN(n19458) );
  NAND2_X1 U22530 ( .A1(n21628), .A2(n19467), .ZN(n19453) );
  OR3_X1 U22531 ( .A1(n19452), .A2(n19451), .A3(n19453), .ZN(n19460) );
  NAND4_X1 U22532 ( .A1(n19456), .A2(n19455), .A3(n19454), .A4(n19453), .ZN(
        n19457) );
  NAND4_X1 U22533 ( .A1(n19459), .A2(n19458), .A3(n19460), .A4(n19457), .ZN(
        P3_U2997) );
  INV_X1 U22534 ( .A(n19577), .ZN(n19462) );
  AND4_X1 U22535 ( .A1(n19462), .A2(n19461), .A3(n19551), .A4(n19460), .ZN(
        P3_U2998) );
  AND2_X1 U22536 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19547), .ZN(
        P3_U2999) );
  AND2_X1 U22537 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19547), .ZN(
        P3_U3000) );
  AND2_X1 U22538 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19547), .ZN(
        P3_U3001) );
  AND2_X1 U22539 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19547), .ZN(
        P3_U3002) );
  AND2_X1 U22540 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19547), .ZN(
        P3_U3003) );
  INV_X1 U22541 ( .A(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21614) );
  NOR2_X1 U22542 ( .A1(n21614), .A2(n19550), .ZN(P3_U3004) );
  AND2_X1 U22543 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19547), .ZN(
        P3_U3005) );
  AND2_X1 U22544 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19547), .ZN(
        P3_U3006) );
  AND2_X1 U22545 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19547), .ZN(
        P3_U3007) );
  AND2_X1 U22546 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19547), .ZN(
        P3_U3008) );
  AND2_X1 U22547 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19547), .ZN(
        P3_U3009) );
  AND2_X1 U22548 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19547), .ZN(
        P3_U3010) );
  AND2_X1 U22549 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19547), .ZN(
        P3_U3011) );
  AND2_X1 U22550 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19547), .ZN(
        P3_U3012) );
  AND2_X1 U22551 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19547), .ZN(
        P3_U3013) );
  AND2_X1 U22552 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19547), .ZN(
        P3_U3014) );
  INV_X1 U22553 ( .A(P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21640) );
  NOR2_X1 U22554 ( .A1(n21640), .A2(n19550), .ZN(P3_U3015) );
  AND2_X1 U22555 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19547), .ZN(
        P3_U3016) );
  AND2_X1 U22556 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19547), .ZN(
        P3_U3017) );
  AND2_X1 U22557 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19547), .ZN(
        P3_U3018) );
  AND2_X1 U22558 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19547), .ZN(
        P3_U3019) );
  AND2_X1 U22559 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19547), .ZN(
        P3_U3020) );
  AND2_X1 U22560 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19547), .ZN(P3_U3021) );
  AND2_X1 U22561 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19547), .ZN(P3_U3022) );
  AND2_X1 U22562 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19547), .ZN(P3_U3023) );
  AND2_X1 U22563 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19547), .ZN(P3_U3024) );
  AND2_X1 U22564 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19547), .ZN(P3_U3025) );
  AND2_X1 U22565 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19547), .ZN(P3_U3026) );
  AND2_X1 U22566 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19547), .ZN(P3_U3027) );
  AND2_X1 U22567 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19547), .ZN(P3_U3028) );
  INV_X1 U22568 ( .A(HOLD), .ZN(n21423) );
  OAI21_X1 U22569 ( .B1(n19463), .B2(n21423), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19464) );
  AOI22_X1 U22570 ( .A1(n19479), .A2(n19480), .B1(n19581), .B2(n19464), .ZN(
        n19466) );
  NAND2_X1 U22571 ( .A1(n19465), .A2(NA), .ZN(n19475) );
  OAI211_X1 U22572 ( .C1(n19468), .C2(n19572), .A(n19466), .B(n19475), .ZN(
        P3_U3029) );
  INV_X1 U22573 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19579) );
  AOI21_X1 U22574 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n19579), .ZN(
        n19470) );
  NAND2_X1 U22575 ( .A1(n19467), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19474) );
  OAI21_X1 U22576 ( .B1(n21423), .B2(n19468), .A(n19474), .ZN(n19469) );
  OAI21_X1 U22577 ( .B1(n19470), .B2(n19469), .A(P3_STATE_REG_0__SCAN_IN), 
        .ZN(n19471) );
  OAI211_X1 U22578 ( .C1(n19581), .C2(n19572), .A(n19569), .B(n19471), .ZN(
        P3_U3030) );
  NOR2_X1 U22579 ( .A1(n19480), .A2(n21423), .ZN(n19473) );
  OAI22_X1 U22580 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19474), .ZN(n19472) );
  OAI22_X1 U22581 ( .A1(n19473), .A2(n19472), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19478) );
  INV_X1 U22582 ( .A(n19474), .ZN(n19476) );
  OAI211_X1 U22583 ( .C1(n19476), .C2(n19479), .A(n19475), .B(
        P3_STATE_REG_2__SCAN_IN), .ZN(n19477) );
  OAI21_X1 U22584 ( .B1(n19479), .B2(n19478), .A(n19477), .ZN(P3_U3031) );
  NAND2_X1 U22585 ( .A1(n19583), .A2(n19480), .ZN(n19534) );
  CLKBUF_X1 U22586 ( .A(n19534), .Z(n19535) );
  OAI222_X1 U22587 ( .A1(n19554), .A2(n19538), .B1(n19481), .B2(n19583), .C1(
        n14113), .C2(n19535), .ZN(P3_U3032) );
  OAI222_X1 U22588 ( .A1(n19534), .A2(n19483), .B1(n19482), .B2(n19583), .C1(
        n14113), .C2(n19538), .ZN(P3_U3033) );
  OAI222_X1 U22589 ( .A1(n19534), .A2(n19485), .B1(n19484), .B2(n19583), .C1(
        n19483), .C2(n19538), .ZN(P3_U3034) );
  OAI222_X1 U22590 ( .A1(n19534), .A2(n19488), .B1(n19486), .B2(n19583), .C1(
        n19485), .C2(n19538), .ZN(P3_U3035) );
  OAI222_X1 U22591 ( .A1(n19488), .A2(n19538), .B1(n19487), .B2(n19583), .C1(
        n14303), .C2(n19535), .ZN(P3_U3036) );
  OAI222_X1 U22592 ( .A1(n19534), .A2(n19490), .B1(n19489), .B2(n19583), .C1(
        n14303), .C2(n19538), .ZN(P3_U3037) );
  OAI222_X1 U22593 ( .A1(n19534), .A2(n14261), .B1(n19491), .B2(n19583), .C1(
        n19490), .C2(n19538), .ZN(P3_U3038) );
  OAI222_X1 U22594 ( .A1(n14261), .A2(n19538), .B1(n19492), .B2(n19583), .C1(
        n19493), .C2(n19535), .ZN(P3_U3039) );
  OAI222_X1 U22595 ( .A1(n19534), .A2(n19495), .B1(n19494), .B2(n19583), .C1(
        n19493), .C2(n19538), .ZN(P3_U3040) );
  OAI222_X1 U22596 ( .A1(n19535), .A2(n19497), .B1(n19496), .B2(n19583), .C1(
        n19495), .C2(n19538), .ZN(P3_U3041) );
  OAI222_X1 U22597 ( .A1(n19535), .A2(n19499), .B1(n19498), .B2(n19583), .C1(
        n19497), .C2(n19538), .ZN(P3_U3042) );
  OAI222_X1 U22598 ( .A1(n19535), .A2(n19501), .B1(n19500), .B2(n19583), .C1(
        n19499), .C2(n19538), .ZN(P3_U3043) );
  OAI222_X1 U22599 ( .A1(n19535), .A2(n19504), .B1(n19502), .B2(n19583), .C1(
        n19501), .C2(n19538), .ZN(P3_U3044) );
  OAI222_X1 U22600 ( .A1(n19504), .A2(n19538), .B1(n19503), .B2(n19583), .C1(
        n19505), .C2(n19535), .ZN(P3_U3045) );
  OAI222_X1 U22601 ( .A1(n19535), .A2(n19507), .B1(n19506), .B2(n19583), .C1(
        n19505), .C2(n19538), .ZN(P3_U3046) );
  OAI222_X1 U22602 ( .A1(n19535), .A2(n19510), .B1(n19508), .B2(n19583), .C1(
        n19507), .C2(n19538), .ZN(P3_U3047) );
  OAI222_X1 U22603 ( .A1(n19510), .A2(n19538), .B1(n19509), .B2(n19583), .C1(
        n19511), .C2(n19535), .ZN(P3_U3048) );
  OAI222_X1 U22604 ( .A1(n19534), .A2(n19514), .B1(n19512), .B2(n19583), .C1(
        n19511), .C2(n19538), .ZN(P3_U3049) );
  OAI222_X1 U22605 ( .A1(n19514), .A2(n19538), .B1(n19513), .B2(n19583), .C1(
        n19515), .C2(n19535), .ZN(P3_U3050) );
  OAI222_X1 U22606 ( .A1(n19534), .A2(n19518), .B1(n19516), .B2(n19583), .C1(
        n19515), .C2(n19538), .ZN(P3_U3051) );
  OAI222_X1 U22607 ( .A1(n19518), .A2(n19538), .B1(n19517), .B2(n19583), .C1(
        n21548), .C2(n19535), .ZN(P3_U3052) );
  INV_X1 U22608 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19521) );
  OAI222_X1 U22609 ( .A1(n19534), .A2(n19521), .B1(n19519), .B2(n19583), .C1(
        n21548), .C2(n19538), .ZN(P3_U3053) );
  OAI222_X1 U22610 ( .A1(n19521), .A2(n19538), .B1(n19520), .B2(n19583), .C1(
        n19522), .C2(n19535), .ZN(P3_U3054) );
  OAI222_X1 U22611 ( .A1(n19534), .A2(n19524), .B1(n19523), .B2(n19583), .C1(
        n19522), .C2(n19538), .ZN(P3_U3055) );
  OAI222_X1 U22612 ( .A1(n19534), .A2(n19526), .B1(n19525), .B2(n19583), .C1(
        n19524), .C2(n19538), .ZN(P3_U3056) );
  OAI222_X1 U22613 ( .A1(n19535), .A2(n19528), .B1(n19527), .B2(n19583), .C1(
        n19526), .C2(n19538), .ZN(P3_U3057) );
  OAI222_X1 U22614 ( .A1(n19535), .A2(n19531), .B1(n19529), .B2(n19583), .C1(
        n19528), .C2(n19538), .ZN(P3_U3058) );
  OAI222_X1 U22615 ( .A1(n19531), .A2(n19538), .B1(n19530), .B2(n19583), .C1(
        n19532), .C2(n19535), .ZN(P3_U3059) );
  OAI222_X1 U22616 ( .A1(n19534), .A2(n19537), .B1(n19533), .B2(n19583), .C1(
        n19532), .C2(n19538), .ZN(P3_U3060) );
  OAI222_X1 U22617 ( .A1(n19538), .A2(n19537), .B1(n21582), .B2(n19583), .C1(
        n19536), .C2(n19535), .ZN(P3_U3061) );
  INV_X1 U22618 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n19539) );
  AOI22_X1 U22619 ( .A1(n19583), .A2(n19540), .B1(n19539), .B2(n19581), .ZN(
        P3_U3274) );
  INV_X1 U22620 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19557) );
  INV_X1 U22621 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n19541) );
  AOI22_X1 U22622 ( .A1(n19583), .A2(n19557), .B1(n19541), .B2(n19581), .ZN(
        P3_U3275) );
  INV_X1 U22623 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n19542) );
  AOI22_X1 U22624 ( .A1(n19583), .A2(n19543), .B1(n19542), .B2(n19581), .ZN(
        P3_U3276) );
  INV_X1 U22625 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19560) );
  INV_X1 U22626 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n19544) );
  AOI22_X1 U22627 ( .A1(n19583), .A2(n19560), .B1(n19544), .B2(n19581), .ZN(
        P3_U3277) );
  INV_X1 U22628 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19546) );
  INV_X1 U22629 ( .A(n19548), .ZN(n19545) );
  AOI21_X1 U22630 ( .B1(n19547), .B2(n19546), .A(n19545), .ZN(P3_U3280) );
  OAI21_X1 U22631 ( .B1(n19550), .B2(n19549), .A(n19548), .ZN(P3_U3281) );
  OAI21_X1 U22632 ( .B1(n19553), .B2(n19552), .A(n19551), .ZN(P3_U3282) );
  AOI21_X1 U22633 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19555) );
  AOI22_X1 U22634 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n19555), .B2(n19554), .ZN(n19558) );
  AOI22_X1 U22635 ( .A1(n19561), .A2(n19558), .B1(n19557), .B2(n19556), .ZN(
        P3_U3292) );
  OAI21_X1 U22636 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n19561), .ZN(n19559) );
  OAI21_X1 U22637 ( .B1(n19561), .B2(n19560), .A(n19559), .ZN(P3_U3293) );
  INV_X1 U22638 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19562) );
  AOI22_X1 U22639 ( .A1(n19583), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19562), 
        .B2(n19581), .ZN(P3_U3294) );
  MUX2_X1 U22640 ( .A(P3_MORE_REG_SCAN_IN), .B(n19564), .S(n19563), .Z(
        P3_U3295) );
  AOI21_X1 U22641 ( .B1(n19565), .B2(n19572), .A(n19586), .ZN(n19566) );
  OAI21_X1 U22642 ( .B1(n19568), .B2(n19567), .A(n19566), .ZN(n19580) );
  AOI21_X1 U22643 ( .B1(n19571), .B2(n19570), .A(n19569), .ZN(n19573) );
  OAI211_X1 U22644 ( .C1(n19574), .C2(n19573), .A(n19572), .B(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n19575) );
  AND2_X1 U22645 ( .A1(n19575), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n19576) );
  OAI21_X1 U22646 ( .B1(n19577), .B2(n19576), .A(n19580), .ZN(n19578) );
  OAI21_X1 U22647 ( .B1(n19580), .B2(n19579), .A(n19578), .ZN(P3_U3296) );
  INV_X1 U22648 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19589) );
  INV_X1 U22649 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n19582) );
  AOI22_X1 U22650 ( .A1(n19583), .A2(n19589), .B1(n19582), .B2(n19581), .ZN(
        P3_U3297) );
  AOI21_X1 U22651 ( .B1(n19584), .B2(n21628), .A(n19586), .ZN(n19590) );
  INV_X1 U22652 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n19585) );
  AOI22_X1 U22653 ( .A1(n19587), .A2(n19586), .B1(n19590), .B2(n19585), .ZN(
        P3_U3298) );
  AOI21_X1 U22654 ( .B1(n19590), .B2(n19589), .A(n19588), .ZN(P3_U3299) );
  INV_X1 U22655 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n19592) );
  NAND2_X1 U22656 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20507), .ZN(n20500) );
  INV_X1 U22657 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19591) );
  NAND2_X1 U22658 ( .A1(n20496), .A2(n19591), .ZN(n20497) );
  OAI21_X1 U22659 ( .B1(n20496), .B2(n19592), .A(n20570), .ZN(P2_U2815) );
  INV_X1 U22660 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19593) );
  NAND2_X1 U22661 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20579), .ZN(n20482) );
  OAI22_X1 U22662 ( .A1(n19594), .A2(n19593), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n20482), .ZN(P2_U2816) );
  AOI21_X1 U22663 ( .B1(n20496), .B2(n20507), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19595) );
  AOI22_X1 U22664 ( .A1(n20618), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19595), 
        .B2(n20619), .ZN(P2_U2817) );
  OAI21_X1 U22665 ( .B1(n20490), .B2(BS16), .A(n20573), .ZN(n20571) );
  OAI21_X1 U22666 ( .B1(n20573), .B2(n19970), .A(n20571), .ZN(P2_U2818) );
  NOR2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21523) );
  AOI211_X1 U22668 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19596) );
  INV_X1 U22669 ( .A(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n21534) );
  INV_X1 U22670 ( .A(P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n21580) );
  AND4_X1 U22671 ( .A1(n21523), .A2(n19596), .A3(n21534), .A4(n21580), .ZN(
        n19604) );
  NOR4_X1 U22672 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_10__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19603) );
  NOR4_X1 U22673 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19602) );
  NOR4_X1 U22674 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19600) );
  NOR4_X1 U22675 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_15__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19599) );
  NOR4_X1 U22676 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19598) );
  NOR4_X1 U22677 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19597) );
  AND4_X1 U22678 ( .A1(n19600), .A2(n19599), .A3(n19598), .A4(n19597), .ZN(
        n19601) );
  NAND4_X1 U22679 ( .A1(n19604), .A2(n19603), .A3(n19602), .A4(n19601), .ZN(
        n19611) );
  NOR2_X1 U22680 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19611), .ZN(n19605) );
  INV_X1 U22681 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20568) );
  AOI22_X1 U22682 ( .A1(n19605), .A2(n19606), .B1(n19611), .B2(n20568), .ZN(
        P2_U2820) );
  INV_X1 U22683 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21542) );
  INV_X1 U22684 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20572) );
  NAND3_X1 U22685 ( .A1(n19606), .A2(n21542), .A3(n20572), .ZN(n19610) );
  INV_X1 U22686 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20566) );
  AOI22_X1 U22687 ( .A1(n19605), .A2(n19610), .B1(n19611), .B2(n20566), .ZN(
        P2_U2821) );
  NAND2_X1 U22688 ( .A1(n19605), .A2(n20572), .ZN(n19609) );
  INV_X1 U22689 ( .A(n19611), .ZN(n19612) );
  OAI21_X1 U22690 ( .B1(n19606), .B2(n20509), .A(n19612), .ZN(n19607) );
  OAI21_X1 U22691 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19612), .A(n19607), 
        .ZN(n19608) );
  OAI221_X1 U22692 ( .B1(n19609), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19609), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19608), .ZN(P2_U2822) );
  INV_X1 U22693 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20564) );
  OAI221_X1 U22694 ( .B1(n19612), .B2(n20564), .C1(n19611), .C2(n19610), .A(
        n19609), .ZN(P2_U2823) );
  NAND2_X1 U22695 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n19616) );
  NAND2_X1 U22696 ( .A1(n19784), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n19615) );
  NAND2_X1 U22697 ( .A1(n19613), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n19614) );
  NAND4_X1 U22698 ( .A1(n19616), .A2(n19701), .A3(n19615), .A4(n19614), .ZN(
        n19617) );
  AOI21_X1 U22699 ( .B1(n19618), .B2(n19736), .A(n19617), .ZN(n19628) );
  NOR2_X1 U22700 ( .A1(n19619), .A2(n19767), .ZN(n19620) );
  AOI21_X1 U22701 ( .B1(n19621), .B2(n19754), .A(n19620), .ZN(n19627) );
  OR2_X1 U22702 ( .A1(n19622), .A2(n19764), .ZN(n19624) );
  NAND2_X1 U22703 ( .A1(n19624), .A2(n19625), .ZN(n19623) );
  OAI211_X1 U22704 ( .C1(n19625), .C2(n19624), .A(n19771), .B(n19623), .ZN(
        n19626) );
  NAND3_X1 U22705 ( .A1(n19628), .A2(n19627), .A3(n19626), .ZN(P2_U2836) );
  NAND2_X1 U22706 ( .A1(n19784), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n19629) );
  OAI211_X1 U22707 ( .C1(n19630), .C2(n19778), .A(n19629), .B(n19701), .ZN(
        n19631) );
  AOI21_X1 U22708 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19777), .A(
        n19631), .ZN(n19632) );
  OAI21_X1 U22709 ( .B1(n19633), .B2(n19782), .A(n19632), .ZN(n19634) );
  INV_X1 U22710 ( .A(n19634), .ZN(n19644) );
  INV_X1 U22711 ( .A(n19635), .ZN(n19636) );
  AOI22_X1 U22712 ( .A1(n19637), .A2(n19754), .B1(n19636), .B2(n19785), .ZN(
        n19643) );
  NAND2_X1 U22713 ( .A1(n19638), .A2(n19790), .ZN(n19640) );
  NAND2_X1 U22714 ( .A1(n19640), .A2(n19641), .ZN(n19639) );
  OAI211_X1 U22715 ( .C1(n19641), .C2(n19640), .A(n19771), .B(n19639), .ZN(
        n19642) );
  NAND3_X1 U22716 ( .A1(n19644), .A2(n19643), .A3(n19642), .ZN(P2_U2837) );
  NAND2_X1 U22717 ( .A1(n19645), .A2(n19790), .ZN(n19646) );
  XNOR2_X1 U22718 ( .A(n19647), .B(n19646), .ZN(n19657) );
  NAND2_X1 U22719 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19650) );
  OAI21_X1 U22720 ( .B1(n19778), .B2(n20533), .A(n19701), .ZN(n19648) );
  INV_X1 U22721 ( .A(n19648), .ZN(n19649) );
  OAI211_X1 U22722 ( .C1(n19651), .C2(n12692), .A(n19650), .B(n19649), .ZN(
        n19652) );
  AOI21_X1 U22723 ( .B1(n19653), .B2(n19736), .A(n19652), .ZN(n19656) );
  AOI22_X1 U22724 ( .A1(n19654), .A2(n19754), .B1(n19803), .B2(n19785), .ZN(
        n19655) );
  OAI211_X1 U22725 ( .C1(n20488), .C2(n19657), .A(n19656), .B(n19655), .ZN(
        P2_U2839) );
  NAND2_X1 U22726 ( .A1(n19784), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n19658) );
  OAI211_X1 U22727 ( .C1(n20531), .C2(n19778), .A(n19658), .B(n19701), .ZN(
        n19659) );
  AOI21_X1 U22728 ( .B1(n19660), .B2(n19736), .A(n19659), .ZN(n19670) );
  NOR2_X1 U22729 ( .A1(n19661), .A2(n19764), .ZN(n19662) );
  XNOR2_X1 U22730 ( .A(n19663), .B(n19662), .ZN(n19668) );
  INV_X1 U22731 ( .A(n19664), .ZN(n19666) );
  OAI22_X1 U22732 ( .A1(n19666), .A2(n19786), .B1(n19665), .B2(n19767), .ZN(
        n19667) );
  AOI21_X1 U22733 ( .B1(n19668), .B2(n19771), .A(n19667), .ZN(n19669) );
  OAI211_X1 U22734 ( .C1(n19671), .C2(n19775), .A(n19670), .B(n19669), .ZN(
        P2_U2840) );
  OAI21_X1 U22735 ( .B1(n19672), .B2(n20488), .A(n19716), .ZN(n19679) );
  INV_X1 U22736 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n19675) );
  OAI21_X1 U22737 ( .B1(n19778), .B2(n20529), .A(n19701), .ZN(n19673) );
  AOI21_X1 U22738 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19784), .A(n19673), .ZN(
        n19674) );
  OAI21_X1 U22739 ( .B1(n19675), .B2(n19775), .A(n19674), .ZN(n19678) );
  NOR2_X1 U22740 ( .A1(n19676), .A2(n19782), .ZN(n19677) );
  AOI211_X1 U22741 ( .C1(n19686), .C2(n19679), .A(n19678), .B(n19677), .ZN(
        n19684) );
  INV_X1 U22742 ( .A(n19680), .ZN(n19681) );
  AOI22_X1 U22743 ( .A1(n19682), .A2(n19754), .B1(n19681), .B2(n19785), .ZN(
        n19683) );
  OAI211_X1 U22744 ( .C1(n19686), .C2(n19685), .A(n19684), .B(n19683), .ZN(
        P2_U2841) );
  INV_X1 U22745 ( .A(n19687), .ZN(n19688) );
  NOR2_X1 U22746 ( .A1(n19764), .A2(n19688), .ZN(n19711) );
  INV_X1 U22747 ( .A(n19711), .ZN(n19689) );
  XNOR2_X1 U22748 ( .A(n19690), .B(n19689), .ZN(n19700) );
  NAND2_X1 U22749 ( .A1(n19784), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n19691) );
  OAI211_X1 U22750 ( .C1(n20526), .C2(n19778), .A(n19691), .B(n19701), .ZN(
        n19692) );
  AOI21_X1 U22751 ( .B1(n19693), .B2(n19736), .A(n19692), .ZN(n19694) );
  INV_X1 U22752 ( .A(n19694), .ZN(n19695) );
  AOI21_X1 U22753 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19777), .A(
        n19695), .ZN(n19699) );
  AOI22_X1 U22754 ( .A1(n19697), .A2(n19754), .B1(n19696), .B2(n19785), .ZN(
        n19698) );
  OAI211_X1 U22755 ( .C1(n20488), .C2(n19700), .A(n19699), .B(n19698), .ZN(
        P2_U2843) );
  NAND2_X1 U22756 ( .A1(n19784), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n19702) );
  OAI211_X1 U22757 ( .C1(n19703), .C2(n19778), .A(n19702), .B(n19701), .ZN(
        n19704) );
  AOI21_X1 U22758 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19777), .A(
        n19704), .ZN(n19705) );
  OAI21_X1 U22759 ( .B1(n19706), .B2(n19782), .A(n19705), .ZN(n19709) );
  NOR2_X1 U22760 ( .A1(n19707), .A2(n19767), .ZN(n19708) );
  AOI211_X1 U22761 ( .C1(n19710), .C2(n19754), .A(n19709), .B(n19708), .ZN(
        n19714) );
  OAI211_X1 U22762 ( .C1(n19712), .C2(n19715), .A(n19771), .B(n19711), .ZN(
        n19713) );
  OAI211_X1 U22763 ( .C1(n19716), .C2(n19715), .A(n19714), .B(n19713), .ZN(
        P2_U2844) );
  NAND2_X1 U22764 ( .A1(n19790), .A2(n19717), .ZN(n19718) );
  XOR2_X1 U22765 ( .A(n19719), .B(n19718), .Z(n19730) );
  OAI21_X1 U22766 ( .B1(n19778), .B2(n20520), .A(n19701), .ZN(n19724) );
  INV_X1 U22767 ( .A(n19720), .ZN(n19722) );
  OAI22_X1 U22768 ( .A1(n19722), .A2(n19782), .B1(n19721), .B2(n19775), .ZN(
        n19723) );
  AOI211_X1 U22769 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19784), .A(n19724), .B(
        n19723), .ZN(n19729) );
  OAI22_X1 U22770 ( .A1(n19726), .A2(n19786), .B1(n19725), .B2(n19767), .ZN(
        n19727) );
  INV_X1 U22771 ( .A(n19727), .ZN(n19728) );
  OAI211_X1 U22772 ( .C1(n20488), .C2(n19730), .A(n19729), .B(n19728), .ZN(
        P2_U2847) );
  NOR2_X1 U22773 ( .A1(n19764), .A2(n19731), .ZN(n19732) );
  XOR2_X1 U22774 ( .A(n19733), .B(n19732), .Z(n19744) );
  NAND2_X1 U22775 ( .A1(n19784), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n19734) );
  OAI211_X1 U22776 ( .C1(n20518), .C2(n19778), .A(n19734), .B(n19701), .ZN(
        n19735) );
  AOI21_X1 U22777 ( .B1(n19737), .B2(n19736), .A(n19735), .ZN(n19738) );
  INV_X1 U22778 ( .A(n19738), .ZN(n19742) );
  OAI22_X1 U22779 ( .A1(n19740), .A2(n19786), .B1(n19739), .B2(n19767), .ZN(
        n19741) );
  AOI211_X1 U22780 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19777), .A(
        n19742), .B(n19741), .ZN(n19743) );
  OAI21_X1 U22781 ( .B1(n20488), .B2(n19744), .A(n19743), .ZN(P2_U2848) );
  NAND2_X1 U22782 ( .A1(n19790), .A2(n19745), .ZN(n19746) );
  XOR2_X1 U22783 ( .A(n19747), .B(n19746), .Z(n19758) );
  OAI21_X1 U22784 ( .B1(n19778), .B2(n20516), .A(n19701), .ZN(n19751) );
  OAI22_X1 U22785 ( .A1(n19749), .A2(n19782), .B1(n19775), .B2(n19748), .ZN(
        n19750) );
  AOI211_X1 U22786 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19784), .A(n19751), .B(
        n19750), .ZN(n19757) );
  INV_X1 U22787 ( .A(n19752), .ZN(n19753) );
  AOI22_X1 U22788 ( .A1(n19755), .A2(n19754), .B1(n19785), .B2(n19753), .ZN(
        n19756) );
  OAI211_X1 U22789 ( .C1(n20488), .C2(n19758), .A(n19757), .B(n19756), .ZN(
        P2_U2849) );
  INV_X1 U22790 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n19776) );
  OAI21_X1 U22791 ( .B1(n19778), .B2(n19759), .A(n19701), .ZN(n19762) );
  NOR2_X1 U22792 ( .A1(n19760), .A2(n19782), .ZN(n19761) );
  AOI211_X1 U22793 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19784), .A(n19762), .B(
        n19761), .ZN(n19774) );
  NOR2_X1 U22794 ( .A1(n19764), .A2(n19763), .ZN(n19765) );
  XNOR2_X1 U22795 ( .A(n19766), .B(n19765), .ZN(n19772) );
  OAI22_X1 U22796 ( .A1(n19769), .A2(n19786), .B1(n19768), .B2(n19767), .ZN(
        n19770) );
  AOI21_X1 U22797 ( .B1(n19772), .B2(n19771), .A(n19770), .ZN(n19773) );
  OAI211_X1 U22798 ( .C1(n19776), .C2(n19775), .A(n19774), .B(n19773), .ZN(
        P2_U2850) );
  NAND2_X1 U22799 ( .A1(n19777), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19781) );
  OAI21_X1 U22800 ( .B1(n19778), .B2(n19915), .A(n19701), .ZN(n19779) );
  INV_X1 U22801 ( .A(n19779), .ZN(n19780) );
  OAI211_X1 U22802 ( .C1(n19782), .C2(n19925), .A(n19781), .B(n19780), .ZN(
        n19783) );
  INV_X1 U22803 ( .A(n19783), .ZN(n19796) );
  INV_X1 U22804 ( .A(n19960), .ZN(n19807) );
  AOI22_X1 U22805 ( .A1(n19807), .A2(n19785), .B1(P2_EBX_REG_4__SCAN_IN), .B2(
        n19784), .ZN(n19795) );
  OAI22_X1 U22806 ( .A1(n19808), .A2(n19787), .B1(n19786), .B2(n19951), .ZN(
        n19788) );
  INV_X1 U22807 ( .A(n19788), .ZN(n19794) );
  AND2_X1 U22808 ( .A1(n19790), .A2(n19789), .ZN(n19792) );
  AOI21_X1 U22809 ( .B1(n19916), .B2(n19792), .A(n20488), .ZN(n19791) );
  OAI21_X1 U22810 ( .B1(n19916), .B2(n19792), .A(n19791), .ZN(n19793) );
  NAND4_X1 U22811 ( .A1(n19796), .A2(n19795), .A3(n19794), .A4(n19793), .ZN(
        P2_U2851) );
  AOI22_X1 U22812 ( .A1(n19798), .A2(n19797), .B1(n19813), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19806) );
  AOI22_X1 U22813 ( .A1(n19800), .A2(BUF1_REG_16__SCAN_IN), .B1(n19799), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19805) );
  INV_X1 U22814 ( .A(n19801), .ZN(n19802) );
  AOI22_X1 U22815 ( .A1(n19803), .A2(n19823), .B1(n19828), .B2(n19802), .ZN(
        n19804) );
  NAND3_X1 U22816 ( .A1(n19806), .A2(n19805), .A3(n19804), .ZN(P2_U2903) );
  AOI22_X1 U22817 ( .A1(n19824), .A2(n20001), .B1(n19823), .B2(n19807), .ZN(
        n19812) );
  XNOR2_X1 U22818 ( .A(n19809), .B(n19808), .ZN(n19810) );
  NAND2_X1 U22819 ( .A1(n19810), .A2(n19828), .ZN(n19811) );
  OAI211_X1 U22820 ( .C1(n19832), .C2(n19895), .A(n19812), .B(n19811), .ZN(
        P2_U2915) );
  AOI22_X1 U22821 ( .A1(n19814), .A2(n19823), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19813), .ZN(n19820) );
  OAI21_X1 U22822 ( .B1(n19817), .B2(n19816), .A(n19815), .ZN(n19818) );
  NAND2_X1 U22823 ( .A1(n19818), .A2(n19828), .ZN(n19819) );
  OAI211_X1 U22824 ( .C1(n19822), .C2(n19821), .A(n19820), .B(n19819), .ZN(
        P2_U2916) );
  INV_X1 U22825 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19899) );
  AOI22_X1 U22826 ( .A1(n19824), .A2(n19989), .B1(n19823), .B2(n20592), .ZN(
        n19831) );
  OAI21_X1 U22827 ( .B1(n19827), .B2(n19826), .A(n19825), .ZN(n19829) );
  NAND2_X1 U22828 ( .A1(n19829), .A2(n19828), .ZN(n19830) );
  OAI211_X1 U22829 ( .C1(n19832), .C2(n19899), .A(n19831), .B(n19830), .ZN(
        P2_U2917) );
  OR2_X1 U22830 ( .A1(n19833), .A2(n20481), .ZN(n19835) );
  NOR2_X1 U22831 ( .A1(n19852), .A2(n19838), .ZN(P2_U2920) );
  INV_X1 U22832 ( .A(n19905), .ZN(n19840) );
  INV_X1 U22833 ( .A(n19871), .ZN(n19850) );
  AOI22_X1 U22834 ( .A1(n19850), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19842) );
  OAI21_X1 U22835 ( .B1(n19852), .B2(n19843), .A(n19842), .ZN(P2_U2921) );
  INV_X1 U22836 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19845) );
  AOI22_X1 U22837 ( .A1(n19903), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n19844) );
  OAI21_X1 U22838 ( .B1(n19845), .B2(n19871), .A(n19844), .ZN(P2_U2922) );
  INV_X1 U22839 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19847) );
  AOI22_X1 U22840 ( .A1(n19903), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n19846) );
  OAI21_X1 U22841 ( .B1(n19847), .B2(n19871), .A(n19846), .ZN(P2_U2923) );
  INV_X1 U22842 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19849) );
  AOI22_X1 U22843 ( .A1(n19903), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n19848) );
  OAI21_X1 U22844 ( .B1(n19849), .B2(n19871), .A(n19848), .ZN(P2_U2924) );
  AOI22_X1 U22845 ( .A1(n19850), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n19851) );
  OAI21_X1 U22846 ( .B1(n19852), .B2(n21644), .A(n19851), .ZN(P2_U2925) );
  INV_X1 U22847 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19854) );
  AOI22_X1 U22848 ( .A1(n19903), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n19853) );
  OAI21_X1 U22849 ( .B1(n19854), .B2(n19871), .A(n19853), .ZN(P2_U2926) );
  INV_X1 U22850 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U22851 ( .A1(n19903), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_8__SCAN_IN), .ZN(n19855) );
  OAI21_X1 U22852 ( .B1(n19856), .B2(n19871), .A(n19855), .ZN(P2_U2927) );
  INV_X1 U22853 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19858) );
  AOI22_X1 U22854 ( .A1(n19903), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n19857) );
  OAI21_X1 U22855 ( .B1(n19858), .B2(n19871), .A(n19857), .ZN(P2_U2928) );
  AOI22_X1 U22856 ( .A1(n19903), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n19859) );
  OAI21_X1 U22857 ( .B1(n19860), .B2(n19871), .A(n19859), .ZN(P2_U2929) );
  INV_X1 U22858 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U22859 ( .A1(n19903), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U22860 ( .B1(n19862), .B2(n19871), .A(n19861), .ZN(P2_U2930) );
  AOI22_X1 U22861 ( .A1(n19903), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U22862 ( .B1(n19864), .B2(n19871), .A(n19863), .ZN(P2_U2931) );
  INV_X1 U22863 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U22864 ( .A1(n19903), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n19865) );
  OAI21_X1 U22865 ( .B1(n19866), .B2(n19871), .A(n19865), .ZN(P2_U2932) );
  AOI22_X1 U22866 ( .A1(n19903), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22867 ( .B1(n21632), .B2(n19871), .A(n19867), .ZN(P2_U2933) );
  INV_X1 U22868 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U22869 ( .A1(n19903), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n19868) );
  OAI21_X1 U22870 ( .B1(n19869), .B2(n19871), .A(n19868), .ZN(P2_U2934) );
  AOI22_X1 U22871 ( .A1(n19903), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n19902), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22872 ( .B1(n21566), .B2(n19871), .A(n19870), .ZN(P2_U2935) );
  AOI22_X1 U22873 ( .A1(n19903), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_15__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U22874 ( .B1(n19873), .B2(n19905), .A(n19872), .ZN(P2_U2936) );
  INV_X1 U22875 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19875) );
  AOI22_X1 U22876 ( .A1(n19903), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22877 ( .B1(n19875), .B2(n19905), .A(n19874), .ZN(P2_U2937) );
  AOI22_X1 U22878 ( .A1(n19903), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22879 ( .B1(n19877), .B2(n19905), .A(n19876), .ZN(P2_U2938) );
  AOI22_X1 U22880 ( .A1(n19903), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19878) );
  OAI21_X1 U22881 ( .B1(n19879), .B2(n19905), .A(n19878), .ZN(P2_U2939) );
  AOI22_X1 U22882 ( .A1(n19903), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n19880) );
  OAI21_X1 U22883 ( .B1(n19881), .B2(n19905), .A(n19880), .ZN(P2_U2940) );
  INV_X1 U22884 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U22885 ( .A1(n19903), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22886 ( .B1(n19883), .B2(n19905), .A(n19882), .ZN(P2_U2941) );
  AOI22_X1 U22887 ( .A1(n19903), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_9__SCAN_IN), .ZN(n19884) );
  OAI21_X1 U22888 ( .B1(n19885), .B2(n19905), .A(n19884), .ZN(P2_U2942) );
  AOI22_X1 U22889 ( .A1(n19903), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_8__SCAN_IN), .ZN(n19886) );
  OAI21_X1 U22890 ( .B1(n19887), .B2(n19905), .A(n19886), .ZN(P2_U2943) );
  AOI22_X1 U22891 ( .A1(n19903), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_7__SCAN_IN), .ZN(n19888) );
  OAI21_X1 U22892 ( .B1(n19889), .B2(n19905), .A(n19888), .ZN(P2_U2944) );
  AOI22_X1 U22893 ( .A1(n19903), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_6__SCAN_IN), .ZN(n19890) );
  OAI21_X1 U22894 ( .B1(n19891), .B2(n19905), .A(n19890), .ZN(P2_U2945) );
  INV_X1 U22895 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U22896 ( .A1(n19903), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n19892) );
  OAI21_X1 U22897 ( .B1(n19893), .B2(n19905), .A(n19892), .ZN(P2_U2946) );
  AOI22_X1 U22898 ( .A1(n19903), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_4__SCAN_IN), .ZN(n19894) );
  OAI21_X1 U22899 ( .B1(n19895), .B2(n19905), .A(n19894), .ZN(P2_U2947) );
  INV_X1 U22900 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U22901 ( .A1(n19903), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_3__SCAN_IN), .ZN(n19896) );
  OAI21_X1 U22902 ( .B1(n19897), .B2(n19905), .A(n19896), .ZN(P2_U2948) );
  AOI22_X1 U22903 ( .A1(n19903), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_2__SCAN_IN), .ZN(n19898) );
  OAI21_X1 U22904 ( .B1(n19899), .B2(n19905), .A(n19898), .ZN(P2_U2949) );
  INV_X1 U22905 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19901) );
  AOI22_X1 U22906 ( .A1(n19903), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19900) );
  OAI21_X1 U22907 ( .B1(n19901), .B2(n19905), .A(n19900), .ZN(P2_U2950) );
  AOI22_X1 U22908 ( .A1(n19903), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n19902), 
        .B2(P2_LWORD_REG_0__SCAN_IN), .ZN(n19904) );
  OAI21_X1 U22909 ( .B1(n12181), .B2(n19905), .A(n19904), .ZN(P2_U2951) );
  AOI22_X1 U22910 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n19907) );
  NAND2_X1 U22911 ( .A1(n19909), .A2(n19906), .ZN(n19911) );
  NAND2_X1 U22912 ( .A1(n19907), .A2(n19911), .ZN(P2_U2962) );
  AOI22_X1 U22913 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U22914 ( .A1(n19909), .A2(n19908), .ZN(n19913) );
  NAND2_X1 U22915 ( .A1(n19910), .A2(n19913), .ZN(P2_U2966) );
  AOI22_X1 U22916 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19912) );
  NAND2_X1 U22917 ( .A1(n19912), .A2(n19911), .ZN(P2_U2977) );
  AOI22_X1 U22918 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n13850), .B1(n13961), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19914) );
  NAND2_X1 U22919 ( .A1(n19914), .A2(n19913), .ZN(P2_U2981) );
  NOR2_X1 U22920 ( .A1(n19701), .A2(n19915), .ZN(n19956) );
  AOI21_X1 U22921 ( .B1(n19917), .B2(n19916), .A(n19956), .ZN(n19933) );
  XNOR2_X1 U22922 ( .A(n19918), .B(n19954), .ZN(n19919) );
  INV_X1 U22923 ( .A(n19920), .ZN(n19921) );
  NAND2_X1 U22924 ( .A1(n19922), .A2(n19921), .ZN(n19923) );
  NAND2_X1 U22925 ( .A1(n19924), .A2(n19923), .ZN(n19927) );
  XNOR2_X1 U22926 ( .A(n19925), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19926) );
  XNOR2_X1 U22927 ( .A(n19927), .B(n19926), .ZN(n19963) );
  NAND2_X1 U22928 ( .A1(n19963), .A2(n19936), .ZN(n19930) );
  OR2_X1 U22929 ( .A1(n19951), .A2(n19928), .ZN(n19929) );
  OAI211_X1 U22930 ( .C1(n19966), .C2(n19941), .A(n19930), .B(n19929), .ZN(
        n19931) );
  INV_X1 U22931 ( .A(n19931), .ZN(n19932) );
  OAI211_X1 U22932 ( .C1(n19934), .C2(n19950), .A(n19933), .B(n19932), .ZN(
        P2_U3010) );
  AND3_X1 U22933 ( .A1(n19937), .A2(n19936), .A3(n19935), .ZN(n19944) );
  INV_X1 U22934 ( .A(n19938), .ZN(n19940) );
  OAI22_X1 U22935 ( .A1(n19942), .A2(n19941), .B1(n19940), .B2(n19939), .ZN(
        n19943) );
  AOI211_X1 U22936 ( .C1(n19946), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        n19948) );
  OAI211_X1 U22937 ( .C1(n19950), .C2(n19949), .A(n19948), .B(n19947), .ZN(
        P2_U3012) );
  INV_X1 U22938 ( .A(n19951), .ZN(n19953) );
  AOI22_X1 U22939 ( .A1(n19955), .A2(n19954), .B1(n19953), .B2(n19952), .ZN(
        n19965) );
  AOI21_X1 U22940 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19957), .A(
        n19956), .ZN(n19958) );
  OAI21_X1 U22941 ( .B1(n19960), .B2(n19959), .A(n19958), .ZN(n19961) );
  AOI21_X1 U22942 ( .B1(n19963), .B2(n19962), .A(n19961), .ZN(n19964) );
  OAI211_X1 U22943 ( .C1(n19967), .C2(n19966), .A(n19965), .B(n19964), .ZN(
        P2_U3042) );
  NOR2_X4 U22944 ( .A1(n20246), .A2(n20049), .ZN(n20044) );
  INV_X1 U22945 ( .A(n20044), .ZN(n19969) );
  AND2_X1 U22946 ( .A1(n20382), .A2(n19969), .ZN(n19971) );
  AND2_X1 U22947 ( .A1(n20382), .A2(n19970), .ZN(n20270) );
  AOI21_X1 U22948 ( .B1(n19972), .B2(n19971), .A(n20270), .ZN(n19974) );
  AOI22_X1 U22949 ( .A1(n19974), .A2(n19973), .B1(n20392), .B2(n19978), .ZN(
        n19975) );
  NAND2_X1 U22950 ( .A1(n20586), .A2(n20594), .ZN(n20084) );
  OR2_X1 U22951 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20084), .ZN(
        n20023) );
  NOR2_X1 U22952 ( .A1(n20023), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20014) );
  INV_X1 U22953 ( .A(n19974), .ZN(n19979) );
  AOI22_X1 U22954 ( .A1(n20436), .A2(n20475), .B1(n20433), .B2(n20014), .ZN(
        n19982) );
  AOI21_X1 U22955 ( .B1(n19976), .B2(n20581), .A(n20382), .ZN(n19977) );
  AOI21_X1 U22956 ( .B1(n19979), .B2(n19978), .A(n19977), .ZN(n19980) );
  OAI21_X1 U22957 ( .B1(n19980), .B2(n20014), .A(n20397), .ZN(n20015) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20435), .ZN(n19981) );
  OAI211_X1 U22959 ( .C1(n20018), .C2(n20401), .A(n19982), .B(n19981), .ZN(
        P2_U3048) );
  NAND2_X1 U22960 ( .A1(n20397), .A2(n19983), .ZN(n20404) );
  OAI22_X2 U22961 ( .A1(n19984), .A2(n20007), .B1(n16018), .B2(n20005), .ZN(
        n20442) );
  NOR2_X2 U22962 ( .A1(n20004), .A2(n19985), .ZN(n20440) );
  AOI22_X1 U22963 ( .A1(n20442), .A2(n20475), .B1(n20440), .B2(n20014), .ZN(
        n19988) );
  OAI22_X2 U22964 ( .A1(n19986), .A2(n20007), .B1(n16076), .B2(n20005), .ZN(
        n20443) );
  AOI22_X1 U22965 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20443), .ZN(n19987) );
  OAI211_X1 U22966 ( .C1(n20018), .C2(n20404), .A(n19988), .B(n19987), .ZN(
        P2_U3049) );
  NAND2_X1 U22967 ( .A1(n20397), .A2(n19989), .ZN(n20407) );
  OAI22_X2 U22968 ( .A1(n19991), .A2(n20007), .B1(n19990), .B2(n20005), .ZN(
        n20450) );
  NOR2_X2 U22969 ( .A1(n20004), .A2(n19992), .ZN(n20447) );
  AOI22_X1 U22970 ( .A1(n20450), .A2(n20475), .B1(n20447), .B2(n20014), .ZN(
        n19994) );
  OAI22_X2 U22971 ( .A1(n21551), .A2(n20007), .B1(n16070), .B2(n20005), .ZN(
        n20449) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20449), .ZN(n19993) );
  OAI211_X1 U22973 ( .C1(n20018), .C2(n20407), .A(n19994), .B(n19993), .ZN(
        P2_U3050) );
  NAND2_X1 U22974 ( .A1(n20397), .A2(n19995), .ZN(n20410) );
  OAI22_X2 U22975 ( .A1(n14536), .A2(n20005), .B1(n19996), .B2(n20007), .ZN(
        n20456) );
  AOI22_X1 U22976 ( .A1(n20456), .A2(n20475), .B1(n9749), .B2(n20014), .ZN(
        n20000) );
  OAI22_X2 U22977 ( .A1(n19998), .A2(n20007), .B1(n16061), .B2(n20005), .ZN(
        n20457) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20457), .ZN(n19999) );
  OAI211_X1 U22979 ( .C1(n20018), .C2(n20410), .A(n20000), .B(n19999), .ZN(
        P2_U3051) );
  NAND2_X1 U22980 ( .A1(n20397), .A2(n20001), .ZN(n20413) );
  OAI22_X2 U22981 ( .A1(n16005), .A2(n20005), .B1(n20002), .B2(n20007), .ZN(
        n20463) );
  NOR2_X2 U22982 ( .A1(n20004), .A2(n20003), .ZN(n20461) );
  AOI22_X1 U22983 ( .A1(n20463), .A2(n20475), .B1(n20461), .B2(n20014), .ZN(
        n20009) );
  OAI22_X2 U22984 ( .A1(n16053), .A2(n20007), .B1(n20006), .B2(n20005), .ZN(
        n20464) );
  AOI22_X1 U22985 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20464), .ZN(n20008) );
  OAI211_X1 U22986 ( .C1(n20018), .C2(n20413), .A(n20009), .B(n20008), .ZN(
        P2_U3052) );
  AOI22_X1 U22987 ( .A1(n20415), .A2(n20475), .B1(n20414), .B2(n20014), .ZN(
        n20011) );
  AOI22_X1 U22988 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20416), .ZN(n20010) );
  OAI211_X1 U22989 ( .C1(n20018), .C2(n20419), .A(n20011), .B(n20010), .ZN(
        P2_U3053) );
  AOI22_X1 U22990 ( .A1(n20421), .A2(n20475), .B1(n20420), .B2(n20014), .ZN(
        n20013) );
  AOI22_X1 U22991 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20422), .ZN(n20012) );
  OAI211_X1 U22992 ( .C1(n20018), .C2(n20425), .A(n20013), .B(n20012), .ZN(
        P2_U3054) );
  AOI22_X1 U22993 ( .A1(n20472), .A2(n20475), .B1(n20468), .B2(n20014), .ZN(
        n20017) );
  AOI22_X1 U22994 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20015), .B1(
        n20044), .B2(n20474), .ZN(n20016) );
  OAI211_X1 U22995 ( .C1(n20018), .C2(n20431), .A(n20017), .B(n20016), .ZN(
        P2_U3055) );
  INV_X1 U22996 ( .A(n20246), .ZN(n20587) );
  NAND2_X1 U22997 ( .A1(n20182), .A2(n20587), .ZN(n20020) );
  NOR2_X1 U22998 ( .A1(n20237), .A2(n20084), .ZN(n20042) );
  AOI211_X1 U22999 ( .C1(n20021), .C2(n20581), .A(n20382), .B(n20042), .ZN(
        n20019) );
  INV_X1 U23000 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U23001 ( .B1(n20021), .B2(n20042), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20022) );
  AOI22_X1 U23002 ( .A1(n20043), .A2(n20434), .B1(n20433), .B2(n20042), .ZN(
        n20025) );
  AOI22_X1 U23003 ( .A1(n20044), .A2(n20436), .B1(n20078), .B2(n20435), .ZN(
        n20024) );
  OAI211_X1 U23004 ( .C1(n20048), .C2(n20026), .A(n20025), .B(n20024), .ZN(
        P2_U3056) );
  AOI22_X1 U23005 ( .A1(n20043), .A2(n20441), .B1(n20440), .B2(n20042), .ZN(
        n20028) );
  AOI22_X1 U23006 ( .A1(n20078), .A2(n20443), .B1(n20044), .B2(n20442), .ZN(
        n20027) );
  OAI211_X1 U23007 ( .C1(n20048), .C2(n12462), .A(n20028), .B(n20027), .ZN(
        P2_U3057) );
  INV_X1 U23008 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n20031) );
  AOI22_X1 U23009 ( .A1(n20043), .A2(n20448), .B1(n20447), .B2(n20042), .ZN(
        n20030) );
  AOI22_X1 U23010 ( .A1(n20044), .A2(n20450), .B1(n20078), .B2(n20449), .ZN(
        n20029) );
  OAI211_X1 U23011 ( .C1(n20048), .C2(n20031), .A(n20030), .B(n20029), .ZN(
        P2_U3058) );
  AOI22_X1 U23012 ( .A1(n20043), .A2(n20455), .B1(n9749), .B2(n20042), .ZN(
        n20033) );
  AOI22_X1 U23013 ( .A1(n20078), .A2(n20457), .B1(n20044), .B2(n20456), .ZN(
        n20032) );
  OAI211_X1 U23014 ( .C1(n20048), .C2(n20034), .A(n20033), .B(n20032), .ZN(
        P2_U3059) );
  INV_X1 U23015 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n20037) );
  AOI22_X1 U23016 ( .A1(n20043), .A2(n20462), .B1(n20461), .B2(n20042), .ZN(
        n20036) );
  AOI22_X1 U23017 ( .A1(n20078), .A2(n20464), .B1(n20044), .B2(n20463), .ZN(
        n20035) );
  OAI211_X1 U23018 ( .C1(n20048), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        P2_U3060) );
  AOI22_X1 U23019 ( .A1(n20043), .A2(n20373), .B1(n20414), .B2(n20042), .ZN(
        n20039) );
  AOI22_X1 U23020 ( .A1(n20044), .A2(n20415), .B1(n20078), .B2(n20416), .ZN(
        n20038) );
  OAI211_X1 U23021 ( .C1(n20048), .C2(n12478), .A(n20039), .B(n20038), .ZN(
        P2_U3061) );
  AOI22_X1 U23022 ( .A1(n20043), .A2(n20376), .B1(n20420), .B2(n20042), .ZN(
        n20041) );
  AOI22_X1 U23023 ( .A1(n20078), .A2(n20422), .B1(n20044), .B2(n20421), .ZN(
        n20040) );
  OAI211_X1 U23024 ( .C1(n20048), .C2(n21585), .A(n20041), .B(n20040), .ZN(
        P2_U3062) );
  INV_X1 U23025 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n20047) );
  AOI22_X1 U23026 ( .A1(n20043), .A2(n20470), .B1(n20468), .B2(n20042), .ZN(
        n20046) );
  AOI22_X1 U23027 ( .A1(n20078), .A2(n20474), .B1(n20044), .B2(n20472), .ZN(
        n20045) );
  OAI211_X1 U23028 ( .C1(n20048), .C2(n20047), .A(n20046), .B(n20045), .ZN(
        P2_U3063) );
  NOR2_X1 U23029 ( .A1(n20057), .A2(n20084), .ZN(n20050) );
  AOI221_X1 U23030 ( .B1(n10452), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n20078), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n20050), .ZN(n20054) );
  AOI21_X1 U23031 ( .B1(n20051), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20052) );
  NOR2_X1 U23032 ( .A1(n20274), .A2(n20084), .ZN(n20076) );
  OAI21_X1 U23033 ( .B1(n20052), .B2(n20076), .A(n20397), .ZN(n20053) );
  INV_X1 U23034 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U23035 ( .B1(n20055), .B2(n20076), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20056) );
  AOI22_X1 U23036 ( .A1(n20077), .A2(n20434), .B1(n20433), .B2(n20076), .ZN(
        n20059) );
  AOI22_X1 U23037 ( .A1(n20078), .A2(n20436), .B1(n10452), .B2(n20435), .ZN(
        n20058) );
  OAI211_X1 U23038 ( .C1(n20082), .C2(n20060), .A(n20059), .B(n20058), .ZN(
        P2_U3064) );
  AOI22_X1 U23039 ( .A1(n20077), .A2(n20441), .B1(n20440), .B2(n20076), .ZN(
        n20062) );
  AOI22_X1 U23040 ( .A1(n10452), .A2(n20443), .B1(n20078), .B2(n20442), .ZN(
        n20061) );
  OAI211_X1 U23041 ( .C1(n20082), .C2(n12460), .A(n20062), .B(n20061), .ZN(
        P2_U3065) );
  INV_X1 U23042 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20065) );
  AOI22_X1 U23043 ( .A1(n20077), .A2(n20448), .B1(n20447), .B2(n20076), .ZN(
        n20064) );
  AOI22_X1 U23044 ( .A1(n20078), .A2(n20450), .B1(n10452), .B2(n20449), .ZN(
        n20063) );
  OAI211_X1 U23045 ( .C1(n20082), .C2(n20065), .A(n20064), .B(n20063), .ZN(
        P2_U3066) );
  AOI22_X1 U23046 ( .A1(n20077), .A2(n20455), .B1(n9749), .B2(n20076), .ZN(
        n20067) );
  AOI22_X1 U23047 ( .A1(n10452), .A2(n20457), .B1(n20078), .B2(n20456), .ZN(
        n20066) );
  OAI211_X1 U23048 ( .C1(n20082), .C2(n12408), .A(n20067), .B(n20066), .ZN(
        P2_U3067) );
  INV_X1 U23049 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20070) );
  AOI22_X1 U23050 ( .A1(n20077), .A2(n20462), .B1(n20461), .B2(n20076), .ZN(
        n20069) );
  AOI22_X1 U23051 ( .A1(n10452), .A2(n20464), .B1(n20078), .B2(n20463), .ZN(
        n20068) );
  OAI211_X1 U23052 ( .C1(n20082), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P2_U3068) );
  AOI22_X1 U23053 ( .A1(n20077), .A2(n20373), .B1(n20414), .B2(n20076), .ZN(
        n20072) );
  AOI22_X1 U23054 ( .A1(n20078), .A2(n20415), .B1(n10452), .B2(n20416), .ZN(
        n20071) );
  OAI211_X1 U23055 ( .C1(n20082), .C2(n12483), .A(n20072), .B(n20071), .ZN(
        P2_U3069) );
  INV_X1 U23056 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n20075) );
  AOI22_X1 U23057 ( .A1(n20077), .A2(n20376), .B1(n20420), .B2(n20076), .ZN(
        n20074) );
  AOI22_X1 U23058 ( .A1(n10452), .A2(n20422), .B1(n20078), .B2(n20421), .ZN(
        n20073) );
  OAI211_X1 U23059 ( .C1(n20082), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        P2_U3070) );
  INV_X1 U23060 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20081) );
  AOI22_X1 U23061 ( .A1(n20077), .A2(n20470), .B1(n20468), .B2(n20076), .ZN(
        n20080) );
  AOI22_X1 U23062 ( .A1(n10452), .A2(n20474), .B1(n20078), .B2(n20472), .ZN(
        n20079) );
  OAI211_X1 U23063 ( .C1(n20082), .C2(n20081), .A(n20080), .B(n20079), .ZN(
        P2_U3071) );
  INV_X1 U23064 ( .A(n20308), .ZN(n20083) );
  AOI21_X1 U23065 ( .B1(n20182), .B2(n20083), .A(n20575), .ZN(n20092) );
  INV_X1 U23066 ( .A(n20084), .ZN(n20085) );
  AND2_X1 U23067 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20085), .ZN(
        n20090) );
  INV_X1 U23068 ( .A(n20109), .ZN(n20086) );
  AOI21_X1 U23069 ( .B1(n20089), .B2(n20086), .A(n20392), .ZN(n20087) );
  AOI22_X1 U23070 ( .A1(n20435), .A2(n20088), .B1(n20433), .B2(n20109), .ZN(
        n20096) );
  AOI21_X1 U23071 ( .B1(n20089), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20094) );
  INV_X1 U23072 ( .A(n20090), .ZN(n20091) );
  NAND2_X1 U23073 ( .A1(n20092), .A2(n20091), .ZN(n20093) );
  OAI211_X1 U23074 ( .C1(n20109), .C2(n20094), .A(n20093), .B(n20397), .ZN(
        n20110) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20110), .B1(
        n10452), .B2(n20436), .ZN(n20095) );
  OAI211_X1 U23076 ( .C1(n20113), .C2(n20401), .A(n20096), .B(n20095), .ZN(
        P2_U3072) );
  AOI22_X1 U23077 ( .A1(n20442), .A2(n10452), .B1(n20109), .B2(n20440), .ZN(
        n20098) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20110), .B1(
        n20088), .B2(n20443), .ZN(n20097) );
  OAI211_X1 U23079 ( .C1(n20113), .C2(n20404), .A(n20098), .B(n20097), .ZN(
        P2_U3073) );
  AOI22_X1 U23080 ( .A1(n20450), .A2(n10452), .B1(n20109), .B2(n20447), .ZN(
        n20100) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20110), .B1(
        n20088), .B2(n20449), .ZN(n20099) );
  OAI211_X1 U23082 ( .C1(n20113), .C2(n20407), .A(n20100), .B(n20099), .ZN(
        P2_U3074) );
  AOI22_X1 U23083 ( .A1(n20457), .A2(n20088), .B1(n20109), .B2(n9749), .ZN(
        n20102) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20110), .B1(
        n10452), .B2(n20456), .ZN(n20101) );
  OAI211_X1 U23085 ( .C1(n20113), .C2(n20410), .A(n20102), .B(n20101), .ZN(
        P2_U3075) );
  AOI22_X1 U23086 ( .A1(n20463), .A2(n10452), .B1(n20109), .B2(n20461), .ZN(
        n20104) );
  AOI22_X1 U23087 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20110), .B1(
        n20088), .B2(n20464), .ZN(n20103) );
  OAI211_X1 U23088 ( .C1(n20113), .C2(n20413), .A(n20104), .B(n20103), .ZN(
        P2_U3076) );
  AOI22_X1 U23089 ( .A1(n20416), .A2(n20088), .B1(n20414), .B2(n20109), .ZN(
        n20106) );
  AOI22_X1 U23090 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20110), .B1(
        n10452), .B2(n20415), .ZN(n20105) );
  OAI211_X1 U23091 ( .C1(n20113), .C2(n20419), .A(n20106), .B(n20105), .ZN(
        P2_U3077) );
  AOI22_X1 U23092 ( .A1(n20422), .A2(n20088), .B1(n20420), .B2(n20109), .ZN(
        n20108) );
  AOI22_X1 U23093 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20110), .B1(
        n10452), .B2(n20421), .ZN(n20107) );
  OAI211_X1 U23094 ( .C1(n20113), .C2(n20425), .A(n20108), .B(n20107), .ZN(
        P2_U3078) );
  AOI22_X1 U23095 ( .A1(n20472), .A2(n10452), .B1(n20468), .B2(n20109), .ZN(
        n20112) );
  AOI22_X1 U23096 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20110), .B1(
        n20088), .B2(n20474), .ZN(n20111) );
  OAI211_X1 U23097 ( .C1(n20113), .C2(n20431), .A(n20112), .B(n20111), .ZN(
        P2_U3079) );
  INV_X1 U23098 ( .A(n20435), .ZN(n20314) );
  NAND3_X1 U23099 ( .A1(n20117), .A2(n20586), .A3(n20581), .ZN(n20116) );
  NOR2_X1 U23100 ( .A1(n20114), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20136) );
  NOR3_X1 U23101 ( .A1(n20115), .A2(n20136), .A3(n20392), .ZN(n20118) );
  AOI22_X1 U23102 ( .A1(n20137), .A2(n20434), .B1(n20433), .B2(n20136), .ZN(
        n20123) );
  OAI21_X1 U23103 ( .B1(n20088), .B2(n20157), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20120) );
  NAND2_X1 U23104 ( .A1(n20117), .A2(n20586), .ZN(n20119) );
  AOI211_X1 U23105 ( .C1(n20120), .C2(n20119), .A(n20183), .B(n20118), .ZN(
        n20121) );
  AOI22_X1 U23106 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20436), .ZN(n20122) );
  OAI211_X1 U23107 ( .C1(n20314), .C2(n16720), .A(n20123), .B(n20122), .ZN(
        P2_U3080) );
  INV_X1 U23108 ( .A(n20443), .ZN(n20317) );
  AOI22_X1 U23109 ( .A1(n20137), .A2(n20441), .B1(n20440), .B2(n20136), .ZN(
        n20125) );
  AOI22_X1 U23110 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20442), .ZN(n20124) );
  OAI211_X1 U23111 ( .C1(n20317), .C2(n16720), .A(n20125), .B(n20124), .ZN(
        P2_U3081) );
  INV_X1 U23112 ( .A(n20449), .ZN(n20320) );
  AOI22_X1 U23113 ( .A1(n20137), .A2(n20448), .B1(n20447), .B2(n20136), .ZN(
        n20127) );
  AOI22_X1 U23114 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20450), .ZN(n20126) );
  OAI211_X1 U23115 ( .C1(n20320), .C2(n16720), .A(n20127), .B(n20126), .ZN(
        P2_U3082) );
  INV_X1 U23116 ( .A(n20457), .ZN(n20323) );
  AOI22_X1 U23117 ( .A1(n20137), .A2(n20455), .B1(n9749), .B2(n20136), .ZN(
        n20129) );
  AOI22_X1 U23118 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20456), .ZN(n20128) );
  OAI211_X1 U23119 ( .C1(n20323), .C2(n16720), .A(n20129), .B(n20128), .ZN(
        P2_U3083) );
  INV_X1 U23120 ( .A(n20464), .ZN(n20326) );
  AOI22_X1 U23121 ( .A1(n20137), .A2(n20462), .B1(n20461), .B2(n20136), .ZN(
        n20131) );
  AOI22_X1 U23122 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20463), .ZN(n20130) );
  OAI211_X1 U23123 ( .C1(n20326), .C2(n16720), .A(n20131), .B(n20130), .ZN(
        P2_U3084) );
  INV_X1 U23124 ( .A(n20416), .ZN(n20329) );
  AOI22_X1 U23125 ( .A1(n20137), .A2(n20373), .B1(n20414), .B2(n20136), .ZN(
        n20133) );
  AOI22_X1 U23126 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20415), .ZN(n20132) );
  OAI211_X1 U23127 ( .C1(n20329), .C2(n16720), .A(n20133), .B(n20132), .ZN(
        P2_U3085) );
  INV_X1 U23128 ( .A(n20422), .ZN(n20332) );
  AOI22_X1 U23129 ( .A1(n20137), .A2(n20376), .B1(n20420), .B2(n20136), .ZN(
        n20135) );
  AOI22_X1 U23130 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20421), .ZN(n20134) );
  OAI211_X1 U23131 ( .C1(n20332), .C2(n16720), .A(n20135), .B(n20134), .ZN(
        P2_U3086) );
  INV_X1 U23132 ( .A(n20474), .ZN(n20340) );
  AOI22_X1 U23133 ( .A1(n20137), .A2(n20470), .B1(n20468), .B2(n20136), .ZN(
        n20140) );
  AOI22_X1 U23134 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20138), .B1(
        n20088), .B2(n20472), .ZN(n20139) );
  OAI211_X1 U23135 ( .C1(n20340), .C2(n16720), .A(n20140), .B(n20139), .ZN(
        P2_U3087) );
  AOI22_X1 U23136 ( .A1(n20442), .A2(n20157), .B1(n20156), .B2(n20440), .ZN(
        n20142) );
  AOI22_X1 U23137 ( .A1(n20441), .A2(n20158), .B1(n10453), .B2(n20443), .ZN(
        n20141) );
  OAI211_X1 U23138 ( .C1(n20162), .C2(n12450), .A(n20142), .B(n20141), .ZN(
        P2_U3089) );
  INV_X1 U23139 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20145) );
  AOI22_X1 U23140 ( .A1(n20450), .A2(n20157), .B1(n20156), .B2(n20447), .ZN(
        n20144) );
  AOI22_X1 U23141 ( .A1(n20448), .A2(n20158), .B1(n10453), .B2(n20449), .ZN(
        n20143) );
  OAI211_X1 U23142 ( .C1(n20162), .C2(n20145), .A(n20144), .B(n20143), .ZN(
        P2_U3090) );
  AOI22_X1 U23143 ( .A1(n20457), .A2(n10453), .B1(n20156), .B2(n9749), .ZN(
        n20147) );
  AOI22_X1 U23144 ( .A1(n20455), .A2(n20158), .B1(n20157), .B2(n20456), .ZN(
        n20146) );
  OAI211_X1 U23145 ( .C1(n20162), .C2(n12414), .A(n20147), .B(n20146), .ZN(
        P2_U3091) );
  INV_X1 U23146 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U23147 ( .A1(n20463), .A2(n20157), .B1(n20156), .B2(n20461), .ZN(
        n20149) );
  AOI22_X1 U23148 ( .A1(n20462), .A2(n20158), .B1(n10453), .B2(n20464), .ZN(
        n20148) );
  OAI211_X1 U23149 ( .C1(n20162), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        P2_U3092) );
  AOI22_X1 U23150 ( .A1(n20415), .A2(n20157), .B1(n20156), .B2(n20414), .ZN(
        n20152) );
  AOI22_X1 U23151 ( .A1(n20373), .A2(n20158), .B1(n10453), .B2(n20416), .ZN(
        n20151) );
  OAI211_X1 U23152 ( .C1(n20162), .C2(n12485), .A(n20152), .B(n20151), .ZN(
        P2_U3093) );
  INV_X1 U23153 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n20155) );
  AOI22_X1 U23154 ( .A1(n20422), .A2(n10453), .B1(n20156), .B2(n20420), .ZN(
        n20154) );
  AOI22_X1 U23155 ( .A1(n20376), .A2(n20158), .B1(n20157), .B2(n20421), .ZN(
        n20153) );
  OAI211_X1 U23156 ( .C1(n20162), .C2(n20155), .A(n20154), .B(n20153), .ZN(
        P2_U3094) );
  INV_X1 U23157 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n20161) );
  AOI22_X1 U23158 ( .A1(n20474), .A2(n10453), .B1(n20156), .B2(n20468), .ZN(
        n20160) );
  AOI22_X1 U23159 ( .A1(n20470), .A2(n20158), .B1(n20157), .B2(n20472), .ZN(
        n20159) );
  OAI211_X1 U23160 ( .C1(n20162), .C2(n20161), .A(n20160), .B(n20159), .ZN(
        P2_U3095) );
  AOI22_X1 U23161 ( .A1(n20174), .A2(n20441), .B1(n20173), .B2(n20440), .ZN(
        n20164) );
  AOI22_X1 U23162 ( .A1(n20202), .A2(n20443), .B1(n10453), .B2(n20442), .ZN(
        n20163) );
  OAI211_X1 U23163 ( .C1(n20177), .C2(n12452), .A(n20164), .B(n20163), .ZN(
        P2_U3097) );
  INV_X1 U23164 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n20167) );
  AOI22_X1 U23165 ( .A1(n20174), .A2(n20448), .B1(n20173), .B2(n20447), .ZN(
        n20166) );
  AOI22_X1 U23166 ( .A1(n10453), .A2(n20450), .B1(n20202), .B2(n20449), .ZN(
        n20165) );
  OAI211_X1 U23167 ( .C1(n20177), .C2(n20167), .A(n20166), .B(n20165), .ZN(
        P2_U3098) );
  AOI22_X1 U23168 ( .A1(n20174), .A2(n20455), .B1(n20173), .B2(n20454), .ZN(
        n20169) );
  AOI22_X1 U23169 ( .A1(n20202), .A2(n20457), .B1(n10453), .B2(n20456), .ZN(
        n20168) );
  OAI211_X1 U23170 ( .C1(n20177), .C2(n12421), .A(n20169), .B(n20168), .ZN(
        P2_U3099) );
  INV_X1 U23171 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n20172) );
  AOI22_X1 U23172 ( .A1(n20174), .A2(n20462), .B1(n20173), .B2(n20461), .ZN(
        n20171) );
  AOI22_X1 U23173 ( .A1(n20202), .A2(n20464), .B1(n10453), .B2(n20463), .ZN(
        n20170) );
  OAI211_X1 U23174 ( .C1(n20177), .C2(n20172), .A(n20171), .B(n20170), .ZN(
        P2_U3100) );
  AOI22_X1 U23175 ( .A1(n20174), .A2(n20373), .B1(n20173), .B2(n20414), .ZN(
        n20176) );
  AOI22_X1 U23176 ( .A1(n10453), .A2(n20415), .B1(n20202), .B2(n20416), .ZN(
        n20175) );
  OAI211_X1 U23177 ( .C1(n20177), .C2(n12490), .A(n20176), .B(n20175), .ZN(
        P2_U3101) );
  NOR3_X1 U23178 ( .A1(n20179), .A2(n20213), .A3(n20392), .ZN(n20184) );
  AOI21_X1 U23179 ( .B1(n20181), .B2(n20581), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20180) );
  AOI22_X1 U23180 ( .A1(n20201), .A2(n20434), .B1(n20433), .B2(n20213), .ZN(
        n20188) );
  AOI21_X1 U23181 ( .B1(n20182), .B2(n20577), .A(n20181), .ZN(n20185) );
  NOR3_X1 U23182 ( .A1(n20185), .A2(n20184), .A3(n20183), .ZN(n20186) );
  AOI22_X1 U23183 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20436), .ZN(n20187) );
  OAI211_X1 U23184 ( .C1(n20314), .C2(n20206), .A(n20188), .B(n20187), .ZN(
        P2_U3104) );
  AOI22_X1 U23185 ( .A1(n20201), .A2(n20441), .B1(n20213), .B2(n20440), .ZN(
        n20190) );
  AOI22_X1 U23186 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20442), .ZN(n20189) );
  OAI211_X1 U23187 ( .C1(n20317), .C2(n20206), .A(n20190), .B(n20189), .ZN(
        P2_U3105) );
  AOI22_X1 U23188 ( .A1(n20201), .A2(n20448), .B1(n20213), .B2(n20447), .ZN(
        n20192) );
  AOI22_X1 U23189 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20450), .ZN(n20191) );
  OAI211_X1 U23190 ( .C1(n20320), .C2(n20206), .A(n20192), .B(n20191), .ZN(
        P2_U3106) );
  AOI22_X1 U23191 ( .A1(n20201), .A2(n20455), .B1(n20213), .B2(n20454), .ZN(
        n20194) );
  AOI22_X1 U23192 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20456), .ZN(n20193) );
  OAI211_X1 U23193 ( .C1(n20323), .C2(n20206), .A(n20194), .B(n20193), .ZN(
        P2_U3107) );
  AOI22_X1 U23194 ( .A1(n20201), .A2(n20462), .B1(n20213), .B2(n20461), .ZN(
        n20196) );
  AOI22_X1 U23195 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20463), .ZN(n20195) );
  OAI211_X1 U23196 ( .C1(n20326), .C2(n20206), .A(n20196), .B(n20195), .ZN(
        P2_U3108) );
  AOI22_X1 U23197 ( .A1(n20201), .A2(n20373), .B1(n20213), .B2(n20414), .ZN(
        n20198) );
  AOI22_X1 U23198 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20415), .ZN(n20197) );
  OAI211_X1 U23199 ( .C1(n20329), .C2(n20206), .A(n20198), .B(n20197), .ZN(
        P2_U3109) );
  AOI22_X1 U23200 ( .A1(n20201), .A2(n20376), .B1(n20420), .B2(n20213), .ZN(
        n20200) );
  AOI22_X1 U23201 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20421), .ZN(n20199) );
  OAI211_X1 U23202 ( .C1(n20332), .C2(n20206), .A(n20200), .B(n20199), .ZN(
        P2_U3110) );
  AOI22_X1 U23203 ( .A1(n20201), .A2(n20470), .B1(n20468), .B2(n20213), .ZN(
        n20205) );
  AOI22_X1 U23204 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20203), .B1(
        n20202), .B2(n20472), .ZN(n20204) );
  OAI211_X1 U23205 ( .C1(n20340), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P2_U3111) );
  NOR2_X4 U23206 ( .A1(n20269), .A2(n20246), .ZN(n20263) );
  NOR3_X1 U23207 ( .A1(n20263), .A2(n10443), .A3(n20575), .ZN(n20207) );
  NOR2_X1 U23208 ( .A1(n20207), .A2(n20270), .ZN(n20214) );
  INV_X1 U23209 ( .A(n20213), .ZN(n20208) );
  NOR2_X1 U23210 ( .A1(n20214), .A2(n20208), .ZN(n20211) );
  NAND2_X1 U23211 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20594), .ZN(
        n20273) );
  NOR2_X1 U23212 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20273), .ZN(
        n20241) );
  NAND2_X1 U23213 ( .A1(n20241), .A2(n20604), .ZN(n20212) );
  OAI21_X1 U23214 ( .B1(n20216), .B2(n20392), .A(n20212), .ZN(n20210) );
  INV_X1 U23215 ( .A(n20214), .ZN(n20209) );
  INV_X1 U23216 ( .A(n20212), .ZN(n20232) );
  AOI22_X1 U23217 ( .A1(n20436), .A2(n10443), .B1(n20433), .B2(n20232), .ZN(
        n20219) );
  NOR2_X1 U23218 ( .A1(n20214), .A2(n20213), .ZN(n20215) );
  AOI211_X1 U23219 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20216), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n20215), .ZN(n20217) );
  OAI21_X1 U23220 ( .B1(n20217), .B2(n20232), .A(n20397), .ZN(n20233) );
  AOI22_X1 U23221 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20233), .B1(
        n20263), .B2(n20435), .ZN(n20218) );
  OAI211_X1 U23222 ( .C1(n20401), .C2(n20236), .A(n20219), .B(n20218), .ZN(
        P2_U3112) );
  AOI22_X1 U23223 ( .A1(n20443), .A2(n20263), .B1(n20232), .B2(n20440), .ZN(
        n20221) );
  AOI22_X1 U23224 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20233), .B1(
        n10443), .B2(n20442), .ZN(n20220) );
  OAI211_X1 U23225 ( .C1(n20236), .C2(n20404), .A(n20221), .B(n20220), .ZN(
        P2_U3113) );
  AOI22_X1 U23226 ( .A1(n20450), .A2(n10443), .B1(n20232), .B2(n20447), .ZN(
        n20223) );
  AOI22_X1 U23227 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20233), .B1(
        n20263), .B2(n20449), .ZN(n20222) );
  OAI211_X1 U23228 ( .C1(n20236), .C2(n20407), .A(n20223), .B(n20222), .ZN(
        P2_U3114) );
  AOI22_X1 U23229 ( .A1(n20457), .A2(n20263), .B1(n20232), .B2(n20454), .ZN(
        n20225) );
  AOI22_X1 U23230 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20233), .B1(
        n10443), .B2(n20456), .ZN(n20224) );
  OAI211_X1 U23231 ( .C1(n20236), .C2(n20410), .A(n20225), .B(n20224), .ZN(
        P2_U3115) );
  AOI22_X1 U23232 ( .A1(n20464), .A2(n20263), .B1(n20232), .B2(n20461), .ZN(
        n20227) );
  AOI22_X1 U23233 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20233), .B1(
        n10443), .B2(n20463), .ZN(n20226) );
  OAI211_X1 U23234 ( .C1(n20236), .C2(n20413), .A(n20227), .B(n20226), .ZN(
        P2_U3116) );
  AOI22_X1 U23235 ( .A1(n20415), .A2(n10443), .B1(n20414), .B2(n20232), .ZN(
        n20229) );
  AOI22_X1 U23236 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20233), .B1(
        n20263), .B2(n20416), .ZN(n20228) );
  OAI211_X1 U23237 ( .C1(n20236), .C2(n20419), .A(n20229), .B(n20228), .ZN(
        P2_U3117) );
  AOI22_X1 U23238 ( .A1(n20422), .A2(n20263), .B1(n20420), .B2(n20232), .ZN(
        n20231) );
  AOI22_X1 U23239 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20233), .B1(
        n10443), .B2(n20421), .ZN(n20230) );
  OAI211_X1 U23240 ( .C1(n20236), .C2(n20425), .A(n20231), .B(n20230), .ZN(
        P2_U3118) );
  AOI22_X1 U23241 ( .A1(n20474), .A2(n20263), .B1(n20468), .B2(n20232), .ZN(
        n20235) );
  AOI22_X1 U23242 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20233), .B1(
        n10443), .B2(n20472), .ZN(n20234) );
  OAI211_X1 U23243 ( .C1(n20236), .C2(n20431), .A(n20235), .B(n20234), .ZN(
        P2_U3119) );
  AOI21_X1 U23244 ( .B1(n20306), .B2(n20587), .A(n20575), .ZN(n20243) );
  OR2_X1 U23245 ( .A1(n20237), .A2(n20273), .ZN(n20239) );
  AOI21_X1 U23246 ( .B1(n20240), .B2(n20239), .A(n20392), .ZN(n20238) );
  INV_X1 U23247 ( .A(n20239), .ZN(n20262) );
  AOI22_X1 U23248 ( .A1(n20436), .A2(n20263), .B1(n20433), .B2(n20262), .ZN(
        n20249) );
  AOI21_X1 U23249 ( .B1(n20240), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20245) );
  INV_X1 U23250 ( .A(n20241), .ZN(n20242) );
  NAND2_X1 U23251 ( .A1(n20243), .A2(n20242), .ZN(n20244) );
  OAI211_X1 U23252 ( .C1(n20262), .C2(n20245), .A(n20244), .B(n20397), .ZN(
        n20264) );
  AOI22_X1 U23253 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20435), .ZN(n20248) );
  OAI211_X1 U23254 ( .C1(n20267), .C2(n20401), .A(n20249), .B(n20248), .ZN(
        P2_U3120) );
  AOI22_X1 U23255 ( .A1(n20442), .A2(n20263), .B1(n20262), .B2(n20440), .ZN(
        n20251) );
  AOI22_X1 U23256 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20443), .ZN(n20250) );
  OAI211_X1 U23257 ( .C1(n20267), .C2(n20404), .A(n20251), .B(n20250), .ZN(
        P2_U3121) );
  AOI22_X1 U23258 ( .A1(n20450), .A2(n20263), .B1(n20262), .B2(n20447), .ZN(
        n20253) );
  AOI22_X1 U23259 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20449), .ZN(n20252) );
  OAI211_X1 U23260 ( .C1(n20267), .C2(n20407), .A(n20253), .B(n20252), .ZN(
        P2_U3122) );
  AOI22_X1 U23261 ( .A1(n20457), .A2(n20296), .B1(n20262), .B2(n20454), .ZN(
        n20255) );
  AOI22_X1 U23262 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20264), .B1(
        n20263), .B2(n20456), .ZN(n20254) );
  OAI211_X1 U23263 ( .C1(n20267), .C2(n20410), .A(n20255), .B(n20254), .ZN(
        P2_U3123) );
  AOI22_X1 U23264 ( .A1(n20464), .A2(n20296), .B1(n20262), .B2(n20461), .ZN(
        n20257) );
  AOI22_X1 U23265 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20264), .B1(
        n20263), .B2(n20463), .ZN(n20256) );
  OAI211_X1 U23266 ( .C1(n20267), .C2(n20413), .A(n20257), .B(n20256), .ZN(
        P2_U3124) );
  AOI22_X1 U23267 ( .A1(n20415), .A2(n20263), .B1(n20414), .B2(n20262), .ZN(
        n20259) );
  AOI22_X1 U23268 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20416), .ZN(n20258) );
  OAI211_X1 U23269 ( .C1(n20267), .C2(n20419), .A(n20259), .B(n20258), .ZN(
        P2_U3125) );
  AOI22_X1 U23270 ( .A1(n20421), .A2(n20263), .B1(n20420), .B2(n20262), .ZN(
        n20261) );
  AOI22_X1 U23271 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20422), .ZN(n20260) );
  OAI211_X1 U23272 ( .C1(n20267), .C2(n20425), .A(n20261), .B(n20260), .ZN(
        P2_U3126) );
  AOI22_X1 U23273 ( .A1(n20472), .A2(n20263), .B1(n20468), .B2(n20262), .ZN(
        n20266) );
  AOI22_X1 U23274 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20264), .B1(
        n20296), .B2(n20474), .ZN(n20265) );
  OAI211_X1 U23275 ( .C1(n20267), .C2(n20431), .A(n20266), .B(n20265), .ZN(
        P2_U3127) );
  INV_X1 U23276 ( .A(n20296), .ZN(n20268) );
  NAND2_X1 U23277 ( .A1(n20268), .A2(n20382), .ZN(n20271) );
  INV_X1 U23278 ( .A(n20270), .ZN(n20385) );
  OAI21_X1 U23279 ( .B1(n20271), .B2(n20335), .A(n20385), .ZN(n20276) );
  INV_X1 U23280 ( .A(n20273), .ZN(n20301) );
  AND2_X1 U23281 ( .A1(n20272), .A2(n20301), .ZN(n20279) );
  NOR2_X1 U23282 ( .A1(n20274), .A2(n20273), .ZN(n20295) );
  INV_X1 U23283 ( .A(n20295), .ZN(n20277) );
  AOI22_X1 U23284 ( .A1(n20435), .A2(n20335), .B1(n20433), .B2(n20295), .ZN(
        n20282) );
  INV_X1 U23285 ( .A(n20276), .ZN(n20280) );
  OAI211_X1 U23286 ( .C1(n20280), .C2(n20279), .A(n20397), .B(n20278), .ZN(
        n20297) );
  AOI22_X1 U23287 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20297), .B1(
        n20296), .B2(n20436), .ZN(n20281) );
  OAI211_X1 U23288 ( .C1(n20300), .C2(n20401), .A(n20282), .B(n20281), .ZN(
        P2_U3128) );
  AOI22_X1 U23289 ( .A1(n20442), .A2(n20296), .B1(n20440), .B2(n20295), .ZN(
        n20284) );
  AOI22_X1 U23290 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20297), .B1(
        n20335), .B2(n20443), .ZN(n20283) );
  OAI211_X1 U23291 ( .C1(n20300), .C2(n20404), .A(n20284), .B(n20283), .ZN(
        P2_U3129) );
  AOI22_X1 U23292 ( .A1(n20450), .A2(n20296), .B1(n20447), .B2(n20295), .ZN(
        n20286) );
  AOI22_X1 U23293 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20297), .B1(
        n20335), .B2(n20449), .ZN(n20285) );
  OAI211_X1 U23294 ( .C1(n20300), .C2(n20407), .A(n20286), .B(n20285), .ZN(
        P2_U3130) );
  AOI22_X1 U23295 ( .A1(n20456), .A2(n20296), .B1(n9749), .B2(n20295), .ZN(
        n20288) );
  AOI22_X1 U23296 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20297), .B1(
        n20335), .B2(n20457), .ZN(n20287) );
  OAI211_X1 U23297 ( .C1(n20300), .C2(n20410), .A(n20288), .B(n20287), .ZN(
        P2_U3131) );
  AOI22_X1 U23298 ( .A1(n20464), .A2(n20335), .B1(n20461), .B2(n20295), .ZN(
        n20290) );
  AOI22_X1 U23299 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20297), .B1(
        n20296), .B2(n20463), .ZN(n20289) );
  OAI211_X1 U23300 ( .C1(n20300), .C2(n20413), .A(n20290), .B(n20289), .ZN(
        P2_U3132) );
  AOI22_X1 U23301 ( .A1(n20416), .A2(n20335), .B1(n20414), .B2(n20295), .ZN(
        n20292) );
  AOI22_X1 U23302 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20297), .B1(
        n20296), .B2(n20415), .ZN(n20291) );
  OAI211_X1 U23303 ( .C1(n20300), .C2(n20419), .A(n20292), .B(n20291), .ZN(
        P2_U3133) );
  AOI22_X1 U23304 ( .A1(n20421), .A2(n20296), .B1(n20420), .B2(n20295), .ZN(
        n20294) );
  AOI22_X1 U23305 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20297), .B1(
        n20335), .B2(n20422), .ZN(n20293) );
  OAI211_X1 U23306 ( .C1(n20300), .C2(n20425), .A(n20294), .B(n20293), .ZN(
        P2_U3134) );
  AOI22_X1 U23307 ( .A1(n20472), .A2(n20296), .B1(n20468), .B2(n20295), .ZN(
        n20299) );
  AOI22_X1 U23308 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20297), .B1(
        n20335), .B2(n20474), .ZN(n20298) );
  OAI211_X1 U23309 ( .C1(n20300), .C2(n20431), .A(n20299), .B(n20298), .ZN(
        P2_U3135) );
  NAND2_X1 U23310 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20301), .ZN(
        n20307) );
  INV_X1 U23311 ( .A(n20305), .ZN(n20303) );
  AND2_X1 U23312 ( .A1(n20302), .A2(n20301), .ZN(n20333) );
  OAI21_X1 U23313 ( .B1(n20303), .B2(n20333), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20304) );
  AOI22_X1 U23314 ( .A1(n20334), .A2(n20434), .B1(n20433), .B2(n20333), .ZN(
        n20313) );
  AOI21_X1 U23315 ( .B1(n20305), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20311) );
  INV_X1 U23316 ( .A(n20306), .ZN(n20309) );
  OAI21_X1 U23317 ( .B1(n20309), .B2(n20308), .A(n20307), .ZN(n20310) );
  OAI211_X1 U23318 ( .C1(n20333), .C2(n20311), .A(n20310), .B(n20397), .ZN(
        n20336) );
  AOI22_X1 U23319 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20436), .ZN(n20312) );
  OAI211_X1 U23320 ( .C1(n20314), .C2(n20339), .A(n20313), .B(n20312), .ZN(
        P2_U3136) );
  AOI22_X1 U23321 ( .A1(n20334), .A2(n20441), .B1(n20440), .B2(n20333), .ZN(
        n20316) );
  AOI22_X1 U23322 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20442), .ZN(n20315) );
  OAI211_X1 U23323 ( .C1(n20317), .C2(n20339), .A(n20316), .B(n20315), .ZN(
        P2_U3137) );
  AOI22_X1 U23324 ( .A1(n20334), .A2(n20448), .B1(n20447), .B2(n20333), .ZN(
        n20319) );
  AOI22_X1 U23325 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20450), .ZN(n20318) );
  OAI211_X1 U23326 ( .C1(n20320), .C2(n20339), .A(n20319), .B(n20318), .ZN(
        P2_U3138) );
  AOI22_X1 U23327 ( .A1(n20334), .A2(n20455), .B1(n9749), .B2(n20333), .ZN(
        n20322) );
  AOI22_X1 U23328 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20456), .ZN(n20321) );
  OAI211_X1 U23329 ( .C1(n20323), .C2(n20339), .A(n20322), .B(n20321), .ZN(
        P2_U3139) );
  AOI22_X1 U23330 ( .A1(n20334), .A2(n20462), .B1(n20461), .B2(n20333), .ZN(
        n20325) );
  AOI22_X1 U23331 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20463), .ZN(n20324) );
  OAI211_X1 U23332 ( .C1(n20326), .C2(n20339), .A(n20325), .B(n20324), .ZN(
        P2_U3140) );
  AOI22_X1 U23333 ( .A1(n20334), .A2(n20373), .B1(n20414), .B2(n20333), .ZN(
        n20328) );
  AOI22_X1 U23334 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20415), .ZN(n20327) );
  OAI211_X1 U23335 ( .C1(n20329), .C2(n20339), .A(n20328), .B(n20327), .ZN(
        P2_U3141) );
  AOI22_X1 U23336 ( .A1(n20334), .A2(n20376), .B1(n20420), .B2(n20333), .ZN(
        n20331) );
  AOI22_X1 U23337 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20421), .ZN(n20330) );
  OAI211_X1 U23338 ( .C1(n20332), .C2(n20339), .A(n20331), .B(n20330), .ZN(
        P2_U3142) );
  AOI22_X1 U23339 ( .A1(n20334), .A2(n20470), .B1(n20468), .B2(n20333), .ZN(
        n20338) );
  AOI22_X1 U23340 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20336), .B1(
        n20335), .B2(n20472), .ZN(n20337) );
  OAI211_X1 U23341 ( .C1(n20340), .C2(n20339), .A(n20338), .B(n20337), .ZN(
        P2_U3143) );
  INV_X1 U23342 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n20343) );
  AOI22_X1 U23343 ( .A1(n20357), .A2(n20434), .B1(n20433), .B2(n20356), .ZN(
        n20342) );
  AOI22_X1 U23344 ( .A1(n20358), .A2(n20436), .B1(n20378), .B2(n20435), .ZN(
        n20341) );
  OAI211_X1 U23345 ( .C1(n20362), .C2(n20343), .A(n20342), .B(n20341), .ZN(
        P2_U3144) );
  AOI22_X1 U23346 ( .A1(n20357), .A2(n20441), .B1(n20356), .B2(n20440), .ZN(
        n20345) );
  AOI22_X1 U23347 ( .A1(n20378), .A2(n20443), .B1(n20358), .B2(n20442), .ZN(
        n20344) );
  OAI211_X1 U23348 ( .C1(n20362), .C2(n12455), .A(n20345), .B(n20344), .ZN(
        P2_U3145) );
  INV_X1 U23349 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20348) );
  AOI22_X1 U23350 ( .A1(n20357), .A2(n20448), .B1(n20356), .B2(n20447), .ZN(
        n20347) );
  AOI22_X1 U23351 ( .A1(n20358), .A2(n20450), .B1(n20378), .B2(n20449), .ZN(
        n20346) );
  OAI211_X1 U23352 ( .C1(n20362), .C2(n20348), .A(n20347), .B(n20346), .ZN(
        P2_U3146) );
  AOI22_X1 U23353 ( .A1(n20357), .A2(n20455), .B1(n20356), .B2(n20454), .ZN(
        n20350) );
  AOI22_X1 U23354 ( .A1(n20378), .A2(n20457), .B1(n20358), .B2(n20456), .ZN(
        n20349) );
  OAI211_X1 U23355 ( .C1(n20362), .C2(n12405), .A(n20350), .B(n20349), .ZN(
        P2_U3147) );
  INV_X1 U23356 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20353) );
  AOI22_X1 U23357 ( .A1(n20357), .A2(n20462), .B1(n20356), .B2(n20461), .ZN(
        n20352) );
  AOI22_X1 U23358 ( .A1(n20378), .A2(n20464), .B1(n20358), .B2(n20463), .ZN(
        n20351) );
  OAI211_X1 U23359 ( .C1(n20362), .C2(n20353), .A(n20352), .B(n20351), .ZN(
        P2_U3148) );
  AOI22_X1 U23360 ( .A1(n20357), .A2(n20373), .B1(n20356), .B2(n20414), .ZN(
        n20355) );
  AOI22_X1 U23361 ( .A1(n20358), .A2(n20415), .B1(n20378), .B2(n20416), .ZN(
        n20354) );
  OAI211_X1 U23362 ( .C1(n20362), .C2(n12474), .A(n20355), .B(n20354), .ZN(
        P2_U3149) );
  INV_X1 U23363 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n20361) );
  AOI22_X1 U23364 ( .A1(n20357), .A2(n20470), .B1(n20468), .B2(n20356), .ZN(
        n20360) );
  AOI22_X1 U23365 ( .A1(n20378), .A2(n20474), .B1(n20358), .B2(n20472), .ZN(
        n20359) );
  OAI211_X1 U23366 ( .C1(n20362), .C2(n20361), .A(n20360), .B(n20359), .ZN(
        P2_U3151) );
  AOI22_X1 U23367 ( .A1(n20377), .A2(n20441), .B1(n20387), .B2(n20440), .ZN(
        n20364) );
  AOI22_X1 U23368 ( .A1(n20427), .A2(n20443), .B1(n20378), .B2(n20442), .ZN(
        n20363) );
  OAI211_X1 U23369 ( .C1(n20381), .C2(n12441), .A(n20364), .B(n20363), .ZN(
        P2_U3153) );
  INV_X1 U23370 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20367) );
  AOI22_X1 U23371 ( .A1(n20377), .A2(n20448), .B1(n20387), .B2(n20447), .ZN(
        n20366) );
  AOI22_X1 U23372 ( .A1(n20378), .A2(n20450), .B1(n20427), .B2(n20449), .ZN(
        n20365) );
  OAI211_X1 U23373 ( .C1(n20381), .C2(n20367), .A(n20366), .B(n20365), .ZN(
        P2_U3154) );
  AOI22_X1 U23374 ( .A1(n20377), .A2(n20455), .B1(n20387), .B2(n20454), .ZN(
        n20369) );
  AOI22_X1 U23375 ( .A1(n20427), .A2(n20457), .B1(n20378), .B2(n20456), .ZN(
        n20368) );
  OAI211_X1 U23376 ( .C1(n20381), .C2(n12398), .A(n20369), .B(n20368), .ZN(
        P2_U3155) );
  AOI22_X1 U23377 ( .A1(n20377), .A2(n20462), .B1(n20387), .B2(n20461), .ZN(
        n20371) );
  AOI22_X1 U23378 ( .A1(n20427), .A2(n20464), .B1(n20378), .B2(n20463), .ZN(
        n20370) );
  OAI211_X1 U23379 ( .C1(n20381), .C2(n20372), .A(n20371), .B(n20370), .ZN(
        P2_U3156) );
  AOI22_X1 U23380 ( .A1(n20377), .A2(n20373), .B1(n20387), .B2(n20414), .ZN(
        n20375) );
  AOI22_X1 U23381 ( .A1(n20378), .A2(n20415), .B1(n20427), .B2(n20416), .ZN(
        n20374) );
  OAI211_X1 U23382 ( .C1(n20381), .C2(n12470), .A(n20375), .B(n20374), .ZN(
        P2_U3157) );
  AOI22_X1 U23383 ( .A1(n20377), .A2(n20376), .B1(n20420), .B2(n20387), .ZN(
        n20380) );
  AOI22_X1 U23384 ( .A1(n20427), .A2(n20422), .B1(n20378), .B2(n20421), .ZN(
        n20379) );
  OAI211_X1 U23385 ( .C1(n20381), .C2(n12510), .A(n20380), .B(n20379), .ZN(
        P2_U3158) );
  NAND3_X1 U23386 ( .A1(n20384), .A2(n20383), .A3(n20382), .ZN(n20386) );
  INV_X1 U23387 ( .A(n20387), .ZN(n20395) );
  AOI22_X1 U23388 ( .A1(n20390), .A2(n20388), .B1(n20392), .B2(n20395), .ZN(
        n20391) );
  AND2_X1 U23389 ( .A1(n20389), .A2(n20604), .ZN(n20426) );
  AOI22_X1 U23390 ( .A1(n20435), .A2(n20473), .B1(n20433), .B2(n20426), .ZN(
        n20400) );
  OAI21_X1 U23391 ( .B1(n20393), .B2(n20392), .A(n20581), .ZN(n20394) );
  AOI21_X1 U23392 ( .B1(n20396), .B2(n20395), .A(n20394), .ZN(n20398) );
  OAI21_X1 U23393 ( .B1(n20398), .B2(n20426), .A(n20397), .ZN(n20428) );
  AOI22_X1 U23394 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20436), .ZN(n20399) );
  OAI211_X1 U23395 ( .C1(n20432), .C2(n20401), .A(n20400), .B(n20399), .ZN(
        P2_U3160) );
  AOI22_X1 U23396 ( .A1(n20442), .A2(n20427), .B1(n20426), .B2(n20440), .ZN(
        n20403) );
  AOI22_X1 U23397 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20428), .B1(
        n20473), .B2(n20443), .ZN(n20402) );
  OAI211_X1 U23398 ( .C1(n20432), .C2(n20404), .A(n20403), .B(n20402), .ZN(
        P2_U3161) );
  AOI22_X1 U23399 ( .A1(n20449), .A2(n20473), .B1(n20426), .B2(n20447), .ZN(
        n20406) );
  AOI22_X1 U23400 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20450), .ZN(n20405) );
  OAI211_X1 U23401 ( .C1(n20432), .C2(n20407), .A(n20406), .B(n20405), .ZN(
        P2_U3162) );
  AOI22_X1 U23402 ( .A1(n20457), .A2(n20473), .B1(n20426), .B2(n20454), .ZN(
        n20409) );
  AOI22_X1 U23403 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20456), .ZN(n20408) );
  OAI211_X1 U23404 ( .C1(n20432), .C2(n20410), .A(n20409), .B(n20408), .ZN(
        P2_U3163) );
  AOI22_X1 U23405 ( .A1(n20464), .A2(n20473), .B1(n20426), .B2(n20461), .ZN(
        n20412) );
  AOI22_X1 U23406 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20463), .ZN(n20411) );
  OAI211_X1 U23407 ( .C1(n20432), .C2(n20413), .A(n20412), .B(n20411), .ZN(
        P2_U3164) );
  AOI22_X1 U23408 ( .A1(n20415), .A2(n20427), .B1(n20426), .B2(n20414), .ZN(
        n20418) );
  AOI22_X1 U23409 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20428), .B1(
        n20473), .B2(n20416), .ZN(n20417) );
  OAI211_X1 U23410 ( .C1(n20432), .C2(n20419), .A(n20418), .B(n20417), .ZN(
        P2_U3165) );
  AOI22_X1 U23411 ( .A1(n20421), .A2(n20427), .B1(n20420), .B2(n20426), .ZN(
        n20424) );
  AOI22_X1 U23412 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20428), .B1(
        n20473), .B2(n20422), .ZN(n20423) );
  OAI211_X1 U23413 ( .C1(n20432), .C2(n20425), .A(n20424), .B(n20423), .ZN(
        P2_U3166) );
  AOI22_X1 U23414 ( .A1(n20474), .A2(n20473), .B1(n20468), .B2(n20426), .ZN(
        n20430) );
  AOI22_X1 U23415 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20428), .B1(
        n20427), .B2(n20472), .ZN(n20429) );
  OAI211_X1 U23416 ( .C1(n20432), .C2(n20431), .A(n20430), .B(n20429), .ZN(
        P2_U3167) );
  INV_X1 U23417 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n20439) );
  AOI22_X1 U23418 ( .A1(n20471), .A2(n20434), .B1(n20469), .B2(n20433), .ZN(
        n20438) );
  AOI22_X1 U23419 ( .A1(n20473), .A2(n20436), .B1(n20475), .B2(n20435), .ZN(
        n20437) );
  OAI211_X1 U23420 ( .C1(n20479), .C2(n20439), .A(n20438), .B(n20437), .ZN(
        P2_U3168) );
  AOI22_X1 U23421 ( .A1(n20471), .A2(n20441), .B1(n20469), .B2(n20440), .ZN(
        n20445) );
  AOI22_X1 U23422 ( .A1(n20475), .A2(n20443), .B1(n20473), .B2(n20442), .ZN(
        n20444) );
  OAI211_X1 U23423 ( .C1(n20479), .C2(n20446), .A(n20445), .B(n20444), .ZN(
        P2_U3169) );
  AOI22_X1 U23424 ( .A1(n20471), .A2(n20448), .B1(n20469), .B2(n20447), .ZN(
        n20452) );
  AOI22_X1 U23425 ( .A1(n20473), .A2(n20450), .B1(n20475), .B2(n20449), .ZN(
        n20451) );
  OAI211_X1 U23426 ( .C1(n20479), .C2(n20453), .A(n20452), .B(n20451), .ZN(
        P2_U3170) );
  INV_X1 U23427 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20460) );
  AOI22_X1 U23428 ( .A1(n20471), .A2(n20455), .B1(n20469), .B2(n20454), .ZN(
        n20459) );
  AOI22_X1 U23429 ( .A1(n20475), .A2(n20457), .B1(n20473), .B2(n20456), .ZN(
        n20458) );
  OAI211_X1 U23430 ( .C1(n20479), .C2(n20460), .A(n20459), .B(n20458), .ZN(
        P2_U3171) );
  INV_X1 U23431 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n20467) );
  AOI22_X1 U23432 ( .A1(n20471), .A2(n20462), .B1(n20469), .B2(n20461), .ZN(
        n20466) );
  AOI22_X1 U23433 ( .A1(n20475), .A2(n20464), .B1(n20473), .B2(n20463), .ZN(
        n20465) );
  OAI211_X1 U23434 ( .C1(n20479), .C2(n20467), .A(n20466), .B(n20465), .ZN(
        P2_U3172) );
  INV_X1 U23435 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20478) );
  AOI22_X1 U23436 ( .A1(n20471), .A2(n20470), .B1(n20469), .B2(n20468), .ZN(
        n20477) );
  AOI22_X1 U23437 ( .A1(n20475), .A2(n20474), .B1(n20473), .B2(n20472), .ZN(
        n20476) );
  OAI211_X1 U23438 ( .C1(n20479), .C2(n20478), .A(n20477), .B(n20476), .ZN(
        P2_U3175) );
  OAI21_X1 U23439 ( .B1(n10291), .B2(n20482), .A(n20481), .ZN(n20486) );
  NAND2_X1 U23440 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n10291), .ZN(n20483) );
  AOI21_X1 U23441 ( .B1(n20487), .B2(n20484), .A(n20483), .ZN(n20485) );
  AOI21_X1 U23442 ( .B1(n20487), .B2(n20486), .A(n20485), .ZN(n20489) );
  NAND2_X1 U23443 ( .A1(n20489), .A2(n20488), .ZN(P2_U3177) );
  AND2_X1 U23444 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20570), .ZN(
        P2_U3179) );
  NOR2_X1 U23445 ( .A1(n21580), .A2(n20573), .ZN(P2_U3180) );
  AND2_X1 U23446 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20570), .ZN(
        P2_U3181) );
  AND2_X1 U23447 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20570), .ZN(
        P2_U3182) );
  AND2_X1 U23448 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20570), .ZN(
        P2_U3183) );
  AND2_X1 U23449 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20570), .ZN(
        P2_U3184) );
  AND2_X1 U23450 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20570), .ZN(
        P2_U3185) );
  AND2_X1 U23451 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20570), .ZN(
        P2_U3186) );
  AND2_X1 U23452 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20570), .ZN(
        P2_U3187) );
  AND2_X1 U23453 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20570), .ZN(
        P2_U3188) );
  AND2_X1 U23454 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20570), .ZN(
        P2_U3189) );
  AND2_X1 U23455 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20570), .ZN(
        P2_U3190) );
  AND2_X1 U23456 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20570), .ZN(
        P2_U3191) );
  AND2_X1 U23457 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20570), .ZN(
        P2_U3192) );
  AND2_X1 U23458 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20570), .ZN(
        P2_U3193) );
  INV_X1 U23459 ( .A(P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21617) );
  NOR2_X1 U23460 ( .A1(n21617), .A2(n20573), .ZN(P2_U3194) );
  AND2_X1 U23461 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20570), .ZN(
        P2_U3195) );
  NOR2_X1 U23462 ( .A1(n21534), .A2(n20573), .ZN(P2_U3196) );
  AND2_X1 U23463 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20570), .ZN(
        P2_U3197) );
  AND2_X1 U23464 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20570), .ZN(
        P2_U3198) );
  AND2_X1 U23465 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20570), .ZN(
        P2_U3199) );
  AND2_X1 U23466 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20570), .ZN(
        P2_U3200) );
  AND2_X1 U23467 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20570), .ZN(P2_U3201) );
  AND2_X1 U23468 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20570), .ZN(P2_U3202) );
  AND2_X1 U23469 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20570), .ZN(P2_U3203) );
  AND2_X1 U23470 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20570), .ZN(P2_U3204) );
  AND2_X1 U23471 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20570), .ZN(P2_U3205) );
  AND2_X1 U23472 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20570), .ZN(P2_U3206) );
  INV_X1 U23473 ( .A(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n21540) );
  NOR2_X1 U23474 ( .A1(n21540), .A2(n20573), .ZN(P2_U3207) );
  AND2_X1 U23475 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20570), .ZN(P2_U3208) );
  AOI21_X1 U23476 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n21423), .A(n20490), .ZN(n20492) );
  INV_X1 U23477 ( .A(NA), .ZN(n21416) );
  OAI21_X1 U23478 ( .B1(n21416), .B2(n20497), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20506) );
  NAND2_X1 U23479 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n10291), .ZN(n20504) );
  NAND3_X1 U23480 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n20504), .ZN(n20491) );
  AOI22_X1 U23481 ( .A1(n20492), .A2(n20619), .B1(n20506), .B2(n20491), .ZN(
        n20493) );
  INV_X1 U23482 ( .A(n20493), .ZN(P2_U3209) );
  INV_X1 U23483 ( .A(n20504), .ZN(n20494) );
  NOR2_X1 U23484 ( .A1(n20495), .A2(n20494), .ZN(n20499) );
  NOR2_X1 U23485 ( .A1(HOLD), .A2(n20496), .ZN(n20505) );
  OAI211_X1 U23486 ( .C1(n20505), .C2(n20507), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n20497), .ZN(n20498) );
  OAI211_X1 U23487 ( .C1(n20500), .C2(n21423), .A(n20499), .B(n20498), .ZN(
        P2_U3210) );
  OAI22_X1 U23488 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20501), .B1(NA), 
        .B2(n20504), .ZN(n20502) );
  OAI211_X1 U23489 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20502), .ZN(n20503) );
  OAI221_X1 U23490 ( .B1(n20506), .B2(n20505), .C1(n20506), .C2(n20504), .A(
        n20503), .ZN(P2_U3211) );
  OAI222_X1 U23491 ( .A1(n20558), .A2(n20509), .B1(n20508), .B2(n20618), .C1(
        n20511), .C2(n20562), .ZN(P2_U3212) );
  OAI222_X1 U23492 ( .A1(n20558), .A2(n20511), .B1(n20510), .B2(n20618), .C1(
        n20513), .C2(n20562), .ZN(P2_U3213) );
  OAI222_X1 U23493 ( .A1(n20558), .A2(n20513), .B1(n20512), .B2(n20618), .C1(
        n19915), .C2(n20562), .ZN(P2_U3214) );
  OAI222_X1 U23494 ( .A1(n20562), .A2(n19759), .B1(n20514), .B2(n20618), .C1(
        n19915), .C2(n20558), .ZN(P2_U3215) );
  OAI222_X1 U23495 ( .A1(n20562), .A2(n20516), .B1(n20515), .B2(n20618), .C1(
        n19759), .C2(n20558), .ZN(P2_U3216) );
  OAI222_X1 U23496 ( .A1(n20562), .A2(n20518), .B1(n20517), .B2(n20618), .C1(
        n20516), .C2(n20558), .ZN(P2_U3217) );
  OAI222_X1 U23497 ( .A1(n20562), .A2(n20520), .B1(n20519), .B2(n20618), .C1(
        n20518), .C2(n20558), .ZN(P2_U3218) );
  OAI222_X1 U23498 ( .A1(n20562), .A2(n16306), .B1(n20521), .B2(n20618), .C1(
        n20520), .C2(n20558), .ZN(P2_U3219) );
  OAI222_X1 U23499 ( .A1(n20562), .A2(n20523), .B1(n20522), .B2(n20618), .C1(
        n16306), .C2(n20558), .ZN(P2_U3220) );
  OAI222_X1 U23500 ( .A1(n20562), .A2(n19703), .B1(n20524), .B2(n20618), .C1(
        n20523), .C2(n20558), .ZN(P2_U3221) );
  OAI222_X1 U23501 ( .A1(n20562), .A2(n20526), .B1(n20525), .B2(n20618), .C1(
        n19703), .C2(n20558), .ZN(P2_U3222) );
  OAI222_X1 U23502 ( .A1(n20562), .A2(n15767), .B1(n20527), .B2(n20618), .C1(
        n20526), .C2(n20558), .ZN(P2_U3223) );
  OAI222_X1 U23503 ( .A1(n20562), .A2(n20529), .B1(n20528), .B2(n20618), .C1(
        n15767), .C2(n20558), .ZN(P2_U3224) );
  OAI222_X1 U23504 ( .A1(n20562), .A2(n20531), .B1(n20530), .B2(n20618), .C1(
        n20529), .C2(n20558), .ZN(P2_U3225) );
  OAI222_X1 U23505 ( .A1(n20562), .A2(n20533), .B1(n20532), .B2(n20618), .C1(
        n20531), .C2(n20558), .ZN(P2_U3226) );
  OAI222_X1 U23506 ( .A1(n20562), .A2(n20535), .B1(n20534), .B2(n20618), .C1(
        n20533), .C2(n20558), .ZN(P2_U3227) );
  OAI222_X1 U23507 ( .A1(n20562), .A2(n19630), .B1(n20536), .B2(n20618), .C1(
        n20535), .C2(n20558), .ZN(P2_U3228) );
  OAI222_X1 U23508 ( .A1(n20562), .A2(n20538), .B1(n20537), .B2(n20618), .C1(
        n19630), .C2(n20558), .ZN(P2_U3229) );
  OAI222_X1 U23509 ( .A1(n20562), .A2(n20540), .B1(n20539), .B2(n20618), .C1(
        n20538), .C2(n20558), .ZN(P2_U3230) );
  OAI222_X1 U23510 ( .A1(n20562), .A2(n20542), .B1(n20541), .B2(n20618), .C1(
        n20540), .C2(n20558), .ZN(P2_U3231) );
  OAI222_X1 U23511 ( .A1(n20562), .A2(n20544), .B1(n20543), .B2(n20618), .C1(
        n20542), .C2(n20558), .ZN(P2_U3232) );
  OAI222_X1 U23512 ( .A1(n20562), .A2(n20546), .B1(n20545), .B2(n20618), .C1(
        n20544), .C2(n20558), .ZN(P2_U3233) );
  OAI222_X1 U23513 ( .A1(n20562), .A2(n20548), .B1(n20547), .B2(n20618), .C1(
        n20546), .C2(n20558), .ZN(P2_U3234) );
  OAI222_X1 U23514 ( .A1(n20562), .A2(n20550), .B1(n20549), .B2(n20618), .C1(
        n20548), .C2(n20558), .ZN(P2_U3235) );
  OAI222_X1 U23515 ( .A1(n20562), .A2(n16142), .B1(n20551), .B2(n20618), .C1(
        n20550), .C2(n20558), .ZN(P2_U3236) );
  OAI222_X1 U23516 ( .A1(n20562), .A2(n20554), .B1(n20552), .B2(n20618), .C1(
        n16142), .C2(n20558), .ZN(P2_U3237) );
  OAI222_X1 U23517 ( .A1(n20558), .A2(n20554), .B1(n20553), .B2(n20618), .C1(
        n16117), .C2(n20562), .ZN(P2_U3238) );
  OAI222_X1 U23518 ( .A1(n20562), .A2(n20556), .B1(n20555), .B2(n20618), .C1(
        n16117), .C2(n20558), .ZN(P2_U3239) );
  OAI222_X1 U23519 ( .A1(n20562), .A2(n20559), .B1(n20557), .B2(n20618), .C1(
        n20556), .C2(n20558), .ZN(P2_U3240) );
  OAI222_X1 U23520 ( .A1(n20562), .A2(n20561), .B1(n20560), .B2(n20618), .C1(
        n20559), .C2(n20558), .ZN(P2_U3241) );
  INV_X1 U23521 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n20563) );
  AOI22_X1 U23522 ( .A1(n20618), .A2(n20564), .B1(n20563), .B2(n20619), .ZN(
        P2_U3585) );
  MUX2_X1 U23523 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n20618), .Z(P2_U3586) );
  INV_X1 U23524 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n20565) );
  AOI22_X1 U23525 ( .A1(n20618), .A2(n20566), .B1(n20565), .B2(n20619), .ZN(
        P2_U3587) );
  INV_X1 U23526 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U23527 ( .A1(n20618), .A2(n20568), .B1(n20567), .B2(n20619), .ZN(
        P2_U3588) );
  INV_X1 U23528 ( .A(n20571), .ZN(n20569) );
  AOI21_X1 U23529 ( .B1(n20570), .B2(n21542), .A(n20569), .ZN(P2_U3591) );
  OAI21_X1 U23530 ( .B1(n20573), .B2(n20572), .A(n20571), .ZN(P2_U3592) );
  NOR3_X1 U23531 ( .A1(n20576), .A2(n20575), .A3(n20574), .ZN(n20584) );
  NAND2_X1 U23532 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20577), .ZN(n20578) );
  OAI21_X1 U23533 ( .B1(n20579), .B2(n20578), .A(n20600), .ZN(n20588) );
  OAI22_X1 U23534 ( .A1(n20582), .A2(n20588), .B1(n20581), .B2(n20580), .ZN(
        n20583) );
  NOR2_X1 U23535 ( .A1(n20584), .A2(n20583), .ZN(n20585) );
  AOI22_X1 U23536 ( .A1(n20605), .A2(n20586), .B1(n20585), .B2(n20602), .ZN(
        P2_U3602) );
  AOI211_X1 U23537 ( .C1(n20590), .C2(n20589), .A(n20588), .B(n20587), .ZN(
        n20591) );
  AOI21_X1 U23538 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20592), .A(n20591), 
        .ZN(n20593) );
  AOI22_X1 U23539 ( .A1(n20605), .A2(n20594), .B1(n20593), .B2(n20602), .ZN(
        P2_U3603) );
  INV_X1 U23540 ( .A(n20595), .ZN(n20598) );
  OAI21_X1 U23541 ( .B1(n20598), .B2(n20597), .A(n20596), .ZN(n20599) );
  AOI21_X1 U23542 ( .B1(n20601), .B2(n20600), .A(n20599), .ZN(n20603) );
  AOI22_X1 U23543 ( .A1(n20605), .A2(n20604), .B1(n20603), .B2(n20602), .ZN(
        P2_U3605) );
  INV_X1 U23544 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20606) );
  AOI22_X1 U23545 ( .A1(n20618), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20606), 
        .B2(n20619), .ZN(P2_U3608) );
  INV_X1 U23546 ( .A(n20607), .ZN(n20613) );
  INV_X1 U23547 ( .A(n20608), .ZN(n20611) );
  OAI21_X1 U23548 ( .B1(n20611), .B2(n20610), .A(n20609), .ZN(n20612) );
  OAI211_X1 U23549 ( .C1(n20615), .C2(n20614), .A(n20613), .B(n20612), .ZN(
        n20617) );
  MUX2_X1 U23550 ( .A(P2_MORE_REG_SCAN_IN), .B(n20617), .S(n20616), .Z(
        P2_U3609) );
  OAI22_X1 U23551 ( .A1(n20619), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20618), .ZN(n20620) );
  INV_X1 U23552 ( .A(n20620), .ZN(P2_U3611) );
  NOR2_X1 U23553 ( .A1(n21418), .A2(n21415), .ZN(n20623) );
  INV_X1 U23554 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20622) );
  NOR2_X4 U23555 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20621), .ZN(n21511) );
  AOI21_X1 U23556 ( .B1(n20623), .B2(n20622), .A(n21511), .ZN(P1_U2802) );
  NAND2_X1 U23557 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20624), .ZN(n20629) );
  INV_X1 U23558 ( .A(n20625), .ZN(n20627) );
  OAI21_X1 U23559 ( .B1(n20627), .B2(n20626), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20628) );
  OAI21_X1 U23560 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20629), .A(n20628), 
        .ZN(P1_U2803) );
  INV_X2 U23561 ( .A(n21511), .ZN(n21495) );
  NOR2_X1 U23562 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21408) );
  OAI21_X1 U23563 ( .B1(n21408), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21495), .ZN(
        n20630) );
  OAI21_X1 U23564 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21495), .A(n20630), 
        .ZN(P1_U2804) );
  OAI21_X1 U23565 ( .B1(BS16), .B2(n21408), .A(n21486), .ZN(n21484) );
  OAI21_X1 U23566 ( .B1(n21486), .B2(n21497), .A(n21484), .ZN(P1_U2805) );
  OAI21_X1 U23567 ( .B1(n20632), .B2(n21646), .A(n20631), .ZN(P1_U2806) );
  NOR4_X1 U23568 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20636) );
  NOR4_X1 U23569 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20635) );
  NOR4_X1 U23570 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20634) );
  NOR4_X1 U23571 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20633) );
  NAND4_X1 U23572 ( .A1(n20636), .A2(n20635), .A3(n20634), .A4(n20633), .ZN(
        n20642) );
  NOR4_X1 U23573 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n20640) );
  AOI211_X1 U23574 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20639) );
  NOR4_X1 U23575 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20638) );
  NOR4_X1 U23576 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20637) );
  NAND4_X1 U23577 ( .A1(n20640), .A2(n20639), .A3(n20638), .A4(n20637), .ZN(
        n20641) );
  NOR2_X1 U23578 ( .A1(n20642), .A2(n20641), .ZN(n21494) );
  INV_X1 U23579 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21479) );
  NOR3_X1 U23580 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20644) );
  OAI21_X1 U23581 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20644), .A(n21494), .ZN(
        n20643) );
  OAI21_X1 U23582 ( .B1(n21494), .B2(n21479), .A(n20643), .ZN(P1_U2807) );
  INV_X1 U23583 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21487) );
  INV_X1 U23584 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21485) );
  AOI21_X1 U23585 ( .B1(n21487), .B2(n21485), .A(n20644), .ZN(n20645) );
  INV_X1 U23586 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21649) );
  INV_X1 U23587 ( .A(n21494), .ZN(n21489) );
  AOI22_X1 U23588 ( .A1(n21494), .A2(n20645), .B1(n21649), .B2(n21489), .ZN(
        P1_U2808) );
  OAI21_X1 U23589 ( .B1(n20646), .B2(n21565), .A(n20688), .ZN(n20647) );
  AOI21_X1 U23590 ( .B1(n20685), .B2(P1_EBX_REG_9__SCAN_IN), .A(n20647), .ZN(
        n20648) );
  OAI21_X1 U23591 ( .B1(n20650), .B2(n20649), .A(n20648), .ZN(n20651) );
  AOI221_X1 U23592 ( .B1(n20653), .B2(P1_REIP_REG_9__SCAN_IN), .C1(n20652), 
        .C2(n21439), .A(n20651), .ZN(n20659) );
  INV_X1 U23593 ( .A(n20654), .ZN(n20657) );
  INV_X1 U23594 ( .A(n20655), .ZN(n20656) );
  AOI22_X1 U23595 ( .A1(n20657), .A2(n13732), .B1(n20656), .B2(n20709), .ZN(
        n20658) );
  NAND2_X1 U23596 ( .A1(n20659), .A2(n20658), .ZN(P1_U2831) );
  AOI21_X1 U23597 ( .B1(n20672), .B2(n20671), .A(n20660), .ZN(n20676) );
  NOR3_X1 U23598 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20687), .A3(n20671), .ZN(
        n20661) );
  AOI211_X1 U23599 ( .C1(n20698), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n20662), .B(n20661), .ZN(n20665) );
  AOI22_X1 U23600 ( .A1(n20705), .A2(n20663), .B1(n20685), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n20664) );
  OAI211_X1 U23601 ( .C1(n20666), .C2(n20691), .A(n20665), .B(n20664), .ZN(
        n20667) );
  AOI21_X1 U23602 ( .B1(n13732), .B2(n20668), .A(n20667), .ZN(n20669) );
  OAI21_X1 U23603 ( .B1(n20676), .B2(n21435), .A(n20669), .ZN(P1_U2833) );
  AND3_X1 U23604 ( .A1(n20672), .A2(n20671), .A3(n20670), .ZN(n20673) );
  AOI21_X1 U23605 ( .B1(n20674), .B2(n20705), .A(n20673), .ZN(n20682) );
  INV_X1 U23606 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21433) );
  NAND2_X1 U23607 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n20675) );
  OAI211_X1 U23608 ( .C1(n21433), .C2(n20676), .A(n20675), .B(n20688), .ZN(
        n20680) );
  NOR2_X1 U23609 ( .A1(n20678), .A2(n20677), .ZN(n20679) );
  AOI211_X1 U23610 ( .C1(n20685), .C2(P1_EBX_REG_6__SCAN_IN), .A(n20680), .B(
        n20679), .ZN(n20681) );
  OAI211_X1 U23611 ( .C1(n20683), .C2(n20691), .A(n20682), .B(n20681), .ZN(
        P1_U2834) );
  INV_X1 U23612 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21429) );
  INV_X1 U23613 ( .A(n20684), .ZN(n20787) );
  AOI22_X1 U23614 ( .A1(n20705), .A2(n20787), .B1(n20685), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n20695) );
  NAND2_X1 U23615 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20686) );
  NOR2_X1 U23616 ( .A1(n20687), .A2(n20686), .ZN(n20697) );
  NAND3_X1 U23617 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20697), .A3(n21429), 
        .ZN(n20689) );
  OAI211_X1 U23618 ( .C1(n20690), .C2(n20701), .A(n20689), .B(n20688), .ZN(
        n20693) );
  OAI211_X1 U23619 ( .C1(n21429), .C2(n20696), .A(n20695), .B(n20694), .ZN(
        P1_U2836) );
  NAND2_X1 U23620 ( .A1(n20697), .A2(n14493), .ZN(n20700) );
  NAND2_X1 U23621 ( .A1(n20698), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n20699) );
  OAI211_X1 U23622 ( .C1(n20702), .C2(n20701), .A(n20700), .B(n20699), .ZN(
        n20703) );
  INV_X1 U23623 ( .A(n20703), .ZN(n20717) );
  INV_X1 U23624 ( .A(n20704), .ZN(n20793) );
  AOI22_X1 U23625 ( .A1(n20705), .A2(n20793), .B1(n20685), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20716) );
  INV_X1 U23626 ( .A(n20706), .ZN(n20711) );
  INV_X1 U23627 ( .A(n20707), .ZN(n20708) );
  AOI22_X1 U23628 ( .A1(n20711), .A2(n20710), .B1(n20709), .B2(n20708), .ZN(
        n20715) );
  OAI21_X1 U23629 ( .B1(n20713), .B2(n20712), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n20714) );
  NAND4_X1 U23630 ( .A1(n20717), .A2(n20716), .A3(n20715), .A4(n20714), .ZN(
        P1_U2837) );
  AOI22_X1 U23631 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20718), .B1(n20737), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20719) );
  OAI21_X1 U23632 ( .B1(n21615), .B2(n20720), .A(n20719), .ZN(P1_U2921) );
  AOI22_X1 U23633 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20721) );
  OAI21_X1 U23634 ( .B1(n21625), .B2(n20740), .A(n20721), .ZN(P1_U2922) );
  AOI22_X1 U23635 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20722) );
  OAI21_X1 U23636 ( .B1(n15184), .B2(n20740), .A(n20722), .ZN(P1_U2923) );
  AOI22_X1 U23637 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20723) );
  OAI21_X1 U23638 ( .B1(n15186), .B2(n20740), .A(n20723), .ZN(P1_U2924) );
  AOI22_X1 U23639 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20724) );
  OAI21_X1 U23640 ( .B1(n15187), .B2(n20740), .A(n20724), .ZN(P1_U2925) );
  AOI22_X1 U23641 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20725) );
  OAI21_X1 U23642 ( .B1(n15190), .B2(n20740), .A(n20725), .ZN(P1_U2926) );
  AOI22_X1 U23643 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20726) );
  OAI21_X1 U23644 ( .B1(n15192), .B2(n20740), .A(n20726), .ZN(P1_U2927) );
  AOI22_X1 U23645 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20727) );
  OAI21_X1 U23646 ( .B1(n20728), .B2(n20740), .A(n20727), .ZN(P1_U2928) );
  AOI22_X1 U23647 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20729) );
  OAI21_X1 U23648 ( .B1(n11031), .B2(n20740), .A(n20729), .ZN(P1_U2929) );
  AOI22_X1 U23649 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20730) );
  OAI21_X1 U23650 ( .B1(n11039), .B2(n20740), .A(n20730), .ZN(P1_U2930) );
  AOI22_X1 U23651 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20731) );
  OAI21_X1 U23652 ( .B1(n11024), .B2(n20740), .A(n20731), .ZN(P1_U2931) );
  AOI22_X1 U23653 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20732) );
  OAI21_X1 U23654 ( .B1(n20733), .B2(n20740), .A(n20732), .ZN(P1_U2932) );
  AOI22_X1 U23655 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20734) );
  OAI21_X1 U23656 ( .B1(n11000), .B2(n20740), .A(n20734), .ZN(P1_U2933) );
  AOI22_X1 U23657 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20735) );
  OAI21_X1 U23658 ( .B1(n10972), .B2(n20740), .A(n20735), .ZN(P1_U2934) );
  AOI22_X1 U23659 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20736) );
  OAI21_X1 U23660 ( .B1(n10980), .B2(n20740), .A(n20736), .ZN(P1_U2935) );
  AOI22_X1 U23661 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20738), .B1(n20737), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20739) );
  OAI21_X1 U23662 ( .B1(n20741), .B2(n20740), .A(n20739), .ZN(P1_U2936) );
  AOI22_X1 U23663 ( .A1(n20770), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20765), .ZN(n20744) );
  INV_X1 U23664 ( .A(n20742), .ZN(n20743) );
  NAND2_X1 U23665 ( .A1(n20757), .A2(n20743), .ZN(n20759) );
  NAND2_X1 U23666 ( .A1(n20744), .A2(n20759), .ZN(P1_U2946) );
  AOI22_X1 U23667 ( .A1(n20770), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20765), .ZN(n20747) );
  INV_X1 U23668 ( .A(n20745), .ZN(n20746) );
  NAND2_X1 U23669 ( .A1(n20757), .A2(n20746), .ZN(n20761) );
  NAND2_X1 U23670 ( .A1(n20747), .A2(n20761), .ZN(P1_U2947) );
  AOI22_X1 U23671 ( .A1(n20770), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20765), .ZN(n20749) );
  NAND2_X1 U23672 ( .A1(n20757), .A2(n20748), .ZN(n20763) );
  NAND2_X1 U23673 ( .A1(n20749), .A2(n20763), .ZN(P1_U2948) );
  AOI22_X1 U23674 ( .A1(n20770), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20765), .ZN(n20752) );
  INV_X1 U23675 ( .A(n20750), .ZN(n20751) );
  NAND2_X1 U23676 ( .A1(n20757), .A2(n20751), .ZN(n20766) );
  NAND2_X1 U23677 ( .A1(n20752), .A2(n20766), .ZN(P1_U2949) );
  AOI22_X1 U23678 ( .A1(n20770), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20765), .ZN(n20755) );
  INV_X1 U23679 ( .A(n20753), .ZN(n20754) );
  NAND2_X1 U23680 ( .A1(n20757), .A2(n20754), .ZN(n20768) );
  NAND2_X1 U23681 ( .A1(n20755), .A2(n20768), .ZN(P1_U2950) );
  AOI22_X1 U23682 ( .A1(n20770), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20765), .ZN(n20758) );
  NAND2_X1 U23683 ( .A1(n20757), .A2(n20756), .ZN(n20771) );
  NAND2_X1 U23684 ( .A1(n20758), .A2(n20771), .ZN(P1_U2951) );
  AOI22_X1 U23685 ( .A1(n20770), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20765), .ZN(n20760) );
  NAND2_X1 U23686 ( .A1(n20760), .A2(n20759), .ZN(P1_U2961) );
  AOI22_X1 U23687 ( .A1(n20770), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20765), .ZN(n20762) );
  NAND2_X1 U23688 ( .A1(n20762), .A2(n20761), .ZN(P1_U2962) );
  AOI22_X1 U23689 ( .A1(n20770), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20765), .ZN(n20764) );
  NAND2_X1 U23690 ( .A1(n20764), .A2(n20763), .ZN(P1_U2963) );
  AOI22_X1 U23691 ( .A1(n20770), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20765), .ZN(n20767) );
  NAND2_X1 U23692 ( .A1(n20767), .A2(n20766), .ZN(P1_U2964) );
  AOI22_X1 U23693 ( .A1(n20770), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20765), .ZN(n20769) );
  NAND2_X1 U23694 ( .A1(n20769), .A2(n20768), .ZN(P1_U2965) );
  AOI22_X1 U23695 ( .A1(n20770), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20765), .ZN(n20772) );
  NAND2_X1 U23696 ( .A1(n20772), .A2(n20771), .ZN(P1_U2966) );
  AOI22_X1 U23697 ( .A1(n20773), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20786), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20782) );
  AOI21_X1 U23698 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20775), .A(
        n20774), .ZN(n20777) );
  XNOR2_X1 U23699 ( .A(n9633), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n20776) );
  XNOR2_X1 U23700 ( .A(n20777), .B(n20776), .ZN(n20788) );
  AOI22_X1 U23701 ( .A1(n20788), .A2(n20780), .B1(n20779), .B2(n9918), .ZN(
        n20781) );
  OAI211_X1 U23702 ( .C1(n20784), .C2(n20783), .A(n20782), .B(n20781), .ZN(
        P1_U2995) );
  OAI21_X1 U23703 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20785), .ZN(n20791) );
  AOI22_X1 U23704 ( .A1(n20801), .A2(n20787), .B1(n20786), .B2(
        P1_REIP_REG_4__SCAN_IN), .ZN(n20790) );
  AOI22_X1 U23705 ( .A1(n20788), .A2(n20795), .B1(
        P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n20794), .ZN(n20789) );
  OAI211_X1 U23706 ( .C1(n20799), .C2(n20791), .A(n20790), .B(n20789), .ZN(
        P1_U3027) );
  AOI21_X1 U23707 ( .B1(n20801), .B2(n20793), .A(n20792), .ZN(n20798) );
  AOI22_X1 U23708 ( .A1(n20796), .A2(n20795), .B1(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n20794), .ZN(n20797) );
  OAI211_X1 U23709 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n20799), .A(
        n20798), .B(n20797), .ZN(P1_U3028) );
  AOI21_X1 U23710 ( .B1(n20801), .B2(n10433), .A(n20800), .ZN(n20816) );
  AND2_X1 U23711 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20804) );
  INV_X1 U23712 ( .A(n20802), .ZN(n20803) );
  AOI21_X1 U23713 ( .B1(n20805), .B2(n20804), .A(n20803), .ZN(n20806) );
  OAI22_X1 U23714 ( .A1(n20808), .A2(n20807), .B1(n20806), .B2(n20812), .ZN(
        n20809) );
  INV_X1 U23715 ( .A(n20809), .ZN(n20815) );
  NAND4_X1 U23716 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20812), .A3(
        n20811), .A4(n20810), .ZN(n20813) );
  NAND4_X1 U23717 ( .A1(n20816), .A2(n20815), .A3(n20814), .A4(n20813), .ZN(
        P1_U3029) );
  NOR2_X1 U23718 ( .A1(n20818), .A2(n20817), .ZN(P1_U3032) );
  AOI22_X2 U23719 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9746), .B1(DATAI_17_), 
        .B2(n9567), .ZN(n21360) );
  AOI22_X1 U23720 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20852), .B1(DATAI_25_), 
        .B2(n20853), .ZN(n21310) );
  NAND2_X1 U23721 ( .A1(n20854), .A2(n20819), .ZN(n21230) );
  OAI22_X1 U23722 ( .A1(n21401), .A2(n21310), .B1(n20855), .B2(n21230), .ZN(
        n20820) );
  INV_X1 U23723 ( .A(n20820), .ZN(n20823) );
  NOR2_X2 U23724 ( .A1(n20821), .A2(n20973), .ZN(n21355) );
  AOI22_X1 U23725 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20859), .B1(
        n21355), .B2(n20858), .ZN(n20822) );
  OAI211_X1 U23726 ( .C1(n21360), .C2(n20888), .A(n20823), .B(n20822), .ZN(
        P1_U3034) );
  AOI22_X1 U23727 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20852), .B1(DATAI_18_), 
        .B2(n20853), .ZN(n21366) );
  AOI22_X2 U23728 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9746), .B1(DATAI_26_), 
        .B2(n9567), .ZN(n21314) );
  NAND2_X1 U23729 ( .A1(n20854), .A2(n20824), .ZN(n21234) );
  OAI22_X1 U23730 ( .A1(n21401), .A2(n21314), .B1(n20855), .B2(n21234), .ZN(
        n20825) );
  INV_X1 U23731 ( .A(n20825), .ZN(n20828) );
  NOR2_X2 U23732 ( .A1(n20973), .A2(n20826), .ZN(n21361) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20859), .B1(
        n21361), .B2(n20858), .ZN(n20827) );
  OAI211_X1 U23734 ( .C1(n21366), .C2(n20888), .A(n20828), .B(n20827), .ZN(
        P1_U3035) );
  AOI22_X1 U23735 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20852), .B1(DATAI_19_), 
        .B2(n20853), .ZN(n21372) );
  AOI22_X2 U23736 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9746), .B1(DATAI_27_), 
        .B2(n9567), .ZN(n21318) );
  NAND2_X1 U23737 ( .A1(n20854), .A2(n10811), .ZN(n21238) );
  OAI22_X1 U23738 ( .A1(n21401), .A2(n21318), .B1(n20855), .B2(n21238), .ZN(
        n20829) );
  INV_X1 U23739 ( .A(n20829), .ZN(n20832) );
  NOR2_X2 U23740 ( .A1(n20973), .A2(n20830), .ZN(n21367) );
  AOI22_X1 U23741 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20859), .B1(
        n21367), .B2(n20858), .ZN(n20831) );
  OAI211_X1 U23742 ( .C1(n21372), .C2(n20888), .A(n20832), .B(n20831), .ZN(
        P1_U3036) );
  AOI22_X2 U23743 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n9746), .B1(DATAI_20_), 
        .B2(n9567), .ZN(n21378) );
  AOI22_X1 U23744 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20852), .B1(DATAI_28_), 
        .B2(n20853), .ZN(n21322) );
  NAND2_X1 U23745 ( .A1(n20854), .A2(n20833), .ZN(n21242) );
  OAI22_X1 U23746 ( .A1(n21401), .A2(n21322), .B1(n20855), .B2(n21242), .ZN(
        n20834) );
  INV_X1 U23747 ( .A(n20834), .ZN(n20837) );
  NOR2_X2 U23748 ( .A1(n20973), .A2(n20835), .ZN(n21373) );
  AOI22_X1 U23749 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20859), .B1(
        n21373), .B2(n20858), .ZN(n20836) );
  OAI211_X1 U23750 ( .C1(n21378), .C2(n20888), .A(n20837), .B(n20836), .ZN(
        P1_U3037) );
  AOI22_X1 U23751 ( .A1(DATAI_21_), .A2(n20853), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20852), .ZN(n21384) );
  AOI22_X2 U23752 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9746), .B1(DATAI_29_), 
        .B2(n9567), .ZN(n21326) );
  NAND2_X1 U23753 ( .A1(n20854), .A2(n20838), .ZN(n21246) );
  OAI22_X1 U23754 ( .A1(n21401), .A2(n21326), .B1(n20855), .B2(n21246), .ZN(
        n20839) );
  INV_X1 U23755 ( .A(n20839), .ZN(n20842) );
  NOR2_X2 U23756 ( .A1(n20973), .A2(n20840), .ZN(n21379) );
  AOI22_X1 U23757 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20859), .B1(
        n21379), .B2(n20858), .ZN(n20841) );
  OAI211_X1 U23758 ( .C1(n21384), .C2(n20888), .A(n20842), .B(n20841), .ZN(
        P1_U3038) );
  AOI22_X2 U23759 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9746), .B1(DATAI_30_), 
        .B2(n9567), .ZN(n21392) );
  OAI22_X1 U23760 ( .A1(n21401), .A2(n21392), .B1(n20855), .B2(n21250), .ZN(
        n20843) );
  INV_X1 U23761 ( .A(n20843), .ZN(n20849) );
  NOR2_X2 U23762 ( .A1(n20973), .A2(n20844), .ZN(n21385) );
  INV_X1 U23763 ( .A(n9746), .ZN(n20847) );
  INV_X1 U23764 ( .A(DATAI_22_), .ZN(n20846) );
  INV_X1 U23765 ( .A(n20853), .ZN(n20845) );
  OAI22_X2 U23766 ( .A1(n16039), .A2(n20847), .B1(n20846), .B2(n20845), .ZN(
        n21387) );
  AOI22_X1 U23767 ( .A1(n21385), .A2(n20858), .B1(n20876), .B2(n21387), .ZN(
        n20848) );
  OAI211_X1 U23768 ( .C1(n20851), .C2(n20850), .A(n20849), .B(n20848), .ZN(
        P1_U3039) );
  AOI22_X1 U23769 ( .A1(DATAI_31_), .A2(n9567), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n9746), .ZN(n21336) );
  NAND2_X1 U23770 ( .A1(n20854), .A2(n10599), .ZN(n21256) );
  OAI22_X1 U23771 ( .A1(n21401), .A2(n9748), .B1(n20855), .B2(n21256), .ZN(
        n20856) );
  INV_X1 U23772 ( .A(n20856), .ZN(n20861) );
  NOR2_X2 U23773 ( .A1(n20973), .A2(n20857), .ZN(n21394) );
  AOI22_X1 U23774 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20859), .B1(
        n21394), .B2(n20858), .ZN(n20860) );
  OAI211_X1 U23775 ( .C1(n21402), .C2(n20888), .A(n20861), .B(n20860), .ZN(
        P1_U3040) );
  INV_X1 U23776 ( .A(n20933), .ZN(n20863) );
  INV_X1 U23777 ( .A(n20862), .ZN(n21266) );
  NOR2_X1 U23778 ( .A1(n21264), .A2(n20864), .ZN(n20883) );
  AOI21_X1 U23779 ( .B1(n20863), .B2(n21266), .A(n20883), .ZN(n20865) );
  OAI22_X1 U23780 ( .A1(n20865), .A2(n21341), .B1(n20864), .B2(n11005), .ZN(
        n20884) );
  AOI22_X1 U23781 ( .A1(n20884), .A2(n21342), .B1(n21343), .B2(n20883), .ZN(
        n20869) );
  INV_X1 U23782 ( .A(n20864), .ZN(n20867) );
  OAI211_X1 U23783 ( .C1(n20930), .C2(n21497), .A(n21349), .B(n20865), .ZN(
        n20866) );
  OAI211_X1 U23784 ( .C1(n21349), .C2(n20867), .A(n21348), .B(n20866), .ZN(
        n20885) );
  INV_X1 U23785 ( .A(n21306), .ZN(n21351) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20885), .B1(
        n20876), .B2(n21351), .ZN(n20868) );
  OAI211_X1 U23787 ( .C1(n21354), .C2(n20920), .A(n20869), .B(n20868), .ZN(
        P1_U3041) );
  AOI22_X1 U23788 ( .A1(n20884), .A2(n21355), .B1(n21356), .B2(n20883), .ZN(
        n20871) );
  INV_X1 U23789 ( .A(n21310), .ZN(n21357) );
  AOI22_X1 U23790 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20885), .B1(
        n20876), .B2(n21357), .ZN(n20870) );
  OAI211_X1 U23791 ( .C1(n21360), .C2(n20920), .A(n20871), .B(n20870), .ZN(
        P1_U3042) );
  AOI22_X1 U23792 ( .A1(n20884), .A2(n21361), .B1(n21362), .B2(n20883), .ZN(
        n20873) );
  INV_X1 U23793 ( .A(n21366), .ZN(n21311) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20885), .B1(
        n20891), .B2(n21311), .ZN(n20872) );
  OAI211_X1 U23795 ( .C1(n21314), .C2(n20888), .A(n20873), .B(n20872), .ZN(
        P1_U3043) );
  AOI22_X1 U23796 ( .A1(n20884), .A2(n21367), .B1(n21368), .B2(n20883), .ZN(
        n20875) );
  INV_X1 U23797 ( .A(n21372), .ZN(n21315) );
  AOI22_X1 U23798 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20885), .B1(
        n20891), .B2(n21315), .ZN(n20874) );
  OAI211_X1 U23799 ( .C1(n21318), .C2(n20888), .A(n20875), .B(n20874), .ZN(
        P1_U3044) );
  AOI22_X1 U23800 ( .A1(n20884), .A2(n21373), .B1(n21374), .B2(n20883), .ZN(
        n20878) );
  INV_X1 U23801 ( .A(n21322), .ZN(n21375) );
  AOI22_X1 U23802 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20885), .B1(
        n20876), .B2(n21375), .ZN(n20877) );
  OAI211_X1 U23803 ( .C1(n21378), .C2(n20920), .A(n20878), .B(n20877), .ZN(
        P1_U3045) );
  AOI22_X1 U23804 ( .A1(n20884), .A2(n21379), .B1(n21380), .B2(n20883), .ZN(
        n20880) );
  INV_X1 U23805 ( .A(n21384), .ZN(n21323) );
  AOI22_X1 U23806 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20885), .B1(
        n20891), .B2(n21323), .ZN(n20879) );
  OAI211_X1 U23807 ( .C1(n21326), .C2(n20888), .A(n20880), .B(n20879), .ZN(
        P1_U3046) );
  AOI22_X1 U23808 ( .A1(n20884), .A2(n21385), .B1(n21386), .B2(n20883), .ZN(
        n20882) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20885), .B1(
        n20891), .B2(n21387), .ZN(n20881) );
  OAI211_X1 U23810 ( .C1(n21392), .C2(n20888), .A(n20882), .B(n20881), .ZN(
        P1_U3047) );
  AOI22_X1 U23811 ( .A1(n20884), .A2(n21394), .B1(n21396), .B2(n20883), .ZN(
        n20887) );
  INV_X1 U23812 ( .A(n21402), .ZN(n21331) );
  AOI22_X1 U23813 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20885), .B1(
        n20891), .B2(n21331), .ZN(n20886) );
  OAI211_X1 U23814 ( .C1(n9748), .C2(n20888), .A(n20887), .B(n20886), .ZN(
        P1_U3048) );
  NAND3_X1 U23815 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n21184), .A3(
        n21143), .ZN(n20938) );
  OR2_X1 U23816 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20938), .ZN(
        n20919) );
  OAI22_X1 U23817 ( .A1(n20962), .A2(n21354), .B1(n20919), .B2(n21217), .ZN(
        n20890) );
  INV_X1 U23818 ( .A(n20890), .ZN(n20900) );
  INV_X1 U23819 ( .A(n20962), .ZN(n20892) );
  OAI21_X1 U23820 ( .B1(n20892), .B2(n20891), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20893) );
  NAND2_X1 U23821 ( .A1(n20893), .A2(n21349), .ZN(n20898) );
  NOR2_X1 U23822 ( .A1(n20933), .A2(n14504), .ZN(n20896) );
  OR2_X1 U23823 ( .A1(n21148), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21029) );
  AND2_X1 U23824 ( .A1(n21029), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21025) );
  AOI211_X1 U23825 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20919), .A(n21025), 
        .B(n20894), .ZN(n20895) );
  INV_X1 U23826 ( .A(n20896), .ZN(n20897) );
  AOI22_X1 U23827 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20923), .B1(
        n21342), .B2(n20922), .ZN(n20899) );
  OAI211_X1 U23828 ( .C1(n21306), .C2(n20920), .A(n20900), .B(n20899), .ZN(
        P1_U3049) );
  OAI22_X1 U23829 ( .A1(n20920), .A2(n21310), .B1(n21230), .B2(n20919), .ZN(
        n20901) );
  INV_X1 U23830 ( .A(n20901), .ZN(n20903) );
  AOI22_X1 U23831 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20923), .B1(
        n21355), .B2(n20922), .ZN(n20902) );
  OAI211_X1 U23832 ( .C1(n21360), .C2(n20962), .A(n20903), .B(n20902), .ZN(
        P1_U3050) );
  OAI22_X1 U23833 ( .A1(n20962), .A2(n21366), .B1(n21234), .B2(n20919), .ZN(
        n20904) );
  INV_X1 U23834 ( .A(n20904), .ZN(n20906) );
  AOI22_X1 U23835 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20923), .B1(
        n21361), .B2(n20922), .ZN(n20905) );
  OAI211_X1 U23836 ( .C1(n21314), .C2(n20920), .A(n20906), .B(n20905), .ZN(
        P1_U3051) );
  OAI22_X1 U23837 ( .A1(n20962), .A2(n21372), .B1(n21238), .B2(n20919), .ZN(
        n20907) );
  INV_X1 U23838 ( .A(n20907), .ZN(n20909) );
  AOI22_X1 U23839 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20923), .B1(
        n21367), .B2(n20922), .ZN(n20908) );
  OAI211_X1 U23840 ( .C1(n21318), .C2(n20920), .A(n20909), .B(n20908), .ZN(
        P1_U3052) );
  OAI22_X1 U23841 ( .A1(n20962), .A2(n21378), .B1(n21242), .B2(n20919), .ZN(
        n20910) );
  INV_X1 U23842 ( .A(n20910), .ZN(n20912) );
  AOI22_X1 U23843 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20923), .B1(
        n21373), .B2(n20922), .ZN(n20911) );
  OAI211_X1 U23844 ( .C1(n21322), .C2(n20920), .A(n20912), .B(n20911), .ZN(
        P1_U3053) );
  OAI22_X1 U23845 ( .A1(n20962), .A2(n21384), .B1(n21246), .B2(n20919), .ZN(
        n20913) );
  INV_X1 U23846 ( .A(n20913), .ZN(n20915) );
  AOI22_X1 U23847 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20923), .B1(
        n21379), .B2(n20922), .ZN(n20914) );
  OAI211_X1 U23848 ( .C1(n21326), .C2(n20920), .A(n20915), .B(n20914), .ZN(
        P1_U3054) );
  INV_X1 U23849 ( .A(n21387), .ZN(n21251) );
  OAI22_X1 U23850 ( .A1(n20962), .A2(n21251), .B1(n21250), .B2(n20919), .ZN(
        n20916) );
  INV_X1 U23851 ( .A(n20916), .ZN(n20918) );
  AOI22_X1 U23852 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20923), .B1(
        n21385), .B2(n20922), .ZN(n20917) );
  OAI211_X1 U23853 ( .C1(n21392), .C2(n20920), .A(n20918), .B(n20917), .ZN(
        P1_U3055) );
  OAI22_X1 U23854 ( .A1(n20920), .A2(n9748), .B1(n21256), .B2(n20919), .ZN(
        n20921) );
  INV_X1 U23855 ( .A(n20921), .ZN(n20925) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20923), .B1(
        n21394), .B2(n20922), .ZN(n20924) );
  OAI211_X1 U23857 ( .C1(n21402), .C2(n20962), .A(n20925), .B(n20924), .ZN(
        P1_U3056) );
  INV_X1 U23858 ( .A(n21185), .ZN(n20927) );
  NAND2_X1 U23859 ( .A1(n20927), .A2(n21184), .ZN(n20961) );
  OAI22_X1 U23860 ( .A1(n20962), .A2(n21306), .B1(n20961), .B2(n21217), .ZN(
        n20928) );
  INV_X1 U23861 ( .A(n20928), .ZN(n20942) );
  AOI21_X1 U23862 ( .B1(n21349), .B2(n20930), .A(n20929), .ZN(n20939) );
  AND2_X1 U23863 ( .A1(n20931), .A2(n10986), .ZN(n21338) );
  INV_X1 U23864 ( .A(n21338), .ZN(n20932) );
  OR2_X1 U23865 ( .A1(n20933), .A2(n20932), .ZN(n20934) );
  INV_X1 U23866 ( .A(n20940), .ZN(n20937) );
  INV_X1 U23867 ( .A(n21348), .ZN(n20935) );
  AOI21_X1 U23868 ( .B1(n21341), .B2(n20938), .A(n20935), .ZN(n20936) );
  AOI22_X1 U23869 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20965), .B1(
        n21342), .B2(n20964), .ZN(n20941) );
  OAI211_X1 U23870 ( .C1(n21354), .C2(n20990), .A(n20942), .B(n20941), .ZN(
        P1_U3057) );
  OAI22_X1 U23871 ( .A1(n20990), .A2(n21360), .B1(n21230), .B2(n20961), .ZN(
        n20943) );
  INV_X1 U23872 ( .A(n20943), .ZN(n20945) );
  AOI22_X1 U23873 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20965), .B1(
        n21355), .B2(n20964), .ZN(n20944) );
  OAI211_X1 U23874 ( .C1(n21310), .C2(n20962), .A(n20945), .B(n20944), .ZN(
        P1_U3058) );
  OAI22_X1 U23875 ( .A1(n20990), .A2(n21366), .B1(n21234), .B2(n20961), .ZN(
        n20946) );
  INV_X1 U23876 ( .A(n20946), .ZN(n20948) );
  AOI22_X1 U23877 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20965), .B1(
        n21361), .B2(n20964), .ZN(n20947) );
  OAI211_X1 U23878 ( .C1(n21314), .C2(n20962), .A(n20948), .B(n20947), .ZN(
        P1_U3059) );
  OAI22_X1 U23879 ( .A1(n20962), .A2(n21318), .B1(n21238), .B2(n20961), .ZN(
        n20949) );
  INV_X1 U23880 ( .A(n20949), .ZN(n20951) );
  AOI22_X1 U23881 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20965), .B1(
        n21367), .B2(n20964), .ZN(n20950) );
  OAI211_X1 U23882 ( .C1(n21372), .C2(n20990), .A(n20951), .B(n20950), .ZN(
        P1_U3060) );
  OAI22_X1 U23883 ( .A1(n20962), .A2(n21322), .B1(n21242), .B2(n20961), .ZN(
        n20952) );
  INV_X1 U23884 ( .A(n20952), .ZN(n20954) );
  AOI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20965), .B1(
        n21373), .B2(n20964), .ZN(n20953) );
  OAI211_X1 U23886 ( .C1(n21378), .C2(n20990), .A(n20954), .B(n20953), .ZN(
        P1_U3061) );
  OAI22_X1 U23887 ( .A1(n20990), .A2(n21384), .B1(n21246), .B2(n20961), .ZN(
        n20955) );
  INV_X1 U23888 ( .A(n20955), .ZN(n20957) );
  AOI22_X1 U23889 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20965), .B1(
        n21379), .B2(n20964), .ZN(n20956) );
  OAI211_X1 U23890 ( .C1(n21326), .C2(n20962), .A(n20957), .B(n20956), .ZN(
        P1_U3062) );
  OAI22_X1 U23891 ( .A1(n20990), .A2(n21251), .B1(n21250), .B2(n20961), .ZN(
        n20958) );
  INV_X1 U23892 ( .A(n20958), .ZN(n20960) );
  AOI22_X1 U23893 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20965), .B1(
        n21385), .B2(n20964), .ZN(n20959) );
  OAI211_X1 U23894 ( .C1(n21392), .C2(n20962), .A(n20960), .B(n20959), .ZN(
        P1_U3063) );
  OAI22_X1 U23895 ( .A1(n20962), .A2(n9748), .B1(n21256), .B2(n20961), .ZN(
        n20963) );
  INV_X1 U23896 ( .A(n20963), .ZN(n20967) );
  AOI22_X1 U23897 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20965), .B1(
        n21394), .B2(n20964), .ZN(n20966) );
  OAI211_X1 U23898 ( .C1(n21402), .C2(n20990), .A(n20967), .B(n20966), .ZN(
        P1_U3064) );
  NAND3_X1 U23899 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n21184), .A3(
        n21216), .ZN(n20997) );
  NOR2_X1 U23900 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20997), .ZN(
        n20992) );
  NOR2_X1 U23901 ( .A1(n13984), .A2(n20968), .ZN(n21061) );
  NAND3_X1 U23902 ( .A1(n21061), .A2(n21349), .A3(n14504), .ZN(n20969) );
  AOI22_X1 U23903 ( .A1(n21343), .A2(n20992), .B1(n21342), .B2(n20991), .ZN(
        n20977) );
  AOI21_X1 U23904 ( .B1(n20990), .B2(n21016), .A(n21497), .ZN(n20971) );
  AOI21_X1 U23905 ( .B1(n21061), .B2(n14504), .A(n20971), .ZN(n20972) );
  NOR2_X1 U23906 ( .A1(n20972), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U23907 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21303), .ZN(n20976) );
  OAI211_X1 U23908 ( .C1(n21306), .C2(n20990), .A(n20977), .B(n20976), .ZN(
        P1_U3065) );
  AOI22_X1 U23909 ( .A1(n21356), .A2(n20992), .B1(n21355), .B2(n20991), .ZN(
        n20979) );
  INV_X1 U23910 ( .A(n20990), .ZN(n20993) );
  AOI22_X1 U23911 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20994), .B1(
        n20993), .B2(n21357), .ZN(n20978) );
  OAI211_X1 U23912 ( .C1(n21360), .C2(n21016), .A(n20979), .B(n20978), .ZN(
        P1_U3066) );
  AOI22_X1 U23913 ( .A1(n21362), .A2(n20992), .B1(n21361), .B2(n20991), .ZN(
        n20981) );
  AOI22_X1 U23914 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21311), .ZN(n20980) );
  OAI211_X1 U23915 ( .C1(n21314), .C2(n20990), .A(n20981), .B(n20980), .ZN(
        P1_U3067) );
  AOI22_X1 U23916 ( .A1(n21368), .A2(n20992), .B1(n21367), .B2(n20991), .ZN(
        n20983) );
  AOI22_X1 U23917 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21315), .ZN(n20982) );
  OAI211_X1 U23918 ( .C1(n21318), .C2(n20990), .A(n20983), .B(n20982), .ZN(
        P1_U3068) );
  AOI22_X1 U23919 ( .A1(n21374), .A2(n20992), .B1(n21373), .B2(n20991), .ZN(
        n20985) );
  INV_X1 U23920 ( .A(n21378), .ZN(n21319) );
  AOI22_X1 U23921 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21319), .ZN(n20984) );
  OAI211_X1 U23922 ( .C1(n21322), .C2(n20990), .A(n20985), .B(n20984), .ZN(
        P1_U3069) );
  AOI22_X1 U23923 ( .A1(n21380), .A2(n20992), .B1(n21379), .B2(n20991), .ZN(
        n20987) );
  AOI22_X1 U23924 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21323), .ZN(n20986) );
  OAI211_X1 U23925 ( .C1(n21326), .C2(n20990), .A(n20987), .B(n20986), .ZN(
        P1_U3070) );
  AOI22_X1 U23926 ( .A1(n21386), .A2(n20992), .B1(n21385), .B2(n20991), .ZN(
        n20989) );
  AOI22_X1 U23927 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20994), .B1(
        n21019), .B2(n21387), .ZN(n20988) );
  OAI211_X1 U23928 ( .C1(n21392), .C2(n20990), .A(n20989), .B(n20988), .ZN(
        P1_U3071) );
  AOI22_X1 U23929 ( .A1(n21396), .A2(n20992), .B1(n21394), .B2(n20991), .ZN(
        n20996) );
  AOI22_X1 U23930 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20994), .B1(
        n20993), .B2(n9747), .ZN(n20995) );
  OAI211_X1 U23931 ( .C1(n21402), .C2(n21016), .A(n20996), .B(n20995), .ZN(
        P1_U3072) );
  NOR2_X1 U23932 ( .A1(n21264), .A2(n20997), .ZN(n21018) );
  AOI21_X1 U23933 ( .B1(n21061), .B2(n21266), .A(n21018), .ZN(n20998) );
  OAI22_X1 U23934 ( .A1(n20998), .A2(n21341), .B1(n20997), .B2(n11005), .ZN(
        n21017) );
  AOI22_X1 U23935 ( .A1(n21343), .A2(n21018), .B1(n21342), .B2(n21017), .ZN(
        n21002) );
  INV_X1 U23936 ( .A(n20997), .ZN(n21000) );
  OAI211_X1 U23937 ( .C1(n21064), .C2(n21497), .A(n21349), .B(n20998), .ZN(
        n20999) );
  OAI211_X1 U23938 ( .C1(n21349), .C2(n21000), .A(n21348), .B(n20999), .ZN(
        n21020) );
  AOI22_X1 U23939 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21351), .ZN(n21001) );
  OAI211_X1 U23940 ( .C1(n21354), .C2(n21058), .A(n21002), .B(n21001), .ZN(
        P1_U3073) );
  AOI22_X1 U23941 ( .A1(n21356), .A2(n21018), .B1(n21355), .B2(n21017), .ZN(
        n21004) );
  AOI22_X1 U23942 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21357), .ZN(n21003) );
  OAI211_X1 U23943 ( .C1(n21360), .C2(n21058), .A(n21004), .B(n21003), .ZN(
        P1_U3074) );
  AOI22_X1 U23944 ( .A1(n21362), .A2(n21018), .B1(n21361), .B2(n21017), .ZN(
        n21006) );
  INV_X1 U23945 ( .A(n21314), .ZN(n21363) );
  AOI22_X1 U23946 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21363), .ZN(n21005) );
  OAI211_X1 U23947 ( .C1(n21366), .C2(n21058), .A(n21006), .B(n21005), .ZN(
        P1_U3075) );
  AOI22_X1 U23948 ( .A1(n21368), .A2(n21018), .B1(n21367), .B2(n21017), .ZN(
        n21008) );
  INV_X1 U23949 ( .A(n21318), .ZN(n21369) );
  AOI22_X1 U23950 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21369), .ZN(n21007) );
  OAI211_X1 U23951 ( .C1(n21372), .C2(n21058), .A(n21008), .B(n21007), .ZN(
        P1_U3076) );
  AOI22_X1 U23952 ( .A1(n21374), .A2(n21018), .B1(n21373), .B2(n21017), .ZN(
        n21010) );
  AOI22_X1 U23953 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n21375), .ZN(n21009) );
  OAI211_X1 U23954 ( .C1(n21378), .C2(n21058), .A(n21010), .B(n21009), .ZN(
        P1_U3077) );
  AOI22_X1 U23955 ( .A1(n21380), .A2(n21018), .B1(n21379), .B2(n21017), .ZN(
        n21012) );
  INV_X1 U23956 ( .A(n21058), .ZN(n21013) );
  AOI22_X1 U23957 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n21020), .B1(
        n21013), .B2(n21323), .ZN(n21011) );
  OAI211_X1 U23958 ( .C1(n21326), .C2(n21016), .A(n21012), .B(n21011), .ZN(
        P1_U3078) );
  AOI22_X1 U23959 ( .A1(n21386), .A2(n21018), .B1(n21385), .B2(n21017), .ZN(
        n21015) );
  AOI22_X1 U23960 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n21020), .B1(
        n21013), .B2(n21387), .ZN(n21014) );
  OAI211_X1 U23961 ( .C1(n21392), .C2(n21016), .A(n21015), .B(n21014), .ZN(
        P1_U3079) );
  AOI22_X1 U23962 ( .A1(n21396), .A2(n21018), .B1(n21394), .B2(n21017), .ZN(
        n21022) );
  AOI22_X1 U23963 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n21020), .B1(
        n21019), .B2(n9747), .ZN(n21021) );
  OAI211_X1 U23964 ( .C1(n21402), .C2(n21058), .A(n21022), .B(n21021), .ZN(
        P1_U3080) );
  INV_X1 U23965 ( .A(n21066), .ZN(n21062) );
  NOR2_X1 U23966 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21062), .ZN(
        n21027) );
  INV_X1 U23967 ( .A(n21027), .ZN(n21052) );
  OAI22_X1 U23968 ( .A1(n21087), .A2(n21354), .B1(n21052), .B2(n21217), .ZN(
        n21023) );
  INV_X1 U23969 ( .A(n21023), .ZN(n21033) );
  NAND3_X1 U23970 ( .A1(n21087), .A2(n21058), .A3(n21349), .ZN(n21024) );
  NAND2_X1 U23971 ( .A1(n21024), .A2(n21219), .ZN(n21028) );
  NAND2_X1 U23972 ( .A1(n21061), .A2(n21292), .ZN(n21030) );
  AOI21_X1 U23973 ( .B1(n21028), .B2(n21030), .A(n21025), .ZN(n21026) );
  INV_X1 U23974 ( .A(n21028), .ZN(n21031) );
  AOI22_X1 U23975 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n21055), .B1(
        n21342), .B2(n21054), .ZN(n21032) );
  OAI211_X1 U23976 ( .C1(n21306), .C2(n21058), .A(n21033), .B(n21032), .ZN(
        P1_U3081) );
  OAI22_X1 U23977 ( .A1(n21058), .A2(n21310), .B1(n21230), .B2(n21052), .ZN(
        n21034) );
  INV_X1 U23978 ( .A(n21034), .ZN(n21036) );
  AOI22_X1 U23979 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n21055), .B1(
        n21355), .B2(n21054), .ZN(n21035) );
  OAI211_X1 U23980 ( .C1(n21360), .C2(n21087), .A(n21036), .B(n21035), .ZN(
        P1_U3082) );
  OAI22_X1 U23981 ( .A1(n21087), .A2(n21366), .B1(n21052), .B2(n21234), .ZN(
        n21037) );
  INV_X1 U23982 ( .A(n21037), .ZN(n21039) );
  AOI22_X1 U23983 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n21055), .B1(
        n21361), .B2(n21054), .ZN(n21038) );
  OAI211_X1 U23984 ( .C1(n21314), .C2(n21058), .A(n21039), .B(n21038), .ZN(
        P1_U3083) );
  OAI22_X1 U23985 ( .A1(n21087), .A2(n21372), .B1(n21238), .B2(n21052), .ZN(
        n21040) );
  INV_X1 U23986 ( .A(n21040), .ZN(n21042) );
  AOI22_X1 U23987 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n21055), .B1(
        n21367), .B2(n21054), .ZN(n21041) );
  OAI211_X1 U23988 ( .C1(n21318), .C2(n21058), .A(n21042), .B(n21041), .ZN(
        P1_U3084) );
  OAI22_X1 U23989 ( .A1(n21087), .A2(n21378), .B1(n21242), .B2(n21052), .ZN(
        n21043) );
  INV_X1 U23990 ( .A(n21043), .ZN(n21045) );
  AOI22_X1 U23991 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n21055), .B1(
        n21373), .B2(n21054), .ZN(n21044) );
  OAI211_X1 U23992 ( .C1(n21322), .C2(n21058), .A(n21045), .B(n21044), .ZN(
        P1_U3085) );
  OAI22_X1 U23993 ( .A1(n21087), .A2(n21384), .B1(n21052), .B2(n21246), .ZN(
        n21046) );
  INV_X1 U23994 ( .A(n21046), .ZN(n21048) );
  AOI22_X1 U23995 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n21055), .B1(
        n21379), .B2(n21054), .ZN(n21047) );
  OAI211_X1 U23996 ( .C1(n21326), .C2(n21058), .A(n21048), .B(n21047), .ZN(
        P1_U3086) );
  OAI22_X1 U23997 ( .A1(n21087), .A2(n21251), .B1(n21250), .B2(n21052), .ZN(
        n21049) );
  INV_X1 U23998 ( .A(n21049), .ZN(n21051) );
  AOI22_X1 U23999 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n21055), .B1(
        n21385), .B2(n21054), .ZN(n21050) );
  OAI211_X1 U24000 ( .C1(n21392), .C2(n21058), .A(n21051), .B(n21050), .ZN(
        P1_U3087) );
  OAI22_X1 U24001 ( .A1(n21087), .A2(n21402), .B1(n21052), .B2(n21256), .ZN(
        n21053) );
  INV_X1 U24002 ( .A(n21053), .ZN(n21057) );
  AOI22_X1 U24003 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n21055), .B1(
        n21394), .B2(n21054), .ZN(n21056) );
  OAI211_X1 U24004 ( .C1(n9748), .C2(n21058), .A(n21057), .B(n21056), .ZN(
        P1_U3088) );
  INV_X1 U24005 ( .A(n21060), .ZN(n21083) );
  AOI21_X1 U24006 ( .B1(n21061), .B2(n21338), .A(n21083), .ZN(n21063) );
  OAI22_X1 U24007 ( .A1(n21063), .A2(n21341), .B1(n21062), .B2(n11005), .ZN(
        n21082) );
  AOI22_X1 U24008 ( .A1(n21343), .A2(n21083), .B1(n21342), .B2(n21082), .ZN(
        n21068) );
  OAI211_X1 U24009 ( .C1(n21346), .C2(n21064), .A(n21349), .B(n21063), .ZN(
        n21065) );
  OAI211_X1 U24010 ( .C1(n21066), .C2(n21349), .A(n21348), .B(n21065), .ZN(
        n21084) );
  AOI22_X1 U24011 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21351), .ZN(n21067) );
  OAI211_X1 U24012 ( .C1(n21354), .C2(n21115), .A(n21068), .B(n21067), .ZN(
        P1_U3089) );
  AOI22_X1 U24013 ( .A1(n21356), .A2(n21083), .B1(n21355), .B2(n21082), .ZN(
        n21070) );
  AOI22_X1 U24014 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21357), .ZN(n21069) );
  OAI211_X1 U24015 ( .C1(n21360), .C2(n21115), .A(n21070), .B(n21069), .ZN(
        P1_U3090) );
  AOI22_X1 U24016 ( .A1(n21362), .A2(n21083), .B1(n21361), .B2(n21082), .ZN(
        n21072) );
  AOI22_X1 U24017 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21363), .ZN(n21071) );
  OAI211_X1 U24018 ( .C1(n21366), .C2(n21115), .A(n21072), .B(n21071), .ZN(
        P1_U3091) );
  AOI22_X1 U24019 ( .A1(n21368), .A2(n21083), .B1(n21367), .B2(n21082), .ZN(
        n21074) );
  AOI22_X1 U24020 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21369), .ZN(n21073) );
  OAI211_X1 U24021 ( .C1(n21372), .C2(n21115), .A(n21074), .B(n21073), .ZN(
        P1_U3092) );
  AOI22_X1 U24022 ( .A1(n21374), .A2(n21083), .B1(n21373), .B2(n21082), .ZN(
        n21076) );
  AOI22_X1 U24023 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21375), .ZN(n21075) );
  OAI211_X1 U24024 ( .C1(n21378), .C2(n21115), .A(n21076), .B(n21075), .ZN(
        P1_U3093) );
  AOI22_X1 U24025 ( .A1(n21380), .A2(n21083), .B1(n21379), .B2(n21082), .ZN(
        n21079) );
  INV_X1 U24026 ( .A(n21326), .ZN(n21381) );
  AOI22_X1 U24027 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n21084), .B1(
        n21077), .B2(n21381), .ZN(n21078) );
  OAI211_X1 U24028 ( .C1(n21384), .C2(n21115), .A(n21079), .B(n21078), .ZN(
        P1_U3094) );
  AOI22_X1 U24029 ( .A1(n21386), .A2(n21083), .B1(n21385), .B2(n21082), .ZN(
        n21081) );
  INV_X1 U24030 ( .A(n21115), .ZN(n21092) );
  AOI22_X1 U24031 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n21084), .B1(
        n21092), .B2(n21387), .ZN(n21080) );
  OAI211_X1 U24032 ( .C1(n21392), .C2(n21087), .A(n21081), .B(n21080), .ZN(
        P1_U3095) );
  AOI22_X1 U24033 ( .A1(n21396), .A2(n21083), .B1(n21394), .B2(n21082), .ZN(
        n21086) );
  AOI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n21084), .B1(
        n21092), .B2(n21331), .ZN(n21085) );
  OAI211_X1 U24035 ( .C1(n9748), .C2(n21087), .A(n21086), .B(n21085), .ZN(
        P1_U3096) );
  NAND3_X1 U24036 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n21143), .A3(
        n21216), .ZN(n21117) );
  NOR2_X1 U24037 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21117), .ZN(
        n21111) );
  AND2_X1 U24038 ( .A1(n21088), .A2(n13984), .ZN(n21186) );
  AOI21_X1 U24039 ( .B1(n21186), .B2(n14504), .A(n21111), .ZN(n21093) );
  INV_X1 U24040 ( .A(n21089), .ZN(n21090) );
  NAND2_X1 U24041 ( .A1(n21090), .A2(n21148), .ZN(n21225) );
  OAI22_X1 U24042 ( .A1(n21093), .A2(n21341), .B1(n21154), .B2(n21225), .ZN(
        n21110) );
  AOI22_X1 U24043 ( .A1(n21343), .A2(n21111), .B1(n21110), .B2(n21342), .ZN(
        n21097) );
  INV_X1 U24044 ( .A(n21215), .ZN(n21091) );
  OAI21_X1 U24045 ( .B1(n21138), .B2(n21092), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21094) );
  NAND2_X1 U24046 ( .A1(n21094), .A2(n21093), .ZN(n21095) );
  AOI22_X1 U24047 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21303), .ZN(n21096) );
  OAI211_X1 U24048 ( .C1(n21306), .C2(n21115), .A(n21097), .B(n21096), .ZN(
        P1_U3097) );
  AOI22_X1 U24049 ( .A1(n21356), .A2(n21111), .B1(n21110), .B2(n21355), .ZN(
        n21099) );
  INV_X1 U24050 ( .A(n21360), .ZN(n21307) );
  AOI22_X1 U24051 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21307), .ZN(n21098) );
  OAI211_X1 U24052 ( .C1(n21310), .C2(n21115), .A(n21099), .B(n21098), .ZN(
        P1_U3098) );
  AOI22_X1 U24053 ( .A1(n21362), .A2(n21111), .B1(n21110), .B2(n21361), .ZN(
        n21101) );
  AOI22_X1 U24054 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21311), .ZN(n21100) );
  OAI211_X1 U24055 ( .C1(n21314), .C2(n21115), .A(n21101), .B(n21100), .ZN(
        P1_U3099) );
  AOI22_X1 U24056 ( .A1(n21368), .A2(n21111), .B1(n21110), .B2(n21367), .ZN(
        n21103) );
  AOI22_X1 U24057 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21315), .ZN(n21102) );
  OAI211_X1 U24058 ( .C1(n21318), .C2(n21115), .A(n21103), .B(n21102), .ZN(
        P1_U3100) );
  AOI22_X1 U24059 ( .A1(n21374), .A2(n21111), .B1(n21110), .B2(n21373), .ZN(
        n21105) );
  AOI22_X1 U24060 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21319), .ZN(n21104) );
  OAI211_X1 U24061 ( .C1(n21322), .C2(n21115), .A(n21105), .B(n21104), .ZN(
        P1_U3101) );
  AOI22_X1 U24062 ( .A1(n21380), .A2(n21111), .B1(n21110), .B2(n21379), .ZN(
        n21107) );
  AOI22_X1 U24063 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21323), .ZN(n21106) );
  OAI211_X1 U24064 ( .C1(n21326), .C2(n21115), .A(n21107), .B(n21106), .ZN(
        P1_U3102) );
  AOI22_X1 U24065 ( .A1(n21386), .A2(n21111), .B1(n21110), .B2(n21385), .ZN(
        n21109) );
  AOI22_X1 U24066 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21387), .ZN(n21108) );
  OAI211_X1 U24067 ( .C1(n21392), .C2(n21115), .A(n21109), .B(n21108), .ZN(
        P1_U3103) );
  AOI22_X1 U24068 ( .A1(n21396), .A2(n21111), .B1(n21110), .B2(n21394), .ZN(
        n21114) );
  AOI22_X1 U24069 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n21112), .B1(
        n21138), .B2(n21331), .ZN(n21113) );
  OAI211_X1 U24070 ( .C1(n9748), .C2(n21115), .A(n21114), .B(n21113), .ZN(
        P1_U3104) );
  INV_X1 U24071 ( .A(n21263), .ZN(n21116) );
  NOR2_X1 U24072 ( .A1(n21264), .A2(n21117), .ZN(n21137) );
  AOI21_X1 U24073 ( .B1(n21186), .B2(n21266), .A(n21137), .ZN(n21118) );
  OAI22_X1 U24074 ( .A1(n21118), .A2(n21341), .B1(n21117), .B2(n11005), .ZN(
        n21136) );
  AOI22_X1 U24075 ( .A1(n21343), .A2(n21137), .B1(n21136), .B2(n21342), .ZN(
        n21122) );
  INV_X1 U24076 ( .A(n21117), .ZN(n21120) );
  OAI211_X1 U24077 ( .C1(n21193), .C2(n21497), .A(n21349), .B(n21118), .ZN(
        n21119) );
  OAI211_X1 U24078 ( .C1(n21349), .C2(n21120), .A(n21348), .B(n21119), .ZN(
        n21139) );
  AOI22_X1 U24079 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n21139), .B1(
        n21138), .B2(n21351), .ZN(n21121) );
  OAI211_X1 U24080 ( .C1(n21354), .C2(n21183), .A(n21122), .B(n21121), .ZN(
        P1_U3105) );
  AOI22_X1 U24081 ( .A1(n21356), .A2(n21137), .B1(n21136), .B2(n21355), .ZN(
        n21124) );
  AOI22_X1 U24082 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n21139), .B1(
        n21145), .B2(n21307), .ZN(n21123) );
  OAI211_X1 U24083 ( .C1(n21310), .C2(n21135), .A(n21124), .B(n21123), .ZN(
        P1_U3106) );
  AOI22_X1 U24084 ( .A1(n21362), .A2(n21137), .B1(n21136), .B2(n21361), .ZN(
        n21126) );
  AOI22_X1 U24085 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n21139), .B1(
        n21145), .B2(n21311), .ZN(n21125) );
  OAI211_X1 U24086 ( .C1(n21314), .C2(n21135), .A(n21126), .B(n21125), .ZN(
        P1_U3107) );
  AOI22_X1 U24087 ( .A1(n21368), .A2(n21137), .B1(n21136), .B2(n21367), .ZN(
        n21128) );
  AOI22_X1 U24088 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n21139), .B1(
        n21145), .B2(n21315), .ZN(n21127) );
  OAI211_X1 U24089 ( .C1(n21318), .C2(n21135), .A(n21128), .B(n21127), .ZN(
        P1_U3108) );
  AOI22_X1 U24090 ( .A1(n21374), .A2(n21137), .B1(n21136), .B2(n21373), .ZN(
        n21130) );
  AOI22_X1 U24091 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n21139), .B1(
        n21138), .B2(n21375), .ZN(n21129) );
  OAI211_X1 U24092 ( .C1(n21378), .C2(n21183), .A(n21130), .B(n21129), .ZN(
        P1_U3109) );
  AOI22_X1 U24093 ( .A1(n21380), .A2(n21137), .B1(n21136), .B2(n21379), .ZN(
        n21132) );
  AOI22_X1 U24094 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n21139), .B1(
        n21145), .B2(n21323), .ZN(n21131) );
  OAI211_X1 U24095 ( .C1(n21326), .C2(n21135), .A(n21132), .B(n21131), .ZN(
        P1_U3110) );
  AOI22_X1 U24096 ( .A1(n21386), .A2(n21137), .B1(n21136), .B2(n21385), .ZN(
        n21134) );
  AOI22_X1 U24097 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n21139), .B1(
        n21145), .B2(n21387), .ZN(n21133) );
  OAI211_X1 U24098 ( .C1(n21392), .C2(n21135), .A(n21134), .B(n21133), .ZN(
        P1_U3111) );
  AOI22_X1 U24099 ( .A1(n21396), .A2(n21137), .B1(n21136), .B2(n21394), .ZN(
        n21141) );
  AOI22_X1 U24100 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n21139), .B1(
        n21138), .B2(n9747), .ZN(n21140) );
  OAI211_X1 U24101 ( .C1(n21402), .C2(n21183), .A(n21141), .B(n21140), .ZN(
        P1_U3112) );
  INV_X1 U24102 ( .A(n21295), .ZN(n21142) );
  NAND3_X1 U24103 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n21143), .ZN(n21187) );
  NOR2_X1 U24104 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21187), .ZN(
        n21150) );
  INV_X1 U24105 ( .A(n21150), .ZN(n21177) );
  OAI22_X1 U24106 ( .A1(n21214), .A2(n21354), .B1(n21177), .B2(n21217), .ZN(
        n21144) );
  INV_X1 U24107 ( .A(n21144), .ZN(n21158) );
  INV_X1 U24108 ( .A(n21214), .ZN(n21146) );
  OAI21_X1 U24109 ( .B1(n21146), .B2(n21145), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21147) );
  NAND2_X1 U24110 ( .A1(n21147), .A2(n21349), .ZN(n21156) );
  AND2_X1 U24111 ( .A1(n21186), .A2(n21292), .ZN(n21153) );
  OR2_X1 U24112 ( .A1(n21148), .A2(n21184), .ZN(n21294) );
  NAND2_X1 U24113 ( .A1(n21294), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21300) );
  OAI211_X1 U24114 ( .C1(n21222), .C2(n21150), .A(n21300), .B(n21149), .ZN(
        n21151) );
  INV_X1 U24115 ( .A(n21151), .ZN(n21152) );
  INV_X1 U24116 ( .A(n21153), .ZN(n21155) );
  AOI22_X1 U24117 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n21180), .B1(
        n21342), .B2(n21179), .ZN(n21157) );
  OAI211_X1 U24118 ( .C1(n21306), .C2(n21183), .A(n21158), .B(n21157), .ZN(
        P1_U3113) );
  OAI22_X1 U24119 ( .A1(n21214), .A2(n21360), .B1(n21177), .B2(n21230), .ZN(
        n21159) );
  INV_X1 U24120 ( .A(n21159), .ZN(n21161) );
  AOI22_X1 U24121 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n21180), .B1(
        n21355), .B2(n21179), .ZN(n21160) );
  OAI211_X1 U24122 ( .C1(n21310), .C2(n21183), .A(n21161), .B(n21160), .ZN(
        P1_U3114) );
  OAI22_X1 U24123 ( .A1(n21214), .A2(n21366), .B1(n21177), .B2(n21234), .ZN(
        n21162) );
  INV_X1 U24124 ( .A(n21162), .ZN(n21164) );
  AOI22_X1 U24125 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n21180), .B1(
        n21361), .B2(n21179), .ZN(n21163) );
  OAI211_X1 U24126 ( .C1(n21314), .C2(n21183), .A(n21164), .B(n21163), .ZN(
        P1_U3115) );
  OAI22_X1 U24127 ( .A1(n21183), .A2(n21318), .B1(n21177), .B2(n21238), .ZN(
        n21165) );
  INV_X1 U24128 ( .A(n21165), .ZN(n21167) );
  AOI22_X1 U24129 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n21180), .B1(
        n21367), .B2(n21179), .ZN(n21166) );
  OAI211_X1 U24130 ( .C1(n21372), .C2(n21214), .A(n21167), .B(n21166), .ZN(
        P1_U3116) );
  OAI22_X1 U24131 ( .A1(n21183), .A2(n21322), .B1(n21177), .B2(n21242), .ZN(
        n21168) );
  INV_X1 U24132 ( .A(n21168), .ZN(n21170) );
  AOI22_X1 U24133 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n21180), .B1(
        n21373), .B2(n21179), .ZN(n21169) );
  OAI211_X1 U24134 ( .C1(n21378), .C2(n21214), .A(n21170), .B(n21169), .ZN(
        P1_U3117) );
  OAI22_X1 U24135 ( .A1(n21214), .A2(n21384), .B1(n21177), .B2(n21246), .ZN(
        n21171) );
  INV_X1 U24136 ( .A(n21171), .ZN(n21173) );
  AOI22_X1 U24137 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n21180), .B1(
        n21379), .B2(n21179), .ZN(n21172) );
  OAI211_X1 U24138 ( .C1(n21326), .C2(n21183), .A(n21173), .B(n21172), .ZN(
        P1_U3118) );
  OAI22_X1 U24139 ( .A1(n21214), .A2(n21251), .B1(n21177), .B2(n21250), .ZN(
        n21174) );
  INV_X1 U24140 ( .A(n21174), .ZN(n21176) );
  AOI22_X1 U24141 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n21180), .B1(
        n21385), .B2(n21179), .ZN(n21175) );
  OAI211_X1 U24142 ( .C1(n21392), .C2(n21183), .A(n21176), .B(n21175), .ZN(
        P1_U3119) );
  OAI22_X1 U24143 ( .A1(n21214), .A2(n21402), .B1(n21177), .B2(n21256), .ZN(
        n21178) );
  INV_X1 U24144 ( .A(n21178), .ZN(n21182) );
  AOI22_X1 U24145 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n21180), .B1(
        n21394), .B2(n21179), .ZN(n21181) );
  OAI211_X1 U24146 ( .C1(n9748), .C2(n21183), .A(n21182), .B(n21181), .ZN(
        P1_U3120) );
  NOR2_X1 U24147 ( .A1(n21185), .A2(n21184), .ZN(n21209) );
  AOI21_X1 U24148 ( .B1(n21186), .B2(n21338), .A(n21209), .ZN(n21188) );
  OAI22_X1 U24149 ( .A1(n21188), .A2(n21341), .B1(n21187), .B2(n11005), .ZN(
        n21208) );
  AOI22_X1 U24150 ( .A1(n21343), .A2(n21209), .B1(n21208), .B2(n21342), .ZN(
        n21195) );
  INV_X1 U24151 ( .A(n21187), .ZN(n21190) );
  OAI211_X1 U24152 ( .C1(n21193), .C2(n21346), .A(n21349), .B(n21188), .ZN(
        n21189) );
  OAI211_X1 U24153 ( .C1(n21349), .C2(n21190), .A(n21348), .B(n21189), .ZN(
        n21211) );
  INV_X1 U24154 ( .A(n21191), .ZN(n21192) );
  AOI22_X1 U24155 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21303), .ZN(n21194) );
  OAI211_X1 U24156 ( .C1(n21306), .C2(n21214), .A(n21195), .B(n21194), .ZN(
        P1_U3121) );
  AOI22_X1 U24157 ( .A1(n21356), .A2(n21209), .B1(n21208), .B2(n21355), .ZN(
        n21197) );
  AOI22_X1 U24158 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21307), .ZN(n21196) );
  OAI211_X1 U24159 ( .C1(n21310), .C2(n21214), .A(n21197), .B(n21196), .ZN(
        P1_U3122) );
  AOI22_X1 U24160 ( .A1(n21362), .A2(n21209), .B1(n21208), .B2(n21361), .ZN(
        n21199) );
  AOI22_X1 U24161 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21311), .ZN(n21198) );
  OAI211_X1 U24162 ( .C1(n21314), .C2(n21214), .A(n21199), .B(n21198), .ZN(
        P1_U3123) );
  AOI22_X1 U24163 ( .A1(n21368), .A2(n21209), .B1(n21208), .B2(n21367), .ZN(
        n21201) );
  AOI22_X1 U24164 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21315), .ZN(n21200) );
  OAI211_X1 U24165 ( .C1(n21318), .C2(n21214), .A(n21201), .B(n21200), .ZN(
        P1_U3124) );
  AOI22_X1 U24166 ( .A1(n21374), .A2(n21209), .B1(n21208), .B2(n21373), .ZN(
        n21203) );
  AOI22_X1 U24167 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21319), .ZN(n21202) );
  OAI211_X1 U24168 ( .C1(n21322), .C2(n21214), .A(n21203), .B(n21202), .ZN(
        P1_U3125) );
  AOI22_X1 U24169 ( .A1(n21380), .A2(n21209), .B1(n21208), .B2(n21379), .ZN(
        n21205) );
  AOI22_X1 U24170 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21323), .ZN(n21204) );
  OAI211_X1 U24171 ( .C1(n21326), .C2(n21214), .A(n21205), .B(n21204), .ZN(
        P1_U3126) );
  AOI22_X1 U24172 ( .A1(n21386), .A2(n21209), .B1(n21208), .B2(n21385), .ZN(
        n21207) );
  AOI22_X1 U24173 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21387), .ZN(n21206) );
  OAI211_X1 U24174 ( .C1(n21392), .C2(n21214), .A(n21207), .B(n21206), .ZN(
        P1_U3127) );
  AOI22_X1 U24175 ( .A1(n21396), .A2(n21209), .B1(n21208), .B2(n21394), .ZN(
        n21213) );
  AOI22_X1 U24176 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n21211), .B1(
        n21210), .B2(n21331), .ZN(n21212) );
  OAI211_X1 U24177 ( .C1(n9748), .C2(n21214), .A(n21213), .B(n21212), .ZN(
        P1_U3128) );
  NAND3_X1 U24178 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n21216), .ZN(n21267) );
  NOR2_X1 U24179 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21267), .ZN(
        n21223) );
  INV_X1 U24180 ( .A(n21223), .ZN(n21255) );
  OAI22_X1 U24181 ( .A1(n21285), .A2(n21354), .B1(n21255), .B2(n21217), .ZN(
        n21218) );
  INV_X1 U24182 ( .A(n21218), .ZN(n21229) );
  NAND3_X1 U24183 ( .A1(n21262), .A2(n21349), .A3(n21285), .ZN(n21220) );
  NAND2_X1 U24184 ( .A1(n21220), .A2(n21219), .ZN(n21224) );
  OR2_X1 U24185 ( .A1(n13984), .A2(n9872), .ZN(n21265) );
  OR2_X1 U24186 ( .A1(n21265), .A2(n21292), .ZN(n21226) );
  AOI22_X1 U24187 ( .A1(n21224), .A2(n21226), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n21225), .ZN(n21221) );
  INV_X1 U24188 ( .A(n21224), .ZN(n21227) );
  AOI22_X1 U24189 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n21259), .B1(
        n21342), .B2(n21258), .ZN(n21228) );
  OAI211_X1 U24190 ( .C1(n21306), .C2(n21262), .A(n21229), .B(n21228), .ZN(
        P1_U3129) );
  OAI22_X1 U24191 ( .A1(n21285), .A2(n21360), .B1(n21230), .B2(n21255), .ZN(
        n21231) );
  INV_X1 U24192 ( .A(n21231), .ZN(n21233) );
  AOI22_X1 U24193 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n21259), .B1(
        n21355), .B2(n21258), .ZN(n21232) );
  OAI211_X1 U24194 ( .C1(n21310), .C2(n21262), .A(n21233), .B(n21232), .ZN(
        P1_U3130) );
  OAI22_X1 U24195 ( .A1(n21285), .A2(n21366), .B1(n21234), .B2(n21255), .ZN(
        n21235) );
  INV_X1 U24196 ( .A(n21235), .ZN(n21237) );
  AOI22_X1 U24197 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n21259), .B1(
        n21361), .B2(n21258), .ZN(n21236) );
  OAI211_X1 U24198 ( .C1(n21314), .C2(n21262), .A(n21237), .B(n21236), .ZN(
        P1_U3131) );
  OAI22_X1 U24199 ( .A1(n21285), .A2(n21372), .B1(n21238), .B2(n21255), .ZN(
        n21239) );
  INV_X1 U24200 ( .A(n21239), .ZN(n21241) );
  AOI22_X1 U24201 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n21259), .B1(
        n21367), .B2(n21258), .ZN(n21240) );
  OAI211_X1 U24202 ( .C1(n21318), .C2(n21262), .A(n21241), .B(n21240), .ZN(
        P1_U3132) );
  OAI22_X1 U24203 ( .A1(n21285), .A2(n21378), .B1(n21242), .B2(n21255), .ZN(
        n21243) );
  INV_X1 U24204 ( .A(n21243), .ZN(n21245) );
  AOI22_X1 U24205 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n21259), .B1(
        n21373), .B2(n21258), .ZN(n21244) );
  OAI211_X1 U24206 ( .C1(n21322), .C2(n21262), .A(n21245), .B(n21244), .ZN(
        P1_U3133) );
  OAI22_X1 U24207 ( .A1(n21285), .A2(n21384), .B1(n21246), .B2(n21255), .ZN(
        n21247) );
  INV_X1 U24208 ( .A(n21247), .ZN(n21249) );
  AOI22_X1 U24209 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n21259), .B1(
        n21379), .B2(n21258), .ZN(n21248) );
  OAI211_X1 U24210 ( .C1(n21326), .C2(n21262), .A(n21249), .B(n21248), .ZN(
        P1_U3134) );
  OAI22_X1 U24211 ( .A1(n21285), .A2(n21251), .B1(n21250), .B2(n21255), .ZN(
        n21252) );
  INV_X1 U24212 ( .A(n21252), .ZN(n21254) );
  AOI22_X1 U24213 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n21259), .B1(
        n21385), .B2(n21258), .ZN(n21253) );
  OAI211_X1 U24214 ( .C1(n21392), .C2(n21262), .A(n21254), .B(n21253), .ZN(
        P1_U3135) );
  OAI22_X1 U24215 ( .A1(n21285), .A2(n21402), .B1(n21256), .B2(n21255), .ZN(
        n21257) );
  INV_X1 U24216 ( .A(n21257), .ZN(n21261) );
  AOI22_X1 U24217 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n21259), .B1(
        n21394), .B2(n21258), .ZN(n21260) );
  OAI211_X1 U24218 ( .C1(n9748), .C2(n21262), .A(n21261), .B(n21260), .ZN(
        P1_U3136) );
  NOR2_X1 U24219 ( .A1(n21264), .A2(n21267), .ZN(n21287) );
  AOI21_X1 U24220 ( .B1(n21339), .B2(n21266), .A(n21287), .ZN(n21268) );
  OAI22_X1 U24221 ( .A1(n21268), .A2(n21341), .B1(n21267), .B2(n11005), .ZN(
        n21286) );
  AOI22_X1 U24222 ( .A1(n21343), .A2(n21287), .B1(n21342), .B2(n21286), .ZN(
        n21272) );
  INV_X1 U24223 ( .A(n21267), .ZN(n21270) );
  OAI211_X1 U24224 ( .C1(n21345), .C2(n21497), .A(n21349), .B(n21268), .ZN(
        n21269) );
  OAI211_X1 U24225 ( .C1(n21349), .C2(n21270), .A(n21348), .B(n21269), .ZN(
        n21289) );
  AOI22_X1 U24226 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21351), .ZN(n21271) );
  OAI211_X1 U24227 ( .C1(n21354), .C2(n21335), .A(n21272), .B(n21271), .ZN(
        P1_U3137) );
  AOI22_X1 U24228 ( .A1(n21356), .A2(n21287), .B1(n21355), .B2(n21286), .ZN(
        n21274) );
  AOI22_X1 U24229 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21357), .ZN(n21273) );
  OAI211_X1 U24230 ( .C1(n21360), .C2(n21335), .A(n21274), .B(n21273), .ZN(
        P1_U3138) );
  AOI22_X1 U24231 ( .A1(n21362), .A2(n21287), .B1(n21361), .B2(n21286), .ZN(
        n21276) );
  AOI22_X1 U24232 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21363), .ZN(n21275) );
  OAI211_X1 U24233 ( .C1(n21366), .C2(n21335), .A(n21276), .B(n21275), .ZN(
        P1_U3139) );
  AOI22_X1 U24234 ( .A1(n21368), .A2(n21287), .B1(n21367), .B2(n21286), .ZN(
        n21278) );
  AOI22_X1 U24235 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21369), .ZN(n21277) );
  OAI211_X1 U24236 ( .C1(n21372), .C2(n21335), .A(n21278), .B(n21277), .ZN(
        P1_U3140) );
  AOI22_X1 U24237 ( .A1(n21374), .A2(n21287), .B1(n21373), .B2(n21286), .ZN(
        n21280) );
  AOI22_X1 U24238 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21375), .ZN(n21279) );
  OAI211_X1 U24239 ( .C1(n21378), .C2(n21335), .A(n21280), .B(n21279), .ZN(
        P1_U3141) );
  AOI22_X1 U24240 ( .A1(n21380), .A2(n21287), .B1(n21379), .B2(n21286), .ZN(
        n21282) );
  AOI22_X1 U24241 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n21381), .ZN(n21281) );
  OAI211_X1 U24242 ( .C1(n21384), .C2(n21335), .A(n21282), .B(n21281), .ZN(
        P1_U3142) );
  AOI22_X1 U24243 ( .A1(n21386), .A2(n21287), .B1(n21385), .B2(n21286), .ZN(
        n21284) );
  INV_X1 U24244 ( .A(n21335), .ZN(n21297) );
  AOI22_X1 U24245 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n21289), .B1(
        n21297), .B2(n21387), .ZN(n21283) );
  OAI211_X1 U24246 ( .C1(n21392), .C2(n21285), .A(n21284), .B(n21283), .ZN(
        P1_U3143) );
  AOI22_X1 U24247 ( .A1(n21396), .A2(n21287), .B1(n21394), .B2(n21286), .ZN(
        n21291) );
  AOI22_X1 U24248 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n21289), .B1(
        n21288), .B2(n9747), .ZN(n21290) );
  OAI211_X1 U24249 ( .C1(n21402), .C2(n21335), .A(n21291), .B(n21290), .ZN(
        P1_U3144) );
  NOR2_X1 U24250 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21340), .ZN(
        n21330) );
  NAND2_X1 U24251 ( .A1(n21339), .A2(n21292), .ZN(n21298) );
  OAI22_X1 U24252 ( .A1(n21298), .A2(n21341), .B1(n21294), .B2(n21293), .ZN(
        n21329) );
  AOI22_X1 U24253 ( .A1(n21343), .A2(n21330), .B1(n21342), .B2(n21329), .ZN(
        n21305) );
  NAND2_X1 U24254 ( .A1(n21296), .A2(n21295), .ZN(n21391) );
  OAI21_X1 U24255 ( .B1(n21397), .B2(n21297), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21299) );
  AOI21_X1 U24256 ( .B1(n21299), .B2(n21298), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21302) );
  AOI22_X1 U24257 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21303), .ZN(n21304) );
  OAI211_X1 U24258 ( .C1(n21306), .C2(n21335), .A(n21305), .B(n21304), .ZN(
        P1_U3145) );
  AOI22_X1 U24259 ( .A1(n21356), .A2(n21330), .B1(n21355), .B2(n21329), .ZN(
        n21309) );
  AOI22_X1 U24260 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21307), .ZN(n21308) );
  OAI211_X1 U24261 ( .C1(n21310), .C2(n21335), .A(n21309), .B(n21308), .ZN(
        P1_U3146) );
  AOI22_X1 U24262 ( .A1(n21362), .A2(n21330), .B1(n21361), .B2(n21329), .ZN(
        n21313) );
  AOI22_X1 U24263 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21311), .ZN(n21312) );
  OAI211_X1 U24264 ( .C1(n21314), .C2(n21335), .A(n21313), .B(n21312), .ZN(
        P1_U3147) );
  AOI22_X1 U24265 ( .A1(n21368), .A2(n21330), .B1(n21367), .B2(n21329), .ZN(
        n21317) );
  AOI22_X1 U24266 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21315), .ZN(n21316) );
  OAI211_X1 U24267 ( .C1(n21318), .C2(n21335), .A(n21317), .B(n21316), .ZN(
        P1_U3148) );
  AOI22_X1 U24268 ( .A1(n21374), .A2(n21330), .B1(n21373), .B2(n21329), .ZN(
        n21321) );
  AOI22_X1 U24269 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21319), .ZN(n21320) );
  OAI211_X1 U24270 ( .C1(n21322), .C2(n21335), .A(n21321), .B(n21320), .ZN(
        P1_U3149) );
  AOI22_X1 U24271 ( .A1(n21380), .A2(n21330), .B1(n21379), .B2(n21329), .ZN(
        n21325) );
  AOI22_X1 U24272 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21323), .ZN(n21324) );
  OAI211_X1 U24273 ( .C1(n21326), .C2(n21335), .A(n21325), .B(n21324), .ZN(
        P1_U3150) );
  AOI22_X1 U24274 ( .A1(n21386), .A2(n21330), .B1(n21385), .B2(n21329), .ZN(
        n21328) );
  AOI22_X1 U24275 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21387), .ZN(n21327) );
  OAI211_X1 U24276 ( .C1(n21392), .C2(n21335), .A(n21328), .B(n21327), .ZN(
        P1_U3151) );
  AOI22_X1 U24277 ( .A1(n21396), .A2(n21330), .B1(n21394), .B2(n21329), .ZN(
        n21334) );
  AOI22_X1 U24278 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n21332), .B1(
        n21397), .B2(n21331), .ZN(n21333) );
  OAI211_X1 U24279 ( .C1(n9748), .C2(n21335), .A(n21334), .B(n21333), .ZN(
        P1_U3152) );
  INV_X1 U24280 ( .A(n21337), .ZN(n21395) );
  AOI21_X1 U24281 ( .B1(n21339), .B2(n21338), .A(n21395), .ZN(n21344) );
  OAI22_X1 U24282 ( .A1(n21344), .A2(n21341), .B1(n21340), .B2(n11005), .ZN(
        n21393) );
  AOI22_X1 U24283 ( .A1(n21343), .A2(n21395), .B1(n21342), .B2(n21393), .ZN(
        n21353) );
  OAI211_X1 U24284 ( .C1(n21346), .C2(n21345), .A(n21349), .B(n21344), .ZN(
        n21347) );
  OAI211_X1 U24285 ( .C1(n21350), .C2(n21349), .A(n21348), .B(n21347), .ZN(
        n21398) );
  AOI22_X1 U24286 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21351), .ZN(n21352) );
  OAI211_X1 U24287 ( .C1(n21354), .C2(n21401), .A(n21353), .B(n21352), .ZN(
        P1_U3153) );
  AOI22_X1 U24288 ( .A1(n21356), .A2(n21395), .B1(n21355), .B2(n21393), .ZN(
        n21359) );
  AOI22_X1 U24289 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21357), .ZN(n21358) );
  OAI211_X1 U24290 ( .C1(n21360), .C2(n21401), .A(n21359), .B(n21358), .ZN(
        P1_U3154) );
  AOI22_X1 U24291 ( .A1(n21362), .A2(n21395), .B1(n21361), .B2(n21393), .ZN(
        n21365) );
  AOI22_X1 U24292 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21363), .ZN(n21364) );
  OAI211_X1 U24293 ( .C1(n21366), .C2(n21401), .A(n21365), .B(n21364), .ZN(
        P1_U3155) );
  AOI22_X1 U24294 ( .A1(n21368), .A2(n21395), .B1(n21367), .B2(n21393), .ZN(
        n21371) );
  AOI22_X1 U24295 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21369), .ZN(n21370) );
  OAI211_X1 U24296 ( .C1(n21372), .C2(n21401), .A(n21371), .B(n21370), .ZN(
        P1_U3156) );
  AOI22_X1 U24297 ( .A1(n21374), .A2(n21395), .B1(n21373), .B2(n21393), .ZN(
        n21377) );
  AOI22_X1 U24298 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21375), .ZN(n21376) );
  OAI211_X1 U24299 ( .C1(n21378), .C2(n21401), .A(n21377), .B(n21376), .ZN(
        P1_U3157) );
  AOI22_X1 U24300 ( .A1(n21380), .A2(n21395), .B1(n21379), .B2(n21393), .ZN(
        n21383) );
  AOI22_X1 U24301 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n21381), .ZN(n21382) );
  OAI211_X1 U24302 ( .C1(n21384), .C2(n21401), .A(n21383), .B(n21382), .ZN(
        P1_U3158) );
  AOI22_X1 U24303 ( .A1(n21386), .A2(n21395), .B1(n21385), .B2(n21393), .ZN(
        n21390) );
  AOI22_X1 U24304 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n21398), .B1(
        n21388), .B2(n21387), .ZN(n21389) );
  OAI211_X1 U24305 ( .C1(n21392), .C2(n21391), .A(n21390), .B(n21389), .ZN(
        P1_U3159) );
  AOI22_X1 U24306 ( .A1(n21396), .A2(n21395), .B1(n21394), .B2(n21393), .ZN(
        n21400) );
  AOI22_X1 U24307 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n21398), .B1(
        n21397), .B2(n9747), .ZN(n21399) );
  OAI211_X1 U24308 ( .C1(n21402), .C2(n21401), .A(n21400), .B(n21399), .ZN(
        P1_U3160) );
  NOR2_X1 U24309 ( .A1(n10276), .A2(n21403), .ZN(n21406) );
  INV_X1 U24310 ( .A(n21404), .ZN(n21405) );
  OAI21_X1 U24311 ( .B1(n21406), .B2(n11005), .A(n21405), .ZN(P1_U3163) );
  INV_X1 U24312 ( .A(n21486), .ZN(n21482) );
  AND2_X1 U24313 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21482), .ZN(
        P1_U3164) );
  AND2_X1 U24314 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21482), .ZN(
        P1_U3165) );
  AND2_X1 U24315 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21482), .ZN(
        P1_U3166) );
  AND2_X1 U24316 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21482), .ZN(
        P1_U3167) );
  AND2_X1 U24317 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21482), .ZN(
        P1_U3168) );
  AND2_X1 U24318 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21482), .ZN(
        P1_U3169) );
  AND2_X1 U24319 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21407), .ZN(
        P1_U3170) );
  AND2_X1 U24320 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21407), .ZN(
        P1_U3171) );
  AND2_X1 U24321 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21407), .ZN(
        P1_U3172) );
  AND2_X1 U24322 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21407), .ZN(
        P1_U3173) );
  AND2_X1 U24323 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21407), .ZN(
        P1_U3174) );
  AND2_X1 U24324 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21407), .ZN(
        P1_U3175) );
  AND2_X1 U24325 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21407), .ZN(
        P1_U3176) );
  AND2_X1 U24326 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21407), .ZN(
        P1_U3177) );
  AND2_X1 U24327 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21407), .ZN(
        P1_U3178) );
  AND2_X1 U24328 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21482), .ZN(
        P1_U3179) );
  INV_X1 U24329 ( .A(P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n21611) );
  NOR2_X1 U24330 ( .A1(n21486), .A2(n21611), .ZN(P1_U3180) );
  AND2_X1 U24331 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21482), .ZN(
        P1_U3181) );
  AND2_X1 U24332 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21482), .ZN(
        P1_U3182) );
  AND2_X1 U24333 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21482), .ZN(
        P1_U3183) );
  AND2_X1 U24334 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21482), .ZN(
        P1_U3184) );
  AND2_X1 U24335 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21482), .ZN(
        P1_U3185) );
  AND2_X1 U24336 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21482), .ZN(P1_U3186) );
  AND2_X1 U24337 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21482), .ZN(P1_U3187) );
  AND2_X1 U24338 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21482), .ZN(P1_U3188) );
  AND2_X1 U24339 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21482), .ZN(P1_U3189) );
  AND2_X1 U24340 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21482), .ZN(P1_U3190) );
  AND2_X1 U24341 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21482), .ZN(P1_U3191) );
  AND2_X1 U24342 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21482), .ZN(P1_U3192) );
  AND2_X1 U24343 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21482), .ZN(P1_U3193) );
  INV_X1 U24344 ( .A(n21418), .ZN(n21413) );
  INV_X1 U24345 ( .A(n21408), .ZN(n21412) );
  OAI21_X1 U24346 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n21416), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21410) );
  OR2_X1 U24347 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21409) );
  OAI221_X1 U24348 ( .B1(n21410), .B2(HOLD), .C1(n21410), .C2(n21409), .A(
        n21495), .ZN(n21411) );
  OAI211_X1 U24349 ( .C1(n21413), .C2(n21419), .A(n21412), .B(n21411), .ZN(
        P1_U3194) );
  AOI221_X1 U24350 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n21415), .C1(n21416), 
        .C2(n21415), .A(n21414), .ZN(n21425) );
  AOI21_X1 U24351 ( .B1(n21417), .B2(n21416), .A(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n21424) );
  OAI21_X1 U24352 ( .B1(NA), .B2(n21419), .A(n21418), .ZN(n21420) );
  OAI211_X1 U24353 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21421), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n21420), .ZN(n21422) );
  OAI22_X1 U24354 ( .A1(n21425), .A2(n21424), .B1(n21423), .B2(n21422), .ZN(
        P1_U3196) );
  NOR2_X1 U24355 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21495), .ZN(n21474) );
  AOI22_X1 U24356 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21474), .ZN(n21426) );
  OAI21_X1 U24357 ( .B1(n21487), .B2(n21472), .A(n21426), .ZN(P1_U3197) );
  INV_X1 U24358 ( .A(n21472), .ZN(n21475) );
  AOI22_X1 U24359 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n21475), .ZN(n21427) );
  OAI21_X1 U24360 ( .B1(n14493), .B2(n21468), .A(n21427), .ZN(P1_U3198) );
  OAI222_X1 U24361 ( .A1(n21472), .A2(n14493), .B1(n21428), .B2(n21511), .C1(
        n21429), .C2(n21468), .ZN(P1_U3199) );
  INV_X1 U24362 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n21631) );
  OAI222_X1 U24363 ( .A1(n21472), .A2(n21429), .B1(n21631), .B2(n21511), .C1(
        n21431), .C2(n21468), .ZN(P1_U3200) );
  INV_X1 U24364 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n21430) );
  OAI222_X1 U24365 ( .A1(n21472), .A2(n21431), .B1(n21430), .B2(n21511), .C1(
        n21433), .C2(n21468), .ZN(P1_U3201) );
  INV_X1 U24366 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n21432) );
  OAI222_X1 U24367 ( .A1(n21472), .A2(n21433), .B1(n21432), .B2(n21511), .C1(
        n21435), .C2(n21468), .ZN(P1_U3202) );
  INV_X1 U24368 ( .A(P1_ADDRESS_REG_6__SCAN_IN), .ZN(n21434) );
  OAI222_X1 U24369 ( .A1(n21472), .A2(n21435), .B1(n21434), .B2(n21511), .C1(
        n21436), .C2(n21468), .ZN(P1_U3203) );
  INV_X1 U24370 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21437) );
  OAI222_X1 U24371 ( .A1(n21468), .A2(n21439), .B1(n21437), .B2(n21511), .C1(
        n21436), .C2(n21472), .ZN(P1_U3204) );
  AOI22_X1 U24372 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21474), .ZN(n21438) );
  OAI21_X1 U24373 ( .B1(n21439), .B2(n21472), .A(n21438), .ZN(P1_U3205) );
  AOI22_X1 U24374 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n21475), .ZN(n21440) );
  OAI21_X1 U24375 ( .B1(n15336), .B2(n21468), .A(n21440), .ZN(P1_U3206) );
  AOI222_X1 U24376 ( .A1(n21475), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n21495), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n21474), .ZN(n21441) );
  INV_X1 U24377 ( .A(n21441), .ZN(P1_U3207) );
  AOI222_X1 U24378 ( .A1(n21475), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n21495), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n21474), .ZN(n21442) );
  INV_X1 U24379 ( .A(n21442), .ZN(P1_U3208) );
  AOI22_X1 U24380 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21474), .ZN(n21443) );
  OAI21_X1 U24381 ( .B1(n21444), .B2(n21472), .A(n21443), .ZN(P1_U3209) );
  AOI22_X1 U24382 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21475), .ZN(n21445) );
  OAI21_X1 U24383 ( .B1(n21447), .B2(n21468), .A(n21445), .ZN(P1_U3210) );
  AOI22_X1 U24384 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n21474), .ZN(n21446) );
  OAI21_X1 U24385 ( .B1(n21447), .B2(n21472), .A(n21446), .ZN(P1_U3211) );
  AOI22_X1 U24386 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21474), .ZN(n21448) );
  OAI21_X1 U24387 ( .B1(n15290), .B2(n21472), .A(n21448), .ZN(P1_U3212) );
  AOI22_X1 U24388 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21475), .ZN(n21449) );
  OAI21_X1 U24389 ( .B1(n21451), .B2(n21468), .A(n21449), .ZN(P1_U3213) );
  AOI22_X1 U24390 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21474), .ZN(n21450) );
  OAI21_X1 U24391 ( .B1(n21451), .B2(n21472), .A(n21450), .ZN(P1_U3214) );
  AOI22_X1 U24392 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n21475), .ZN(n21452) );
  OAI21_X1 U24393 ( .B1(n21454), .B2(n21468), .A(n21452), .ZN(P1_U3215) );
  INV_X1 U24394 ( .A(P1_ADDRESS_REG_19__SCAN_IN), .ZN(n21453) );
  OAI222_X1 U24395 ( .A1(n21472), .A2(n21454), .B1(n21453), .B2(n21511), .C1(
        n21456), .C2(n21468), .ZN(P1_U3216) );
  INV_X1 U24396 ( .A(P1_ADDRESS_REG_20__SCAN_IN), .ZN(n21455) );
  OAI222_X1 U24397 ( .A1(n21472), .A2(n21456), .B1(n21455), .B2(n21511), .C1(
        n21458), .C2(n21468), .ZN(P1_U3217) );
  AOI22_X1 U24398 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21474), .ZN(n21457) );
  OAI21_X1 U24399 ( .B1(n21458), .B2(n21472), .A(n21457), .ZN(P1_U3218) );
  AOI22_X1 U24400 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n21495), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n21475), .ZN(n21459) );
  OAI21_X1 U24401 ( .B1(n21461), .B2(n21468), .A(n21459), .ZN(P1_U3219) );
  INV_X1 U24402 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n21460) );
  OAI222_X1 U24403 ( .A1(n21472), .A2(n21461), .B1(n21460), .B2(n21511), .C1(
        n21462), .C2(n21468), .ZN(P1_U3220) );
  INV_X1 U24404 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n21463) );
  OAI222_X1 U24405 ( .A1(n21468), .A2(n21465), .B1(n21463), .B2(n21511), .C1(
        n21462), .C2(n21472), .ZN(P1_U3221) );
  INV_X1 U24406 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n21464) );
  OAI222_X1 U24407 ( .A1(n21472), .A2(n21465), .B1(n21464), .B2(n21511), .C1(
        n21467), .C2(n21468), .ZN(P1_U3222) );
  INV_X1 U24408 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n21466) );
  OAI222_X1 U24409 ( .A1(n21472), .A2(n21467), .B1(n21466), .B2(n21511), .C1(
        n21471), .C2(n21468), .ZN(P1_U3223) );
  INV_X1 U24410 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n21470) );
  OAI222_X1 U24411 ( .A1(n21472), .A2(n21471), .B1(n21470), .B2(n21511), .C1(
        n21469), .C2(n21468), .ZN(P1_U3224) );
  AOI222_X1 U24412 ( .A1(n21474), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21495), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n21475), .ZN(n21473) );
  INV_X1 U24413 ( .A(n21473), .ZN(P1_U3225) );
  AOI222_X1 U24414 ( .A1(n21475), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21495), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n21474), .ZN(n21476) );
  INV_X1 U24415 ( .A(n21476), .ZN(P1_U3226) );
  INV_X1 U24416 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n21563) );
  AOI22_X1 U24417 ( .A1(n21511), .A2(n21649), .B1(n21563), .B2(n21495), .ZN(
        P1_U3458) );
  INV_X1 U24418 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21490) );
  INV_X1 U24419 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n21477) );
  AOI22_X1 U24420 ( .A1(n21511), .A2(n21490), .B1(n21477), .B2(n21495), .ZN(
        P1_U3459) );
  INV_X1 U24421 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n21478) );
  AOI22_X1 U24422 ( .A1(n21511), .A2(n21479), .B1(n21478), .B2(n21495), .ZN(
        P1_U3460) );
  INV_X1 U24423 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21493) );
  INV_X1 U24424 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n21480) );
  AOI22_X1 U24425 ( .A1(n21511), .A2(n21493), .B1(n21480), .B2(n21495), .ZN(
        P1_U3461) );
  INV_X1 U24426 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21483) );
  INV_X1 U24427 ( .A(n21484), .ZN(n21481) );
  AOI21_X1 U24428 ( .B1(n21483), .B2(n21482), .A(n21481), .ZN(P1_U3464) );
  OAI21_X1 U24429 ( .B1(n21486), .B2(n21485), .A(n21484), .ZN(P1_U3465) );
  AOI21_X1 U24430 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n21488) );
  AOI22_X1 U24431 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n21488), .B2(n21487), .ZN(n21491) );
  AOI22_X1 U24432 ( .A1(n21494), .A2(n21491), .B1(n21490), .B2(n21489), .ZN(
        P1_U3481) );
  OAI21_X1 U24433 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n21494), .ZN(n21492) );
  OAI21_X1 U24434 ( .B1(n21494), .B2(n21493), .A(n21492), .ZN(P1_U3482) );
  AOI22_X1 U24435 ( .A1(n21511), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21496), 
        .B2(n21495), .ZN(P1_U3483) );
  OAI22_X1 U24436 ( .A1(n21500), .A2(n21499), .B1(n21498), .B2(n21497), .ZN(
        n21502) );
  NOR2_X1 U24437 ( .A1(n21501), .A2(n11005), .ZN(n21507) );
  AND2_X1 U24438 ( .A1(n21502), .A2(n21507), .ZN(n21504) );
  OAI21_X1 U24439 ( .B1(n21504), .B2(n10276), .A(n21503), .ZN(n21510) );
  AOI211_X1 U24440 ( .C1(n21508), .C2(n21507), .A(n21506), .B(n21505), .ZN(
        n21509) );
  MUX2_X1 U24441 ( .A(n21510), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21509), 
        .Z(P1_U3485) );
  MUX2_X1 U24442 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(P1_MEMORYFETCH_REG_SCAN_IN), 
        .S(n21511), .Z(P1_U3486) );
  NAND4_X1 U24443 ( .A1(P1_BE_N_REG_3__SCAN_IN), .A2(n21566), .A3(n15142), 
        .A4(n21551), .ZN(n21521) );
  NAND4_X1 U24444 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(P3_DATAO_REG_25__SCAN_IN), 
        .A3(n21565), .A4(n21572), .ZN(n21520) );
  NOR4_X1 U24445 ( .A1(BUF2_REG_30__SCAN_IN), .A2(P1_EAX_REG_21__SCAN_IN), 
        .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(n21571), .ZN(n21513) );
  NOR2_X1 U24446 ( .A1(BUF1_REG_7__SCAN_IN), .A2(P2_LWORD_REG_14__SCAN_IN), 
        .ZN(n21512) );
  NAND4_X1 U24447 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n21513), .A3(
        P3_ADDRESS_REG_29__SCAN_IN), .A4(n21512), .ZN(n21519) );
  NOR4_X1 U24448 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(
        P3_DATAO_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        n21644), .ZN(n21517) );
  INV_X1 U24449 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n21650) );
  NOR4_X1 U24450 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n21650), .A3(n21647), .A4(
        n21649), .ZN(n21516) );
  NOR4_X1 U24451 ( .A1(P1_ADDRESS_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n21625), .A4(n21630), .ZN(
        n21515) );
  NOR4_X1 U24452 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(
        P2_EAX_REG_18__SCAN_IN), .A3(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A4(
        n21628), .ZN(n21514) );
  NAND4_X1 U24453 ( .A1(n21517), .A2(n21516), .A3(n21515), .A4(n21514), .ZN(
        n21518) );
  NOR4_X1 U24454 ( .A1(n21521), .A2(n21520), .A3(n21519), .A4(n21518), .ZN(
        n21662) );
  NOR4_X1 U24455 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__3__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), 
        .A4(n21612), .ZN(n21532) );
  INV_X1 U24456 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n21598) );
  NOR4_X1 U24457 ( .A1(P2_UWORD_REG_9__SCAN_IN), .A2(P3_LWORD_REG_0__SCAN_IN), 
        .A3(n21598), .A4(n16031), .ZN(n21531) );
  NOR4_X1 U24458 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_26__SCAN_IN), .A3(n21618), .A4(n21615), .ZN(n21530)
         );
  NOR4_X1 U24459 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        BUF2_REG_10__SCAN_IN), .A3(P1_UWORD_REG_2__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21522) );
  NAND4_X1 U24460 ( .A1(DATAI_27_), .A2(P2_DATAWIDTH_REG_14__SCAN_IN), .A3(
        n21523), .A4(n21522), .ZN(n21528) );
  AND4_X1 U24461 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_1__5__SCAN_IN), .A3(P1_EAX_REG_23__SCAN_IN), .A4(
        n21554), .ZN(n21524) );
  NAND4_X1 U24462 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n21549), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A4(n21524), .ZN(n21525) );
  NOR3_X1 U24463 ( .A1(n21525), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_14__SCAN_IN), .ZN(n21526) );
  NAND4_X1 U24464 ( .A1(n21526), .A2(n21552), .A3(P3_REIP_REG_22__SCAN_IN), 
        .A4(BUF1_REG_10__SCAN_IN), .ZN(n21527) );
  NOR2_X1 U24465 ( .A1(n21528), .A2(n21527), .ZN(n21529) );
  AND4_X1 U24466 ( .A1(n21532), .A2(n21531), .A3(n21530), .A4(n21529), .ZN(
        n21661) );
  AOI22_X1 U24467 ( .A1(n15126), .A2(keyinput27), .B1(keyinput61), .B2(n21534), 
        .ZN(n21533) );
  OAI221_X1 U24468 ( .B1(n15126), .B2(keyinput27), .C1(n21534), .C2(keyinput61), .A(n21533), .ZN(n21546) );
  INV_X1 U24469 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n21537) );
  AOI22_X1 U24470 ( .A1(n21537), .A2(keyinput29), .B1(n21536), .B2(keyinput16), 
        .ZN(n21535) );
  OAI221_X1 U24471 ( .B1(n21537), .B2(keyinput29), .C1(n21536), .C2(keyinput16), .A(n21535), .ZN(n21545) );
  AOI22_X1 U24472 ( .A1(n21540), .A2(keyinput31), .B1(n21539), .B2(keyinput34), 
        .ZN(n21538) );
  OAI221_X1 U24473 ( .B1(n21540), .B2(keyinput31), .C1(n21539), .C2(keyinput34), .A(n21538), .ZN(n21544) );
  AOI22_X1 U24474 ( .A1(n21542), .A2(keyinput52), .B1(n10557), .B2(keyinput33), 
        .ZN(n21541) );
  OAI221_X1 U24475 ( .B1(n21542), .B2(keyinput52), .C1(n10557), .C2(keyinput33), .A(n21541), .ZN(n21543) );
  NOR4_X1 U24476 ( .A1(n21546), .A2(n21545), .A3(n21544), .A4(n21543), .ZN(
        n21594) );
  AOI22_X1 U24477 ( .A1(n21549), .A2(keyinput41), .B1(keyinput59), .B2(n21548), 
        .ZN(n21547) );
  OAI221_X1 U24478 ( .B1(n21549), .B2(keyinput41), .C1(n21548), .C2(keyinput59), .A(n21547), .ZN(n21561) );
  AOI22_X1 U24479 ( .A1(n21552), .A2(keyinput18), .B1(n21551), .B2(keyinput45), 
        .ZN(n21550) );
  OAI221_X1 U24480 ( .B1(n21552), .B2(keyinput18), .C1(n21551), .C2(keyinput45), .A(n21550), .ZN(n21560) );
  AOI22_X1 U24481 ( .A1(n11415), .A2(keyinput28), .B1(n21554), .B2(keyinput21), 
        .ZN(n21553) );
  OAI221_X1 U24482 ( .B1(n11415), .B2(keyinput28), .C1(n21554), .C2(keyinput21), .A(n21553), .ZN(n21559) );
  XOR2_X1 U24483 ( .A(n21555), .B(keyinput24), .Z(n21557) );
  XNOR2_X1 U24484 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B(keyinput38), 
        .ZN(n21556) );
  NAND2_X1 U24485 ( .A1(n21557), .A2(n21556), .ZN(n21558) );
  NOR4_X1 U24486 ( .A1(n21561), .A2(n21560), .A3(n21559), .A4(n21558), .ZN(
        n21593) );
  AOI22_X1 U24487 ( .A1(n21563), .A2(keyinput13), .B1(n15142), .B2(keyinput50), 
        .ZN(n21562) );
  OAI221_X1 U24488 ( .B1(n21563), .B2(keyinput13), .C1(n15142), .C2(keyinput50), .A(n21562), .ZN(n21576) );
  AOI22_X1 U24489 ( .A1(n21566), .A2(keyinput56), .B1(keyinput44), .B2(n21565), 
        .ZN(n21564) );
  OAI221_X1 U24490 ( .B1(n21566), .B2(keyinput56), .C1(n21565), .C2(keyinput44), .A(n21564), .ZN(n21575) );
  INV_X1 U24491 ( .A(P1_EAX_REG_31__SCAN_IN), .ZN(n21569) );
  INV_X1 U24492 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n21568) );
  AOI22_X1 U24493 ( .A1(n21569), .A2(keyinput32), .B1(keyinput1), .B2(n21568), 
        .ZN(n21567) );
  OAI221_X1 U24494 ( .B1(n21569), .B2(keyinput32), .C1(n21568), .C2(keyinput1), 
        .A(n21567), .ZN(n21574) );
  AOI22_X1 U24495 ( .A1(n21572), .A2(keyinput12), .B1(keyinput4), .B2(n21571), 
        .ZN(n21570) );
  OAI221_X1 U24496 ( .B1(n21572), .B2(keyinput12), .C1(n21571), .C2(keyinput4), 
        .A(n21570), .ZN(n21573) );
  NOR4_X1 U24497 ( .A1(n21576), .A2(n21575), .A3(n21574), .A4(n21573), .ZN(
        n21592) );
  AOI22_X1 U24498 ( .A1(n15155), .A2(keyinput62), .B1(n14609), .B2(keyinput39), 
        .ZN(n21577) );
  OAI221_X1 U24499 ( .B1(n15155), .B2(keyinput62), .C1(n14609), .C2(keyinput39), .A(n21577), .ZN(n21590) );
  INV_X1 U24500 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n21579) );
  AOI22_X1 U24501 ( .A1(n21580), .A2(keyinput49), .B1(n21579), .B2(keyinput23), 
        .ZN(n21578) );
  OAI221_X1 U24502 ( .B1(n21580), .B2(keyinput49), .C1(n21579), .C2(keyinput23), .A(n21578), .ZN(n21589) );
  AOI22_X1 U24503 ( .A1(n21583), .A2(keyinput36), .B1(keyinput17), .B2(n21582), 
        .ZN(n21581) );
  OAI221_X1 U24504 ( .B1(n21583), .B2(keyinput36), .C1(n21582), .C2(keyinput17), .A(n21581), .ZN(n21588) );
  INV_X1 U24505 ( .A(P3_EAX_REG_31__SCAN_IN), .ZN(n21586) );
  AOI22_X1 U24506 ( .A1(n21586), .A2(keyinput53), .B1(n21585), .B2(keyinput8), 
        .ZN(n21584) );
  OAI221_X1 U24507 ( .B1(n21586), .B2(keyinput53), .C1(n21585), .C2(keyinput8), 
        .A(n21584), .ZN(n21587) );
  NOR4_X1 U24508 ( .A1(n21590), .A2(n21589), .A3(n21588), .A4(n21587), .ZN(
        n21591) );
  NAND4_X1 U24509 ( .A1(n21594), .A2(n21593), .A3(n21592), .A4(n21591), .ZN(
        n21660) );
  AOI22_X1 U24510 ( .A1(n21596), .A2(keyinput15), .B1(n17237), .B2(keyinput37), 
        .ZN(n21595) );
  OAI221_X1 U24511 ( .B1(n21596), .B2(keyinput15), .C1(n17237), .C2(keyinput37), .A(n21595), .ZN(n21607) );
  INV_X1 U24512 ( .A(P3_LWORD_REG_0__SCAN_IN), .ZN(n21599) );
  AOI22_X1 U24513 ( .A1(n21599), .A2(keyinput6), .B1(n21598), .B2(keyinput43), 
        .ZN(n21597) );
  OAI221_X1 U24514 ( .B1(n21599), .B2(keyinput6), .C1(n21598), .C2(keyinput43), 
        .A(n21597), .ZN(n21606) );
  INV_X1 U24515 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n21601) );
  AOI22_X1 U24516 ( .A1(n16031), .A2(keyinput30), .B1(keyinput48), .B2(n21601), 
        .ZN(n21600) );
  OAI221_X1 U24517 ( .B1(n16031), .B2(keyinput30), .C1(n21601), .C2(keyinput48), .A(n21600), .ZN(n21605) );
  XOR2_X1 U24518 ( .A(n12697), .B(keyinput35), .Z(n21603) );
  XNOR2_X1 U24519 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput26), .ZN(
        n21602) );
  NAND2_X1 U24520 ( .A1(n21603), .A2(n21602), .ZN(n21604) );
  NOR4_X1 U24521 ( .A1(n21607), .A2(n21606), .A3(n21605), .A4(n21604), .ZN(
        n21658) );
  AOI22_X1 U24522 ( .A1(n21609), .A2(keyinput7), .B1(n11024), .B2(keyinput25), 
        .ZN(n21608) );
  OAI221_X1 U24523 ( .B1(n21609), .B2(keyinput7), .C1(n11024), .C2(keyinput25), 
        .A(n21608), .ZN(n21622) );
  AOI22_X1 U24524 ( .A1(n21612), .A2(keyinput20), .B1(keyinput46), .B2(n21611), 
        .ZN(n21610) );
  OAI221_X1 U24525 ( .B1(n21612), .B2(keyinput20), .C1(n21611), .C2(keyinput46), .A(n21610), .ZN(n21621) );
  AOI22_X1 U24526 ( .A1(n21615), .A2(keyinput60), .B1(keyinput5), .B2(n21614), 
        .ZN(n21613) );
  OAI221_X1 U24527 ( .B1(n21615), .B2(keyinput60), .C1(n21614), .C2(keyinput5), 
        .A(n21613), .ZN(n21620) );
  AOI22_X1 U24528 ( .A1(n21618), .A2(keyinput51), .B1(keyinput10), .B2(n21617), 
        .ZN(n21616) );
  OAI221_X1 U24529 ( .B1(n21618), .B2(keyinput51), .C1(n21617), .C2(keyinput10), .A(n21616), .ZN(n21619) );
  NOR4_X1 U24530 ( .A1(n21622), .A2(n21621), .A3(n21620), .A4(n21619), .ZN(
        n21657) );
  AOI22_X1 U24531 ( .A1(n21625), .A2(keyinput58), .B1(keyinput3), .B2(n21624), 
        .ZN(n21623) );
  OAI221_X1 U24532 ( .B1(n21625), .B2(keyinput58), .C1(n21624), .C2(keyinput3), 
        .A(n21623), .ZN(n21638) );
  INV_X1 U24533 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21627) );
  AOI22_X1 U24534 ( .A1(n21628), .A2(keyinput55), .B1(n21627), .B2(keyinput40), 
        .ZN(n21626) );
  OAI221_X1 U24535 ( .B1(n21628), .B2(keyinput55), .C1(n21627), .C2(keyinput40), .A(n21626), .ZN(n21637) );
  AOI22_X1 U24536 ( .A1(n21631), .A2(keyinput0), .B1(n21630), .B2(keyinput2), 
        .ZN(n21629) );
  OAI221_X1 U24537 ( .B1(n21631), .B2(keyinput0), .C1(n21630), .C2(keyinput2), 
        .A(n21629), .ZN(n21636) );
  XOR2_X1 U24538 ( .A(n21632), .B(keyinput19), .Z(n21634) );
  XNOR2_X1 U24539 ( .A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B(keyinput63), .ZN(
        n21633) );
  NAND2_X1 U24540 ( .A1(n21634), .A2(n21633), .ZN(n21635) );
  NOR4_X1 U24541 ( .A1(n21638), .A2(n21637), .A3(n21636), .A4(n21635), .ZN(
        n21656) );
  AOI22_X1 U24542 ( .A1(n21641), .A2(keyinput14), .B1(keyinput57), .B2(n21640), 
        .ZN(n21639) );
  OAI221_X1 U24543 ( .B1(n21641), .B2(keyinput14), .C1(n21640), .C2(keyinput57), .A(n21639), .ZN(n21654) );
  INV_X1 U24544 ( .A(P3_DATAO_REG_20__SCAN_IN), .ZN(n21643) );
  AOI22_X1 U24545 ( .A1(n21644), .A2(keyinput22), .B1(keyinput9), .B2(n21643), 
        .ZN(n21642) );
  OAI221_X1 U24546 ( .B1(n21644), .B2(keyinput22), .C1(n21643), .C2(keyinput9), 
        .A(n21642), .ZN(n21653) );
  AOI22_X1 U24547 ( .A1(n21647), .A2(keyinput54), .B1(keyinput11), .B2(n21646), 
        .ZN(n21645) );
  OAI221_X1 U24548 ( .B1(n21647), .B2(keyinput54), .C1(n21646), .C2(keyinput11), .A(n21645), .ZN(n21652) );
  AOI22_X1 U24549 ( .A1(n21650), .A2(keyinput42), .B1(keyinput47), .B2(n21649), 
        .ZN(n21648) );
  OAI221_X1 U24550 ( .B1(n21650), .B2(keyinput42), .C1(n21649), .C2(keyinput47), .A(n21648), .ZN(n21651) );
  NOR4_X1 U24551 ( .A1(n21654), .A2(n21653), .A3(n21652), .A4(n21651), .ZN(
        n21655) );
  NAND4_X1 U24552 ( .A1(n21658), .A2(n21657), .A3(n21656), .A4(n21655), .ZN(
        n21659) );
  AOI211_X1 U24553 ( .C1(n21662), .C2(n21661), .A(n21660), .B(n21659), .ZN(
        n21676) );
  AOI22_X1 U24554 ( .A1(n21666), .A2(n21665), .B1(n21664), .B2(n21663), .ZN(
        n21667) );
  INV_X1 U24555 ( .A(n21667), .ZN(n21673) );
  OAI22_X1 U24556 ( .A1(n21671), .A2(n21670), .B1(n21669), .B2(n21668), .ZN(
        n21672) );
  AOI211_X1 U24557 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n21674), .A(
        n21673), .B(n21672), .ZN(n21675) );
  XNOR2_X1 U24558 ( .A(n21676), .B(n21675), .ZN(P3_U2891) );
  NOR2_X2 U13063 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10136) );
  CLKBUF_X1 U11093 ( .A(n12932), .Z(n12951) );
  AND2_X1 U12159 ( .A1(n9761), .A2(n13580), .ZN(n13663) );
  CLKBUF_X2 U12544 ( .A(n18046), .Z(n9570) );
  CLKBUF_X1 U12545 ( .A(n19565), .Z(n18374) );
  CLKBUF_X1 U12965 ( .A(n18417), .Z(n18424) );
endmodule

