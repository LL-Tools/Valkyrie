

module b15_C_gen_AntiSAT_k_256_9 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3445, U3446, U3447, U3448, U3213, U3212, 
        U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, U3203, U3202, 
        U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, U3193, U3192, 
        U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, U3183, U3182, 
        U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, U3175, U3174, 
        U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, U3165, U3164, 
        U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, U3155, U3154, 
        U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, U3146, U3145, 
        U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, U3136, U3135, 
        U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, U3126, U3125, 
        U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, U3116, U3115, 
        U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, U3106, U3105, 
        U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, U3096, U3095, 
        U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, U3086, U3085, 
        U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, U3076, U3075, 
        U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, U3066, U3065, 
        U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, U3056, U3055, 
        U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, U3046, U3045, 
        U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, U3036, U3035, 
        U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, U3026, U3025, 
        U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, U3460, U3461, 
        U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, U3015, U3014, 
        U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, U3005, U3004, 
        U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, U2995, U2994, 
        U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, U2985, U2984, 
        U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, U2975, U2974, 
        U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, U2965, U2964, 
        U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, U2955, U2954, 
        U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, U2945, U2944, 
        U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, U2935, U2934, 
        U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, U2925, U2924, 
        U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, U2915, U2914, 
        U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, U2905, U2904, 
        U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, U2895, U2894, 
        U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, U2885, U2884, 
        U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, U2875, U2874, 
        U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, U2865, U2864, 
        U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, U2855, U2854, 
        U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, U2845, U2844, 
        U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, U2835, U2834, 
        U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, U2825, U2824, 
        U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, U2815, U2814, 
        U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, U2805, U2804, 
        U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, U2795, U3468, 
        U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, U3473, U2790, 
        U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput_f0, keyinput_f1,
         keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6,
         keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11,
         keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16,
         keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21,
         keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26,
         keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31,
         keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36,
         keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41,
         keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46,
         keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51,
         keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56,
         keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61,
         keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66,
         keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71,
         keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76,
         keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81,
         keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86,
         keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91,
         keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96,
         keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131;

  AND2_X1 U3601 ( .A1(n5636), .A2(n3233), .ZN(n5573) );
  INV_X4 U3602 ( .A(n5944), .ZN(n6356) );
  CLKBUF_X1 U3605 ( .A(n3386), .Z(n4058) );
  BUF_X2 U3606 ( .A(n3500), .Z(n4202) );
  CLKBUF_X2 U3607 ( .A(n3471), .Z(n4235) );
  CLKBUF_X2 U3608 ( .A(n3350), .Z(n4237) );
  INV_X2 U3609 ( .A(n4287), .ZN(n3446) );
  NAND2_X1 U3610 ( .A1(n3413), .A2(n3373), .ZN(n3422) );
  INV_X1 U3611 ( .A(n3373), .ZN(n3384) );
  CLKBUF_X2 U3612 ( .A(n4719), .Z(n3172) );
  CLKBUF_X2 U3613 ( .A(n4120), .Z(n3170) );
  BUF_X2 U3614 ( .A(n3363), .Z(n3167) );
  INV_X4 U3615 ( .A(n3400), .ZN(n4125) );
  AND2_X1 U3616 ( .A1(n3289), .A2(n3290), .ZN(n3173) );
  CLKBUF_X3 U3617 ( .A(n4120), .Z(n3171) );
  INV_X1 U3618 ( .A(n3383), .ZN(n3711) );
  AND2_X1 U3619 ( .A1(n3791), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4714)
         );
  AND4_X1 U3620 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  NAND2_X1 U3621 ( .A1(n3768), .A2(n3446), .ZN(n3717) );
  NAND2_X1 U3622 ( .A1(n5410), .A2(n5411), .ZN(n3684) );
  CLKBUF_X3 U3623 ( .A(n4719), .Z(n3155) );
  NOR2_X1 U3624 ( .A1(n4434), .A2(n4437), .ZN(n5802) );
  AOI221_X1 U3625 ( .B1(REIP_REG_23__SCAN_IN), .B2(n6075), .C1(n6074), .C2(
        n6075), .A(n6073), .ZN(n6076) );
  INV_X1 U3626 ( .A(n6294), .ZN(n6279) );
  NAND2_X2 U3627 ( .A1(n3253), .A2(n3252), .ZN(n5410) );
  NOR2_X2 U3628 ( .A1(n6382), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3564)
         );
  NAND2_X2 U3629 ( .A1(n3563), .A2(n3562), .ZN(n6382) );
  NOR2_X1 U3630 ( .A1(n5793), .A2(n5775), .ZN(n5787) );
  NAND2_X2 U3631 ( .A1(n3370), .A2(n3369), .ZN(n3432) );
  NAND2_X2 U3632 ( .A1(n3384), .A2(n3417), .ZN(n4285) );
  NAND2_X4 U3633 ( .A1(n3296), .A2(n3295), .ZN(n3417) );
  BUF_X1 U3634 ( .A(n3391), .Z(n3153) );
  BUF_X4 U3635 ( .A(n3391), .Z(n3154) );
  OR2_X2 U3636 ( .A1(n5546), .A2(n4502), .ZN(n6072) );
  CLKBUF_X3 U3637 ( .A(n4719), .Z(n3156) );
  NOR2_X4 U3638 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3290) );
  CLKBUF_X1 U3639 ( .A(n4218), .Z(n5519) );
  NAND2_X1 U3640 ( .A1(n5585), .A2(n5680), .ZN(n5570) );
  CLKBUF_X2 U3641 ( .A(n3775), .Z(n4747) );
  INV_X1 U3642 ( .A(n4899), .ZN(n3230) );
  NAND2_X1 U3643 ( .A1(n3485), .A2(n3486), .ZN(n3530) );
  CLKBUF_X1 U3644 ( .A(n3463), .Z(n3161) );
  NAND2_X1 U3645 ( .A1(n4403), .A2(n3446), .ZN(n4739) );
  AND2_X2 U3646 ( .A1(n4295), .A2(n4560), .ZN(n4378) );
  INV_X4 U3647 ( .A(n4324), .ZN(n4295) );
  BUF_X1 U3648 ( .A(n3537), .Z(n3164) );
  BUF_X1 U3649 ( .A(n3413), .Z(n3773) );
  AND2_X1 U3650 ( .A1(n3714), .A2(n3383), .ZN(n3709) );
  INV_X1 U3651 ( .A(n3417), .ZN(n3413) );
  BUF_X1 U3652 ( .A(n4287), .Z(n4801) );
  INV_X2 U3653 ( .A(n4286), .ZN(n3768) );
  BUF_X2 U3655 ( .A(n3332), .Z(n3158) );
  CLKBUF_X2 U3656 ( .A(n3173), .Z(n3174) );
  AND2_X2 U3657 ( .A1(n4714), .A2(n3288), .ZN(n3363) );
  AND2_X2 U3658 ( .A1(n4715), .A2(n3289), .ZN(n3332) );
  AND2_X1 U3659 ( .A1(n4714), .A2(n4582), .ZN(n4719) );
  BUF_X2 U3660 ( .A(n3345), .Z(n4242) );
  NAND2_X2 U3661 ( .A1(n4582), .A2(n4733), .ZN(n3400) );
  AND2_X2 U3662 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4582) );
  INV_X2 U3663 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4728) );
  NOR2_X1 U3665 ( .A1(n5794), .A2(n5795), .ZN(n5793) );
  OR2_X1 U3666 ( .A1(n5519), .A2(n4219), .ZN(n4220) );
  NOR2_X1 U3667 ( .A1(n4262), .A2(n4274), .ZN(n4266) );
  NAND2_X1 U3668 ( .A1(n4218), .A2(n4219), .ZN(n4262) );
  CLKBUF_X1 U3669 ( .A(n5544), .Z(n5670) );
  CLKBUF_X1 U3670 ( .A(n4500), .Z(n5546) );
  CLKBUF_X1 U3671 ( .A(n5585), .Z(n5586) );
  NAND2_X2 U3672 ( .A1(n5734), .A2(n3921), .ZN(n5705) );
  AND2_X1 U3673 ( .A1(n4393), .A2(n4392), .ZN(n4394) );
  INV_X1 U3674 ( .A(n4423), .ZN(n3228) );
  NOR2_X1 U3675 ( .A1(n3691), .A2(n3210), .ZN(n3209) );
  NOR2_X1 U3676 ( .A1(n5448), .A2(n3240), .ZN(n3239) );
  NOR2_X1 U3677 ( .A1(n3244), .A2(n3243), .ZN(n3242) );
  INV_X1 U3678 ( .A(n5448), .ZN(n3241) );
  OR2_X1 U3679 ( .A1(n3667), .A2(n3666), .ZN(n3673) );
  NAND2_X1 U3680 ( .A1(n3187), .A2(n5425), .ZN(n3245) );
  AOI21_X1 U3681 ( .B1(n3822), .B2(n3944), .A(n3821), .ZN(n5135) );
  OR2_X1 U3682 ( .A1(n5774), .A2(n3685), .ZN(n6354) );
  XNOR2_X1 U3683 ( .A(n3628), .B(n3638), .ZN(n3806) );
  CLKBUF_X1 U3684 ( .A(n5025), .Z(n5406) );
  XNOR2_X1 U3685 ( .A(n3665), .B(n3664), .ZN(n3822) );
  AND2_X1 U3686 ( .A1(n3790), .A2(n3789), .ZN(n4759) );
  NAND2_X1 U3687 ( .A1(n3650), .A2(n3649), .ZN(n3665) );
  INV_X1 U3688 ( .A(n3652), .ZN(n3650) );
  NAND2_X1 U3689 ( .A1(n3592), .A2(n3591), .ZN(n3593) );
  XNOR2_X1 U3690 ( .A(n3636), .B(n3637), .ZN(n3805) );
  CLKBUF_X1 U3691 ( .A(n4781), .Z(n4782) );
  AND2_X1 U3692 ( .A1(n4640), .A2(n4641), .ZN(n3787) );
  OAI21_X1 U3693 ( .B1(n5969), .B2(n3666), .A(n3547), .ZN(n4550) );
  NAND2_X2 U3694 ( .A1(n3544), .A2(n3543), .ZN(n5969) );
  NAND2_X2 U3695 ( .A1(n5738), .A2(n4709), .ZN(n6086) );
  NAND2_X2 U3696 ( .A1(n6307), .A2(n3357), .ZN(n5704) );
  NAND2_X1 U3697 ( .A1(n3199), .A2(n3202), .ZN(n3544) );
  CLKBUF_X1 U3698 ( .A(n3781), .Z(n4752) );
  NOR2_X1 U3699 ( .A1(n6720), .A2(n6321), .ZN(n6350) );
  NAND2_X1 U3700 ( .A1(n4882), .A2(n4883), .ZN(n4881) );
  NOR2_X2 U3701 ( .A1(n4766), .A2(n4767), .ZN(n4882) );
  NAND2_X1 U3702 ( .A1(n4770), .A2(n4769), .ZN(n4766) );
  AND2_X1 U3703 ( .A1(n4301), .A2(n3219), .ZN(n4770) );
  NOR2_X1 U3704 ( .A1(n5136), .A2(n3232), .ZN(n3231) );
  OAI211_X1 U3705 ( .C1(n4395), .C2(n3449), .A(n4739), .B(n4456), .ZN(n3450)
         );
  NAND2_X1 U3706 ( .A1(n4560), .A2(n4324), .ZN(n4375) );
  OAI211_X1 U3707 ( .C1(n3753), .C2(n3515), .A(n3514), .B(n3513), .ZN(n3542)
         );
  AND2_X1 U3708 ( .A1(n3537), .A2(n3711), .ZN(n4470) );
  NAND2_X1 U3709 ( .A1(n4280), .A2(n4286), .ZN(n4368) );
  AND2_X2 U3710 ( .A1(n3446), .A2(n4286), .ZN(n4462) );
  AND2_X1 U3711 ( .A1(n4286), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3714) );
  INV_X1 U3712 ( .A(n3432), .ZN(n3439) );
  OR2_X1 U3713 ( .A1(n3510), .A2(n3509), .ZN(n3676) );
  OR2_X1 U3714 ( .A1(n3499), .A2(n3498), .ZN(n3556) );
  NOR2_X1 U3715 ( .A1(n3323), .A2(n3322), .ZN(n3330) );
  OR2_X2 U3716 ( .A1(n3342), .A2(n3341), .ZN(n3385) );
  AND4_X1 U3717 ( .A1(n3362), .A2(n3361), .A3(n3360), .A4(n3359), .ZN(n3370)
         );
  AND4_X1 U3718 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3296)
         );
  AND4_X1 U3719 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3295)
         );
  AND4_X1 U3720 ( .A1(n3399), .A2(n3398), .A3(n3397), .A4(n3396), .ZN(n3407)
         );
  AND4_X1 U3721 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3306)
         );
  AND4_X1 U3722 ( .A1(n3377), .A2(n3376), .A3(n3375), .A4(n3374), .ZN(n3382)
         );
  AND4_X1 U3723 ( .A1(n3390), .A2(n3389), .A3(n3388), .A4(n3387), .ZN(n3409)
         );
  AND4_X1 U3724 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3408)
         );
  AND4_X1 U3725 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  NAND2_X2 U3726 ( .A1(n7129), .A2(n6814), .ZN(n6694) );
  NAND2_X2 U3727 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7129), .ZN(n6696) );
  NOR2_X1 U3728 ( .A1(n5839), .A2(n7100), .ZN(n6517) );
  AND4_X1 U3729 ( .A1(n3405), .A2(n3404), .A3(n3403), .A4(n3402), .ZN(n3406)
         );
  AND4_X1 U3730 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3317)
         );
  AND2_X1 U3731 ( .A1(n3280), .A2(n3279), .ZN(n3286) );
  AOI22_X1 U3732 ( .A1(n4719), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3292) );
  AND4_X1 U3733 ( .A1(n3315), .A2(n3314), .A3(n3313), .A4(n3312), .ZN(n3316)
         );
  BUF_X2 U3734 ( .A(n3154), .Z(n4088) );
  BUF_X2 U3735 ( .A(n3332), .Z(n3175) );
  CLKBUF_X3 U3736 ( .A(n3332), .Z(n3176) );
  AND2_X2 U3737 ( .A1(n6659), .A2(n4753), .ZN(n6720) );
  AND2_X2 U3738 ( .A1(n3288), .A2(n4733), .ZN(n3391) );
  AND2_X2 U3739 ( .A1(n4728), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4715)
         );
  AND2_X2 U3740 ( .A1(n4583), .A2(n3290), .ZN(n4120) );
  AND2_X2 U3741 ( .A1(n3290), .A2(n4582), .ZN(n3350) );
  AND2_X2 U3742 ( .A1(n4733), .A2(n4583), .ZN(n3386) );
  AND2_X2 U3743 ( .A1(n3281), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3288)
         );
  OR2_X1 U3744 ( .A1(n5587), .A2(n5694), .ZN(n3159) );
  OR2_X1 U3745 ( .A1(n5693), .A2(n5694), .ZN(n5584) );
  OR2_X1 U3746 ( .A1(n5851), .A2(n6274), .ZN(n3160) );
  NAND2_X1 U3747 ( .A1(n3160), .A2(n3224), .ZN(U2796) );
  XNOR2_X1 U3748 ( .A(n3228), .B(n4424), .ZN(n5851) );
  AND2_X1 U3749 ( .A1(n5712), .A2(n4408), .ZN(n3185) );
  XNOR2_X1 U3750 ( .A(n4266), .B(n4265), .ZN(n5712) );
  AND2_X1 U3751 ( .A1(n3282), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3289)
         );
  AND2_X1 U3752 ( .A1(n3288), .A2(n3290), .ZN(n3177) );
  AND2_X1 U3753 ( .A1(n3288), .A2(n3290), .ZN(n3178) );
  AND2_X1 U3754 ( .A1(n4715), .A2(n4583), .ZN(n3162) );
  INV_X1 U3755 ( .A(n3400), .ZN(n3163) );
  AND4_X1 U3756 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3329)
         );
  NAND2_X1 U3757 ( .A1(n4772), .A2(n4773), .ZN(n4774) );
  AND2_X2 U3758 ( .A1(n4715), .A2(n3288), .ZN(n3500) );
  AND2_X1 U3759 ( .A1(n3373), .A2(n4287), .ZN(n3537) );
  AND2_X1 U3760 ( .A1(n4715), .A2(n4582), .ZN(n3165) );
  AND2_X4 U3761 ( .A1(n4715), .A2(n4582), .ZN(n3166) );
  NAND2_X2 U3762 ( .A1(n3586), .A2(n3585), .ZN(n5314) );
  AND2_X1 U3764 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U3765 ( .A1(n3214), .A2(n5314), .ZN(n3636) );
  INV_X2 U3766 ( .A(n3774), .ZN(n3772) );
  NAND2_X1 U3767 ( .A1(n3798), .A2(n3797), .ZN(n4765) );
  OAI21_X1 U3768 ( .B1(n3444), .B2(n3419), .A(n3768), .ZN(n3420) );
  OAI21_X1 U3769 ( .B1(n3416), .B2(n3415), .A(n3414), .ZN(n3444) );
  INV_X2 U3770 ( .A(n5544), .ZN(n4142) );
  BUF_X4 U3771 ( .A(n3363), .Z(n3168) );
  INV_X2 U3772 ( .A(n3442), .ZN(n3418) );
  AOI21_X2 U3773 ( .B1(n5477), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5476), 
        .ZN(n5478) );
  NOR2_X2 U3774 ( .A1(n5754), .A2(n5846), .ZN(n5477) );
  NOR2_X1 U3775 ( .A1(n3185), .A2(n3225), .ZN(n3224) );
  CLKBUF_X1 U3776 ( .A(n3282), .Z(n3169) );
  AND2_X1 U3777 ( .A1(n3773), .A2(n3383), .ZN(n3415) );
  AND2_X4 U3778 ( .A1(n4733), .A2(n3289), .ZN(n3364) );
  NOR2_X2 U3779 ( .A1(n5134), .A2(n5135), .ZN(n5246) );
  NOR2_X2 U3780 ( .A1(n3445), .A2(n3444), .ZN(n4403) );
  AND2_X1 U3781 ( .A1(n3289), .A2(n3290), .ZN(n3344) );
  OR2_X1 U3782 ( .A1(n3552), .A2(n3551), .ZN(n3205) );
  XNOR2_X1 U3784 ( .A(n4262), .B(n4274), .ZN(n5492) );
  NAND2_X1 U3785 ( .A1(n4262), .A2(n4220), .ZN(n5503) );
  XNOR2_X1 U3786 ( .A(n3554), .B(n3553), .ZN(n3775) );
  NOR2_X4 U3787 ( .A1(n4277), .A2(n3440), .ZN(n4442) );
  AND2_X4 U3788 ( .A1(n4715), .A2(n4583), .ZN(n3331) );
  NOR2_X4 U3789 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4583) );
  AND2_X4 U3790 ( .A1(n3288), .A2(n3290), .ZN(n3324) );
  NOR2_X1 U3791 ( .A1(n3678), .A2(n3677), .ZN(n3679) );
  NAND2_X1 U3792 ( .A1(n3214), .A2(n3213), .ZN(n3652) );
  AND2_X1 U3793 ( .A1(n5314), .A2(n3277), .ZN(n3213) );
  NOR2_X1 U3794 ( .A1(n5608), .A2(n3238), .ZN(n3237) );
  INV_X1 U3795 ( .A(n5620), .ZN(n3238) );
  INV_X1 U3796 ( .A(n3431), .ZN(n4280) );
  INV_X1 U3797 ( .A(n3416), .ZN(n3371) );
  OR2_X1 U3798 ( .A1(n4286), .A2(n6659), .ZN(n3573) );
  OR2_X1 U3799 ( .A1(n3383), .A2(n6659), .ZN(n3574) );
  AOI21_X1 U3800 ( .B1(n6487), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3750), 
        .ZN(n3757) );
  INV_X1 U3801 ( .A(n3709), .ZN(n3753) );
  AOI21_X1 U3802 ( .B1(n3431), .B2(n3422), .A(n4390), .ZN(n3414) );
  NOR2_X1 U3803 ( .A1(n4584), .A2(n6659), .ZN(n4213) );
  AND2_X1 U3804 ( .A1(n5436), .A2(n5431), .ZN(n3266) );
  NAND2_X1 U3805 ( .A1(n5418), .A2(n3264), .ZN(n3921) );
  AND2_X1 U3806 ( .A1(n3266), .A2(n3265), .ZN(n3264) );
  NOR2_X1 U3807 ( .A1(n3191), .A2(n3207), .ZN(n3206) );
  INV_X1 U3808 ( .A(n3690), .ZN(n3207) );
  AND2_X1 U3809 ( .A1(n4368), .A2(n4324), .ZN(n4382) );
  NAND2_X1 U3810 ( .A1(n5621), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5009) );
  NAND2_X1 U3811 ( .A1(n4512), .A2(n4518), .ZN(n4533) );
  OR3_X1 U3812 ( .A1(n6356), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n3702), 
        .ZN(n4230) );
  NOR2_X1 U3813 ( .A1(n5944), .A2(n5759), .ZN(n3705) );
  NOR2_X1 U3814 ( .A1(n4914), .A2(n4731), .ZN(n4407) );
  INV_X1 U3815 ( .A(n5836), .ZN(n6380) );
  NOR2_X1 U3816 ( .A1(n3469), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U3817 ( .A1(n3469), .A2(n6659), .ZN(n3248) );
  NAND2_X1 U3818 ( .A1(n4285), .A2(n3439), .ZN(n3416) );
  NAND2_X1 U3819 ( .A1(n3607), .A2(n3606), .ZN(n3637) );
  INV_X1 U3820 ( .A(n4470), .ZN(n3678) );
  AND2_X1 U3821 ( .A1(n4279), .A2(n4278), .ZN(n4448) );
  NAND2_X1 U3822 ( .A1(n3709), .A2(n3164), .ZN(n3756) );
  AOI21_X1 U3823 ( .B1(n3202), .B2(n3201), .A(n3186), .ZN(n3200) );
  OAI211_X1 U3824 ( .C1(n3753), .C2(n3529), .A(n3528), .B(n3527), .ZN(n3551)
         );
  OAI21_X1 U3825 ( .B1(n4577), .B2(STATE2_REG_0__SCAN_IN), .A(n3533), .ZN(
        n3554) );
  NOR2_X1 U3826 ( .A1(n3274), .A2(n3273), .ZN(n3272) );
  INV_X1 U3827 ( .A(n3275), .ZN(n3273) );
  INV_X1 U3828 ( .A(n5531), .ZN(n3274) );
  NOR2_X1 U3829 ( .A1(n5556), .A2(n5571), .ZN(n3268) );
  NAND2_X1 U3830 ( .A1(n3262), .A2(n5706), .ZN(n3261) );
  INV_X1 U3831 ( .A(n5632), .ZN(n3262) );
  NOR2_X1 U3832 ( .A1(n4367), .A2(n5663), .ZN(n3223) );
  NAND2_X1 U3833 ( .A1(n3249), .A2(n3209), .ZN(n3208) );
  INV_X1 U3834 ( .A(n3689), .ZN(n3210) );
  INV_X1 U3835 ( .A(n5361), .ZN(n3229) );
  NAND2_X1 U3836 ( .A1(n4298), .A2(n4297), .ZN(n4301) );
  NOR2_X1 U3837 ( .A1(n3766), .A2(n3769), .ZN(n4459) );
  NAND2_X1 U3838 ( .A1(n3574), .A2(n3573), .ZN(n3762) );
  OR2_X1 U3839 ( .A1(n3752), .A2(n3751), .ZN(n4397) );
  NOR2_X1 U3840 ( .A1(n4353), .A2(n3235), .ZN(n3233) );
  OR2_X1 U3841 ( .A1(n5486), .A2(n4116), .ZN(n4260) );
  INV_X1 U3842 ( .A(n5570), .ZN(n3269) );
  OR2_X1 U3843 ( .A1(n3266), .A2(n3265), .ZN(n3263) );
  NOR2_X1 U3844 ( .A1(n3886), .A2(n6232), .ZN(n3902) );
  AND2_X1 U3845 ( .A1(n3811), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3833)
         );
  NAND2_X1 U3846 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n3802), .ZN(n3810)
         );
  AOI21_X1 U3847 ( .B1(n3242), .B2(n3239), .A(n3198), .ZN(n3215) );
  NAND2_X1 U3848 ( .A1(n3242), .A2(n3241), .ZN(n3216) );
  INV_X1 U3849 ( .A(n3684), .ZN(n3217) );
  NAND2_X1 U3850 ( .A1(n4455), .A2(n4454), .ZN(n4484) );
  XNOR2_X1 U3851 ( .A(n3595), .B(n5314), .ZN(n4781) );
  OR2_X1 U3852 ( .A1(n5059), .A2(n4747), .ZN(n5066) );
  INV_X1 U3853 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6613) );
  INV_X1 U3854 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6487) );
  INV_X1 U3855 ( .A(n4822), .ZN(n6012) );
  NAND2_X1 U3856 ( .A1(n3781), .A2(n3541), .ZN(n3199) );
  AND2_X1 U3857 ( .A1(n4731), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3765) );
  NAND2_X1 U3858 ( .A1(n3227), .A2(n4427), .ZN(n3226) );
  NAND2_X1 U3859 ( .A1(n4433), .A2(REIP_REG_31__SCAN_IN), .ZN(n3227) );
  OR3_X1 U3860 ( .A1(n6717), .A2(n6648), .A3(n4406), .ZN(n5621) );
  INV_X1 U3861 ( .A(n6270), .ZN(n6288) );
  XNOR2_X1 U3862 ( .A(n4270), .B(n4269), .ZN(n4914) );
  OR2_X1 U3863 ( .A1(n4268), .A2(n4267), .ZN(n4270) );
  NAND2_X1 U3864 ( .A1(n6364), .A2(n4221), .ZN(n5836) );
  XNOR2_X1 U3865 ( .A(n4234), .B(n4233), .ZN(n5855) );
  AND2_X1 U3866 ( .A1(n6118), .A2(n5845), .ZN(n6110) );
  AND2_X1 U3867 ( .A1(n5916), .A2(n5925), .ZN(n5912) );
  INV_X1 U3868 ( .A(n6455), .ZN(n6474) );
  INV_X1 U3869 ( .A(n5969), .ZN(n5316) );
  CLKBUF_X1 U3870 ( .A(n4711), .Z(n4712) );
  AND2_X1 U3871 ( .A1(n6639), .A2(n6638), .ZN(n6656) );
  OAI21_X1 U3872 ( .B1(n3753), .B2(n3620), .A(n3627), .ZN(n3638) );
  AOI21_X1 U3873 ( .B1(n3418), .B2(n3417), .A(n3439), .ZN(n3419) );
  AND2_X1 U3874 ( .A1(n3748), .A2(n3747), .ZN(n3750) );
  XNOR2_X1 U3875 ( .A(n3484), .B(n3483), .ZN(n3257) );
  NAND2_X1 U3876 ( .A1(n3554), .A2(n3205), .ZN(n3535) );
  AND2_X1 U3877 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3464) );
  OR2_X1 U3878 ( .A1(n3400), .A2(n3307), .ZN(n3308) );
  OR2_X1 U3879 ( .A1(n3584), .A2(n3583), .ZN(n3608) );
  INV_X1 U3880 ( .A(n3574), .ZN(n3532) );
  INV_X1 U3881 ( .A(n5592), .ZN(n3236) );
  INV_X1 U3882 ( .A(n5520), .ZN(n3271) );
  NOR2_X1 U3883 ( .A1(n5660), .A2(n5669), .ZN(n3275) );
  INV_X1 U3884 ( .A(n3268), .ZN(n3267) );
  INV_X1 U3885 ( .A(n4501), .ZN(n3270) );
  INV_X1 U3886 ( .A(n4213), .ZN(n4256) );
  INV_X1 U3887 ( .A(n3907), .ZN(n3265) );
  AOI21_X1 U3888 ( .B1(n4264), .B2(EAX_REG_13__SCAN_IN), .A(n3906), .ZN(n3907)
         );
  NAND2_X1 U3889 ( .A1(n5636), .A2(n3237), .ZN(n5610) );
  INV_X1 U3890 ( .A(n3245), .ZN(n3240) );
  INV_X1 U3891 ( .A(n3675), .ZN(n3255) );
  INV_X1 U3892 ( .A(n5253), .ZN(n3232) );
  NAND2_X1 U3894 ( .A1(n3460), .A2(n3458), .ZN(n3531) );
  NAND2_X1 U3895 ( .A1(n3457), .A2(n3456), .ZN(n3458) );
  NAND2_X1 U3896 ( .A1(n4470), .A2(n3431), .ZN(n4579) );
  AND3_X1 U3897 ( .A1(n4275), .A2(n4448), .A3(n4284), .ZN(n4581) );
  XNOR2_X1 U3898 ( .A(n3552), .B(n3551), .ZN(n3553) );
  XNOR2_X1 U3899 ( .A(n3256), .B(n3257), .ZN(n3774) );
  INV_X1 U3900 ( .A(n3536), .ZN(n3256) );
  NAND2_X1 U3901 ( .A1(n3572), .A2(n3571), .ZN(n4818) );
  INV_X1 U3902 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6623) );
  INV_X1 U3903 ( .A(n4935), .ZN(n5263) );
  AOI22_X1 U3904 ( .A1(n3173), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3366) );
  AOI21_X1 U3905 ( .B1(n3386), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n3358), 
        .ZN(n3359) );
  AOI21_X1 U3906 ( .B1(n3176), .B2(INSTQUEUE_REG_10__3__SCAN_IN), .A(n3343), 
        .ZN(n3347) );
  AND2_X1 U3907 ( .A1(n4719), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U3908 ( .A1(n4125), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U3909 ( .A1(n3350), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U3910 ( .A1(n3165), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U3911 ( .A1(n3363), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3283) );
  AOI22_X1 U3912 ( .A1(n3500), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3153), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3284) );
  OAI21_X1 U3913 ( .B1(n6723), .B2(n4753), .A(n6646), .ZN(n4796) );
  AND2_X1 U3914 ( .A1(n4730), .A2(n4729), .ZN(n6624) );
  AND2_X1 U3915 ( .A1(n3768), .A2(n3417), .ZN(n3443) );
  AND2_X1 U3916 ( .A1(n4380), .A2(n4379), .ZN(n5522) );
  NOR2_X1 U3917 ( .A1(n3222), .A2(n5533), .ZN(n3221) );
  INV_X1 U3918 ( .A(n3223), .ZN(n3222) );
  AND2_X1 U3919 ( .A1(n4359), .A2(n4358), .ZN(n5560) );
  NAND2_X1 U3920 ( .A1(n5573), .A2(n4356), .ZN(n5574) );
  NAND2_X1 U3921 ( .A1(n5636), .A2(n5620), .ZN(n5619) );
  NAND2_X1 U3922 ( .A1(n3220), .A2(n4560), .ZN(n3219) );
  AND2_X1 U3923 ( .A1(n4512), .A2(n4511), .ZN(n6321) );
  INV_X1 U3924 ( .A(n4706), .ZN(n4660) );
  OR2_X1 U3925 ( .A1(n4259), .A2(n4258), .ZN(n4268) );
  AOI22_X1 U3926 ( .A1(n4217), .A2(n4216), .B1(n4404), .B2(n5511), .ZN(n4219)
         );
  AND2_X1 U3927 ( .A1(n4181), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4182)
         );
  NAND2_X1 U3928 ( .A1(n4182), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4259)
         );
  AOI22_X1 U3929 ( .A1(n4180), .A2(n4179), .B1(n4404), .B2(n5752), .ZN(n5531)
         );
  OR2_X1 U3930 ( .A1(n4158), .A2(n5766), .ZN(n4160) );
  NOR2_X1 U3931 ( .A1(n4160), .A2(n4159), .ZN(n4181) );
  INV_X1 U3932 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4503) );
  NAND2_X1 U3933 ( .A1(n4071), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4114)
         );
  NOR2_X1 U3934 ( .A1(n4018), .A2(n5599), .ZN(n4019) );
  NAND2_X1 U3935 ( .A1(n4019), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4069)
         );
  NOR2_X1 U3936 ( .A1(n3984), .A2(n5606), .ZN(n3985) );
  NAND2_X1 U3937 ( .A1(n3965), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3984)
         );
  NOR2_X1 U3938 ( .A1(n3952), .A2(n5635), .ZN(n3965) );
  NOR2_X1 U3939 ( .A1(n3261), .A2(n3260), .ZN(n3259) );
  INV_X1 U3940 ( .A(n5617), .ZN(n3260) );
  AND3_X1 U3941 ( .A1(n3951), .A2(n3950), .A3(n3949), .ZN(n5632) );
  INV_X1 U3942 ( .A(n5705), .ZN(n3258) );
  AND2_X1 U3943 ( .A1(n3902), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3903)
         );
  NAND2_X1 U3944 ( .A1(n3903), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3947)
         );
  NAND2_X1 U3945 ( .A1(n3901), .A2(n3900), .ZN(n5436) );
  NAND2_X1 U3946 ( .A1(n3872), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3886)
         );
  NOR2_X1 U3947 ( .A1(n3857), .A2(n3856), .ZN(n3872) );
  INV_X1 U3948 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3856) );
  CLKBUF_X1 U3949 ( .A(n5418), .Z(n5419) );
  NAND2_X1 U3950 ( .A1(n3838), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3857)
         );
  INV_X1 U3951 ( .A(n5359), .ZN(n3854) );
  CLKBUF_X1 U3952 ( .A(n5247), .Z(n5248) );
  NOR2_X1 U3953 ( .A1(n3810), .A2(n4922), .ZN(n3811) );
  AOI21_X1 U3954 ( .B1(n3817), .B2(n3944), .A(n3816), .ZN(n5131) );
  AOI21_X1 U3955 ( .B1(n3805), .B2(n3944), .A(n3804), .ZN(n4878) );
  NOR2_X1 U3956 ( .A1(n3792), .A2(n4776), .ZN(n3802) );
  INV_X1 U3957 ( .A(n3796), .ZN(n3797) );
  NAND2_X1 U3958 ( .A1(n4781), .A2(n3944), .ZN(n3798) );
  NAND2_X1 U3959 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3792) );
  AND2_X1 U3960 ( .A1(n4459), .A2(n3771), .ZN(n4520) );
  NAND2_X1 U3961 ( .A1(n5549), .A2(n3223), .ZN(n5665) );
  AND2_X1 U3962 ( .A1(n5774), .A2(n5927), .ZN(n5775) );
  OAI21_X1 U3963 ( .B1(n4435), .B2(n6123), .A(n6356), .ZN(n4436) );
  NOR2_X1 U3964 ( .A1(n3192), .A2(n3251), .ZN(n3250) );
  INV_X1 U3965 ( .A(n3687), .ZN(n3251) );
  NAND2_X1 U3966 ( .A1(n6155), .A2(n5708), .ZN(n5707) );
  NOR2_X2 U3967 ( .A1(n5438), .A2(n6156), .ZN(n6155) );
  NAND2_X1 U3968 ( .A1(n6354), .A2(n3218), .ZN(n3244) );
  NOR2_X1 U3969 ( .A1(n5412), .A2(n3245), .ZN(n3243) );
  NAND2_X1 U3970 ( .A1(n5944), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U3971 ( .A1(n3230), .A2(n3181), .ZN(n6230) );
  AND2_X1 U3972 ( .A1(n3180), .A2(n5421), .ZN(n3181) );
  NOR2_X1 U3973 ( .A1(n4899), .A2(n5136), .ZN(n5252) );
  NOR2_X2 U3974 ( .A1(n4881), .A2(n4857), .ZN(n4900) );
  AND2_X1 U3975 ( .A1(n4581), .A2(n4447), .ZN(n4609) );
  INV_X1 U3976 ( .A(n6433), .ZN(n6471) );
  XNOR2_X1 U3977 ( .A(n4301), .B(n4551), .ZN(n4642) );
  INV_X1 U3978 ( .A(n4382), .ZN(n4552) );
  OR2_X1 U3979 ( .A1(n3422), .A2(n3767), .ZN(n4584) );
  OR2_X1 U3980 ( .A1(n3764), .A2(n3763), .ZN(n4587) );
  AOI21_X1 U3981 ( .B1(n3761), .B2(n3760), .A(n3759), .ZN(n3764) );
  OR3_X1 U3982 ( .A1(n4782), .A2(n5139), .A3(n4747), .ZN(n5145) );
  NAND2_X1 U3983 ( .A1(n6659), .A2(n4796), .ZN(n4935) );
  NAND2_X1 U3984 ( .A1(n4782), .A2(n3772), .ZN(n5059) );
  AND2_X1 U3985 ( .A1(n6709), .A2(n4796), .ZN(n4841) );
  OR2_X1 U3986 ( .A1(n3772), .A2(n5024), .ZN(n5971) );
  NOR2_X1 U3987 ( .A1(n6009), .A2(n5316), .ZN(n5317) );
  INV_X1 U3988 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4731) );
  OR2_X1 U3989 ( .A1(n5009), .A2(n4411), .ZN(n6272) );
  INV_X1 U3990 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5635) );
  INV_X1 U3991 ( .A(n6285), .ZN(n6258) );
  AND2_X1 U3992 ( .A1(n4914), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4915) );
  OR2_X1 U3993 ( .A1(n5009), .A2(n4919), .ZN(n6270) );
  AND2_X1 U3994 ( .A1(n4913), .A2(n6212), .ZN(n5305) );
  INV_X1 U3995 ( .A(n5709), .ZN(n6303) );
  INV_X1 U3996 ( .A(n6086), .ZN(n6315) );
  INV_X1 U3997 ( .A(n5738), .ZN(n6317) );
  AND2_X1 U3998 ( .A1(n5738), .A2(n4710), .ZN(n6318) );
  NAND2_X1 U3999 ( .A1(n4706), .A2(n4705), .ZN(n5738) );
  OAI21_X1 U4000 ( .B1(n4704), .B2(n4703), .A(n6657), .ZN(n4705) );
  NOR2_X2 U4001 ( .A1(n6314), .A2(n6318), .ZN(n5739) );
  BUF_X1 U4002 ( .A(n6350), .Z(n6341) );
  NAND2_X1 U4003 ( .A1(n3269), .A2(n4053), .ZN(n5557) );
  INV_X1 U4004 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4776) );
  INV_X1 U4005 ( .A(n6390), .ZN(n6360) );
  INV_X1 U4006 ( .A(n5959), .ZN(n6403) );
  AND2_X1 U4007 ( .A1(n3703), .A2(n5858), .ZN(n3211) );
  NAND2_X1 U4008 ( .A1(n5459), .A2(n6471), .ZN(n5959) );
  NAND2_X1 U4009 ( .A1(n5741), .A2(n3703), .ZN(n3212) );
  NOR2_X1 U4010 ( .A1(n6128), .A2(n4481), .ZN(n6118) );
  NAND2_X1 U4011 ( .A1(n5424), .A2(n5425), .ZN(n6355) );
  NAND2_X1 U4012 ( .A1(n5365), .A2(n5364), .ZN(n5363) );
  NAND2_X1 U4013 ( .A1(n5239), .A2(n3675), .ZN(n5365) );
  NAND2_X1 U4014 ( .A1(n4484), .A2(n4463), .ZN(n6448) );
  NOR2_X1 U4015 ( .A1(n4731), .A2(n4510), .ZN(n4753) );
  AND2_X1 U4016 ( .A1(n4747), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4787) );
  INV_X1 U4017 ( .A(n6496), .ZN(n6015) );
  OR2_X1 U4018 ( .A1(n4587), .A2(n6166), .ZN(n6646) );
  INV_X1 U4019 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U4020 ( .A1(n4823), .A2(n6012), .ZN(n4848) );
  AND2_X1 U4021 ( .A1(n6491), .A2(n6490), .ZN(n6544) );
  OAI21_X1 U4022 ( .B1(n5100), .B2(n5102), .A(n5099), .ZN(n5124) );
  OAI211_X1 U4023 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4510), .A(n5375), .B(n5268), .ZN(n5291) );
  AOI22_X1 U4024 ( .A1(n5267), .A2(n5264), .B1(n6488), .B2(n5262), .ZN(n5297)
         );
  NAND2_X1 U4025 ( .A1(n4938), .A2(n4937), .ZN(n4964) );
  INV_X1 U4026 ( .A(n5231), .ZN(n6492) );
  INV_X1 U4027 ( .A(n5212), .ZN(n6514) );
  INV_X1 U4028 ( .A(n6566), .ZN(n6526) );
  INV_X1 U4029 ( .A(n6596), .ZN(n6532) );
  INV_X1 U4030 ( .A(n6573), .ZN(n6537) );
  OAI211_X1 U4031 ( .C1(n6015), .C2(n6014), .A(n6013), .B(n6012), .ZN(n6043)
         );
  INV_X1 U4032 ( .A(n6606), .ZN(n6543) );
  AND2_X1 U4033 ( .A1(n4745), .A2(n6635), .ZN(n6649) );
  AND2_X1 U4034 ( .A1(n6645), .A2(n6644), .ZN(n6710) );
  OR2_X1 U4035 ( .A1(n4409), .A2(STATE_REG_0__SCAN_IN), .ZN(n6673) );
  INV_X1 U4036 ( .A(STATE_REG_1__SCAN_IN), .ZN(n7000) );
  OR2_X1 U4037 ( .A1(n4432), .A2(n3226), .ZN(n3225) );
  OR2_X1 U4038 ( .A1(n5857), .A2(n5709), .ZN(n4393) );
  OAI21_X1 U4039 ( .B1(n5855), .B2(n6364), .A(n4273), .ZN(U2955) );
  AND2_X1 U4040 ( .A1(n4496), .A2(n3276), .ZN(n4497) );
  NAND2_X2 U4041 ( .A1(n3330), .A2(n3329), .ZN(n3383) );
  NAND2_X1 U4042 ( .A1(n4854), .A2(n4855), .ZN(n4856) );
  OR2_X2 U4043 ( .A1(n3356), .A2(n3355), .ZN(n3431) );
  AND2_X1 U4044 ( .A1(n3269), .A2(n3268), .ZN(n3179) );
  AND2_X1 U4045 ( .A1(n3231), .A2(n3229), .ZN(n3180) );
  NOR2_X1 U4046 ( .A1(n3258), .A2(n3261), .ZN(n5616) );
  AND2_X1 U4047 ( .A1(n4435), .A2(n3195), .ZN(n4434) );
  INV_X1 U4048 ( .A(n3541), .ZN(n3201) );
  NAND2_X1 U4049 ( .A1(n4285), .A2(n3711), .ZN(n3442) );
  OAI21_X1 U4050 ( .B1(n3470), .B2(n3469), .A(n3566), .ZN(n4608) );
  BUF_X1 U4051 ( .A(n3364), .Z(n4236) );
  AND2_X1 U4052 ( .A1(n3230), .A2(n3180), .ZN(n3182) );
  INV_X1 U4053 ( .A(n3935), .ZN(n3944) );
  NAND2_X1 U4054 ( .A1(n3208), .A2(n3690), .ZN(n5817) );
  NAND2_X1 U4055 ( .A1(n3468), .A2(n3467), .ZN(n3469) );
  AND4_X1 U4056 ( .A1(n3381), .A2(n3380), .A3(n3379), .A4(n3378), .ZN(n3183)
         );
  NAND2_X1 U4057 ( .A1(n3208), .A2(n3206), .ZN(n4435) );
  NAND2_X1 U4058 ( .A1(n3688), .A2(n3687), .ZN(n5832) );
  OR2_X1 U4059 ( .A1(n5503), .A2(n5839), .ZN(n3184) );
  NAND2_X1 U4060 ( .A1(n4435), .A2(n3694), .ZN(n5809) );
  BUF_X1 U4061 ( .A(n3704), .Z(n5741) );
  AND2_X1 U4062 ( .A1(n3532), .A2(n3676), .ZN(n3186) );
  INV_X1 U4063 ( .A(n3203), .ZN(n3202) );
  NAND2_X1 U4064 ( .A1(n3204), .A2(n3542), .ZN(n3203) );
  NAND2_X1 U4065 ( .A1(n5774), .A2(n3686), .ZN(n3187) );
  AND2_X1 U4066 ( .A1(n3683), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3188)
         );
  OR2_X1 U4067 ( .A1(n3587), .A2(n3574), .ZN(n3189) );
  AND2_X1 U4068 ( .A1(n3287), .A2(n4718), .ZN(n3345) );
  INV_X1 U4069 ( .A(n4293), .ZN(n4560) );
  OR2_X1 U4070 ( .A1(n3357), .A2(n4510), .ZN(n3190) );
  AND2_X1 U4071 ( .A1(n5418), .A2(n5431), .ZN(n5432) );
  INV_X1 U4072 ( .A(n4747), .ZN(n5024) );
  NAND2_X1 U4073 ( .A1(n5549), .A2(n5672), .ZN(n5662) );
  NOR2_X1 U4074 ( .A1(n5535), .A2(n5522), .ZN(n4383) );
  OAI21_X1 U4075 ( .B1(n3217), .B2(n3216), .A(n3215), .ZN(n6106) );
  OAI21_X1 U4076 ( .B1(n3684), .B2(n3245), .A(n3242), .ZN(n5447) );
  NAND2_X1 U4077 ( .A1(n3249), .A2(n3689), .ZN(n5824) );
  NOR2_X1 U4078 ( .A1(n5574), .A2(n5560), .ZN(n4360) );
  NAND2_X1 U4079 ( .A1(n3684), .A2(n5412), .ZN(n5424) );
  AND2_X1 U4080 ( .A1(n5774), .A2(n3692), .ZN(n3191) );
  AND2_X1 U4081 ( .A1(n5774), .A2(n5833), .ZN(n3192) );
  INV_X1 U4082 ( .A(n5669), .ZN(n4141) );
  NOR2_X1 U4083 ( .A1(n5559), .A2(n4465), .ZN(n4464) );
  INV_X1 U4084 ( .A(n3235), .ZN(n3234) );
  NAND2_X1 U4085 ( .A1(n3237), .A2(n3236), .ZN(n3235) );
  OR2_X1 U4086 ( .A1(n3270), .A2(n3267), .ZN(n3193) );
  AND2_X1 U4087 ( .A1(n4464), .A2(n5551), .ZN(n5549) );
  AND2_X1 U4088 ( .A1(n3272), .A2(n3271), .ZN(n3194) );
  AND2_X1 U4089 ( .A1(n3694), .A2(n6123), .ZN(n3195) );
  INV_X1 U4090 ( .A(n4404), .ZN(n4116) );
  NAND2_X1 U4091 ( .A1(n3230), .A2(n3231), .ZN(n5251) );
  AND2_X1 U4092 ( .A1(n5636), .A2(n3234), .ZN(n3196) );
  NAND2_X1 U4093 ( .A1(n4405), .A2(n4404), .ZN(n3197) );
  INV_X1 U4094 ( .A(n4115), .ZN(n4263) );
  AND2_X1 U4095 ( .A1(n5774), .A2(n5466), .ZN(n3198) );
  AOI21_X1 U4096 ( .B1(n3774), .B2(n3944), .A(n4263), .ZN(n4760) );
  INV_X2 U4097 ( .A(n5839), .ZN(n6385) );
  AND2_X1 U4098 ( .A1(n4300), .A2(n4299), .ZN(n4551) );
  INV_X1 U4099 ( .A(n4551), .ZN(n3220) );
  INV_X1 U4100 ( .A(n3385), .ZN(n4390) );
  OR2_X1 U4101 ( .A1(n6665), .A2(n6496), .ZN(n5839) );
  OAI21_X2 U4102 ( .B1(n3781), .B2(n3203), .A(n3200), .ZN(n3552) );
  NAND2_X1 U4103 ( .A1(n3541), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3204) );
  XNOR2_X1 U4104 ( .A(n3530), .B(n3531), .ZN(n4577) );
  AND2_X2 U4105 ( .A1(n5741), .A2(n3211), .ZN(n5476) );
  NAND2_X1 U4106 ( .A1(n3707), .A2(n3212), .ZN(n3708) );
  INV_X1 U4107 ( .A(n3595), .ZN(n3214) );
  NAND2_X2 U4108 ( .A1(n3665), .A2(n3679), .ZN(n5774) );
  NAND3_X1 U4109 ( .A1(n3665), .A2(n3817), .A3(n3164), .ZN(n3659) );
  NAND2_X1 U4110 ( .A1(n5549), .A2(n3221), .ZN(n5535) );
  NAND2_X1 U4111 ( .A1(n3470), .A2(n3247), .ZN(n3246) );
  NAND2_X1 U4112 ( .A1(n3470), .A2(n3469), .ZN(n3566) );
  OAI211_X1 U4113 ( .C1(n3470), .C2(n3248), .A(n3246), .B(n3189), .ZN(n3484)
         );
  NAND2_X1 U4114 ( .A1(n3688), .A2(n3250), .ZN(n3249) );
  NAND2_X1 U4115 ( .A1(n5238), .A2(n5240), .ZN(n5239) );
  AOI21_X1 U4116 ( .B1(n3255), .B2(n5364), .A(n3188), .ZN(n3252) );
  NAND2_X1 U4117 ( .A1(n5238), .A2(n3254), .ZN(n3253) );
  AND2_X1 U4118 ( .A1(n5240), .A2(n5364), .ZN(n3254) );
  NAND2_X1 U4119 ( .A1(n4759), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U4120 ( .A1(n3257), .A2(n3536), .ZN(n3595) );
  NAND3_X1 U4121 ( .A1(n4854), .A2(n3818), .A3(n4855), .ZN(n5134) );
  NAND2_X1 U4122 ( .A1(n5705), .A2(n3259), .ZN(n5603) );
  NAND2_X1 U4123 ( .A1(n5705), .A2(n5706), .ZN(n5631) );
  INV_X1 U4124 ( .A(n5603), .ZN(n3983) );
  OAI211_X1 U4125 ( .C1(n5418), .C2(n3265), .A(n3921), .B(n3263), .ZN(n5735)
         );
  NOR2_X2 U4126 ( .A1(n5570), .A2(n3193), .ZN(n4500) );
  NAND2_X1 U4127 ( .A1(n4142), .A2(n3272), .ZN(n5518) );
  AND2_X1 U4128 ( .A1(n4142), .A2(n3275), .ZN(n5530) );
  NAND2_X1 U4129 ( .A1(n4142), .A2(n4141), .ZN(n5659) );
  AND2_X2 U4130 ( .A1(n4142), .A2(n3194), .ZN(n4218) );
  INV_X1 U4131 ( .A(n3787), .ZN(n4639) );
  NAND2_X1 U4132 ( .A1(n3163), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3279)
         );
  AOI22_X1 U4133 ( .A1(n3178), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3163), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3303) );
  XNOR2_X1 U4134 ( .A(n3566), .B(n4818), .ZN(n4711) );
  OR2_X1 U4135 ( .A1(n5912), .A2(n4495), .ZN(n3276) );
  INV_X1 U4136 ( .A(READY_N), .ZN(n6719) );
  NAND2_X1 U4137 ( .A1(n3773), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3935) );
  AND2_X1 U4138 ( .A1(n4290), .A2(n6657), .ZN(n6307) );
  AND2_X1 U4139 ( .A1(n3638), .A2(n3637), .ZN(n3277) );
  AND2_X1 U4140 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4141 ( .A1(n6166), .A2(n4510), .ZN(n6496) );
  INV_X1 U4142 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6209) );
  INV_X1 U4143 ( .A(n6700), .ZN(n7128) );
  INV_X1 U4144 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4233) );
  NAND2_X1 U4145 ( .A1(n4512), .A2(n4520), .ZN(n6364) );
  INV_X1 U4146 ( .A(n6364), .ZN(n6386) );
  AND2_X1 U4147 ( .A1(n3165), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3358) );
  OR2_X1 U4148 ( .A1(n3605), .A2(n3604), .ZN(n3654) );
  OR2_X1 U4149 ( .A1(n3481), .A2(n3480), .ZN(n3482) );
  AOI22_X1 U4150 ( .A1(n4125), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3365) );
  INV_X1 U4151 ( .A(n5604), .ZN(n3982) );
  OR2_X1 U4152 ( .A1(n3626), .A2(n3625), .ZN(n3653) );
  INV_X1 U4153 ( .A(n3482), .ZN(n3587) );
  AOI22_X1 U4154 ( .A1(n3709), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3526), 
        .B2(n3482), .ZN(n3483) );
  OR2_X1 U4155 ( .A1(n3455), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3456)
         );
  INV_X1 U4156 ( .A(n3486), .ZN(n3487) );
  AND2_X1 U4157 ( .A1(n6613), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3730)
         );
  OR2_X1 U4158 ( .A1(n4154), .A2(n4153), .ZN(n4165) );
  INV_X1 U4159 ( .A(n5736), .ZN(n3919) );
  INV_X1 U4160 ( .A(n5131), .ZN(n3818) );
  OR2_X1 U4161 ( .A1(n3648), .A2(n3647), .ZN(n3669) );
  OR2_X1 U4162 ( .A1(n3525), .A2(n3524), .ZN(n3555) );
  INV_X1 U4163 ( .A(n3756), .ZN(n3758) );
  INV_X1 U4164 ( .A(n4069), .ZN(n4070) );
  INV_X1 U4165 ( .A(n5571), .ZN(n4053) );
  OR2_X1 U4166 ( .A1(n3947), .A2(n6209), .ZN(n3952) );
  OR2_X1 U4167 ( .A1(n6356), .A2(n5833), .ZN(n3689) );
  AND2_X1 U4168 ( .A1(n3568), .A2(n6045), .ZN(n4975) );
  INV_X1 U4169 ( .A(n4403), .ZN(n4479) );
  AND2_X1 U4170 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4070), .ZN(n4071)
         );
  AND2_X1 U4171 ( .A1(n3833), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3838)
         );
  AND2_X1 U4172 ( .A1(n4396), .A2(n3762), .ZN(n3763) );
  AND2_X1 U4173 ( .A1(n6485), .A2(n5021), .ZN(n5380) );
  INV_X1 U4174 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6618) );
  AND2_X1 U4175 ( .A1(n5060), .A2(n6015), .ZN(n5063) );
  INV_X1 U4176 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4159) );
  INV_X1 U4177 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5599) );
  INV_X1 U4178 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5606) );
  INV_X1 U4179 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6232) );
  INV_X1 U4180 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4922) );
  INV_X1 U4181 ( .A(n6307), .ZN(n4391) );
  NOR2_X1 U4182 ( .A1(n4114), .A2(n4503), .ZN(n4138) );
  XNOR2_X1 U4183 ( .A(n3593), .B(n6463), .ZN(n4773) );
  OR2_X1 U4184 ( .A1(n5921), .A2(n5902), .ZN(n5916) );
  AND2_X1 U4185 ( .A1(n4348), .A2(n4347), .ZN(n5592) );
  AND2_X1 U4186 ( .A1(n6143), .A2(n4904), .ZN(n5459) );
  OR2_X1 U4187 ( .A1(n4225), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6454) );
  INV_X1 U4188 ( .A(n6616), .ZN(n4742) );
  OR2_X1 U4189 ( .A1(n4824), .A2(n5969), .ZN(n6495) );
  OR2_X1 U4190 ( .A1(n5066), .A2(n5969), .ZN(n5269) );
  OR2_X1 U4191 ( .A1(n3542), .A2(n3201), .ZN(n3543) );
  OR3_X1 U4192 ( .A1(n3772), .A2(n5970), .A3(n4747), .ZN(n5185) );
  INV_X1 U4193 ( .A(n5314), .ZN(n5970) );
  INV_X1 U4194 ( .A(n5320), .ZN(n6014) );
  INV_X1 U4195 ( .A(n4462), .ZN(n6722) );
  INV_X1 U4196 ( .A(n6212), .ZN(n4408) );
  INV_X1 U4197 ( .A(n6274), .ZN(n6286) );
  INV_X1 U4198 ( .A(n6272), .ZN(n6247) );
  AND2_X1 U4199 ( .A1(n5621), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6285) );
  AND2_X1 U4200 ( .A1(n5621), .A2(n4915), .ZN(n6294) );
  NAND2_X1 U4201 ( .A1(n3985), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4018)
         );
  AND2_X1 U4202 ( .A1(n5734), .A2(n5737), .ZN(n6300) );
  NOR2_X1 U4203 ( .A1(n4587), .A2(n6655), .ZN(n4512) );
  AND2_X1 U4204 ( .A1(n4491), .A2(n4490), .ZN(n6126) );
  AND2_X1 U4205 ( .A1(n4484), .A2(n4609), .ZN(n6433) );
  AND2_X1 U4206 ( .A1(n3550), .A2(n3562), .ZN(n4644) );
  INV_X1 U4207 ( .A(n6448), .ZN(n6467) );
  NOR2_X1 U4208 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n5499) );
  OAI21_X1 U4209 ( .B1(n5977), .B2(n5980), .A(n5976), .ZN(n6002) );
  NOR2_X1 U4210 ( .A1(n5145), .A2(n5316), .ZN(n5972) );
  OAI221_X1 U4211 ( .B1(n5377), .B2(n6166), .C1(n5377), .C2(n5376), .A(n5375), 
        .ZN(n5402) );
  OAI211_X1 U4212 ( .C1(n6015), .C2(n5031), .A(n5030), .B(n6012), .ZN(n5055)
         );
  INV_X1 U4213 ( .A(n6495), .ZN(n6547) );
  NOR2_X1 U4214 ( .A1(n5066), .A2(n5316), .ZN(n5095) );
  INV_X1 U4215 ( .A(n5269), .ZN(n5294) );
  INV_X1 U4216 ( .A(n6558), .ZN(n6510) );
  INV_X1 U4217 ( .A(n6569), .ZN(n6528) );
  INV_X1 U4218 ( .A(n6611), .ZN(n6548) );
  AND2_X1 U4219 ( .A1(n3765), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6657) );
  INV_X1 U4220 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6814) );
  NAND2_X1 U4221 ( .A1(n4533), .A2(n4528), .ZN(n6717) );
  INV_X1 U4222 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6659) );
  OR2_X1 U4223 ( .A1(n4161), .A2(n4181), .ZN(n6059) );
  NAND2_X1 U4224 ( .A1(n5621), .A2(n4407), .ZN(n6212) );
  OR2_X1 U4225 ( .A1(n5009), .A2(n4425), .ZN(n6274) );
  NAND2_X1 U4226 ( .A1(n4390), .A2(n6307), .ZN(n5709) );
  INV_X1 U4227 ( .A(n5454), .ZN(n5473) );
  INV_X1 U4228 ( .A(n6321), .ZN(n6352) );
  OR3_X1 U4229 ( .A1(n4533), .A2(n3446), .A3(READY_N), .ZN(n4706) );
  NAND2_X1 U4230 ( .A1(n5836), .A2(n4224), .ZN(n6390) );
  AND2_X1 U4231 ( .A1(n5912), .A2(n5844), .ZN(n6117) );
  NAND2_X1 U4232 ( .A1(n4484), .A2(n4461), .ZN(n6455) );
  INV_X1 U4233 ( .A(n6483), .ZN(n4786) );
  INV_X1 U4234 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6169) );
  INV_X1 U4235 ( .A(n5972), .ZN(n6008) );
  OR2_X1 U4236 ( .A1(n5145), .A2(n5969), .ZN(n5409) );
  AOI22_X1 U4237 ( .A1(n5029), .A2(n5023), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5031), .ZN(n5058) );
  INV_X1 U4238 ( .A(n4819), .ZN(n4853) );
  OR2_X1 U4239 ( .A1(n4863), .A2(n5316), .ZN(n6585) );
  INV_X1 U4240 ( .A(n5095), .ZN(n5130) );
  INV_X1 U4241 ( .A(n6589), .ZN(n6521) );
  INV_X1 U4242 ( .A(n6555), .ZN(n6508) );
  OR3_X1 U4243 ( .A1(n5059), .A2(n5316), .A3(n5024), .ZN(n6610) );
  OR3_X1 U4244 ( .A1(n5059), .A2(n5024), .A3(n5969), .ZN(n6603) );
  INV_X1 U4245 ( .A(n5317), .ZN(n6050) );
  INV_X1 U4246 ( .A(n6657), .ZN(n6655) );
  INV_X1 U4247 ( .A(n6707), .ZN(n6703) );
  NOR2_X1 U4248 ( .A1(STATE_REG_0__SCAN_IN), .A2(n7000), .ZN(n6700) );
  OAI21_X1 U4249 ( .B1(n5492), .B2(n5704), .A(n4394), .ZN(U2829) );
  INV_X1 U4250 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3281) );
  INV_X1 U4251 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3282) );
  NOR2_X1 U4252 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3287) );
  AOI22_X1 U4253 ( .A1(n3173), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3294) );
  AND2_X2 U4254 ( .A1(n4714), .A2(n4583), .ZN(n3471) );
  AOI22_X1 U4255 ( .A1(n3471), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4256 ( .A1(n3162), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4257 ( .A1(n3332), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3162), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4258 ( .A1(n3471), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4259 ( .A1(n4719), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4260 ( .A1(n3154), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3297) );
  AOI22_X1 U4261 ( .A1(n3344), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4120), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4262 ( .A1(n3165), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4263 ( .A1(n3500), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3301) );
  NAND2_X1 U4264 ( .A1(n3165), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3311)
         );
  NAND2_X1 U4265 ( .A1(n3350), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4266 ( .A1(n3386), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3309)
         );
  INV_X1 U4267 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3307) );
  NAND2_X1 U4268 ( .A1(n3500), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4269 ( .A1(n3363), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3314) );
  NAND2_X1 U4270 ( .A1(n3154), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3313)
         );
  NAND2_X1 U4271 ( .A1(n3364), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3312)
         );
  NAND2_X1 U4272 ( .A1(n3317), .A2(n3316), .ZN(n3323) );
  NAND2_X1 U4273 ( .A1(n3162), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4274 ( .A1(n3344), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3320) );
  NAND2_X1 U4275 ( .A1(n3171), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3319) );
  NAND2_X1 U4276 ( .A1(n3345), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3318) );
  NAND4_X1 U4277 ( .A1(n3321), .A2(n3320), .A3(n3319), .A4(n3318), .ZN(n3322)
         );
  NAND2_X1 U4278 ( .A1(n3471), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3328) );
  NAND2_X1 U4279 ( .A1(n3156), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3327) );
  NAND2_X1 U4280 ( .A1(n3176), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4281 ( .A1(n3324), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3325) );
  AOI22_X1 U4282 ( .A1(n3173), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4283 ( .A1(n3331), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4284 ( .A1(n3471), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4285 ( .A1(n3156), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4286 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3342)
         );
  AOI22_X1 U4287 ( .A1(n3363), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4288 ( .A1(n3500), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4289 ( .A1(n3166), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4290 ( .A1(n4125), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3350), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4291 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3341)
         );
  AOI22_X1 U4292 ( .A1(n3471), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3349) );
  AOI22_X1 U4293 ( .A1(n3331), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3348) );
  AOI22_X1 U4294 ( .A1(n3344), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3346) );
  NAND4_X1 U4295 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3356)
         );
  AOI22_X1 U4296 ( .A1(n3168), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4297 ( .A1(n3500), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4298 ( .A1(n3166), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3352) );
  NAND4_X1 U4299 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3355)
         );
  OAI211_X1 U4300 ( .C1(n3422), .C2(n3383), .A(n3357), .B(n3431), .ZN(n3429)
         );
  INV_X1 U4301 ( .A(n3429), .ZN(n3372) );
  AOI22_X1 U4302 ( .A1(n3500), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4303 ( .A1(n3155), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U4304 ( .A1(n3471), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4305 ( .A1(n3167), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4306 ( .A1(n3331), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4307 ( .A1(n3372), .A2(n3371), .ZN(n3766) );
  INV_X1 U4308 ( .A(n3766), .ZN(n3412) );
  AOI22_X1 U4309 ( .A1(n3500), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4310 ( .A1(n3350), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3376) );
  AOI22_X1 U4311 ( .A1(n3166), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4312 ( .A1(n3168), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4313 ( .A1(n3172), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4314 ( .A1(n3471), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4315 ( .A1(n3331), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4316 ( .A1(n3344), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3345), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3378) );
  NAND2_X2 U4317 ( .A1(n3382), .A2(n3183), .ZN(n4287) );
  NAND2_X1 U4318 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6681) );
  OAI21_X1 U4319 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n6681), .ZN(n4409) );
  NAND2_X1 U4320 ( .A1(n3446), .A2(n4409), .ZN(n3441) );
  NAND2_X1 U4321 ( .A1(n3441), .A2(n3384), .ZN(n3411) );
  NAND2_X2 U4322 ( .A1(n3418), .A2(n3385), .ZN(n4277) );
  NAND2_X1 U4323 ( .A1(n3168), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3390) );
  NAND2_X1 U4324 ( .A1(n3500), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3389) );
  NAND2_X1 U4325 ( .A1(n3158), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3388)
         );
  NAND2_X1 U4326 ( .A1(n3386), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3387)
         );
  NAND2_X1 U4327 ( .A1(n3154), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3395)
         );
  NAND2_X1 U4328 ( .A1(n3162), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3394) );
  NAND2_X1 U4329 ( .A1(n3324), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3393) );
  NAND2_X1 U4330 ( .A1(n3173), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3392) );
  NAND2_X1 U4331 ( .A1(n3155), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3399) );
  NAND2_X1 U4332 ( .A1(n3471), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3398) );
  NAND2_X1 U4333 ( .A1(n3166), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3397)
         );
  NAND2_X1 U4334 ( .A1(n3345), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4335 ( .A1(n3364), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3405)
         );
  NAND2_X1 U4336 ( .A1(n3171), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3404) );
  NAND2_X1 U4337 ( .A1(n3350), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3403) );
  INV_X1 U4338 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3401) );
  OR2_X1 U4339 ( .A1(n3400), .A2(n3401), .ZN(n3402) );
  NAND4_X4 U4340 ( .A1(n3409), .A2(n3408), .A3(n3407), .A4(n3406), .ZN(n4286)
         );
  NAND2_X1 U4341 ( .A1(n4277), .A2(n4462), .ZN(n3410) );
  NAND4_X1 U4342 ( .A1(n3412), .A2(n4579), .A3(n3411), .A4(n3410), .ZN(n3421)
         );
  NAND2_X1 U4343 ( .A1(n3768), .A2(n4801), .ZN(n5008) );
  NAND2_X1 U4344 ( .A1(n3420), .A2(n5008), .ZN(n3428) );
  OAI21_X1 U4345 ( .B1(n3421), .B2(n3428), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3424) );
  NAND2_X1 U4346 ( .A1(n3709), .A2(n3422), .ZN(n3423) );
  NAND2_X1 U4347 ( .A1(n3424), .A2(n3423), .ZN(n3463) );
  NAND2_X1 U4348 ( .A1(n3463), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U4349 ( .A1(n5499), .A2(n6659), .ZN(n4225) );
  MUX2_X1 U4350 ( .A(n3765), .B(n4225), .S(n6613), .Z(n3425) );
  NAND2_X1 U4351 ( .A1(n3426), .A2(n3425), .ZN(n3485) );
  INV_X1 U4352 ( .A(n3422), .ZN(n3427) );
  NOR2_X1 U4353 ( .A1(n4277), .A2(n3427), .ZN(n4276) );
  AND2_X1 U4354 ( .A1(n4276), .A2(n3431), .ZN(n3438) );
  NAND2_X1 U4355 ( .A1(n3428), .A2(n3678), .ZN(n4275) );
  AND2_X1 U4356 ( .A1(n3442), .A2(n3422), .ZN(n3430) );
  OR2_X1 U4357 ( .A1(n3430), .A2(n3429), .ZN(n3436) );
  NAND2_X1 U4358 ( .A1(n3439), .A2(n4280), .ZN(n4282) );
  AND2_X1 U4359 ( .A1(n5499), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6658) );
  INV_X1 U4360 ( .A(n6658), .ZN(n3433) );
  AOI21_X1 U4361 ( .B1(n4286), .B2(n3432), .A(n3433), .ZN(n3434) );
  OAI211_X1 U4362 ( .C1(n3417), .C2(n4282), .A(n4579), .B(n3434), .ZN(n3435)
         );
  AOI21_X1 U4363 ( .B1(n4801), .B2(n3436), .A(n3435), .ZN(n3437) );
  OAI211_X1 U4364 ( .C1(n3438), .C2(n6722), .A(n4275), .B(n3437), .ZN(n3486)
         );
  INV_X1 U4365 ( .A(n3530), .ZN(n3459) );
  NAND2_X1 U4366 ( .A1(n3463), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3452) );
  NAND3_X1 U4367 ( .A1(n4446), .A2(n3384), .A3(n3431), .ZN(n3440) );
  NAND2_X1 U4368 ( .A1(n4442), .A2(n4286), .ZN(n4395) );
  INV_X1 U4369 ( .A(n3441), .ZN(n3449) );
  NAND2_X1 U4370 ( .A1(n3418), .A2(n3443), .ZN(n3445) );
  INV_X1 U4371 ( .A(n3717), .ZN(n4458) );
  INV_X1 U4372 ( .A(n4282), .ZN(n4468) );
  NAND3_X1 U4373 ( .A1(n4458), .A2(n4468), .A3(n3384), .ZN(n4467) );
  INV_X1 U4374 ( .A(n4467), .ZN(n3448) );
  NAND2_X1 U4375 ( .A1(n3417), .A2(n3385), .ZN(n4707) );
  INV_X1 U4376 ( .A(n4707), .ZN(n3447) );
  NAND2_X1 U4377 ( .A1(n3448), .A2(n3447), .ZN(n4456) );
  NAND2_X1 U4378 ( .A1(n3450), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3453) );
  INV_X1 U4379 ( .A(n4225), .ZN(n3570) );
  XNOR2_X1 U4380 ( .A(n6613), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6488)
         );
  INV_X1 U4381 ( .A(n3765), .ZN(n3569) );
  AND2_X1 U4382 ( .A1(n3569), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3451)
         );
  AOI21_X1 U4383 ( .B1(n3570), .B2(n6488), .A(n3451), .ZN(n3454) );
  NAND3_X1 U4384 ( .A1(n3452), .A2(n3453), .A3(n3454), .ZN(n3460) );
  INV_X1 U4385 ( .A(n3453), .ZN(n3457) );
  INV_X1 U4386 ( .A(n3454), .ZN(n3455) );
  NOR2_X1 U4387 ( .A1(n3459), .A2(n3531), .ZN(n3462) );
  INV_X1 U4388 ( .A(n3460), .ZN(n3461) );
  NOR2_X2 U4389 ( .A1(n3462), .A2(n3461), .ZN(n3470) );
  NAND2_X1 U4390 ( .A1(n3161), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3468) );
  NAND2_X1 U4391 ( .A1(n3464), .A2(n6623), .ZN(n5022) );
  INV_X1 U4392 ( .A(n3464), .ZN(n3465) );
  NAND2_X1 U4393 ( .A1(n3465), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3466) );
  NAND2_X1 U4394 ( .A1(n5022), .A2(n3466), .ZN(n4941) );
  AOI22_X1 U4395 ( .A1(n3570), .A2(n4941), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3569), .ZN(n3467) );
  AOI22_X1 U4396 ( .A1(n3156), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4397 ( .A1(n4235), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4398 ( .A1(n3331), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3473) );
  AOI22_X1 U4399 ( .A1(n3174), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3472) );
  NAND4_X1 U4400 ( .A1(n3475), .A2(n3474), .A3(n3473), .A4(n3472), .ZN(n3481)
         );
  AOI22_X1 U4401 ( .A1(n4202), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4402 ( .A1(n3168), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U4403 ( .A1(n3166), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4404 ( .A1(n4237), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3476) );
  NAND4_X1 U4405 ( .A1(n3479), .A2(n3478), .A3(n3477), .A4(n3476), .ZN(n3480)
         );
  INV_X1 U4406 ( .A(n3573), .ZN(n3526) );
  INV_X1 U4407 ( .A(n3485), .ZN(n3488) );
  NAND2_X1 U4408 ( .A1(n3488), .A2(n3487), .ZN(n3489) );
  NAND2_X1 U4409 ( .A1(n3489), .A2(n3530), .ZN(n3781) );
  AOI22_X1 U4410 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4202), .B1(n3158), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4411 ( .A1(n3156), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3492) );
  AOI22_X1 U4412 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n3364), .B1(n3170), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U4413 ( .A1(n4235), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        INSTQUEUE_REG_7__0__SCAN_IN), .B2(n4242), .ZN(n3490) );
  NAND4_X1 U4414 ( .A1(n3493), .A2(n3492), .A3(n3491), .A4(n3490), .ZN(n3499)
         );
  AOI22_X1 U4415 ( .A1(n4088), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4416 ( .A1(n3166), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4417 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3167), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4418 ( .A1(n3174), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3494) );
  NAND4_X1 U4419 ( .A1(n3497), .A2(n3496), .A3(n3495), .A4(n3494), .ZN(n3498)
         );
  INV_X1 U4420 ( .A(n3556), .ZN(n3511) );
  AOI22_X1 U4421 ( .A1(n4202), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3504) );
  AOI22_X1 U4422 ( .A1(n3172), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3173), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3503) );
  AOI22_X1 U4423 ( .A1(n3158), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U4424 ( .A1(n4235), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3501) );
  NAND4_X1 U4425 ( .A1(n3504), .A2(n3503), .A3(n3502), .A4(n3501), .ZN(n3510)
         );
  AOI22_X1 U4426 ( .A1(n3168), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4427 ( .A1(n3331), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4428 ( .A1(n3166), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3506) );
  AOI22_X1 U4429 ( .A1(n4237), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3505) );
  NAND4_X1 U4430 ( .A1(n3508), .A2(n3507), .A3(n3506), .A4(n3505), .ZN(n3509)
         );
  XNOR2_X1 U4431 ( .A(n3511), .B(n3676), .ZN(n3512) );
  NAND2_X1 U4432 ( .A1(n3512), .A2(n3532), .ZN(n3541) );
  INV_X1 U4433 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3515) );
  AOI21_X1 U4434 ( .B1(n3711), .B2(n3676), .A(n6659), .ZN(n3514) );
  NAND2_X1 U4435 ( .A1(n3768), .A2(n3556), .ZN(n3513) );
  INV_X1 U4436 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4437 ( .A1(n3167), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4438 ( .A1(n3331), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4439 ( .A1(n4088), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3517) );
  AOI22_X1 U4440 ( .A1(n4235), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3516) );
  NAND4_X1 U4441 ( .A1(n3519), .A2(n3518), .A3(n3517), .A4(n3516), .ZN(n3525)
         );
  AOI22_X1 U4442 ( .A1(n4202), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4443 ( .A1(n3171), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3522) );
  AOI22_X1 U4444 ( .A1(n3175), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3521) );
  AOI22_X1 U4445 ( .A1(n3172), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3520) );
  NAND4_X1 U4446 ( .A1(n3523), .A2(n3522), .A3(n3521), .A4(n3520), .ZN(n3524)
         );
  NAND2_X1 U4447 ( .A1(n3526), .A2(n3555), .ZN(n3528) );
  INV_X1 U4448 ( .A(n3676), .ZN(n3680) );
  NAND2_X1 U4449 ( .A1(n3532), .A2(n3680), .ZN(n3527) );
  NAND2_X1 U4450 ( .A1(n3532), .A2(n3555), .ZN(n3533) );
  NAND2_X1 U4451 ( .A1(n3552), .A2(n3551), .ZN(n3534) );
  NAND2_X1 U4452 ( .A1(n3535), .A2(n3534), .ZN(n3536) );
  INV_X1 U4453 ( .A(n3164), .ZN(n3666) );
  OR2_X1 U4454 ( .A1(n3772), .A2(n3666), .ZN(n3540) );
  NAND2_X1 U4455 ( .A1(n3555), .A2(n3556), .ZN(n3588) );
  XNOR2_X1 U4456 ( .A(n3588), .B(n3587), .ZN(n3538) );
  AND2_X1 U4457 ( .A1(n3768), .A2(n3431), .ZN(n4469) );
  AOI21_X1 U4458 ( .B1(n3538), .B2(n4462), .A(n4469), .ZN(n3539) );
  AND2_X2 U4459 ( .A1(n3540), .A2(n3539), .ZN(n6381) );
  INV_X1 U4460 ( .A(n4469), .ZN(n3545) );
  OAI21_X1 U4461 ( .B1(n6722), .B2(n3556), .A(n3545), .ZN(n3546) );
  INV_X1 U4462 ( .A(n3546), .ZN(n3547) );
  NAND2_X1 U4463 ( .A1(n4550), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3548)
         );
  INV_X1 U4464 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U4465 ( .A1(n3548), .A2(n4902), .ZN(n3550) );
  AND2_X1 U4466 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U4467 ( .A1(n4550), .A2(n3549), .ZN(n3562) );
  NAND2_X1 U4468 ( .A1(n4747), .A2(n3164), .ZN(n3561) );
  OAI21_X1 U4469 ( .B1(n3556), .B2(n3555), .A(n3588), .ZN(n3557) );
  INV_X1 U4470 ( .A(n3557), .ZN(n3559) );
  NAND3_X1 U4471 ( .A1(n4446), .A2(n3373), .A3(n3431), .ZN(n3558) );
  AOI21_X1 U4472 ( .B1(n3559), .B2(n4462), .A(n3558), .ZN(n3560) );
  NAND2_X1 U4473 ( .A1(n3561), .A2(n3560), .ZN(n4645) );
  NAND2_X1 U4474 ( .A1(n4644), .A2(n4645), .ZN(n3563) );
  NAND2_X1 U4475 ( .A1(n6382), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3565)
         );
  AOI21_X2 U4476 ( .B1(n6381), .B2(n3565), .A(n3564), .ZN(n4772) );
  NAND2_X1 U4477 ( .A1(n3161), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3572) );
  NAND3_X1 U4478 ( .A1(n6487), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6484) );
  INV_X1 U4479 ( .A(n6484), .ZN(n3567) );
  NAND2_X1 U4480 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3567), .ZN(n6577) );
  NAND2_X1 U4481 ( .A1(n6487), .A2(n6577), .ZN(n3568) );
  NAND3_X1 U4482 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5320) );
  NAND2_X1 U4483 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6014), .ZN(n6045) );
  AOI22_X1 U4484 ( .A1(n3570), .A2(n4975), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3569), .ZN(n3571) );
  NAND2_X1 U4485 ( .A1(n4711), .A2(n6659), .ZN(n3586) );
  AOI22_X1 U4486 ( .A1(n3167), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4487 ( .A1(n4202), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3577) );
  AOI22_X1 U4488 ( .A1(n3331), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4489 ( .A1(n4058), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3575) );
  NAND4_X1 U4490 ( .A1(n3578), .A2(n3577), .A3(n3576), .A4(n3575), .ZN(n3584)
         );
  AOI22_X1 U4491 ( .A1(n4235), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3582) );
  AOI22_X1 U4492 ( .A1(n3172), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4493 ( .A1(n3171), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4494 ( .A1(n3176), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3579) );
  NAND4_X1 U4495 ( .A1(n3582), .A2(n3581), .A3(n3580), .A4(n3579), .ZN(n3583)
         );
  AOI22_X1 U4496 ( .A1(n3709), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3762), 
        .B2(n3608), .ZN(n3585) );
  NAND2_X1 U4497 ( .A1(n4781), .A2(n3164), .ZN(n3592) );
  NAND2_X1 U4498 ( .A1(n3588), .A2(n3587), .ZN(n3609) );
  INV_X1 U4499 ( .A(n3608), .ZN(n3589) );
  XNOR2_X1 U4500 ( .A(n3609), .B(n3589), .ZN(n3590) );
  NAND2_X1 U4501 ( .A1(n3590), .A2(n4462), .ZN(n3591) );
  INV_X1 U4502 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U4503 ( .A1(n3593), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3594)
         );
  NAND2_X1 U4504 ( .A1(n4774), .A2(n3594), .ZN(n6372) );
  NAND2_X1 U4505 ( .A1(n3709), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3607) );
  AOI22_X1 U4506 ( .A1(n3167), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4507 ( .A1(n4202), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4508 ( .A1(n4235), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4509 ( .A1(n3156), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4510 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3605)
         );
  AOI22_X1 U4511 ( .A1(n3166), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3603) );
  AOI22_X1 U4512 ( .A1(n4236), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3602) );
  AOI22_X1 U4513 ( .A1(n3176), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3601) );
  AOI22_X1 U4514 ( .A1(n3331), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3600) );
  NAND4_X1 U4515 ( .A1(n3603), .A2(n3602), .A3(n3601), .A4(n3600), .ZN(n3604)
         );
  NAND2_X1 U4516 ( .A1(n3762), .A2(n3654), .ZN(n3606) );
  NAND2_X1 U4517 ( .A1(n3805), .A2(n3164), .ZN(n3612) );
  NAND2_X1 U4518 ( .A1(n3609), .A2(n3608), .ZN(n3656) );
  XNOR2_X1 U4519 ( .A(n3656), .B(n3654), .ZN(n3610) );
  NAND2_X1 U4520 ( .A1(n3610), .A2(n4462), .ZN(n3611) );
  NAND2_X1 U4521 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  INV_X1 U4522 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6453) );
  XNOR2_X1 U4523 ( .A(n3613), .B(n6453), .ZN(n6371) );
  NAND2_X1 U4524 ( .A1(n6372), .A2(n6371), .ZN(n6374) );
  NAND2_X1 U4525 ( .A1(n3613), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3614)
         );
  NAND2_X1 U4526 ( .A1(n6374), .A2(n3614), .ZN(n4888) );
  INV_X1 U4527 ( .A(n3636), .ZN(n3615) );
  NAND2_X1 U4528 ( .A1(n3615), .A2(n3637), .ZN(n3628) );
  AOI22_X1 U4529 ( .A1(n3155), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4530 ( .A1(n4235), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3618) );
  AOI22_X1 U4531 ( .A1(n3331), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3617) );
  AOI22_X1 U4532 ( .A1(n3174), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3616) );
  NAND4_X1 U4533 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3626)
         );
  AOI22_X1 U4534 ( .A1(n4202), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4535 ( .A1(n3168), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3623) );
  AOI22_X1 U4536 ( .A1(n3166), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3622) );
  INV_X1 U4537 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4538 ( .A1(n4237), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3621) );
  NAND4_X1 U4539 ( .A1(n3624), .A2(n3623), .A3(n3622), .A4(n3621), .ZN(n3625)
         );
  NAND2_X1 U4540 ( .A1(n3762), .A2(n3653), .ZN(n3627) );
  NAND2_X1 U4541 ( .A1(n3806), .A2(n3164), .ZN(n3633) );
  INV_X1 U4542 ( .A(n3656), .ZN(n3629) );
  NAND2_X1 U4543 ( .A1(n3629), .A2(n3654), .ZN(n3630) );
  XNOR2_X1 U4544 ( .A(n3630), .B(n3653), .ZN(n3631) );
  NAND2_X1 U4545 ( .A1(n3631), .A2(n4462), .ZN(n3632) );
  NAND2_X1 U4546 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  INV_X1 U4547 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4476) );
  XNOR2_X1 U4548 ( .A(n3634), .B(n4476), .ZN(n4890) );
  NAND2_X1 U4549 ( .A1(n4888), .A2(n4890), .ZN(n4889) );
  NAND2_X1 U4550 ( .A1(n3634), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3635)
         );
  NAND2_X1 U4551 ( .A1(n4889), .A2(n3635), .ZN(n4898) );
  AOI22_X1 U4552 ( .A1(n3172), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4553 ( .A1(n4235), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4554 ( .A1(n3331), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4555 ( .A1(n3174), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3639) );
  NAND4_X1 U4556 ( .A1(n3642), .A2(n3641), .A3(n3640), .A4(n3639), .ZN(n3648)
         );
  AOI22_X1 U4557 ( .A1(n4202), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3646) );
  AOI22_X1 U4558 ( .A1(n3168), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3645) );
  AOI22_X1 U4559 ( .A1(n3166), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4560 ( .A1(n4237), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3643) );
  NAND4_X1 U4561 ( .A1(n3646), .A2(n3645), .A3(n3644), .A4(n3643), .ZN(n3647)
         );
  AOI22_X1 U4562 ( .A1(n3709), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3762), 
        .B2(n3669), .ZN(n3651) );
  INV_X1 U4563 ( .A(n3651), .ZN(n3649) );
  NAND2_X1 U4564 ( .A1(n3652), .A2(n3651), .ZN(n3817) );
  NAND2_X1 U4565 ( .A1(n3654), .A2(n3653), .ZN(n3655) );
  OR2_X1 U4566 ( .A1(n3656), .A2(n3655), .ZN(n3668) );
  XNOR2_X1 U4567 ( .A(n3668), .B(n3669), .ZN(n3657) );
  NAND2_X1 U4568 ( .A1(n3657), .A2(n4462), .ZN(n3658) );
  NAND2_X1 U4569 ( .A1(n3659), .A2(n3658), .ZN(n3660) );
  INV_X1 U4570 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4475) );
  XNOR2_X1 U4571 ( .A(n3660), .B(n4475), .ZN(n4897) );
  NAND2_X1 U4572 ( .A1(n4898), .A2(n4897), .ZN(n4896) );
  NAND2_X1 U4573 ( .A1(n3660), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3661)
         );
  NAND2_X1 U4574 ( .A1(n4896), .A2(n3661), .ZN(n5238) );
  INV_X1 U4575 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3663) );
  NAND2_X1 U4576 ( .A1(n3762), .A2(n3676), .ZN(n3662) );
  OAI21_X1 U4577 ( .B1(n3753), .B2(n3663), .A(n3662), .ZN(n3664) );
  INV_X1 U4578 ( .A(n3822), .ZN(n3667) );
  INV_X1 U4579 ( .A(n3668), .ZN(n3670) );
  NAND2_X1 U4580 ( .A1(n3670), .A2(n3669), .ZN(n3681) );
  XNOR2_X1 U4581 ( .A(n3681), .B(n3676), .ZN(n3671) );
  NAND2_X1 U4582 ( .A1(n3671), .A2(n4462), .ZN(n3672) );
  NAND2_X1 U4583 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  INV_X1 U4584 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6430) );
  XNOR2_X1 U4585 ( .A(n3674), .B(n6430), .ZN(n5240) );
  NAND2_X1 U4586 ( .A1(n3674), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3675)
         );
  NAND2_X1 U4587 ( .A1(n3676), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3677) );
  OR3_X1 U4588 ( .A1(n3681), .A2(n3680), .A3(n6722), .ZN(n3682) );
  NAND2_X1 U4589 ( .A1(n5774), .A2(n3682), .ZN(n3683) );
  INV_X1 U4590 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6421) );
  XNOR2_X1 U4591 ( .A(n3683), .B(n6421), .ZN(n5364) );
  INV_X1 U4592 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U4593 ( .A1(n5774), .A2(n6398), .ZN(n5411) );
  OR2_X1 U4594 ( .A1(n5774), .A2(n6398), .ZN(n5412) );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3685) );
  NAND2_X1 U4596 ( .A1(n5774), .A2(n3685), .ZN(n5425) );
  INV_X1 U4597 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3686) );
  INV_X1 U4598 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5466) );
  NOR2_X1 U4599 ( .A1(n6356), .A2(n5466), .ZN(n5448) );
  XNOR2_X1 U4600 ( .A(n6356), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6107)
         );
  NAND2_X1 U4601 ( .A1(n6106), .A2(n6107), .ZN(n3688) );
  NAND2_X1 U4602 ( .A1(n5774), .A2(n6142), .ZN(n3687) );
  INV_X1 U4603 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5833) );
  INV_X1 U4604 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6140) );
  NOR2_X1 U4605 ( .A1(n6356), .A2(n6140), .ZN(n3691) );
  NAND2_X1 U4606 ( .A1(n5774), .A2(n6140), .ZN(n3690) );
  AND2_X1 U4607 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4492) );
  NAND2_X1 U4608 ( .A1(n4492), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3692) );
  INV_X1 U4609 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5953) );
  INV_X1 U4610 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5951) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6127) );
  AND3_X1 U4612 ( .A1(n5953), .A2(n5951), .A3(n6127), .ZN(n3693) );
  OR2_X1 U4613 ( .A1(n5774), .A2(n3693), .ZN(n3694) );
  NOR2_X1 U4614 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3695) );
  INV_X1 U4615 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4495) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5940) );
  INV_X1 U4617 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5903) );
  AND4_X1 U4618 ( .A1(n3695), .A2(n4495), .A3(n5940), .A4(n5903), .ZN(n3696)
         );
  NAND2_X1 U4619 ( .A1(n4434), .A2(n3696), .ZN(n3699) );
  AND2_X1 U4620 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5902) );
  AND2_X1 U4621 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5935) );
  AND2_X1 U4622 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5842) );
  AND3_X1 U4623 ( .A1(n5902), .A2(n5935), .A3(n5842), .ZN(n5845) );
  NAND2_X1 U4624 ( .A1(n5809), .A2(n5845), .ZN(n3697) );
  NAND2_X1 U4625 ( .A1(n3697), .A2(n6356), .ZN(n3698) );
  NAND2_X1 U4626 ( .A1(n3699), .A2(n3698), .ZN(n5742) );
  XNOR2_X1 U4627 ( .A(n6356), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5768)
         );
  NAND2_X1 U4628 ( .A1(n5742), .A2(n5768), .ZN(n4228) );
  INV_X1 U4629 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6116) );
  NAND2_X1 U4630 ( .A1(n5774), .A2(n6116), .ZN(n3700) );
  NAND2_X1 U4631 ( .A1(n4228), .A2(n3700), .ZN(n3704) );
  INV_X1 U4632 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n3701) );
  INV_X1 U4633 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U4634 ( .A1(n3701), .A2(n5892), .ZN(n3702) );
  INV_X1 U4635 ( .A(n4230), .ZN(n3703) );
  INV_X1 U4636 ( .A(n3704), .ZN(n3706) );
  INV_X1 U4637 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U4638 ( .A1(n3706), .A2(n3705), .ZN(n5754) );
  NAND2_X1 U4639 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5846) );
  INV_X1 U4640 ( .A(n5477), .ZN(n3707) );
  XNOR2_X1 U4641 ( .A(n3708), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5875)
         );
  XNOR2_X1 U4642 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3729) );
  INV_X1 U4643 ( .A(n3729), .ZN(n3710) );
  XNOR2_X1 U4644 ( .A(n3710), .B(n3730), .ZN(n4399) );
  NAND2_X1 U4645 ( .A1(n3711), .A2(n3373), .ZN(n3770) );
  INV_X1 U4646 ( .A(n3730), .ZN(n3713) );
  NAND2_X1 U4647 ( .A1(n3169), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4648 ( .A1(n3713), .A2(n3712), .ZN(n3720) );
  INV_X1 U4649 ( .A(n3720), .ZN(n3716) );
  INV_X1 U4650 ( .A(n3714), .ZN(n3715) );
  AOI21_X1 U4651 ( .B1(n3770), .B2(n3716), .A(n3715), .ZN(n3724) );
  NAND2_X1 U4652 ( .A1(n3446), .A2(n3373), .ZN(n3718) );
  NAND2_X1 U4653 ( .A1(n3717), .A2(n3718), .ZN(n3737) );
  AOI21_X1 U4654 ( .B1(n3762), .B2(n4801), .A(n3384), .ZN(n3725) );
  INV_X1 U4655 ( .A(n4399), .ZN(n3719) );
  NAND2_X1 U4656 ( .A1(n3725), .A2(n3719), .ZN(n3723) );
  INV_X1 U4657 ( .A(n3762), .ZN(n3721) );
  OAI21_X1 U4658 ( .B1(n3721), .B2(n3720), .A(n3756), .ZN(n3722) );
  OAI211_X1 U4659 ( .C1(n3724), .C2(n3737), .A(n3723), .B(n3722), .ZN(n3728)
         );
  INV_X1 U4660 ( .A(n3725), .ZN(n3726) );
  NAND3_X1 U4661 ( .A1(n3726), .A2(STATE2_REG_0__SCAN_IN), .A3(n4399), .ZN(
        n3727) );
  OAI211_X1 U4662 ( .C1(n3756), .C2(n4399), .A(n3728), .B(n3727), .ZN(n3735)
         );
  NAND2_X1 U4663 ( .A1(n3730), .A2(n3729), .ZN(n3732) );
  NAND2_X1 U4664 ( .A1(n6618), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3731) );
  NAND2_X1 U4665 ( .A1(n3732), .A2(n3731), .ZN(n3743) );
  XNOR2_X1 U4666 ( .A(n4728), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3741)
         );
  XNOR2_X1 U4667 ( .A(n3743), .B(n3741), .ZN(n4400) );
  INV_X1 U4668 ( .A(n3737), .ZN(n3733) );
  NAND2_X1 U4669 ( .A1(n3762), .A2(n4400), .ZN(n3736) );
  OAI211_X1 U4670 ( .C1(n4400), .C2(n3753), .A(n3733), .B(n3736), .ZN(n3734)
         );
  NAND2_X1 U4671 ( .A1(n3735), .A2(n3734), .ZN(n3740) );
  INV_X1 U4672 ( .A(n3736), .ZN(n3738) );
  NAND2_X1 U4673 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  NAND2_X1 U4674 ( .A1(n3740), .A2(n3739), .ZN(n3755) );
  INV_X1 U4675 ( .A(n3741), .ZN(n3742) );
  NAND2_X1 U4676 ( .A1(n3743), .A2(n3742), .ZN(n3745) );
  NAND2_X1 U4677 ( .A1(n6623), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3744) );
  NAND2_X1 U4678 ( .A1(n3745), .A2(n3744), .ZN(n3748) );
  XNOR2_X1 U4679 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4680 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3757), .ZN(n3746) );
  NOR2_X1 U4681 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n3746), .ZN(n3752)
         );
  NOR2_X1 U4682 ( .A1(n3748), .A2(n3747), .ZN(n3749) );
  OR2_X1 U4683 ( .A1(n3750), .A2(n3749), .ZN(n3751) );
  NAND2_X1 U4684 ( .A1(n4397), .A2(n3753), .ZN(n3754) );
  NAND2_X1 U4685 ( .A1(n3755), .A2(n3754), .ZN(n3761) );
  AOI22_X1 U4686 ( .A1(n4397), .A2(n3758), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6659), .ZN(n3760) );
  OAI222_X1 U4687 ( .A1(n6169), .A2(n3757), .B1(n6169), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3757), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4396) );
  AND2_X1 U4688 ( .A1(n4396), .A2(n3758), .ZN(n3759) );
  NAND2_X1 U4689 ( .A1(n3383), .A2(n3357), .ZN(n3767) );
  AND2_X1 U4690 ( .A1(n4584), .A2(n3768), .ZN(n3769) );
  INV_X1 U4691 ( .A(n3770), .ZN(n3771) );
  INV_X2 U4692 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U4693 ( .A1(n4510), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4115) );
  NAND2_X1 U4694 ( .A1(n3775), .A2(n3944), .ZN(n3780) );
  NAND2_X1 U4695 ( .A1(n3447), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U4696 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3777)
         );
  INV_X2 U4697 ( .A(n3190), .ZN(n4264) );
  NAND2_X1 U4698 ( .A1(n4264), .A2(EAX_REG_1__SCAN_IN), .ZN(n3776) );
  OAI211_X1 U4699 ( .C1(n3801), .C2(n3281), .A(n3777), .B(n3776), .ZN(n3778)
         );
  INV_X1 U4700 ( .A(n3778), .ZN(n3779) );
  NAND2_X1 U4701 ( .A1(n3780), .A2(n3779), .ZN(n4640) );
  NOR2_X4 U4702 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4404) );
  AOI21_X1 U4703 ( .B1(n5969), .B2(n3773), .A(n4510), .ZN(n4627) );
  OR2_X1 U4704 ( .A1(n4752), .A2(n3935), .ZN(n3783) );
  AOI22_X1 U4705 ( .A1(n4264), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4510), .ZN(n3782) );
  OAI211_X1 U4706 ( .C1(n3801), .C2(n3169), .A(n3783), .B(n3782), .ZN(n4626)
         );
  MUX2_X1 U4707 ( .A(n4404), .B(n4627), .S(n4626), .Z(n4641) );
  OAI21_X1 U4708 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3792), .ZN(n6389) );
  AOI22_X1 U4709 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4404), 
        .B2(n6389), .ZN(n3785) );
  NAND2_X1 U4710 ( .A1(n4264), .A2(EAX_REG_2__SCAN_IN), .ZN(n3784) );
  OAI211_X1 U4711 ( .C1(n3801), .C2(n4728), .A(n3785), .B(n3784), .ZN(n3788)
         );
  NAND2_X1 U4712 ( .A1(n3787), .A2(n3788), .ZN(n3786) );
  NAND2_X1 U4713 ( .A1(n4760), .A2(n3786), .ZN(n3790) );
  INV_X1 U4714 ( .A(n3788), .ZN(n4761) );
  NAND2_X1 U4715 ( .A1(n4639), .A2(n4761), .ZN(n3789) );
  AOI21_X1 U4716 ( .B1(n4776), .B2(n3792), .A(n3802), .ZN(n6295) );
  OAI22_X1 U4717 ( .A1(n6295), .A2(n4116), .B1(n4115), .B2(n4776), .ZN(n3793)
         );
  INV_X1 U4718 ( .A(n3793), .ZN(n3795) );
  NAND2_X1 U4719 ( .A1(n4264), .A2(EAX_REG_3__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4720 ( .C1(n3801), .C2(n3791), .A(n3795), .B(n3794), .ZN(n3796)
         );
  NAND2_X1 U4721 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4722 ( .A1(n4264), .A2(EAX_REG_4__SCAN_IN), .ZN(n3799) );
  OAI211_X1 U4723 ( .C1(n3801), .C2(n6169), .A(n3800), .B(n3799), .ZN(n3803)
         );
  OAI21_X1 U4724 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3802), .A(n3810), 
        .ZN(n6379) );
  MUX2_X1 U4725 ( .A(n3803), .B(n6379), .S(n4404), .Z(n3804) );
  NOR2_X2 U4726 ( .A1(n4764), .A2(n4878), .ZN(n4854) );
  NAND2_X1 U4727 ( .A1(n3806), .A2(n3944), .ZN(n3809) );
  XNOR2_X1 U4728 ( .A(n3810), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n4929) );
  OAI22_X1 U4729 ( .A1(n4929), .A2(n4116), .B1(n4115), .B2(n4922), .ZN(n3807)
         );
  AOI21_X1 U4730 ( .B1(n4264), .B2(EAX_REG_5__SCAN_IN), .A(n3807), .ZN(n3808)
         );
  NAND2_X1 U4731 ( .A1(n3809), .A2(n3808), .ZN(n4855) );
  NOR2_X1 U4732 ( .A1(n3811), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3812)
         );
  OR2_X1 U4733 ( .A1(n3833), .A2(n3812), .ZN(n6370) );
  INV_X1 U4734 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3814) );
  INV_X1 U4735 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3813) );
  OAI22_X1 U4736 ( .A1(n3190), .A2(n3814), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3813), .ZN(n3815) );
  MUX2_X1 U4737 ( .A(n6370), .B(n3815), .S(n4116), .Z(n3816) );
  INV_X1 U4738 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3820) );
  XNOR2_X1 U4739 ( .A(n3833), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5242) );
  AOI22_X1 U4740 ( .A1(n5242), .A2(n4404), .B1(n4263), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3819) );
  OAI21_X1 U4741 ( .B1(n3190), .B2(n3820), .A(n3819), .ZN(n3821) );
  AOI22_X1 U4742 ( .A1(n3158), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4743 ( .A1(n3324), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4744 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3364), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4745 ( .A1(n3172), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3823) );
  NAND4_X1 U4746 ( .A1(n3826), .A2(n3825), .A3(n3824), .A4(n3823), .ZN(n3832)
         );
  AOI22_X1 U4747 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4235), .B1(n3331), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4748 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3167), .B1(n3166), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4749 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n4202), .B1(n4088), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4750 ( .A1(n3171), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3827) );
  NAND4_X1 U4751 ( .A1(n3830), .A2(n3829), .A3(n3828), .A4(n3827), .ZN(n3831)
         );
  OAI21_X1 U4752 ( .B1(n3832), .B2(n3831), .A(n3944), .ZN(n3837) );
  NAND2_X1 U4753 ( .A1(n4264), .A2(EAX_REG_8__SCAN_IN), .ZN(n3836) );
  XNOR2_X1 U4754 ( .A(n3838), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U4755 ( .A1(n5367), .A2(n4404), .ZN(n3835) );
  NAND2_X1 U4756 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3834)
         );
  NAND4_X1 U4757 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n5249)
         );
  NAND2_X1 U4758 ( .A1(n5246), .A2(n5249), .ZN(n5247) );
  INV_X1 U4759 ( .A(n5247), .ZN(n3855) );
  XNOR2_X1 U4760 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3857), .ZN(n6244) );
  INV_X1 U4761 ( .A(n6244), .ZN(n3853) );
  AOI22_X1 U4762 ( .A1(n3155), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4763 ( .A1(n4088), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4764 ( .A1(n3166), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4765 ( .A1(n4235), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4766 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4767 ( .A1(n3168), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4768 ( .A1(n3324), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4769 ( .A1(n4058), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4770 ( .A1(n3176), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4771 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  OAI21_X1 U4772 ( .B1(n3848), .B2(n3847), .A(n3944), .ZN(n3851) );
  NAND2_X1 U4773 ( .A1(n4264), .A2(EAX_REG_9__SCAN_IN), .ZN(n3850) );
  NAND2_X1 U4774 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3849)
         );
  NAND3_X1 U4775 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(n3852) );
  AOI21_X1 U4776 ( .B1(n3853), .B2(n4404), .A(n3852), .ZN(n5359) );
  NAND2_X1 U4777 ( .A1(n3855), .A2(n3854), .ZN(n5358) );
  XNOR2_X1 U4778 ( .A(n3872), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5644)
         );
  AOI22_X1 U4779 ( .A1(n3331), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4780 ( .A1(n4202), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4781 ( .A1(n3168), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4782 ( .A1(n4235), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4783 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3867)
         );
  AOI22_X1 U4784 ( .A1(n3155), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4785 ( .A1(n3174), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4786 ( .A1(n3166), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4787 ( .A1(n4237), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4788 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3866)
         );
  OAI21_X1 U4789 ( .B1(n3867), .B2(n3866), .A(n3944), .ZN(n3870) );
  NAND2_X1 U4790 ( .A1(n4264), .A2(EAX_REG_10__SCAN_IN), .ZN(n3869) );
  NAND2_X1 U4791 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3868)
         );
  NAND3_X1 U4792 ( .A1(n3870), .A2(n3869), .A3(n3868), .ZN(n3871) );
  AOI21_X1 U4793 ( .B1(n5644), .B2(n4404), .A(n3871), .ZN(n5420) );
  NOR2_X2 U4794 ( .A1(n5358), .A2(n5420), .ZN(n5418) );
  XNOR2_X1 U4795 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3886), .ZN(n6359)
         );
  AOI22_X1 U4796 ( .A1(n3166), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4797 ( .A1(n4202), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4798 ( .A1(n3167), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4799 ( .A1(n3175), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3873) );
  NAND4_X1 U4800 ( .A1(n3876), .A2(n3875), .A3(n3874), .A4(n3873), .ZN(n3882)
         );
  AOI22_X1 U4801 ( .A1(n3331), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4802 ( .A1(n4235), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4803 ( .A1(n4088), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4804 ( .A1(n3156), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3877) );
  NAND4_X1 U4805 ( .A1(n3880), .A2(n3879), .A3(n3878), .A4(n3877), .ZN(n3881)
         );
  OR2_X1 U4806 ( .A1(n3882), .A2(n3881), .ZN(n3883) );
  AOI22_X1 U4807 ( .A1(n3944), .A2(n3883), .B1(n4263), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3885) );
  NAND2_X1 U4808 ( .A1(n4264), .A2(EAX_REG_11__SCAN_IN), .ZN(n3884) );
  OAI211_X1 U4809 ( .C1(n6359), .C2(n4116), .A(n3885), .B(n3884), .ZN(n5431)
         );
  XNOR2_X1 U4810 ( .A(n3902), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5452)
         );
  NAND2_X1 U4811 ( .A1(n5452), .A2(n4404), .ZN(n3901) );
  AOI22_X1 U4812 ( .A1(n3178), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4813 ( .A1(n3168), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4814 ( .A1(n3166), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4815 ( .A1(n4235), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4816 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3896)
         );
  AOI22_X1 U4817 ( .A1(n3156), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4818 ( .A1(n4202), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4819 ( .A1(n3331), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4820 ( .A1(n4237), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3891) );
  NAND4_X1 U4821 ( .A1(n3894), .A2(n3893), .A3(n3892), .A4(n3891), .ZN(n3895)
         );
  OAI21_X1 U4822 ( .B1(n3896), .B2(n3895), .A(n3944), .ZN(n3899) );
  NAND2_X1 U4823 ( .A1(n4264), .A2(EAX_REG_12__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U4824 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3897)
         );
  AND3_X1 U4825 ( .A1(n3899), .A2(n3898), .A3(n3897), .ZN(n3900) );
  INV_X1 U4826 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3905) );
  OAI21_X1 U4827 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3903), .A(n3947), 
        .ZN(n6226) );
  NAND2_X1 U4828 ( .A1(n6226), .A2(n4404), .ZN(n3904) );
  OAI21_X1 U4829 ( .B1(n3905), .B2(n4115), .A(n3904), .ZN(n3906) );
  INV_X1 U4830 ( .A(n5735), .ZN(n3920) );
  AOI22_X1 U4831 ( .A1(n3155), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4832 ( .A1(n3167), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4833 ( .A1(n4202), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4834 ( .A1(n3171), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3908) );
  NAND4_X1 U4835 ( .A1(n3911), .A2(n3910), .A3(n3909), .A4(n3908), .ZN(n3917)
         );
  AOI22_X1 U4836 ( .A1(n4235), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4837 ( .A1(n3176), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3914) );
  AOI22_X1 U4838 ( .A1(n4237), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4839 ( .A1(n4088), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3912) );
  NAND4_X1 U4840 ( .A1(n3915), .A2(n3914), .A3(n3913), .A4(n3912), .ZN(n3916)
         );
  OR2_X1 U4841 ( .A1(n3917), .A2(n3916), .ZN(n3918) );
  NAND2_X1 U4842 ( .A1(n3944), .A2(n3918), .ZN(n5736) );
  NAND2_X1 U4843 ( .A1(n3920), .A2(n3919), .ZN(n5734) );
  AOI22_X1 U4844 ( .A1(n3176), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4845 ( .A1(n3168), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4846 ( .A1(n4236), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4847 ( .A1(n3166), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4848 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3931)
         );
  AOI22_X1 U4849 ( .A1(n3324), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4850 ( .A1(n3156), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4851 ( .A1(n4202), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4852 ( .A1(n4235), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4853 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  NOR2_X1 U4854 ( .A1(n3931), .A2(n3930), .ZN(n3934) );
  XNOR2_X1 U4855 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3947), .ZN(n5838)
         );
  INV_X1 U4856 ( .A(n5838), .ZN(n6211) );
  AOI22_X1 U4857 ( .A1(n4263), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n4404), 
        .B2(n6211), .ZN(n3933) );
  NAND2_X1 U4858 ( .A1(n4264), .A2(EAX_REG_14__SCAN_IN), .ZN(n3932) );
  OAI211_X1 U4859 ( .C1(n3935), .C2(n3934), .A(n3933), .B(n3932), .ZN(n5706)
         );
  AOI22_X1 U4860 ( .A1(n3168), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4861 ( .A1(n4202), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4862 ( .A1(n3172), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4863 ( .A1(n3331), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4864 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3946)
         );
  AOI22_X1 U4865 ( .A1(n4235), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4866 ( .A1(n3158), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4867 ( .A1(n3166), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4868 ( .A1(n3170), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4869 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3945)
         );
  OAI21_X1 U4870 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n3951) );
  NAND2_X1 U4871 ( .A1(n4264), .A2(EAX_REG_15__SCAN_IN), .ZN(n3950) );
  INV_X1 U4872 ( .A(n3952), .ZN(n3948) );
  XNOR2_X1 U4873 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3948), .ZN(n5827)
         );
  AOI22_X1 U4874 ( .A1(n4404), .A2(n5827), .B1(n4263), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3949) );
  INV_X1 U4875 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5627) );
  XNOR2_X1 U4876 ( .A(n5627), .B(n3965), .ZN(n5819) );
  AOI22_X1 U4877 ( .A1(n4264), .A2(EAX_REG_16__SCAN_IN), .B1(n4263), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4878 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3177), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4879 ( .A1(n4088), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4880 ( .A1(n3167), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4881 ( .A1(n3170), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3953) );
  NAND4_X1 U4882 ( .A1(n3956), .A2(n3955), .A3(n3954), .A4(n3953), .ZN(n3962)
         );
  AOI22_X1 U4883 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n4235), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4884 ( .A1(n3156), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3158), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4885 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n4202), .B1(n3166), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4886 ( .A1(n4237), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4887 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3961)
         );
  OAI21_X1 U4888 ( .B1(n3962), .B2(n3961), .A(n4213), .ZN(n3963) );
  OAI211_X1 U4889 ( .C1(n5819), .C2(n4116), .A(n3964), .B(n3963), .ZN(n5617)
         );
  XNOR2_X1 U4890 ( .A(n3984), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6103)
         );
  NAND2_X1 U4891 ( .A1(n6103), .A2(n4404), .ZN(n3981) );
  AOI22_X1 U4892 ( .A1(n4235), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4893 ( .A1(n3158), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4894 ( .A1(n3324), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4895 ( .A1(n3172), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4896 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3977)
         );
  AOI22_X1 U4897 ( .A1(n3166), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4898 ( .A1(n3174), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4899 ( .A1(n4202), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3971)
         );
  AOI21_X1 U4900 ( .B1(n4242), .B2(INSTQUEUE_REG_9__1__SCAN_IN), .A(n4404), 
        .ZN(n3970) );
  AND2_X1 U4901 ( .A1(n3971), .A2(n3970), .ZN(n3973) );
  AOI22_X1 U4902 ( .A1(n3168), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3972) );
  NAND4_X1 U4903 ( .A1(n3975), .A2(n3974), .A3(n3973), .A4(n3972), .ZN(n3976)
         );
  NAND2_X1 U4904 ( .A1(n4256), .A2(n4116), .ZN(n4046) );
  OAI21_X1 U4905 ( .B1(n3977), .B2(n3976), .A(n4046), .ZN(n3979) );
  AOI22_X1 U4906 ( .A1(n4264), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4510), .ZN(n3978) );
  NAND2_X1 U4907 ( .A1(n3979), .A2(n3978), .ZN(n3980) );
  NAND2_X1 U4908 ( .A1(n3981), .A2(n3980), .ZN(n5604) );
  NAND2_X1 U4909 ( .A1(n3983), .A2(n3982), .ZN(n5693) );
  OR2_X1 U4910 ( .A1(n3985), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3986)
         );
  NAND2_X1 U4911 ( .A1(n3986), .A2(n4018), .ZN(n6207) );
  AOI22_X1 U4912 ( .A1(n3172), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4913 ( .A1(n4202), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4914 ( .A1(n3166), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4915 ( .A1(n3177), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U4916 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3996)
         );
  AOI22_X1 U4917 ( .A1(n3176), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4918 ( .A1(n3171), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4919 ( .A1(n3168), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4920 ( .A1(n4235), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4921 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n3995)
         );
  NOR2_X1 U4922 ( .A1(n3996), .A2(n3995), .ZN(n3997) );
  NOR2_X1 U4923 ( .A1(n4256), .A2(n3997), .ZN(n4001) );
  INV_X1 U4924 ( .A(EAX_REG_18__SCAN_IN), .ZN(n3999) );
  NAND2_X1 U4925 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n3998)
         );
  OAI211_X1 U4926 ( .C1(n3190), .C2(n3999), .A(n4116), .B(n3998), .ZN(n4000)
         );
  OAI22_X1 U4927 ( .A1(n6207), .A2(n4116), .B1(n4001), .B2(n4000), .ZN(n5694)
         );
  AOI22_X1 U4928 ( .A1(n3172), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3167), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4929 ( .A1(n4235), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4930 ( .A1(n3331), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4931 ( .A1(n4088), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4002) );
  NAND4_X1 U4932 ( .A1(n4005), .A2(n4004), .A3(n4003), .A4(n4002), .ZN(n4013)
         );
  AOI22_X1 U4933 ( .A1(n3175), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4934 ( .A1(n3177), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4935 ( .A1(n3364), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4009) );
  NAND2_X1 U4936 ( .A1(n4202), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4007)
         );
  AOI21_X1 U4937 ( .B1(n4242), .B2(INSTQUEUE_REG_9__3__SCAN_IN), .A(n4404), 
        .ZN(n4006) );
  AND2_X1 U4938 ( .A1(n4007), .A2(n4006), .ZN(n4008) );
  NAND4_X1 U4939 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4012)
         );
  OAI21_X1 U4940 ( .B1(n4013), .B2(n4012), .A(n4046), .ZN(n4015) );
  AOI22_X1 U4941 ( .A1(n4264), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4510), .ZN(n4014) );
  NAND2_X1 U4942 ( .A1(n4015), .A2(n4014), .ZN(n4017) );
  XNOR2_X1 U4943 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .B(n4018), .ZN(n5588)
         );
  NAND2_X1 U4944 ( .A1(n4404), .A2(n5588), .ZN(n4016) );
  NAND2_X1 U4945 ( .A1(n4017), .A2(n4016), .ZN(n5587) );
  NOR2_X2 U4946 ( .A1(n3159), .A2(n5693), .ZN(n5585) );
  OR2_X1 U4947 ( .A1(n4019), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4020)
         );
  NAND2_X1 U4948 ( .A1(n4020), .A2(n4069), .ZN(n5806) );
  INV_X1 U4949 ( .A(n5806), .ZN(n6080) );
  AOI22_X1 U4950 ( .A1(n4235), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4951 ( .A1(n3176), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4952 ( .A1(n3167), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4953 ( .A1(n3166), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U4954 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4030)
         );
  AOI22_X1 U4955 ( .A1(n3331), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4028) );
  AOI22_X1 U4956 ( .A1(n3156), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4957 ( .A1(n3171), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4958 ( .A1(n4202), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4025) );
  NAND4_X1 U4959 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4029)
         );
  OR2_X1 U4960 ( .A1(n4030), .A2(n4029), .ZN(n4034) );
  INV_X1 U4961 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4032) );
  NAND2_X1 U4962 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4031)
         );
  OAI211_X1 U4963 ( .C1(n3190), .C2(n4032), .A(n4116), .B(n4031), .ZN(n4033)
         );
  AOI21_X1 U4964 ( .B1(n4213), .B2(n4034), .A(n4033), .ZN(n4035) );
  AOI21_X1 U4965 ( .B1(n6080), .B2(n4404), .A(n4035), .ZN(n5680) );
  AOI22_X1 U4966 ( .A1(n3175), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4967 ( .A1(n4088), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4038) );
  AOI22_X1 U4968 ( .A1(n4235), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4969 ( .A1(n4202), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4036) );
  NAND4_X1 U4970 ( .A1(n4039), .A2(n4038), .A3(n4037), .A4(n4036), .ZN(n4048)
         );
  AOI22_X1 U4971 ( .A1(n3168), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4972 ( .A1(n3156), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4973 ( .A1(n3331), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4043) );
  NAND2_X1 U4974 ( .A1(n3364), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4041) );
  AOI21_X1 U4975 ( .B1(n4242), .B2(INSTQUEUE_REG_9__5__SCAN_IN), .A(n4404), 
        .ZN(n4040) );
  AND2_X1 U4976 ( .A1(n4041), .A2(n4040), .ZN(n4042) );
  NAND4_X1 U4977 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4047)
         );
  OAI21_X1 U4978 ( .B1(n4048), .B2(n4047), .A(n4046), .ZN(n4050) );
  AOI22_X1 U4979 ( .A1(n4264), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n4510), .ZN(n4049) );
  NAND2_X1 U4980 ( .A1(n4050), .A2(n4049), .ZN(n4052) );
  XNOR2_X1 U4981 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4069), .ZN(n5798)
         );
  NAND2_X1 U4982 ( .A1(n4404), .A2(n5798), .ZN(n4051) );
  NAND2_X1 U4983 ( .A1(n4052), .A2(n4051), .ZN(n5571) );
  AOI22_X1 U4984 ( .A1(n3167), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3166), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4985 ( .A1(n4202), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4986 ( .A1(n3331), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4987 ( .A1(n3156), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4054) );
  NAND4_X1 U4988 ( .A1(n4057), .A2(n4056), .A3(n4055), .A4(n4054), .ZN(n4064)
         );
  AOI22_X1 U4989 ( .A1(n3158), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4990 ( .A1(n4088), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4991 ( .A1(n4235), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U4992 ( .A1(n3324), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U4993 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  NOR2_X1 U4994 ( .A1(n4064), .A2(n4063), .ZN(n4068) );
  NAND2_X1 U4995 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4065)
         );
  NAND2_X1 U4996 ( .A1(n4116), .A2(n4065), .ZN(n4066) );
  AOI21_X1 U4997 ( .B1(n4264), .B2(EAX_REG_22__SCAN_IN), .A(n4066), .ZN(n4067)
         );
  OAI21_X1 U4998 ( .B1(n4256), .B2(n4068), .A(n4067), .ZN(n4073) );
  OAI21_X1 U4999 ( .B1(n4071), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4114), 
        .ZN(n5790) );
  OR2_X1 U5000 ( .A1(n5790), .A2(n4116), .ZN(n4072) );
  NAND2_X1 U5001 ( .A1(n4073), .A2(n4072), .ZN(n5556) );
  AOI22_X1 U5002 ( .A1(n4235), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5003 ( .A1(n3155), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5004 ( .A1(n4088), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5005 ( .A1(n4058), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5006 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4083)
         );
  AOI22_X1 U5007 ( .A1(n3167), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5008 ( .A1(n3175), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5009 ( .A1(n3171), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5010 ( .A1(n3166), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4078) );
  NAND4_X1 U5011 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .ZN(n4082)
         );
  NOR2_X1 U5012 ( .A1(n4083), .A2(n4082), .ZN(n4101) );
  AOI22_X1 U5013 ( .A1(n3168), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4202), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5014 ( .A1(n3155), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4086) );
  AOI22_X1 U5015 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n3170), .B1(n4058), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5016 ( .A1(n4235), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4084) );
  NAND4_X1 U5017 ( .A1(n4087), .A2(n4086), .A3(n4085), .A4(n4084), .ZN(n4094)
         );
  AOI22_X1 U5018 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n3324), .B1(n3331), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4092) );
  AOI22_X1 U5019 ( .A1(n4088), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5020 ( .A1(n3166), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5021 ( .A1(n3158), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4089) );
  NAND4_X1 U5022 ( .A1(n4092), .A2(n4091), .A3(n4090), .A4(n4089), .ZN(n4093)
         );
  NOR2_X1 U5023 ( .A1(n4094), .A2(n4093), .ZN(n4100) );
  XOR2_X1 U5024 ( .A(n4101), .B(n4100), .Z(n4095) );
  NAND2_X1 U5025 ( .A1(n4095), .A2(n4213), .ZN(n4099) );
  OAI21_X1 U5026 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4503), .A(n4116), .ZN(
        n4096) );
  AOI21_X1 U5027 ( .B1(n4264), .B2(EAX_REG_23__SCAN_IN), .A(n4096), .ZN(n4098)
         );
  XNOR2_X1 U5028 ( .A(n4114), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6069)
         );
  AND2_X1 U5029 ( .A1(n6069), .A2(n4404), .ZN(n4097) );
  AOI21_X1 U5030 ( .B1(n4099), .B2(n4098), .A(n4097), .ZN(n4501) );
  NOR2_X1 U5031 ( .A1(n4101), .A2(n4100), .ZN(n4133) );
  AOI22_X1 U5032 ( .A1(n3172), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5033 ( .A1(n4235), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5034 ( .A1(n3331), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5035 ( .A1(n3174), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U5036 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4111)
         );
  AOI22_X1 U5037 ( .A1(n4202), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5038 ( .A1(n3167), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5039 ( .A1(n3166), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U5040 ( .A1(n4237), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U5041 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4110)
         );
  OR2_X1 U5042 ( .A1(n4111), .A2(n4110), .ZN(n4132) );
  INV_X1 U5043 ( .A(n4132), .ZN(n4112) );
  XNOR2_X1 U5044 ( .A(n4133), .B(n4112), .ZN(n4113) );
  NAND2_X1 U5045 ( .A1(n4113), .A2(n4213), .ZN(n4119) );
  INV_X1 U5046 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5780) );
  XNOR2_X1 U5047 ( .A(n4138), .B(n5780), .ZN(n5784) );
  OAI22_X1 U5048 ( .A1(n5784), .A2(n4116), .B1(n5780), .B2(n4115), .ZN(n4117)
         );
  AOI21_X1 U5049 ( .B1(n4264), .B2(EAX_REG_24__SCAN_IN), .A(n4117), .ZN(n4118)
         );
  NAND2_X1 U5050 ( .A1(n4119), .A2(n4118), .ZN(n5545) );
  NAND2_X1 U5051 ( .A1(n4500), .A2(n5545), .ZN(n5544) );
  AOI22_X1 U5052 ( .A1(n3155), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3175), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5053 ( .A1(n4235), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5054 ( .A1(n3331), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4122) );
  AOI22_X1 U5055 ( .A1(n3174), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4121) );
  NAND4_X1 U5056 ( .A1(n4124), .A2(n4123), .A3(n4122), .A4(n4121), .ZN(n4131)
         );
  AOI22_X1 U5057 ( .A1(n4202), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5058 ( .A1(n3168), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U5059 ( .A1(n3166), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U5060 ( .A1(n4237), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4126) );
  NAND4_X1 U5061 ( .A1(n4129), .A2(n4128), .A3(n4127), .A4(n4126), .ZN(n4130)
         );
  NOR2_X1 U5062 ( .A1(n4131), .A2(n4130), .ZN(n4144) );
  NAND2_X1 U5063 ( .A1(n4133), .A2(n4132), .ZN(n4143) );
  XOR2_X1 U5064 ( .A(n4144), .B(n4143), .Z(n4134) );
  NAND2_X1 U5065 ( .A1(n4134), .A2(n4213), .ZN(n4137) );
  INV_X1 U5066 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5766) );
  OAI21_X1 U5067 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5766), .A(n4116), .ZN(
        n4135) );
  AOI21_X1 U5068 ( .B1(n4264), .B2(EAX_REG_25__SCAN_IN), .A(n4135), .ZN(n4136)
         );
  NAND2_X1 U5069 ( .A1(n4137), .A2(n4136), .ZN(n4140) );
  NAND2_X1 U5070 ( .A1(n4138), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4158)
         );
  XNOR2_X1 U5071 ( .A(n4158), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6061)
         );
  NAND2_X1 U5072 ( .A1(n6061), .A2(n4404), .ZN(n4139) );
  NAND2_X1 U5073 ( .A1(n4140), .A2(n4139), .ZN(n5669) );
  NOR2_X1 U5074 ( .A1(n4144), .A2(n4143), .ZN(n4166) );
  AOI22_X1 U5075 ( .A1(n3155), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5076 ( .A1(n4235), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3178), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5077 ( .A1(n3331), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3171), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5078 ( .A1(n3174), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U5079 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4154)
         );
  AOI22_X1 U5080 ( .A1(n4202), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5081 ( .A1(n3168), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5082 ( .A1(n3166), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5083 ( .A1(n4237), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4149) );
  NAND4_X1 U5084 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  XNOR2_X1 U5085 ( .A(n4166), .B(n4165), .ZN(n4157) );
  OAI21_X1 U5086 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4159), .A(n4116), .ZN(
        n4155) );
  AOI21_X1 U5087 ( .B1(n4264), .B2(EAX_REG_26__SCAN_IN), .A(n4155), .ZN(n4156)
         );
  OAI21_X1 U5088 ( .B1(n4157), .B2(n4256), .A(n4156), .ZN(n4164) );
  AND2_X1 U5089 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  INV_X1 U5090 ( .A(n6059), .ZN(n4162) );
  NAND2_X1 U5091 ( .A1(n4162), .A2(n4404), .ZN(n4163) );
  NAND2_X1 U5092 ( .A1(n4164), .A2(n4163), .ZN(n5660) );
  NAND2_X1 U5093 ( .A1(n4166), .A2(n4165), .ZN(n4184) );
  AOI22_X1 U5094 ( .A1(n4235), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U5095 ( .A1(n4202), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4169) );
  AOI22_X1 U5096 ( .A1(n3166), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5097 ( .A1(n4237), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4167) );
  NAND4_X1 U5098 ( .A1(n4170), .A2(n4169), .A3(n4168), .A4(n4167), .ZN(n4176)
         );
  AOI22_X1 U5099 ( .A1(n3155), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5100 ( .A1(n3177), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4173) );
  AOI22_X1 U5101 ( .A1(n3167), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4058), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5102 ( .A1(n3171), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4171) );
  NAND4_X1 U5103 ( .A1(n4174), .A2(n4173), .A3(n4172), .A4(n4171), .ZN(n4175)
         );
  NOR2_X1 U5104 ( .A1(n4176), .A2(n4175), .ZN(n4185) );
  XOR2_X1 U5105 ( .A(n4184), .B(n4185), .Z(n4177) );
  NAND2_X1 U5106 ( .A1(n4177), .A2(n4213), .ZN(n4180) );
  INV_X1 U5107 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5750) );
  NOR2_X1 U5108 ( .A1(n5750), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4178) );
  AOI211_X1 U5109 ( .C1(n4264), .C2(EAX_REG_27__SCAN_IN), .A(n4404), .B(n4178), 
        .ZN(n4179) );
  XOR2_X1 U5110 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .B(n4181), .Z(n5752) );
  OR2_X1 U5111 ( .A1(n4182), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4183)
         );
  NAND2_X1 U5112 ( .A1(n4259), .A2(n4183), .ZN(n5746) );
  NOR2_X1 U5113 ( .A1(n4185), .A2(n4184), .ZN(n4201) );
  AOI22_X1 U5114 ( .A1(n3155), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3176), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4189) );
  AOI22_X1 U5115 ( .A1(n4235), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4188) );
  AOI22_X1 U5116 ( .A1(n3331), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3170), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5117 ( .A1(n3174), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4186) );
  NAND4_X1 U5118 ( .A1(n4189), .A2(n4188), .A3(n4187), .A4(n4186), .ZN(n4195)
         );
  AOI22_X1 U5119 ( .A1(n4202), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4088), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4193) );
  AOI22_X1 U5120 ( .A1(n3168), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4192) );
  AOI22_X1 U5121 ( .A1(n3166), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4191) );
  AOI22_X1 U5122 ( .A1(n4237), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4190) );
  NAND4_X1 U5123 ( .A1(n4193), .A2(n4192), .A3(n4191), .A4(n4190), .ZN(n4194)
         );
  OR2_X1 U5124 ( .A1(n4195), .A2(n4194), .ZN(n4200) );
  XNOR2_X1 U5125 ( .A(n4201), .B(n4200), .ZN(n4198) );
  AOI21_X1 U5126 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4510), .A(n4404), 
        .ZN(n4197) );
  NAND2_X1 U5127 ( .A1(n4264), .A2(EAX_REG_28__SCAN_IN), .ZN(n4196) );
  OAI211_X1 U5128 ( .C1(n4198), .C2(n4256), .A(n4197), .B(n4196), .ZN(n4199)
         );
  OAI21_X1 U5129 ( .B1(n4116), .B2(n5746), .A(n4199), .ZN(n5520) );
  NAND2_X1 U5130 ( .A1(n4201), .A2(n4200), .ZN(n4249) );
  AOI22_X1 U5131 ( .A1(n4235), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5132 ( .A1(n4202), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5133 ( .A1(n3172), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4204) );
  AOI22_X1 U5134 ( .A1(n3386), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4203) );
  NAND4_X1 U5135 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n4212)
         );
  AOI22_X1 U5136 ( .A1(n3158), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4210) );
  AOI22_X1 U5137 ( .A1(n3166), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3324), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4209) );
  AOI22_X1 U5138 ( .A1(n3168), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3364), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4208) );
  AOI22_X1 U5139 ( .A1(n3171), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4207) );
  NAND4_X1 U5140 ( .A1(n4210), .A2(n4209), .A3(n4208), .A4(n4207), .ZN(n4211)
         );
  NOR2_X1 U5141 ( .A1(n4212), .A2(n4211), .ZN(n4250) );
  XOR2_X1 U5142 ( .A(n4249), .B(n4250), .Z(n4214) );
  NAND2_X1 U5143 ( .A1(n4214), .A2(n4213), .ZN(n4217) );
  INV_X1 U5144 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4258) );
  NOR2_X1 U5145 ( .A1(n4258), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4215) );
  AOI211_X1 U5146 ( .C1(n4264), .C2(EAX_REG_29__SCAN_IN), .A(n4404), .B(n4215), 
        .ZN(n4216) );
  XNOR2_X1 U5147 ( .A(n4259), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5511)
         );
  AND2_X1 U5148 ( .A1(n6659), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4405) );
  NAND2_X1 U5149 ( .A1(n4405), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6665) );
  NAND2_X1 U5150 ( .A1(n4225), .A2(n6496), .ZN(n6718) );
  NAND2_X1 U5151 ( .A1(n6718), .A2(n6659), .ZN(n4221) );
  NAND2_X1 U5152 ( .A1(n6659), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4223) );
  INV_X1 U5153 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6177) );
  NAND2_X1 U5154 ( .A1(n6177), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4222) );
  AND2_X1 U5155 ( .A1(n4223), .A2(n4222), .ZN(n4628) );
  INV_X1 U5156 ( .A(n4628), .ZN(n4224) );
  INV_X2 U5157 ( .A(n6454), .ZN(n6476) );
  NAND2_X1 U5158 ( .A1(n6476), .A2(REIP_REG_29__SCAN_IN), .ZN(n5868) );
  OAI21_X1 U5159 ( .B1(n5836), .B2(n4258), .A(n5868), .ZN(n4226) );
  AOI21_X1 U5160 ( .B1(n5511), .B2(n6360), .A(n4226), .ZN(n4227) );
  OAI211_X1 U5161 ( .C1(n5875), .C2(n6364), .A(n3184), .B(n4227), .ZN(U2957)
         );
  AND2_X1 U5162 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5847) );
  INV_X1 U5164 ( .A(n4229), .ZN(n4232) );
  NOR3_X1 U5165 ( .A1(n4230), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4231) );
  AOI22_X1 U5166 ( .A1(n5477), .A2(n5847), .B1(n4232), .B2(n4231), .ZN(n4234)
         );
  AOI22_X1 U5167 ( .A1(n4235), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5168 ( .A1(n4202), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3154), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4240) );
  AOI22_X1 U5169 ( .A1(n3166), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4239) );
  AOI22_X1 U5170 ( .A1(n3178), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4238) );
  NAND4_X1 U5171 ( .A1(n4241), .A2(n4240), .A3(n4239), .A4(n4238), .ZN(n4248)
         );
  AOI22_X1 U5172 ( .A1(n3158), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3174), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4246) );
  AOI22_X1 U5173 ( .A1(n3167), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3386), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4245) );
  AOI22_X1 U5174 ( .A1(n3170), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4242), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4244) );
  AOI22_X1 U5175 ( .A1(n3156), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4125), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4243) );
  NAND4_X1 U5176 ( .A1(n4246), .A2(n4245), .A3(n4244), .A4(n4243), .ZN(n4247)
         );
  NOR2_X1 U5177 ( .A1(n4248), .A2(n4247), .ZN(n4252) );
  NOR2_X1 U5178 ( .A1(n4250), .A2(n4249), .ZN(n4251) );
  XOR2_X1 U5179 ( .A(n4252), .B(n4251), .Z(n4257) );
  NAND2_X1 U5180 ( .A1(n4510), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4253)
         );
  NAND2_X1 U5181 ( .A1(n4116), .A2(n4253), .ZN(n4254) );
  AOI21_X1 U5182 ( .B1(n4264), .B2(EAX_REG_30__SCAN_IN), .A(n4254), .ZN(n4255)
         );
  OAI21_X1 U5183 ( .B1(n4257), .B2(n4256), .A(n4255), .ZN(n4261) );
  INV_X1 U5184 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4267) );
  XNOR2_X1 U5185 ( .A(n4268), .B(n4267), .ZN(n5486) );
  NAND2_X1 U5186 ( .A1(n4261), .A2(n4260), .ZN(n4274) );
  AOI22_X1 U5187 ( .A1(n4264), .A2(EAX_REG_31__SCAN_IN), .B1(n4263), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4265) );
  INV_X1 U5188 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4269) );
  INV_X1 U5189 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6872) );
  NOR2_X1 U5190 ( .A1(n6454), .A2(n6872), .ZN(n5848) );
  AOI21_X1 U5191 ( .B1(n6380), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5848), 
        .ZN(n4271) );
  OAI21_X1 U5192 ( .B1(n6390), .B2(n4914), .A(n4271), .ZN(n4272) );
  AOI21_X1 U5193 ( .B1(n5712), .B2(n6385), .A(n4272), .ZN(n4273) );
  OR2_X1 U5194 ( .A1(n4276), .A2(n6722), .ZN(n4279) );
  NAND3_X1 U5195 ( .A1(n4277), .A2(n4286), .A3(n3422), .ZN(n4278) );
  NAND2_X2 U5196 ( .A1(n3431), .A2(n4287), .ZN(n4324) );
  OAI21_X1 U5197 ( .B1(n4707), .B2(n4286), .A(n3432), .ZN(n4281) );
  OAI21_X1 U5198 ( .B1(n4282), .B2(n5008), .A(n4281), .ZN(n4283) );
  AOI21_X1 U5199 ( .B1(n3766), .B2(n4552), .A(n4283), .ZN(n4284) );
  NOR2_X1 U5200 ( .A1(n4584), .A2(n3446), .ZN(n4447) );
  NAND2_X1 U5201 ( .A1(n4609), .A2(n4587), .ZN(n4568) );
  INV_X1 U5202 ( .A(n4285), .ZN(n4288) );
  NAND2_X1 U5203 ( .A1(n4287), .A2(n4286), .ZN(n4293) );
  NOR2_X1 U5204 ( .A1(n3357), .A2(n3383), .ZN(n4701) );
  NAND4_X1 U5205 ( .A1(n4468), .A2(n4288), .A3(n4560), .A4(n4701), .ZN(n4289)
         );
  NAND2_X1 U5206 ( .A1(n4568), .A2(n4289), .ZN(n4290) );
  NAND2_X1 U5207 ( .A1(n4295), .A2(EBX_REG_9__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5208 ( .A1(n4382), .A2(n6398), .ZN(n4291) );
  OAI211_X1 U5209 ( .C1(EBX_REG_9__SCAN_IN), .C2(n4375), .A(n4292), .B(n4291), 
        .ZN(n5361) );
  NAND2_X1 U5210 ( .A1(n4368), .A2(n4902), .ZN(n4294) );
  OAI211_X1 U5211 ( .C1(n3157), .C2(EBX_REG_1__SCAN_IN), .A(n4294), .B(n4324), 
        .ZN(n4298) );
  INV_X1 U5212 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4296) );
  NAND2_X1 U5213 ( .A1(n4378), .A2(n4296), .ZN(n4297) );
  NAND2_X1 U5214 ( .A1(n4368), .A2(EBX_REG_0__SCAN_IN), .ZN(n4300) );
  INV_X1 U5215 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5298) );
  NAND2_X1 U5216 ( .A1(n4324), .A2(n5298), .ZN(n4299) );
  OR2_X1 U5217 ( .A1(n4560), .A2(n4368), .ZN(n4341) );
  INV_X1 U5218 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U5219 ( .A1(n4378), .A2(n5306), .ZN(n4304) );
  OR2_X1 U5220 ( .A1(n4368), .A2(n5306), .ZN(n4303) );
  NAND2_X1 U5221 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n3157), .ZN(n4302)
         );
  NAND4_X1 U5222 ( .A1(n4341), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4769)
         );
  NAND2_X1 U5223 ( .A1(n4295), .A2(EBX_REG_3__SCAN_IN), .ZN(n4306) );
  NAND2_X1 U5224 ( .A1(n4382), .A2(n6463), .ZN(n4305) );
  OAI211_X1 U5225 ( .C1(EBX_REG_3__SCAN_IN), .C2(n4375), .A(n4306), .B(n4305), 
        .ZN(n4767) );
  INV_X1 U5226 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U5227 ( .A1(n4378), .A2(n6269), .ZN(n4309) );
  NAND2_X1 U5228 ( .A1(n4368), .A2(n6453), .ZN(n4307) );
  OAI211_X1 U5229 ( .C1(n3157), .C2(EBX_REG_4__SCAN_IN), .A(n4307), .B(n4324), 
        .ZN(n4308) );
  NAND2_X1 U5230 ( .A1(n4309), .A2(n4308), .ZN(n4883) );
  INV_X1 U5231 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4311) );
  INV_X1 U5232 ( .A(n4375), .ZN(n4315) );
  AOI22_X1 U5233 ( .A1(n4315), .A2(n4311), .B1(n4382), .B2(n4476), .ZN(n4310)
         );
  OAI21_X1 U5234 ( .B1(n4324), .B2(n4311), .A(n4310), .ZN(n4857) );
  INV_X1 U5235 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U5236 ( .A1(n4378), .A2(n6252), .ZN(n4314) );
  NAND2_X1 U5237 ( .A1(n4368), .A2(n4475), .ZN(n4312) );
  OAI211_X1 U5238 ( .C1(n3157), .C2(EBX_REG_6__SCAN_IN), .A(n4312), .B(n4324), 
        .ZN(n4313) );
  NAND2_X1 U5239 ( .A1(n4314), .A2(n4313), .ZN(n4901) );
  NAND2_X1 U5240 ( .A1(n4900), .A2(n4901), .ZN(n4899) );
  INV_X1 U5241 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4317) );
  AOI22_X1 U5242 ( .A1(n4315), .A2(n4317), .B1(n4382), .B2(n6430), .ZN(n4316)
         );
  OAI21_X1 U5243 ( .B1(n4317), .B2(n4324), .A(n4316), .ZN(n5136) );
  INV_X1 U5244 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U5245 ( .A1(n4378), .A2(n5355), .ZN(n4320) );
  NAND2_X1 U5246 ( .A1(n4368), .A2(n6421), .ZN(n4318) );
  OAI211_X1 U5247 ( .C1(n3157), .C2(EBX_REG_8__SCAN_IN), .A(n4318), .B(n4324), 
        .ZN(n4319) );
  NAND2_X1 U5248 ( .A1(n4320), .A2(n4319), .ZN(n5253) );
  INV_X1 U5249 ( .A(n4378), .ZN(n4418) );
  INV_X1 U5250 ( .A(n4368), .ZN(n4376) );
  INV_X1 U5251 ( .A(n4341), .ZN(n4321) );
  AOI21_X1 U5252 ( .B1(n4376), .B2(EBX_REG_10__SCAN_IN), .A(n4321), .ZN(n4323)
         );
  NAND2_X1 U5253 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n3157), .ZN(n4322) );
  OAI211_X1 U5254 ( .C1(EBX_REG_10__SCAN_IN), .C2(n4418), .A(n4323), .B(n4322), 
        .ZN(n5421) );
  NAND2_X1 U5255 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4325) );
  OAI211_X1 U5256 ( .C1(n3157), .C2(EBX_REG_11__SCAN_IN), .A(n4368), .B(n4325), 
        .ZN(n4326) );
  OAI21_X1 U5257 ( .B1(n4375), .B2(EBX_REG_11__SCAN_IN), .A(n4326), .ZN(n6231)
         );
  NOR2_X2 U5258 ( .A1(n6230), .A2(n6231), .ZN(n6229) );
  INV_X1 U5259 ( .A(EBX_REG_12__SCAN_IN), .ZN(n4327) );
  NAND2_X1 U5260 ( .A1(n4378), .A2(n4327), .ZN(n4330) );
  OR2_X1 U5261 ( .A1(n4368), .A2(n4327), .ZN(n4329) );
  NAND2_X1 U5262 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n3157), .ZN(n4328) );
  NAND4_X1 U5263 ( .A1(n4341), .A2(n4330), .A3(n4329), .A4(n4328), .ZN(n5439)
         );
  NAND2_X1 U5264 ( .A1(n6229), .A2(n5439), .ZN(n5438) );
  NAND2_X1 U5265 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4331) );
  OAI211_X1 U5266 ( .C1(n3157), .C2(EBX_REG_13__SCAN_IN), .A(n4368), .B(n4331), 
        .ZN(n4332) );
  OAI21_X1 U5267 ( .B1(n4375), .B2(EBX_REG_13__SCAN_IN), .A(n4332), .ZN(n6156)
         );
  INV_X1 U5268 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U5269 ( .A1(n4378), .A2(n5710), .ZN(n4335) );
  OR2_X1 U5270 ( .A1(n4368), .A2(n5710), .ZN(n4334) );
  NAND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n3157), .ZN(n4333) );
  NAND4_X1 U5272 ( .A1(n4341), .A2(n4335), .A3(n4334), .A4(n4333), .ZN(n5708)
         );
  INV_X1 U5273 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U5274 ( .A1(n4560), .A2(n5633), .ZN(n4336) );
  OAI211_X1 U5275 ( .C1(n4295), .C2(n6140), .A(n4368), .B(n4336), .ZN(n4337)
         );
  OAI21_X1 U5276 ( .B1(n4375), .B2(EBX_REG_15__SCAN_IN), .A(n4337), .ZN(n5637)
         );
  NOR2_X4 U5277 ( .A1(n5707), .A2(n5637), .ZN(n5636) );
  INV_X1 U5278 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U5279 ( .A1(n4378), .A2(n5702), .ZN(n4340) );
  OR2_X1 U5280 ( .A1(n4368), .A2(n5702), .ZN(n4339) );
  NAND2_X1 U5281 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n3157), .ZN(n4338) );
  NAND4_X1 U5282 ( .A1(n4341), .A2(n4340), .A3(n4339), .A4(n4338), .ZN(n5620)
         );
  NAND2_X1 U5283 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4342) );
  OAI211_X1 U5284 ( .C1(n3157), .C2(EBX_REG_17__SCAN_IN), .A(n4368), .B(n4342), 
        .ZN(n4343) );
  OAI21_X1 U5285 ( .B1(n4375), .B2(EBX_REG_17__SCAN_IN), .A(n4343), .ZN(n5608)
         );
  INV_X1 U5286 ( .A(EBX_REG_19__SCAN_IN), .ZN(n4344) );
  NAND2_X1 U5287 ( .A1(n4378), .A2(n4344), .ZN(n4348) );
  INV_X1 U5288 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6123) );
  NAND2_X1 U5289 ( .A1(n4368), .A2(n6123), .ZN(n4346) );
  NAND2_X1 U5290 ( .A1(n4560), .A2(n4344), .ZN(n4345) );
  NAND3_X1 U5291 ( .A1(n4346), .A2(n4324), .A3(n4345), .ZN(n4347) );
  NOR2_X1 U5292 ( .A1(n3157), .A2(EBX_REG_20__SCAN_IN), .ZN(n4349) );
  AOI21_X1 U5293 ( .B1(n4382), .B2(n5940), .A(n4349), .ZN(n5684) );
  OR2_X1 U5294 ( .A1(n4552), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4350)
         );
  INV_X1 U5295 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U5296 ( .A1(n4560), .A2(n5697), .ZN(n5589) );
  NAND2_X1 U5297 ( .A1(n4350), .A2(n5589), .ZN(n5681) );
  NAND2_X1 U5298 ( .A1(n4295), .A2(EBX_REG_20__SCAN_IN), .ZN(n4352) );
  NAND2_X1 U5299 ( .A1(n5681), .A2(n4324), .ZN(n4351) );
  OAI211_X1 U5300 ( .C1(n5684), .C2(n5681), .A(n4352), .B(n4351), .ZN(n4353)
         );
  OR2_X1 U5301 ( .A1(n4552), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4355)
         );
  NAND2_X1 U5302 ( .A1(n4295), .A2(EBX_REG_21__SCAN_IN), .ZN(n4354) );
  OAI211_X1 U5303 ( .C1(n4375), .C2(EBX_REG_21__SCAN_IN), .A(n4355), .B(n4354), 
        .ZN(n5576) );
  INV_X1 U5304 ( .A(n5576), .ZN(n4356) );
  AOI22_X1 U5305 ( .A1(n4376), .A2(EBX_REG_22__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3157), .ZN(n4359) );
  INV_X1 U5306 ( .A(EBX_REG_22__SCAN_IN), .ZN(n4357) );
  NAND2_X1 U5307 ( .A1(n4378), .A2(n4357), .ZN(n4358) );
  INV_X1 U5308 ( .A(n4360), .ZN(n5559) );
  NAND2_X1 U5309 ( .A1(n4324), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4361) );
  OAI211_X1 U5310 ( .C1(n3157), .C2(EBX_REG_23__SCAN_IN), .A(n4368), .B(n4361), 
        .ZN(n4362) );
  OAI21_X1 U5311 ( .B1(n4375), .B2(EBX_REG_23__SCAN_IN), .A(n4362), .ZN(n4465)
         );
  NAND2_X1 U5312 ( .A1(n3157), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4364) );
  NAND2_X1 U5313 ( .A1(n4376), .A2(EBX_REG_24__SCAN_IN), .ZN(n4363) );
  OAI211_X1 U5314 ( .C1(n4418), .C2(EBX_REG_24__SCAN_IN), .A(n4364), .B(n4363), 
        .ZN(n5551) );
  OR2_X1 U5315 ( .A1(n4552), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4366)
         );
  NAND2_X1 U5316 ( .A1(n4295), .A2(EBX_REG_25__SCAN_IN), .ZN(n4365) );
  OAI211_X1 U5317 ( .C1(n4375), .C2(EBX_REG_25__SCAN_IN), .A(n4366), .B(n4365), 
        .ZN(n4367) );
  INV_X1 U5318 ( .A(n4367), .ZN(n5672) );
  INV_X1 U5319 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U5320 ( .A1(n4378), .A2(n5666), .ZN(n4372) );
  NAND2_X1 U5321 ( .A1(n4368), .A2(n5759), .ZN(n4370) );
  NAND2_X1 U5322 ( .A1(n4560), .A2(n5666), .ZN(n4369) );
  NAND3_X1 U5323 ( .A1(n4370), .A2(n4324), .A3(n4369), .ZN(n4371) );
  AND2_X1 U5324 ( .A1(n4372), .A2(n4371), .ZN(n5663) );
  OR2_X1 U5325 ( .A1(n4552), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4374)
         );
  NAND2_X1 U5326 ( .A1(n4295), .A2(EBX_REG_27__SCAN_IN), .ZN(n4373) );
  OAI211_X1 U5327 ( .C1(n4375), .C2(EBX_REG_27__SCAN_IN), .A(n4374), .B(n4373), 
        .ZN(n5533) );
  AOI22_X1 U5328 ( .A1(n4376), .A2(EBX_REG_28__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n3157), .ZN(n4380) );
  INV_X1 U5329 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4377) );
  NAND2_X1 U5330 ( .A1(n4378), .A2(n4377), .ZN(n4379) );
  INV_X1 U5331 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5858) );
  NOR2_X1 U5332 ( .A1(n3157), .A2(EBX_REG_29__SCAN_IN), .ZN(n4381) );
  AOI21_X1 U5333 ( .B1(n4382), .B2(n5858), .A(n4381), .ZN(n5506) );
  NAND2_X1 U5334 ( .A1(n4383), .A2(n5506), .ZN(n4417) );
  AND2_X1 U5335 ( .A1(n4417), .A2(n4324), .ZN(n4421) );
  NAND2_X1 U5336 ( .A1(n4417), .A2(n4383), .ZN(n4386) );
  AND2_X1 U5337 ( .A1(n3157), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4384)
         );
  AOI21_X1 U5338 ( .B1(n4552), .B2(EBX_REG_30__SCAN_IN), .A(n4384), .ZN(n4422)
         );
  INV_X1 U5339 ( .A(n4422), .ZN(n4385) );
  NAND2_X1 U5340 ( .A1(n4386), .A2(n4385), .ZN(n4387) );
  OR2_X1 U5341 ( .A1(n4421), .A2(n4387), .ZN(n4389) );
  OAI211_X1 U5342 ( .C1(n4383), .C2(n4324), .A(n4417), .B(n4422), .ZN(n4388)
         );
  NAND2_X1 U5343 ( .A1(n4389), .A2(n4388), .ZN(n5857) );
  NAND2_X1 U5344 ( .A1(n4391), .A2(EBX_REG_30__SCAN_IN), .ZN(n4392) );
  INV_X1 U5345 ( .A(n4395), .ZN(n4518) );
  INV_X1 U5346 ( .A(n4396), .ZN(n4402) );
  INV_X1 U5347 ( .A(n4397), .ZN(n4398) );
  NAND3_X1 U5348 ( .A1(n4400), .A2(n4399), .A3(n4398), .ZN(n4401) );
  NAND2_X1 U5349 ( .A1(n4402), .A2(n4401), .ZN(n4521) );
  NOR2_X1 U5350 ( .A1(n4521), .A2(n4479), .ZN(n4515) );
  NAND2_X1 U5351 ( .A1(n4515), .A2(n6657), .ZN(n4528) );
  NAND2_X1 U5352 ( .A1(n4731), .A2(n4510), .ZN(n6663) );
  NOR3_X1 U5353 ( .A1(n6659), .A2(n6166), .A3(n6663), .ZN(n6648) );
  NAND2_X1 U5354 ( .A1(n3197), .A2(n6454), .ZN(n4406) );
  NAND2_X1 U5355 ( .A1(n3446), .A2(n6673), .ZN(n4443) );
  NAND2_X1 U5356 ( .A1(n6719), .A2(n6177), .ZN(n4916) );
  INV_X1 U5357 ( .A(n4916), .ZN(n4410) );
  NAND3_X1 U5358 ( .A1(n4443), .A2(n4286), .A3(n4410), .ZN(n4411) );
  INV_X1 U5359 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U5360 ( .A1(n6272), .A2(n5621), .ZN(n6263) );
  INV_X1 U5361 ( .A(n6263), .ZN(n4413) );
  INV_X1 U5362 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6695) );
  INV_X1 U5363 ( .A(REIP_REG_22__SCAN_IN), .ZN(n7068) );
  INV_X1 U5364 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6868) );
  NOR3_X1 U5365 ( .A1(n6695), .A2(n7068), .A3(n6868), .ZN(n4412) );
  NAND3_X1 U5366 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n4429) );
  INV_X1 U5367 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6755) );
  INV_X1 U5368 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6691) );
  INV_X1 U5369 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6689) );
  INV_X1 U5370 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6688) );
  INV_X1 U5371 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6687) );
  INV_X1 U5372 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6685) );
  INV_X1 U5373 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6684) );
  NAND3_X1 U5374 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6271) );
  NOR2_X1 U5375 ( .A1(n6684), .A2(n6271), .ZN(n4924) );
  NAND2_X1 U5376 ( .A1(REIP_REG_5__SCAN_IN), .A2(n4924), .ZN(n5181) );
  NOR2_X1 U5377 ( .A1(n6685), .A2(n5181), .ZN(n5177) );
  NAND2_X1 U5378 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5177), .ZN(n5250) );
  NOR2_X1 U5379 ( .A1(n6687), .A2(n5250), .ZN(n6246) );
  NAND2_X1 U5380 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6246), .ZN(n5651) );
  NOR3_X1 U5381 ( .A1(n6689), .A2(n6688), .A3(n5651), .ZN(n5440) );
  NAND4_X1 U5382 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5440), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5622) );
  NOR2_X1 U5383 ( .A1(n6691), .A2(n5622), .ZN(n5625) );
  NAND2_X1 U5384 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5625), .ZN(n5605) );
  NOR2_X1 U5385 ( .A1(n6755), .A2(n5605), .ZN(n4428) );
  NAND2_X1 U5386 ( .A1(n5621), .A2(n4428), .ZN(n5594) );
  OAI21_X1 U5387 ( .B1(n4429), .B2(n5594), .A(n6263), .ZN(n6084) );
  OAI21_X1 U5388 ( .B1(n4413), .B2(n4412), .A(n6084), .ZN(n6075) );
  NAND3_X1 U5389 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4430) );
  AND2_X1 U5390 ( .A1(n6263), .A2(n4430), .ZN(n4414) );
  NOR2_X1 U5391 ( .A1(n6075), .A2(n4414), .ZN(n6053) );
  NAND2_X1 U5392 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4415) );
  NAND2_X1 U5393 ( .A1(n6247), .A2(n4415), .ZN(n4416) );
  NAND2_X1 U5394 ( .A1(n6053), .A2(n4416), .ZN(n5528) );
  AOI21_X1 U5395 ( .B1(n6247), .B2(n6860), .A(n5528), .ZN(n5483) );
  OAI21_X1 U5396 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6272), .A(n5483), .ZN(n4433) );
  OAI22_X1 U5397 ( .A1(n4552), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n3157), .ZN(n4424) );
  OR2_X1 U5398 ( .A1(n4417), .A2(n4295), .ZN(n4420) );
  NOR2_X1 U5399 ( .A1(n4418), .A2(EBX_REG_29__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U5400 ( .A1(n4383), .A2(n5505), .ZN(n4419) );
  NAND2_X1 U5401 ( .A1(n4420), .A2(n4419), .ZN(n5504) );
  AOI21_X1 U5402 ( .B1(n4422), .B2(n5504), .A(n4421), .ZN(n4423) );
  NAND3_X1 U5403 ( .A1(n4560), .A2(EBX_REG_31__SCAN_IN), .A3(n4916), .ZN(n4425) );
  INV_X1 U5404 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5502) );
  OR2_X1 U5405 ( .A1(n6673), .A2(n4916), .ZN(n6642) );
  NAND2_X1 U5406 ( .A1(n4462), .A2(n6642), .ZN(n4918) );
  NOR3_X1 U5407 ( .A1(n5009), .A2(n5502), .A3(n4918), .ZN(n4426) );
  AOI21_X1 U5408 ( .B1(n6285), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n4426), 
        .ZN(n4427) );
  NAND2_X1 U5409 ( .A1(n6247), .A2(n4428), .ZN(n5595) );
  NOR2_X1 U5410 ( .A1(n5595), .A2(n4429), .ZN(n5562) );
  NAND2_X1 U5411 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5562), .ZN(n5566) );
  NOR2_X1 U5412 ( .A1(n7068), .A2(n5566), .ZN(n6074) );
  NAND2_X1 U5413 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6074), .ZN(n6051) );
  INV_X1 U5414 ( .A(n4430), .ZN(n5538) );
  NAND2_X1 U5415 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5538), .ZN(n4431) );
  NOR2_X1 U5416 ( .A1(n6051), .A2(n4431), .ZN(n5521) );
  NAND2_X1 U5417 ( .A1(n5521), .A2(REIP_REG_28__SCAN_IN), .ZN(n5514) );
  INV_X1 U5418 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6861) );
  NOR4_X1 U5419 ( .A1(n5514), .A2(REIP_REG_31__SCAN_IN), .A3(n6861), .A4(n6860), .ZN(n4432) );
  INV_X1 U5420 ( .A(n4436), .ZN(n4437) );
  XNOR2_X1 U5421 ( .A(n6356), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5801)
         );
  NAND2_X1 U5422 ( .A1(n5802), .A2(n5801), .ZN(n4439) );
  NAND2_X1 U5423 ( .A1(n5902), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4440) );
  OR2_X1 U5424 ( .A1(n6356), .A2(n5940), .ZN(n4438) );
  NAND2_X1 U5425 ( .A1(n4439), .A2(n4438), .ZN(n5794) );
  INV_X1 U5426 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5927) );
  XNOR2_X1 U5427 ( .A(n6356), .B(n5927), .ZN(n5795) );
  NOR2_X1 U5428 ( .A1(n6356), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5786)
         );
  NAND2_X1 U5429 ( .A1(n5793), .A2(n5786), .ZN(n5772) );
  OAI21_X1 U5430 ( .B1(n4439), .B2(n4440), .A(n5772), .ZN(n4441) );
  XNOR2_X1 U5431 ( .A(n4441), .B(n4495), .ZN(n4499) );
  NAND3_X1 U5432 ( .A1(n4442), .A2(n4443), .A3(n6719), .ZN(n4444) );
  NAND3_X1 U5433 ( .A1(n4444), .A2(n4286), .A3(n4707), .ZN(n4445) );
  NAND3_X1 U5434 ( .A1(n4512), .A2(n4446), .A3(n4445), .ZN(n4455) );
  NAND2_X1 U5435 ( .A1(n4587), .A2(n4447), .ZN(n4452) );
  NAND2_X1 U5436 ( .A1(n4448), .A2(n4459), .ZN(n4449) );
  NAND2_X1 U5437 ( .A1(n4449), .A2(n4479), .ZN(n4566) );
  NAND2_X1 U5438 ( .A1(n4801), .A2(n6673), .ZN(n4450) );
  NOR2_X1 U5439 ( .A1(READY_N), .A2(n4521), .ZN(n4571) );
  NAND3_X1 U5440 ( .A1(n4450), .A2(n4571), .A3(n3432), .ZN(n4451) );
  NAND3_X1 U5441 ( .A1(n4452), .A2(n4566), .A3(n4451), .ZN(n4453) );
  NAND2_X1 U5442 ( .A1(n4453), .A2(n6657), .ZN(n4454) );
  INV_X1 U5443 ( .A(n4520), .ZN(n6633) );
  INV_X1 U5444 ( .A(n4456), .ZN(n4457) );
  AOI22_X1 U5445 ( .A1(n4442), .A2(n4560), .B1(n4457), .B2(n3383), .ZN(n4460)
         );
  NAND2_X1 U5446 ( .A1(n4459), .A2(n4458), .ZN(n4610) );
  NAND4_X1 U5447 ( .A1(n6633), .A2(n4460), .A3(n4739), .A4(n4610), .ZN(n4461)
         );
  NAND2_X1 U5448 ( .A1(n4499), .A2(n6474), .ZN(n4498) );
  NAND2_X1 U5449 ( .A1(n4442), .A2(n4462), .ZN(n6643) );
  OAI21_X1 U5450 ( .B1(n4456), .B2(n3383), .A(n6643), .ZN(n4463) );
  AND2_X1 U5451 ( .A1(n5559), .A2(n4465), .ZN(n4466) );
  NOR2_X1 U5452 ( .A1(n4464), .A2(n4466), .ZN(n6070) );
  NOR2_X1 U5453 ( .A1(n6454), .A2(n6695), .ZN(n4505) );
  NOR2_X1 U5454 ( .A1(n3686), .A2(n5466), .ZN(n6146) );
  AND2_X1 U5455 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6146), .ZN(n6144)
         );
  NAND2_X1 U5456 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6144), .ZN(n6134) );
  NAND2_X1 U5457 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5957) );
  NOR2_X1 U5458 ( .A1(n6134), .A2(n5957), .ZN(n4487) );
  NOR2_X1 U5459 ( .A1(n6430), .A2(n6421), .ZN(n6402) );
  INV_X1 U5460 ( .A(n6402), .ZN(n6418) );
  NOR3_X1 U5461 ( .A1(n6398), .A2(n3685), .A3(n6418), .ZN(n5461) );
  INV_X1 U5462 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U5463 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U5464 ( .A1(n6477), .A2(n6472), .ZN(n6444) );
  AND3_X1 U5465 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6444), .ZN(n6432) );
  NAND2_X1 U5466 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6432), .ZN(n4907)
         );
  NOR2_X1 U5467 ( .A1(n4475), .A2(n4907), .ZN(n5457) );
  NAND2_X1 U5468 ( .A1(n5461), .A2(n5457), .ZN(n4488) );
  INV_X1 U5469 ( .A(n4488), .ZN(n4478) );
  INV_X1 U5470 ( .A(n4584), .ZN(n5493) );
  NAND2_X1 U5471 ( .A1(n5493), .A2(n4468), .ZN(n4720) );
  NAND2_X1 U5472 ( .A1(n4470), .A2(n4469), .ZN(n4471) );
  OAI211_X1 U5473 ( .C1(n4467), .C2(n3417), .A(n4720), .B(n4471), .ZN(n4472)
         );
  INV_X1 U5474 ( .A(n4472), .ZN(n4473) );
  NAND2_X1 U5475 ( .A1(n4581), .A2(n4473), .ZN(n4474) );
  NAND2_X1 U5476 ( .A1(n4484), .A2(n4474), .ZN(n4904) );
  INV_X1 U5477 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4903) );
  NAND4_X1 U5478 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(INSTADDRPOINTER_REG_3__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6436) );
  NOR3_X1 U5479 ( .A1(n4476), .A2(n4475), .A3(n6436), .ZN(n5458) );
  AND2_X1 U5480 ( .A1(n5458), .A2(n5461), .ZN(n4485) );
  INV_X1 U5481 ( .A(n4485), .ZN(n4477) );
  NOR3_X1 U5482 ( .A1(n4904), .A2(n4903), .A3(n4477), .ZN(n5456) );
  AOI21_X1 U5483 ( .B1(n4478), .B2(n6433), .A(n5456), .ZN(n6148) );
  NOR2_X1 U5484 ( .A1(n4479), .A2(n3446), .ZN(n4723) );
  NAND2_X1 U5485 ( .A1(n4484), .A2(n4723), .ZN(n6143) );
  INV_X1 U5486 ( .A(n6143), .ZN(n4480) );
  NAND2_X1 U5487 ( .A1(n4480), .A2(n4485), .ZN(n5464) );
  NAND2_X1 U5488 ( .A1(n6148), .A2(n5464), .ZN(n6392) );
  NAND2_X1 U5489 ( .A1(n4487), .A2(n6392), .ZN(n6128) );
  INV_X1 U5490 ( .A(n4492), .ZN(n4481) );
  NAND2_X1 U5491 ( .A1(n6118), .A2(n5935), .ZN(n5921) );
  INV_X1 U5492 ( .A(n5902), .ZN(n4482) );
  NOR3_X1 U5493 ( .A1(n5921), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n4482), 
        .ZN(n4483) );
  AOI211_X1 U5494 ( .C1(n6467), .C2(n6070), .A(n4505), .B(n4483), .ZN(n4496)
         );
  INV_X1 U5495 ( .A(n4904), .ZN(n4557) );
  NOR2_X1 U5496 ( .A1(n4484), .A2(n6476), .ZN(n4649) );
  AOI21_X1 U5497 ( .B1(n4903), .B2(n4557), .A(n4649), .ZN(n5462) );
  OAI221_X1 U5498 ( .B1(n5459), .B2(n4485), .C1(n5459), .C2(n4487), .A(n5462), 
        .ZN(n4486) );
  INV_X1 U5499 ( .A(n4486), .ZN(n4491) );
  INV_X1 U5500 ( .A(n4487), .ZN(n4489) );
  OAI21_X1 U5501 ( .B1(n4489), .B2(n4488), .A(n6433), .ZN(n4490) );
  NAND2_X1 U5502 ( .A1(n5935), .A2(n4492), .ZN(n4493) );
  NAND2_X1 U5503 ( .A1(n5959), .A2(n4493), .ZN(n4494) );
  AND2_X1 U5504 ( .A1(n6126), .A2(n4494), .ZN(n5925) );
  NAND2_X1 U5505 ( .A1(n4498), .A2(n4497), .ZN(U2995) );
  NAND2_X1 U5506 ( .A1(n4499), .A2(n6386), .ZN(n4509) );
  NOR2_X1 U5507 ( .A1(n3179), .A2(n4501), .ZN(n4502) );
  NOR2_X1 U5508 ( .A1(n5836), .A2(n4503), .ZN(n4504) );
  AOI211_X1 U5509 ( .C1(n6360), .C2(n6069), .A(n4505), .B(n4504), .ZN(n4506)
         );
  OAI21_X1 U5510 ( .B1(n6072), .B2(n5839), .A(n4506), .ZN(n4507) );
  INV_X1 U5511 ( .A(n4507), .ZN(n4508) );
  NAND2_X1 U5512 ( .A1(n4509), .A2(n4508), .ZN(U2963) );
  INV_X1 U5513 ( .A(n4723), .ZN(n5498) );
  AOI21_X1 U5514 ( .B1(n5498), .B2(n6643), .A(n6673), .ZN(n4511) );
  AND2_X1 U5515 ( .A1(n6341), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U5516 ( .A(n4528), .ZN(n4514) );
  INV_X1 U5517 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6832) );
  OR2_X1 U5518 ( .A1(n6496), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U5519 ( .A1(n4533), .A2(n6173), .ZN(n4527) );
  INV_X1 U5520 ( .A(n4527), .ZN(n4513) );
  OAI21_X1 U5521 ( .B1(n4514), .B2(n6832), .A(n4513), .ZN(U2788) );
  NAND2_X1 U5522 ( .A1(n4587), .A2(n3717), .ZN(n4517) );
  OR2_X1 U5523 ( .A1(n4515), .A2(n4518), .ZN(n4516) );
  NAND2_X1 U5524 ( .A1(n4517), .A2(n4516), .ZN(n6171) );
  NAND2_X1 U5525 ( .A1(n6722), .A2(n5008), .ZN(n4530) );
  AOI21_X1 U5526 ( .B1(n4530), .B2(n6673), .A(READY_N), .ZN(n6721) );
  NOR2_X1 U5527 ( .A1(n6171), .A2(n6721), .ZN(n6631) );
  OR2_X1 U5528 ( .A1(n6631), .A2(n6655), .ZN(n6178) );
  INV_X1 U5529 ( .A(n4610), .ZN(n4519) );
  OR3_X1 U5530 ( .A1(n4520), .A2(n4519), .A3(n4518), .ZN(n4522) );
  AOI22_X1 U5531 ( .A1(n4587), .A2(n4522), .B1(n4403), .B2(n4521), .ZN(n4525)
         );
  INV_X1 U5532 ( .A(n4587), .ZN(n4523) );
  NAND2_X1 U5533 ( .A1(n4523), .A2(n4609), .ZN(n4524) );
  AND2_X1 U5534 ( .A1(n4525), .A2(n4524), .ZN(n6634) );
  NAND2_X1 U5535 ( .A1(n6178), .A2(MORE_REG_SCAN_IN), .ZN(n4526) );
  OAI21_X1 U5536 ( .B1(n6178), .B2(n6634), .A(n4526), .ZN(U3471) );
  NOR2_X1 U5537 ( .A1(n4527), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4529) );
  AND2_X1 U5538 ( .A1(n4529), .A2(n4528), .ZN(n4531) );
  OAI22_X1 U5539 ( .A1(n4531), .A2(n4530), .B1(n4529), .B2(n6717), .ZN(U3474)
         );
  INV_X1 U5540 ( .A(n4533), .ZN(n4532) );
  NAND2_X1 U5541 ( .A1(n4532), .A2(n3446), .ZN(n4592) );
  INV_X1 U5542 ( .A(EAX_REG_15__SCAN_IN), .ZN(n4535) );
  INV_X1 U5543 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4534) );
  AOI21_X1 U5544 ( .B1(n4801), .B2(READY_N), .A(n4533), .ZN(n4591) );
  INV_X1 U5545 ( .A(DATAI_15_), .ZN(n6829) );
  OAI222_X1 U5546 ( .A1(n4592), .A2(n4535), .B1(n4534), .B2(n4591), .C1(n4706), 
        .C2(n6829), .ZN(U2954) );
  INV_X1 U5547 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4537) );
  NAND2_X1 U5548 ( .A1(n6321), .A2(n4286), .ZN(n4694) );
  AOI22_X1 U5549 ( .A1(n6720), .A2(UWORD_REG_9__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4536) );
  OAI21_X1 U5550 ( .B1(n4537), .B2(n4694), .A(n4536), .ZN(U2898) );
  INV_X1 U5551 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4539) );
  AOI22_X1 U5552 ( .A1(n6720), .A2(UWORD_REG_10__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4538) );
  OAI21_X1 U5553 ( .B1(n4539), .B2(n4694), .A(n4538), .ZN(U2897) );
  INV_X1 U5554 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4541) );
  AOI22_X1 U5555 ( .A1(n6720), .A2(UWORD_REG_8__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4540) );
  OAI21_X1 U5556 ( .B1(n4541), .B2(n4694), .A(n4540), .ZN(U2899) );
  INV_X1 U5557 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4543) );
  AOI22_X1 U5558 ( .A1(n6720), .A2(UWORD_REG_12__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4542) );
  OAI21_X1 U5559 ( .B1(n4543), .B2(n4694), .A(n4542), .ZN(U2895) );
  INV_X1 U5560 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4545) );
  AOI22_X1 U5561 ( .A1(n6720), .A2(UWORD_REG_13__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4544) );
  OAI21_X1 U5562 ( .B1(n4545), .B2(n4694), .A(n4544), .ZN(U2894) );
  INV_X1 U5563 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4547) );
  AOI22_X1 U5564 ( .A1(n6720), .A2(UWORD_REG_11__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4546) );
  OAI21_X1 U5565 ( .B1(n4547), .B2(n4694), .A(n4546), .ZN(U2896) );
  INV_X1 U5566 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4549) );
  AOI22_X1 U5567 ( .A1(n6720), .A2(UWORD_REG_14__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4548) );
  OAI21_X1 U5568 ( .B1(n4549), .B2(n4694), .A(n4548), .ZN(U2893) );
  XNOR2_X1 U5569 ( .A(n4550), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4629)
         );
  OAI21_X1 U5570 ( .B1(n4552), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3220), 
        .ZN(n5300) );
  INV_X1 U5571 ( .A(n5300), .ZN(n4556) );
  INV_X1 U5572 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4553) );
  NOR2_X1 U5573 ( .A1(n6454), .A2(n4553), .ZN(n4631) );
  INV_X1 U5574 ( .A(n4649), .ZN(n4554) );
  AOI21_X1 U5575 ( .B1(n4554), .B2(n6143), .A(n4903), .ZN(n4555) );
  AOI211_X1 U5576 ( .C1(n6467), .C2(n4556), .A(n4631), .B(n4555), .ZN(n4559)
         );
  NOR2_X1 U5577 ( .A1(n4557), .A2(n6433), .ZN(n6145) );
  NOR2_X1 U5578 ( .A1(n6145), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4650)
         );
  INV_X1 U5579 ( .A(n4650), .ZN(n4558) );
  OAI211_X1 U5580 ( .C1(n4629), .C2(n6455), .A(n4559), .B(n4558), .ZN(U3018)
         );
  NOR2_X1 U5581 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6166), .ZN(n6709) );
  INV_X1 U5582 ( .A(n6673), .ZN(n4561) );
  NAND2_X1 U5583 ( .A1(n4723), .A2(n4561), .ZN(n4563) );
  OAI21_X1 U5584 ( .B1(n4561), .B2(n4560), .A(n4442), .ZN(n4562) );
  NAND2_X1 U5585 ( .A1(n4563), .A2(n4562), .ZN(n4564) );
  NAND2_X1 U5586 ( .A1(n4564), .A2(n6719), .ZN(n4569) );
  OR2_X1 U5587 ( .A1(n5008), .A2(n3432), .ZN(n4565) );
  AND2_X1 U5588 ( .A1(n4566), .A2(n4565), .ZN(n4567) );
  OAI211_X1 U5589 ( .C1(n4587), .C2(n4569), .A(n4568), .B(n4567), .ZN(n4570)
         );
  INV_X1 U5590 ( .A(n4570), .ZN(n4576) );
  OR2_X1 U5591 ( .A1(n4587), .A2(n4610), .ZN(n4574) );
  INV_X1 U5592 ( .A(n4739), .ZN(n4572) );
  NAND2_X1 U5593 ( .A1(n4572), .A2(n4571), .ZN(n4573) );
  NAND2_X1 U5594 ( .A1(n4574), .A2(n4573), .ZN(n4704) );
  INV_X1 U5595 ( .A(n4704), .ZN(n4575) );
  NAND2_X1 U5596 ( .A1(n4576), .A2(n4575), .ZN(n6616) );
  NAND2_X1 U5597 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4753), .ZN(n6662) );
  INV_X1 U5598 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6179) );
  OAI22_X1 U5599 ( .A1(n4742), .A2(n6655), .B1(n6662), .B2(n6179), .ZN(n6165)
         );
  NOR2_X1 U5600 ( .A1(n6709), .A2(n6165), .ZN(n5967) );
  INV_X1 U5601 ( .A(n4442), .ZN(n4578) );
  AND4_X1 U5602 ( .A1(n4739), .A2(n4579), .A3(n4578), .A4(n4467), .ZN(n4580)
         );
  AND2_X1 U5603 ( .A1(n4581), .A2(n4580), .ZN(n4713) );
  NOR3_X1 U5604 ( .A1(n4584), .A2(n4582), .A3(n4583), .ZN(n4585) );
  AOI21_X1 U5605 ( .B1(n4723), .B2(n3281), .A(n4585), .ZN(n4586) );
  OAI21_X1 U5606 ( .B1(n4577), .B2(n4713), .A(n4586), .ZN(n6617) );
  NOR2_X1 U5607 ( .A1(n4731), .A2(n4903), .ZN(n4618) );
  AOI22_X1 U5608 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n4233), .B2(n4902), .ZN(n4619)
         );
  INV_X1 U5609 ( .A(n4619), .ZN(n4588) );
  INV_X1 U5610 ( .A(n4583), .ZN(n4737) );
  NOR2_X1 U5611 ( .A1(n6646), .A2(n4582), .ZN(n4623) );
  AOI222_X1 U5612 ( .A1(n6617), .A2(n5499), .B1(n4618), .B2(n4588), .C1(n4737), 
        .C2(n4623), .ZN(n4590) );
  NAND2_X1 U5613 ( .A1(n5967), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4589) );
  OAI21_X1 U5614 ( .B1(n5967), .B2(n4590), .A(n4589), .ZN(U3460) );
  INV_X2 U5615 ( .A(n4591), .ZN(n4674) );
  INV_X2 U5616 ( .A(n4592), .ZN(n4653) );
  AOI22_X1 U5617 ( .A1(n4674), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n4653), .ZN(n4593) );
  NAND2_X1 U5618 ( .A1(n4660), .A2(DATAI_0_), .ZN(n4670) );
  NAND2_X1 U5619 ( .A1(n4593), .A2(n4670), .ZN(U2924) );
  AOI22_X1 U5620 ( .A1(n4674), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n4653), .ZN(n4594) );
  NAND2_X1 U5621 ( .A1(n4660), .A2(DATAI_10_), .ZN(n4595) );
  NAND2_X1 U5622 ( .A1(n4594), .A2(n4595), .ZN(U2949) );
  AOI22_X1 U5623 ( .A1(n4674), .A2(UWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_26__SCAN_IN), .B2(n4653), .ZN(n4596) );
  NAND2_X1 U5624 ( .A1(n4596), .A2(n4595), .ZN(U2934) );
  AOI22_X1 U5625 ( .A1(n4674), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4653), .ZN(n4597) );
  NAND2_X1 U5626 ( .A1(n4660), .A2(DATAI_11_), .ZN(n4637) );
  NAND2_X1 U5627 ( .A1(n4597), .A2(n4637), .ZN(U2950) );
  AOI22_X1 U5628 ( .A1(n4674), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4653), .ZN(n4598) );
  NAND2_X1 U5629 ( .A1(n4660), .A2(DATAI_5_), .ZN(n4656) );
  NAND2_X1 U5630 ( .A1(n4598), .A2(n4656), .ZN(U2929) );
  AOI22_X1 U5631 ( .A1(n4674), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n4653), .ZN(n4599) );
  NAND2_X1 U5632 ( .A1(n4660), .A2(DATAI_9_), .ZN(n4635) );
  NAND2_X1 U5633 ( .A1(n4599), .A2(n4635), .ZN(U2948) );
  AOI22_X1 U5634 ( .A1(n4674), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4653), .ZN(n4600) );
  NAND2_X1 U5635 ( .A1(n4660), .A2(DATAI_6_), .ZN(n4672) );
  NAND2_X1 U5636 ( .A1(n4600), .A2(n4672), .ZN(U2930) );
  AOI22_X1 U5637 ( .A1(n4674), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n4653), .ZN(n4601) );
  NAND2_X1 U5638 ( .A1(n4660), .A2(DATAI_2_), .ZN(n4658) );
  NAND2_X1 U5639 ( .A1(n4601), .A2(n4658), .ZN(U2926) );
  AOI22_X1 U5640 ( .A1(n4674), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4653), .ZN(n4602) );
  NAND2_X1 U5641 ( .A1(n4660), .A2(DATAI_4_), .ZN(n4668) );
  NAND2_X1 U5642 ( .A1(n4602), .A2(n4668), .ZN(U2928) );
  AOI22_X1 U5643 ( .A1(n4674), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n4653), .ZN(n4603) );
  NAND2_X1 U5644 ( .A1(n4660), .A2(DATAI_1_), .ZN(n4654) );
  NAND2_X1 U5645 ( .A1(n4603), .A2(n4654), .ZN(U2925) );
  AOI22_X1 U5646 ( .A1(n4674), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4653), .ZN(n4604) );
  NAND2_X1 U5647 ( .A1(n4660), .A2(DATAI_7_), .ZN(n4664) );
  NAND2_X1 U5648 ( .A1(n4604), .A2(n4664), .ZN(U2931) );
  AOI22_X1 U5649 ( .A1(n4674), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4653), .ZN(n4605) );
  NAND2_X1 U5650 ( .A1(n4660), .A2(DATAI_3_), .ZN(n4666) );
  NAND2_X1 U5651 ( .A1(n4605), .A2(n4666), .ZN(U2927) );
  AOI22_X1 U5652 ( .A1(n4674), .A2(UWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_24__SCAN_IN), .B2(n4653), .ZN(n4606) );
  INV_X1 U5653 ( .A(DATAI_8_), .ZN(n5353) );
  OR2_X1 U5654 ( .A1(n4706), .A2(n5353), .ZN(n4679) );
  NAND2_X1 U5655 ( .A1(n4606), .A2(n4679), .ZN(U2932) );
  AOI22_X1 U5656 ( .A1(n4674), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n4653), .ZN(n4607) );
  INV_X1 U5657 ( .A(DATAI_12_), .ZN(n5446) );
  OR2_X1 U5658 ( .A1(n4706), .A2(n5446), .ZN(n4677) );
  NAND2_X1 U5659 ( .A1(n4607), .A2(n4677), .ZN(U2951) );
  INV_X1 U5660 ( .A(n5967), .ZN(n6170) );
  OR2_X1 U5661 ( .A1(n4608), .A2(n4713), .ZN(n4617) );
  INV_X1 U5662 ( .A(n4609), .ZN(n4611) );
  NAND2_X1 U5663 ( .A1(n4611), .A2(n4610), .ZN(n4716) );
  XNOR2_X1 U5664 ( .A(n4582), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4615)
         );
  XNOR2_X1 U5665 ( .A(n3281), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4612)
         );
  NAND2_X1 U5666 ( .A1(n4723), .A2(n4612), .ZN(n4613) );
  OAI21_X1 U5667 ( .B1(n4615), .B2(n4720), .A(n4613), .ZN(n4614) );
  AOI21_X1 U5668 ( .B1(n4716), .B2(n4615), .A(n4614), .ZN(n4616) );
  AND2_X1 U5669 ( .A1(n4617), .A2(n4616), .ZN(n4727) );
  INV_X1 U5670 ( .A(n5499), .ZN(n5965) );
  NAND2_X1 U5671 ( .A1(n4619), .A2(n4618), .ZN(n4621) );
  INV_X1 U5672 ( .A(n6646), .ZN(n5496) );
  NAND3_X1 U5673 ( .A1(n5496), .A2(n4582), .A3(n4728), .ZN(n4620) );
  OAI211_X1 U5674 ( .C1(n4727), .C2(n5965), .A(n4621), .B(n4620), .ZN(n4622)
         );
  NAND2_X1 U5675 ( .A1(n6170), .A2(n4622), .ZN(n4625) );
  OAI21_X1 U5676 ( .B1(n5967), .B2(n4623), .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), 
        .ZN(n4624) );
  NAND2_X1 U5677 ( .A1(n4625), .A2(n4624), .ZN(U3459) );
  XNOR2_X1 U5678 ( .A(n4627), .B(n4626), .ZN(n5304) );
  NAND2_X1 U5679 ( .A1(n4628), .A2(n5836), .ZN(n4632) );
  NOR2_X1 U5680 ( .A1(n4629), .A2(n6364), .ZN(n4630) );
  AOI211_X1 U5681 ( .C1(PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n4632), .A(n4631), 
        .B(n4630), .ZN(n4633) );
  OAI21_X1 U5682 ( .B1(n5304), .B2(n5839), .A(n4633), .ZN(U2986) );
  AOI22_X1 U5683 ( .A1(n4674), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4653), .ZN(n4634) );
  NAND2_X1 U5684 ( .A1(n4660), .A2(DATAI_14_), .ZN(n4662) );
  NAND2_X1 U5685 ( .A1(n4634), .A2(n4662), .ZN(U2953) );
  AOI22_X1 U5686 ( .A1(n4674), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n4653), .ZN(n4636) );
  NAND2_X1 U5687 ( .A1(n4636), .A2(n4635), .ZN(U2933) );
  AOI22_X1 U5688 ( .A1(n4674), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4653), .ZN(n4638) );
  NAND2_X1 U5689 ( .A1(n4638), .A2(n4637), .ZN(U2935) );
  OAI21_X1 U5690 ( .B1(n4641), .B2(n4640), .A(n4639), .ZN(n5017) );
  XNOR2_X1 U5691 ( .A(n4642), .B(n3157), .ZN(n4648) );
  AOI22_X1 U5692 ( .A1(n6303), .A2(n4648), .B1(n4391), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4643) );
  OAI21_X1 U5693 ( .B1(n5017), .B2(n5704), .A(n4643), .ZN(U2858) );
  OAI222_X1 U5694 ( .A1(n5300), .A2(n5709), .B1(n6307), .B2(n5298), .C1(n5704), 
        .C2(n5304), .ZN(U2859) );
  XNOR2_X1 U5695 ( .A(n4645), .B(n4644), .ZN(n4700) );
  NAND2_X1 U5696 ( .A1(n6476), .A2(REIP_REG_1__SCAN_IN), .ZN(n4696) );
  INV_X1 U5697 ( .A(n4696), .ZN(n4647) );
  AOI211_X1 U5698 ( .C1(n4903), .C2(n6143), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .B(n6403), .ZN(n4646) );
  AOI211_X1 U5699 ( .C1(n6467), .C2(n4648), .A(n4647), .B(n4646), .ZN(n4652)
         );
  OAI21_X1 U5700 ( .B1(n4650), .B2(n4649), .A(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .ZN(n4651) );
  OAI211_X1 U5701 ( .C1(n4700), .C2(n6455), .A(n4652), .B(n4651), .ZN(U3017)
         );
  AOI22_X1 U5702 ( .A1(n4674), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4653), .ZN(n4655) );
  NAND2_X1 U5703 ( .A1(n4655), .A2(n4654), .ZN(U2940) );
  AOI22_X1 U5704 ( .A1(n4674), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4653), .ZN(n4657) );
  NAND2_X1 U5705 ( .A1(n4657), .A2(n4656), .ZN(U2944) );
  AOI22_X1 U5706 ( .A1(n4674), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4653), .ZN(n4659) );
  NAND2_X1 U5707 ( .A1(n4659), .A2(n4658), .ZN(U2941) );
  AOI22_X1 U5708 ( .A1(n4674), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n4653), .ZN(n4661) );
  NAND2_X1 U5709 ( .A1(n4660), .A2(DATAI_13_), .ZN(n4675) );
  NAND2_X1 U5710 ( .A1(n4661), .A2(n4675), .ZN(U2937) );
  AOI22_X1 U5711 ( .A1(n4674), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4653), .ZN(n4663) );
  NAND2_X1 U5712 ( .A1(n4663), .A2(n4662), .ZN(U2938) );
  AOI22_X1 U5713 ( .A1(n4674), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4653), .ZN(n4665) );
  NAND2_X1 U5714 ( .A1(n4665), .A2(n4664), .ZN(U2946) );
  AOI22_X1 U5715 ( .A1(n4674), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4653), .ZN(n4667) );
  NAND2_X1 U5716 ( .A1(n4667), .A2(n4666), .ZN(U2942) );
  AOI22_X1 U5717 ( .A1(n4674), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4653), .ZN(n4669) );
  NAND2_X1 U5718 ( .A1(n4669), .A2(n4668), .ZN(U2943) );
  AOI22_X1 U5719 ( .A1(n4674), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4653), .ZN(n4671) );
  NAND2_X1 U5720 ( .A1(n4671), .A2(n4670), .ZN(U2939) );
  AOI22_X1 U5721 ( .A1(n4674), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4653), .ZN(n4673) );
  NAND2_X1 U5722 ( .A1(n4673), .A2(n4672), .ZN(U2945) );
  AOI22_X1 U5723 ( .A1(n4674), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n4653), .ZN(n4676) );
  NAND2_X1 U5724 ( .A1(n4676), .A2(n4675), .ZN(U2952) );
  AOI22_X1 U5725 ( .A1(n4674), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n4653), .ZN(n4678) );
  NAND2_X1 U5726 ( .A1(n4678), .A2(n4677), .ZN(U2936) );
  AOI22_X1 U5727 ( .A1(n4674), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n4653), .ZN(n4680) );
  NAND2_X1 U5728 ( .A1(n4680), .A2(n4679), .ZN(U2947) );
  INV_X1 U5729 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4682) );
  AOI22_X1 U5730 ( .A1(n6720), .A2(UWORD_REG_6__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4681) );
  OAI21_X1 U5731 ( .B1(n4682), .B2(n4694), .A(n4681), .ZN(U2901) );
  INV_X1 U5732 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4684) );
  AOI22_X1 U5733 ( .A1(n6720), .A2(UWORD_REG_7__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4683) );
  OAI21_X1 U5734 ( .B1(n4684), .B2(n4694), .A(n4683), .ZN(U2900) );
  AOI22_X1 U5735 ( .A1(n6720), .A2(UWORD_REG_4__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4685) );
  OAI21_X1 U5736 ( .B1(n4032), .B2(n4694), .A(n4685), .ZN(U2903) );
  INV_X1 U5737 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4687) );
  AOI22_X1 U5738 ( .A1(n6720), .A2(UWORD_REG_5__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4686) );
  OAI21_X1 U5739 ( .B1(n4687), .B2(n4694), .A(n4686), .ZN(U2902) );
  AOI22_X1 U5740 ( .A1(n6720), .A2(UWORD_REG_2__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4688) );
  OAI21_X1 U5741 ( .B1(n3999), .B2(n4694), .A(n4688), .ZN(U2905) );
  INV_X1 U5742 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4690) );
  AOI22_X1 U5743 ( .A1(n6720), .A2(UWORD_REG_3__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4689) );
  OAI21_X1 U5744 ( .B1(n4690), .B2(n4694), .A(n4689), .ZN(U2904) );
  INV_X1 U5745 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4692) );
  AOI22_X1 U5746 ( .A1(n6720), .A2(UWORD_REG_0__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4691) );
  OAI21_X1 U5747 ( .B1(n4692), .B2(n4694), .A(n4691), .ZN(U2907) );
  INV_X1 U5748 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4695) );
  AOI22_X1 U5749 ( .A1(n6720), .A2(UWORD_REG_1__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4693) );
  OAI21_X1 U5750 ( .B1(n4695), .B2(n4694), .A(n4693), .ZN(U2906) );
  INV_X1 U5751 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5012) );
  OAI21_X1 U5752 ( .B1(n5836), .B2(n5012), .A(n4696), .ZN(n4698) );
  NOR2_X1 U5753 ( .A1(n5017), .A2(n5839), .ZN(n4697) );
  AOI211_X1 U5754 ( .C1(n6360), .C2(n5012), .A(n4698), .B(n4697), .ZN(n4699)
         );
  OAI21_X1 U5755 ( .B1(n4700), .B2(n6364), .A(n4699), .ZN(U2985) );
  NAND2_X1 U5756 ( .A1(n4701), .A2(n3417), .ZN(n4702) );
  NOR2_X1 U5757 ( .A1(n4467), .A2(n4702), .ZN(n4703) );
  AND2_X1 U5758 ( .A1(n3384), .A2(n3357), .ZN(n4710) );
  INV_X1 U5759 ( .A(n4710), .ZN(n4708) );
  AND2_X1 U5760 ( .A1(n4708), .A2(n4707), .ZN(n4709) );
  AND2_X1 U5761 ( .A1(n5738), .A2(n3447), .ZN(n6314) );
  INV_X1 U5762 ( .A(DATAI_1_), .ZN(n6843) );
  INV_X1 U5763 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6349) );
  OAI222_X1 U5764 ( .A1(n5017), .A2(n6086), .B1(n5739), .B2(n6843), .C1(n5738), 
        .C2(n6349), .ZN(U2890) );
  INV_X1 U5765 ( .A(n4713), .ZN(n5494) );
  MUX2_X1 U5766 ( .A(n4715), .B(n3791), .S(n4582), .Z(n4717) );
  OAI21_X1 U5767 ( .B1(n4714), .B2(n4717), .A(n4716), .ZN(n4725) );
  XNOR2_X1 U5768 ( .A(n4718), .B(n3791), .ZN(n4722) );
  OAI21_X1 U5769 ( .B1(n3155), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3400), 
        .ZN(n5964) );
  NOR2_X1 U5770 ( .A1(n4720), .A2(n5964), .ZN(n4721) );
  AOI21_X1 U5771 ( .B1(n4723), .B2(n4722), .A(n4721), .ZN(n4724) );
  NAND2_X1 U5772 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  AOI21_X1 U5773 ( .B1(n4712), .B2(n5494), .A(n4726), .ZN(n5966) );
  MUX2_X1 U5774 ( .A(n3791), .B(n5966), .S(n6616), .Z(n6625) );
  INV_X1 U5775 ( .A(n6625), .ZN(n4732) );
  NAND2_X1 U5776 ( .A1(n4727), .A2(n6616), .ZN(n4730) );
  NAND2_X1 U5777 ( .A1(n4742), .A2(n4728), .ZN(n4729) );
  NAND3_X1 U5778 ( .A1(n4732), .A2(n6624), .A3(n4731), .ZN(n4736) );
  AND2_X1 U5779 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6179), .ZN(n4734) );
  NAND2_X1 U5780 ( .A1(n4733), .A2(n4734), .ZN(n4735) );
  NAND2_X1 U5781 ( .A1(n4736), .A2(n4735), .ZN(n6637) );
  NAND2_X1 U5782 ( .A1(n6637), .A2(n4737), .ZN(n4745) );
  INV_X1 U5783 ( .A(n4818), .ZN(n4972) );
  OR2_X1 U5784 ( .A1(n3566), .A2(n4972), .ZN(n4738) );
  XNOR2_X1 U5785 ( .A(n4738), .B(n6169), .ZN(n6266) );
  INV_X1 U5786 ( .A(n6266), .ZN(n4741) );
  NOR2_X1 U5787 ( .A1(n4739), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4740) );
  NAND2_X1 U5788 ( .A1(n4741), .A2(n4740), .ZN(n6164) );
  MUX2_X1 U5789 ( .A(n4742), .B(n6179), .S(STATE2_REG_1__SCAN_IN), .Z(n4743)
         );
  NAND2_X1 U5790 ( .A1(n4743), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4744) );
  AND2_X1 U5791 ( .A1(n6164), .A2(n4744), .ZN(n6635) );
  AND2_X1 U5792 ( .A1(n6649), .A2(n6179), .ZN(n4746) );
  INV_X1 U5793 ( .A(n6663), .ZN(n6723) );
  OAI21_X1 U5794 ( .B1(n4746), .B2(n6662), .A(n4935), .ZN(n6483) );
  XNOR2_X1 U5795 ( .A(n3772), .B(n4787), .ZN(n4749) );
  INV_X1 U5796 ( .A(n4608), .ZN(n4748) );
  NAND2_X1 U5797 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6166), .ZN(n4783) );
  AOI22_X1 U5798 ( .A1(n4749), .A2(n6015), .B1(n4748), .B2(n4783), .ZN(n4751)
         );
  NAND2_X1 U5799 ( .A1(n4786), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4750) );
  OAI21_X1 U5800 ( .B1(n4786), .B2(n4751), .A(n4750), .ZN(U3463) );
  INV_X1 U5801 ( .A(n4752), .ZN(n5495) );
  AOI222_X1 U5802 ( .A1(n6649), .A2(n4753), .B1(n5495), .B2(n4783), .C1(n5316), 
        .C2(n6015), .ZN(n4755) );
  NAND2_X1 U5803 ( .A1(n4786), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4754) );
  OAI21_X1 U5804 ( .B1(n4786), .B2(n4755), .A(n4754), .ZN(U3465) );
  INV_X1 U5805 ( .A(n4577), .ZN(n5010) );
  AOI211_X1 U5806 ( .C1(n5024), .C2(n6177), .A(n6496), .B(n4787), .ZN(n4756)
         );
  AOI21_X1 U5807 ( .B1(n5010), .B2(n4783), .A(n4756), .ZN(n4758) );
  NAND2_X1 U5808 ( .A1(n4786), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4757) );
  OAI21_X1 U5809 ( .B1(n4786), .B2(n4758), .A(n4757), .ZN(U3464) );
  INV_X1 U5810 ( .A(n4759), .ZN(n4763) );
  NAND3_X1 U5811 ( .A1(n4760), .A2(n4761), .A3(n4639), .ZN(n4762) );
  AND2_X1 U5812 ( .A1(n4763), .A2(n4762), .ZN(n6384) );
  INV_X1 U5813 ( .A(n6384), .ZN(n4771) );
  INV_X1 U5814 ( .A(DATAI_2_), .ZN(n4809) );
  INV_X1 U5815 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6347) );
  OAI222_X1 U5816 ( .A1(n4771), .A2(n6086), .B1(n5739), .B2(n4809), .C1(n5738), 
        .C2(n6347), .ZN(U2889) );
  CLKBUF_X1 U5817 ( .A(n4764), .Z(n4880) );
  OAI21_X1 U5818 ( .B1(n4759), .B2(n4765), .A(n4880), .ZN(n6282) );
  AOI21_X1 U5819 ( .B1(n4767), .B2(n4766), .A(n4882), .ZN(n6460) );
  AOI22_X1 U5820 ( .A1(n6303), .A2(n6460), .B1(EBX_REG_3__SCAN_IN), .B2(n4391), 
        .ZN(n4768) );
  OAI21_X1 U5821 ( .B1(n6282), .B2(n5704), .A(n4768), .ZN(U2856) );
  XNOR2_X1 U5822 ( .A(n4770), .B(n4769), .ZN(n6465) );
  OAI222_X1 U5823 ( .A1(n5704), .A2(n4771), .B1(n5306), .B2(n6307), .C1(n5709), 
        .C2(n6465), .ZN(U2857) );
  NOR2_X1 U5824 ( .A1(n4773), .A2(n4772), .ZN(n6457) );
  INV_X1 U5825 ( .A(n4774), .ZN(n6456) );
  OR3_X1 U5826 ( .A1(n6457), .A2(n6456), .A3(n6364), .ZN(n4779) );
  INV_X1 U5827 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4775) );
  OAI22_X1 U5828 ( .A1(n5836), .A2(n4776), .B1(n6454), .B2(n4775), .ZN(n4777)
         );
  AOI21_X1 U5829 ( .B1(n6360), .B2(n6295), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5830 ( .C1(n6282), .C2(n5839), .A(n4779), .B(n4778), .ZN(U2983)
         );
  INV_X1 U5831 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6353) );
  INV_X1 U5832 ( .A(DATAI_0_), .ZN(n7084) );
  OAI222_X1 U5833 ( .A1(n6086), .A2(n5304), .B1(n5738), .B2(n6353), .C1(n7084), 
        .C2(n5739), .ZN(U2891) );
  NOR2_X1 U5834 ( .A1(n3772), .A2(n5314), .ZN(n4817) );
  NAND2_X1 U5835 ( .A1(n4817), .A2(n4787), .ZN(n4859) );
  INV_X1 U5836 ( .A(n5185), .ZN(n4780) );
  NAND2_X1 U5837 ( .A1(n4780), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5194) );
  NAND3_X1 U5838 ( .A1(n4859), .A2(n5194), .A3(n5059), .ZN(n5019) );
  NOR2_X1 U5839 ( .A1(n6496), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6499) );
  AOI222_X1 U5840 ( .A1(n5019), .A2(n6015), .B1(n4712), .B2(n4783), .C1(n4782), 
        .C2(n6499), .ZN(n4785) );
  NAND2_X1 U5841 ( .A1(n4786), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U5842 ( .B1(n4786), .B2(n4785), .A(n4784), .ZN(U3462) );
  INV_X1 U5843 ( .A(n4787), .ZN(n5018) );
  OR2_X1 U5844 ( .A1(n5059), .A2(n5018), .ZN(n4788) );
  NAND2_X1 U5845 ( .A1(n4788), .A2(n6015), .ZN(n4795) );
  AND2_X1 U5846 ( .A1(n4608), .A2(n5010), .ZN(n5021) );
  AND2_X1 U5847 ( .A1(n5021), .A2(n4712), .ZN(n5264) );
  NOR2_X1 U5848 ( .A1(n5022), .A2(n6487), .ZN(n4797) );
  AOI21_X1 U5849 ( .B1(n5264), .B2(n5495), .A(n4797), .ZN(n4792) );
  OR2_X1 U5850 ( .A1(n4795), .A2(n4792), .ZN(n4791) );
  NAND3_X1 U5851 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6623), .ZN(n5265) );
  INV_X1 U5852 ( .A(n5265), .ZN(n4789) );
  NAND2_X1 U5853 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4789), .ZN(n4790) );
  NAND2_X1 U5854 ( .A1(n4791), .A2(n4790), .ZN(n6605) );
  INV_X1 U5855 ( .A(n6605), .ZN(n4816) );
  INV_X1 U5856 ( .A(DATAI_6_), .ZN(n7103) );
  NOR2_X1 U5857 ( .A1(n7103), .A2(n4935), .ZN(n6573) );
  INV_X1 U5858 ( .A(n4792), .ZN(n4794) );
  OAI21_X1 U5859 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6166), .A(n5263), 
        .ZN(n4822) );
  AOI21_X1 U5860 ( .B1(n5265), .B2(n6496), .A(n4822), .ZN(n4793) );
  OAI21_X1 U5861 ( .B1(n4795), .B2(n4794), .A(n4793), .ZN(n6607) );
  NAND2_X1 U5862 ( .A1(n6385), .A2(DATAI_30_), .ZN(n6576) );
  NOR2_X1 U5863 ( .A1(n6610), .A2(n6576), .ZN(n4799) );
  NAND2_X1 U5864 ( .A1(n6385), .A2(DATAI_22_), .ZN(n6542) );
  NAND2_X1 U5865 ( .A1(n4841), .A2(n3417), .ZN(n6570) );
  INV_X1 U5866 ( .A(n4797), .ZN(n6600) );
  OAI22_X1 U5867 ( .A1(n6603), .A2(n6542), .B1(n6570), .B2(n6600), .ZN(n4798)
         );
  AOI211_X1 U5868 ( .C1(n6607), .C2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4799), 
        .B(n4798), .ZN(n4800) );
  OAI21_X1 U5869 ( .B1(n4816), .B2(n6537), .A(n4800), .ZN(U3114) );
  NOR2_X1 U5870 ( .A1(n6843), .A2(n4935), .ZN(n6555) );
  NAND2_X1 U5871 ( .A1(n6385), .A2(DATAI_25_), .ZN(n6558) );
  NOR2_X1 U5872 ( .A1(n6610), .A2(n6558), .ZN(n4803) );
  NAND2_X1 U5873 ( .A1(n6385), .A2(DATAI_17_), .ZN(n6513) );
  NAND2_X1 U5874 ( .A1(n4841), .A2(n4801), .ZN(n6552) );
  OAI22_X1 U5875 ( .A1(n6603), .A2(n6513), .B1(n6552), .B2(n6600), .ZN(n4802)
         );
  AOI211_X1 U5876 ( .C1(n6607), .C2(INSTQUEUE_REG_11__1__SCAN_IN), .A(n4803), 
        .B(n4802), .ZN(n4804) );
  OAI21_X1 U5877 ( .B1(n4816), .B2(n6508), .A(n4804), .ZN(U3109) );
  NOR2_X1 U5878 ( .A1(n7084), .A2(n4935), .ZN(n5231) );
  INV_X1 U5879 ( .A(DATAI_24_), .ZN(n4805) );
  NOR2_X1 U5880 ( .A1(n5839), .A2(n4805), .ZN(n6504) );
  INV_X1 U5881 ( .A(n6504), .ZN(n6021) );
  NOR2_X1 U5882 ( .A1(n6610), .A2(n6021), .ZN(n4807) );
  NAND2_X1 U5883 ( .A1(n6385), .A2(DATAI_16_), .ZN(n6507) );
  NAND2_X1 U5884 ( .A1(n4841), .A2(n4286), .ZN(n6493) );
  OAI22_X1 U5885 ( .A1(n6603), .A2(n6507), .B1(n6493), .B2(n6600), .ZN(n4806)
         );
  AOI211_X1 U5886 ( .C1(n6607), .C2(INSTQUEUE_REG_11__0__SCAN_IN), .A(n4807), 
        .B(n4806), .ZN(n4808) );
  OAI21_X1 U5887 ( .B1(n4816), .B2(n6492), .A(n4808), .ZN(U3108) );
  NOR2_X1 U5888 ( .A1(n4809), .A2(n4935), .ZN(n5212) );
  INV_X1 U5889 ( .A(n6517), .ZN(n6029) );
  NOR2_X1 U5890 ( .A1(n6610), .A2(n6029), .ZN(n4811) );
  NAND2_X1 U5891 ( .A1(n6385), .A2(DATAI_18_), .ZN(n6520) );
  NAND2_X1 U5892 ( .A1(n4841), .A2(n3432), .ZN(n6515) );
  OAI22_X1 U5893 ( .A1(n6603), .A2(n6520), .B1(n6515), .B2(n6600), .ZN(n4810)
         );
  AOI211_X1 U5894 ( .C1(n6607), .C2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4811), 
        .B(n4810), .ZN(n4812) );
  OAI21_X1 U5895 ( .B1(n4816), .B2(n6514), .A(n4812), .ZN(U3110) );
  INV_X1 U5896 ( .A(DATAI_4_), .ZN(n6780) );
  NOR2_X1 U5897 ( .A1(n6780), .A2(n4935), .ZN(n6566) );
  NAND2_X1 U5898 ( .A1(n6385), .A2(DATAI_28_), .ZN(n6569) );
  NOR2_X1 U5899 ( .A1(n6610), .A2(n6569), .ZN(n4814) );
  NAND2_X1 U5900 ( .A1(n6385), .A2(DATAI_20_), .ZN(n6531) );
  NAND2_X1 U5901 ( .A1(n4841), .A2(n3383), .ZN(n6563) );
  OAI22_X1 U5902 ( .A1(n6603), .A2(n6531), .B1(n6563), .B2(n6600), .ZN(n4813)
         );
  AOI211_X1 U5903 ( .C1(n6607), .C2(INSTQUEUE_REG_11__4__SCAN_IN), .A(n4814), 
        .B(n4813), .ZN(n4815) );
  OAI21_X1 U5904 ( .B1(n4816), .B2(n6526), .A(n4815), .ZN(U3112) );
  INV_X1 U5905 ( .A(DATAI_3_), .ZN(n7074) );
  INV_X1 U5906 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6345) );
  OAI222_X1 U5907 ( .A1(n6282), .A2(n6086), .B1(n5739), .B2(n7074), .C1(n5738), 
        .C2(n6345), .ZN(U2888) );
  NAND2_X1 U5908 ( .A1(n4817), .A2(n5024), .ZN(n4824) );
  OAI21_X1 U5909 ( .B1(n4824), .B2(n6177), .A(n6015), .ZN(n4971) );
  NOR2_X1 U5910 ( .A1(n4608), .A2(n5010), .ZN(n5187) );
  NOR2_X1 U5911 ( .A1(n4752), .A2(n4818), .ZN(n4860) );
  NAND2_X1 U5912 ( .A1(n6618), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5189) );
  OR2_X1 U5913 ( .A1(n5189), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4974)
         );
  NOR2_X1 U5914 ( .A1(n6613), .A2(n4974), .ZN(n4825) );
  AOI21_X1 U5915 ( .B1(n5187), .B2(n4860), .A(n4825), .ZN(n4820) );
  OAI22_X1 U5916 ( .A1(n4971), .A2(n4820), .B1(n4974), .B2(n4510), .ZN(n4819)
         );
  INV_X1 U5917 ( .A(DATAI_5_), .ZN(n4886) );
  NOR2_X1 U5918 ( .A1(n4886), .A2(n4935), .ZN(n6596) );
  INV_X1 U5919 ( .A(n4971), .ZN(n4821) );
  AOI22_X1 U5920 ( .A1(n4821), .A2(n4820), .B1(n4974), .B2(n6496), .ZN(n4823)
         );
  NAND2_X1 U5921 ( .A1(n4848), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4828) );
  NAND2_X1 U5922 ( .A1(n6385), .A2(DATAI_29_), .ZN(n6599) );
  INV_X1 U5923 ( .A(n6599), .ZN(n6534) );
  NOR2_X2 U5924 ( .A1(n4824), .A2(n5316), .ZN(n5005) );
  NAND2_X1 U5925 ( .A1(n6385), .A2(DATAI_21_), .ZN(n6594) );
  NAND2_X1 U5926 ( .A1(n4841), .A2(n3373), .ZN(n6593) );
  INV_X1 U5927 ( .A(n4825), .ZN(n4849) );
  OAI22_X1 U5928 ( .A1(n6495), .A2(n6594), .B1(n6593), .B2(n4849), .ZN(n4826)
         );
  AOI21_X1 U5929 ( .B1(n6534), .B2(n5005), .A(n4826), .ZN(n4827) );
  OAI211_X1 U5930 ( .C1(n4853), .C2(n6532), .A(n4828), .B(n4827), .ZN(U3065)
         );
  NAND2_X1 U5931 ( .A1(n4848), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4831) );
  OAI22_X1 U5932 ( .A1(n6495), .A2(n6531), .B1(n6563), .B2(n4849), .ZN(n4829)
         );
  AOI21_X1 U5933 ( .B1(n6528), .B2(n5005), .A(n4829), .ZN(n4830) );
  OAI211_X1 U5934 ( .C1(n4853), .C2(n6526), .A(n4831), .B(n4830), .ZN(U3064)
         );
  NOR2_X1 U5935 ( .A1(n7074), .A2(n4935), .ZN(n6589) );
  NAND2_X1 U5936 ( .A1(n4848), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4834) );
  NAND2_X1 U5937 ( .A1(n6385), .A2(DATAI_27_), .ZN(n6592) );
  INV_X1 U5938 ( .A(n6592), .ZN(n6523) );
  NAND2_X1 U5939 ( .A1(n6385), .A2(DATAI_19_), .ZN(n6587) );
  NAND2_X1 U5940 ( .A1(n4841), .A2(n3431), .ZN(n6586) );
  OAI22_X1 U5941 ( .A1(n6495), .A2(n6587), .B1(n6586), .B2(n4849), .ZN(n4832)
         );
  AOI21_X1 U5942 ( .B1(n6523), .B2(n5005), .A(n4832), .ZN(n4833) );
  OAI211_X1 U5943 ( .C1(n4853), .C2(n6521), .A(n4834), .B(n4833), .ZN(U3063)
         );
  NAND2_X1 U5944 ( .A1(n4848), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4837) );
  OAI22_X1 U5945 ( .A1(n6495), .A2(n6513), .B1(n6552), .B2(n4849), .ZN(n4835)
         );
  AOI21_X1 U5946 ( .B1(n6510), .B2(n5005), .A(n4835), .ZN(n4836) );
  OAI211_X1 U5947 ( .C1(n4853), .C2(n6508), .A(n4837), .B(n4836), .ZN(U3061)
         );
  NAND2_X1 U5948 ( .A1(n4848), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4840) );
  OAI22_X1 U5949 ( .A1(n6495), .A2(n6520), .B1(n6515), .B2(n4849), .ZN(n4838)
         );
  AOI21_X1 U5950 ( .B1(n6517), .B2(n5005), .A(n4838), .ZN(n4839) );
  OAI211_X1 U5951 ( .C1(n4853), .C2(n6514), .A(n4840), .B(n4839), .ZN(U3062)
         );
  INV_X1 U5952 ( .A(DATAI_7_), .ZN(n7065) );
  NOR2_X1 U5953 ( .A1(n7065), .A2(n4935), .ZN(n6606) );
  NAND2_X1 U5954 ( .A1(n4848), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4844) );
  NAND2_X1 U5955 ( .A1(n6385), .A2(DATAI_31_), .ZN(n6611) );
  NAND2_X1 U5956 ( .A1(n6385), .A2(DATAI_23_), .ZN(n6602) );
  NAND2_X1 U5957 ( .A1(n4841), .A2(n3357), .ZN(n6601) );
  OAI22_X1 U5958 ( .A1(n6495), .A2(n6602), .B1(n6601), .B2(n4849), .ZN(n4842)
         );
  AOI21_X1 U5959 ( .B1(n6548), .B2(n5005), .A(n4842), .ZN(n4843) );
  OAI211_X1 U5960 ( .C1(n4853), .C2(n6543), .A(n4844), .B(n4843), .ZN(U3067)
         );
  NAND2_X1 U5961 ( .A1(n4848), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U5962 ( .A1(n6495), .A2(n6507), .B1(n6493), .B2(n4849), .ZN(n4845)
         );
  AOI21_X1 U5963 ( .B1(n6504), .B2(n5005), .A(n4845), .ZN(n4846) );
  OAI211_X1 U5964 ( .C1(n4853), .C2(n6492), .A(n4847), .B(n4846), .ZN(U3060)
         );
  NAND2_X1 U5965 ( .A1(n4848), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4852) );
  INV_X1 U5966 ( .A(n6576), .ZN(n6539) );
  OAI22_X1 U5967 ( .A1(n6495), .A2(n6542), .B1(n6570), .B2(n4849), .ZN(n4850)
         );
  AOI21_X1 U5968 ( .B1(n6539), .B2(n5005), .A(n4850), .ZN(n4851) );
  OAI211_X1 U5969 ( .C1(n4853), .C2(n6537), .A(n4852), .B(n4851), .ZN(U3066)
         );
  OAI21_X1 U5970 ( .B1(n4854), .B2(n4855), .A(n4856), .ZN(n4931) );
  AOI21_X1 U5971 ( .B1(n4857), .B2(n4881), .A(n4900), .ZN(n6435) );
  AOI22_X1 U5972 ( .A1(n6303), .A2(n6435), .B1(EBX_REG_5__SCAN_IN), .B2(n4391), 
        .ZN(n4858) );
  OAI21_X1 U5973 ( .B1(n4931), .B2(n5704), .A(n4858), .ZN(U2854) );
  NAND2_X1 U5974 ( .A1(n4859), .A2(n6015), .ZN(n4866) );
  OR2_X1 U5975 ( .A1(n4608), .A2(n4577), .ZN(n6498) );
  INV_X1 U5976 ( .A(n4860), .ZN(n4861) );
  OAI21_X1 U5977 ( .B1(n6498), .B2(n4861), .A(n6577), .ZN(n4867) );
  INV_X1 U5978 ( .A(n4867), .ZN(n4862) );
  OAI22_X1 U5979 ( .A1(n4866), .A2(n4862), .B1(n6484), .B2(n4510), .ZN(n6581)
         );
  INV_X1 U5980 ( .A(n6581), .ZN(n4877) );
  OR2_X1 U5981 ( .A1(n5971), .A2(n5314), .ZN(n4863) );
  INV_X1 U5982 ( .A(n6585), .ZN(n6497) );
  NOR2_X2 U5983 ( .A1(n4863), .A2(n5969), .ZN(n6580) );
  INV_X1 U5984 ( .A(n6580), .ZN(n4873) );
  OAI22_X1 U5985 ( .A1(n4873), .A2(n6520), .B1(n6577), .B2(n6515), .ZN(n4864)
         );
  AOI21_X1 U5986 ( .B1(n6517), .B2(n6497), .A(n4864), .ZN(n4869) );
  NAND2_X1 U5987 ( .A1(n6496), .A2(n6484), .ZN(n4865) );
  OAI211_X1 U5988 ( .C1(n4867), .C2(n4866), .A(n6012), .B(n4865), .ZN(n6582)
         );
  NAND2_X1 U5989 ( .A1(n6582), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4868) );
  OAI211_X1 U5990 ( .C1(n4877), .C2(n6514), .A(n4869), .B(n4868), .ZN(U3078)
         );
  OAI22_X1 U5991 ( .A1(n4873), .A2(n6507), .B1(n6577), .B2(n6493), .ZN(n4870)
         );
  AOI21_X1 U5992 ( .B1(n6504), .B2(n6497), .A(n4870), .ZN(n4872) );
  NAND2_X1 U5993 ( .A1(n6582), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4871) );
  OAI211_X1 U5994 ( .C1(n4877), .C2(n6492), .A(n4872), .B(n4871), .ZN(U3076)
         );
  OAI22_X1 U5995 ( .A1(n4873), .A2(n6594), .B1(n6577), .B2(n6593), .ZN(n4874)
         );
  AOI21_X1 U5996 ( .B1(n6534), .B2(n6497), .A(n4874), .ZN(n4876) );
  NAND2_X1 U5997 ( .A1(n6582), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4875) );
  OAI211_X1 U5998 ( .C1(n4877), .C2(n6532), .A(n4876), .B(n4875), .ZN(U3081)
         );
  INV_X1 U5999 ( .A(n4878), .ZN(n4879) );
  XNOR2_X1 U6000 ( .A(n4880), .B(n4879), .ZN(n6375) );
  INV_X1 U6001 ( .A(n5704), .ZN(n6304) );
  OAI21_X1 U6002 ( .B1(n4883), .B2(n4882), .A(n4881), .ZN(n6447) );
  OAI22_X1 U6003 ( .A1(n5709), .A2(n6447), .B1(n6307), .B2(n6269), .ZN(n4884)
         );
  AOI21_X1 U6004 ( .B1(n6375), .B2(n6304), .A(n4884), .ZN(n4885) );
  INV_X1 U6005 ( .A(n4885), .ZN(U2855) );
  INV_X1 U6006 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6340) );
  OAI222_X1 U6007 ( .A1(n4931), .A2(n6086), .B1(n5739), .B2(n4886), .C1(n5738), 
        .C2(n6340), .ZN(U2886) );
  INV_X1 U6008 ( .A(n6375), .ZN(n4887) );
  INV_X1 U6009 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6343) );
  OAI222_X1 U6010 ( .A1(n6086), .A2(n4887), .B1(n5738), .B2(n6343), .C1(n6780), 
        .C2(n5739), .ZN(U2887) );
  OAI21_X1 U6011 ( .B1(n4888), .B2(n4890), .A(n4889), .ZN(n4891) );
  INV_X1 U6012 ( .A(n4891), .ZN(n6438) );
  NAND2_X1 U6013 ( .A1(n6438), .A2(n6386), .ZN(n4895) );
  INV_X1 U6014 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4892) );
  NOR2_X1 U6015 ( .A1(n6454), .A2(n4892), .ZN(n6434) );
  NOR2_X1 U6016 ( .A1(n5836), .A2(n4922), .ZN(n4893) );
  AOI211_X1 U6017 ( .C1(n6360), .C2(n4929), .A(n6434), .B(n4893), .ZN(n4894)
         );
  OAI211_X1 U6018 ( .C1(n5839), .C2(n4931), .A(n4895), .B(n4894), .ZN(U2981)
         );
  OAI21_X1 U6019 ( .B1(n4898), .B2(n4897), .A(n4896), .ZN(n6365) );
  OAI21_X1 U6020 ( .B1(n4901), .B2(n4900), .A(n4899), .ZN(n6256) );
  NOR2_X1 U6021 ( .A1(n6448), .A2(n6256), .ZN(n4911) );
  NOR2_X1 U6022 ( .A1(n6477), .A2(n4902), .ZN(n4906) );
  OR2_X1 U6023 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  NAND2_X1 U6024 ( .A1(n4905), .A2(n6143), .ZN(n6478) );
  AOI21_X1 U6025 ( .B1(n4906), .B2(n6478), .A(n6433), .ZN(n6443) );
  NOR2_X1 U6026 ( .A1(n4907), .A2(n6443), .ZN(n4909) );
  OAI21_X1 U6027 ( .B1(n5459), .B2(n4906), .A(n5462), .ZN(n6469) );
  AOI21_X1 U6028 ( .B1(n4907), .B2(n5959), .A(n6469), .ZN(n6442) );
  INV_X1 U6029 ( .A(n6442), .ZN(n4908) );
  MUX2_X1 U6030 ( .A(n4909), .B(n4908), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4910) );
  AOI211_X1 U6031 ( .C1(n6476), .C2(REIP_REG_6__SCAN_IN), .A(n4911), .B(n4910), 
        .ZN(n4912) );
  OAI21_X1 U6032 ( .B1(n6455), .B2(n6365), .A(n4912), .ZN(U3012) );
  OR2_X1 U6033 ( .A1(n5009), .A2(n3717), .ZN(n4913) );
  NAND3_X1 U6034 ( .A1(n4286), .A2(n4916), .A3(n5502), .ZN(n4917) );
  AND2_X1 U6035 ( .A1(n4918), .A2(n4917), .ZN(n4919) );
  AOI22_X1 U6036 ( .A1(n6286), .A2(n6435), .B1(n6288), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4921) );
  INV_X1 U6037 ( .A(n6173), .ZN(n4920) );
  NAND2_X1 U6038 ( .A1(n5621), .A2(n4920), .ZN(n6257) );
  OAI211_X1 U6039 ( .C1(n6258), .C2(n4922), .A(n4921), .B(n6257), .ZN(n4928)
         );
  INV_X1 U6040 ( .A(n5181), .ZN(n4923) );
  OAI21_X1 U6041 ( .B1(n6272), .B2(n4923), .A(n5621), .ZN(n6255) );
  INV_X1 U6042 ( .A(n6255), .ZN(n4926) );
  AOI21_X1 U6043 ( .B1(n6247), .B2(n4924), .A(REIP_REG_5__SCAN_IN), .ZN(n4925)
         );
  NOR2_X1 U6044 ( .A1(n4926), .A2(n4925), .ZN(n4927) );
  AOI211_X1 U6045 ( .C1(n6294), .C2(n4929), .A(n4928), .B(n4927), .ZN(n4930)
         );
  OAI21_X1 U6046 ( .B1(n4931), .B2(n5305), .A(n4930), .ZN(U2822) );
  INV_X1 U6047 ( .A(n6603), .ZN(n4932) );
  NOR2_X2 U6048 ( .A1(n5185), .A2(n5316), .ZN(n5229) );
  NOR3_X1 U6049 ( .A1(n4932), .A2(n5229), .A3(n6496), .ZN(n4933) );
  NAND2_X1 U6050 ( .A1(n5187), .A2(n4712), .ZN(n4939) );
  OAI21_X1 U6051 ( .B1(n4933), .B2(n6499), .A(n4939), .ZN(n4938) );
  NOR2_X1 U6052 ( .A1(n6487), .A2(n5189), .ZN(n5196) );
  NAND2_X1 U6053 ( .A1(n6613), .A2(n5196), .ZN(n4966) );
  INV_X1 U6054 ( .A(n4975), .ZN(n4934) );
  OR2_X1 U6055 ( .A1(n4934), .A2(n6488), .ZN(n4940) );
  AOI21_X1 U6056 ( .B1(n4940), .B2(STATE2_REG_2__SCAN_IN), .A(n4935), .ZN(
        n4936) );
  INV_X1 U6057 ( .A(n4936), .ZN(n5098) );
  NOR2_X1 U6058 ( .A1(n4941), .A2(n4510), .ZN(n5979) );
  AOI211_X1 U6059 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4966), .A(n5098), .B(
        n5979), .ZN(n4937) );
  NAND2_X1 U6060 ( .A1(n4964), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4945)
         );
  INV_X1 U6061 ( .A(n6513), .ZN(n6554) );
  INV_X1 U6062 ( .A(n4939), .ZN(n4942) );
  INV_X1 U6063 ( .A(n4940), .ZN(n5101) );
  AND2_X1 U6064 ( .A1(n4941), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6489) );
  AOI22_X1 U6065 ( .A1(n4942), .A2(n6015), .B1(n5101), .B2(n6489), .ZN(n4965)
         );
  OAI22_X1 U6066 ( .A1(n6552), .A2(n4966), .B1(n4965), .B2(n6508), .ZN(n4943)
         );
  AOI21_X1 U6067 ( .B1(n6554), .B2(n5229), .A(n4943), .ZN(n4944) );
  OAI211_X1 U6068 ( .C1(n6603), .C2(n6558), .A(n4945), .B(n4944), .ZN(U3117)
         );
  NAND2_X1 U6069 ( .A1(n4964), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4948)
         );
  INV_X1 U6070 ( .A(n6531), .ZN(n6565) );
  OAI22_X1 U6071 ( .A1(n6563), .A2(n4966), .B1(n4965), .B2(n6526), .ZN(n4946)
         );
  AOI21_X1 U6072 ( .B1(n6565), .B2(n5229), .A(n4946), .ZN(n4947) );
  OAI211_X1 U6073 ( .C1(n6603), .C2(n6569), .A(n4948), .B(n4947), .ZN(U3120)
         );
  NAND2_X1 U6074 ( .A1(n4964), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4951)
         );
  INV_X1 U6075 ( .A(n6507), .ZN(n6018) );
  OAI22_X1 U6076 ( .A1(n6493), .A2(n4966), .B1(n4965), .B2(n6492), .ZN(n4949)
         );
  AOI21_X1 U6077 ( .B1(n6018), .B2(n5229), .A(n4949), .ZN(n4950) );
  OAI211_X1 U6078 ( .C1(n6603), .C2(n6021), .A(n4951), .B(n4950), .ZN(U3116)
         );
  NAND2_X1 U6079 ( .A1(n4964), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4954)
         );
  INV_X1 U6080 ( .A(n6594), .ZN(n6037) );
  OAI22_X1 U6081 ( .A1(n6593), .A2(n4966), .B1(n4965), .B2(n6532), .ZN(n4952)
         );
  AOI21_X1 U6082 ( .B1(n6037), .B2(n5229), .A(n4952), .ZN(n4953) );
  OAI211_X1 U6083 ( .C1(n6603), .C2(n6599), .A(n4954), .B(n4953), .ZN(U3121)
         );
  NAND2_X1 U6084 ( .A1(n4964), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4957)
         );
  INV_X1 U6085 ( .A(n6542), .ZN(n6572) );
  OAI22_X1 U6086 ( .A1(n6570), .A2(n4966), .B1(n4965), .B2(n6537), .ZN(n4955)
         );
  AOI21_X1 U6087 ( .B1(n6572), .B2(n5229), .A(n4955), .ZN(n4956) );
  OAI211_X1 U6088 ( .C1(n6603), .C2(n6576), .A(n4957), .B(n4956), .ZN(U3122)
         );
  NAND2_X1 U6089 ( .A1(n4964), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4960)
         );
  INV_X1 U6090 ( .A(n6602), .ZN(n6579) );
  OAI22_X1 U6091 ( .A1(n6601), .A2(n4966), .B1(n4965), .B2(n6543), .ZN(n4958)
         );
  AOI21_X1 U6092 ( .B1(n6579), .B2(n5229), .A(n4958), .ZN(n4959) );
  OAI211_X1 U6093 ( .C1(n6603), .C2(n6611), .A(n4960), .B(n4959), .ZN(U3123)
         );
  NAND2_X1 U6094 ( .A1(n4964), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4963)
         );
  INV_X1 U6095 ( .A(n6587), .ZN(n6560) );
  OAI22_X1 U6096 ( .A1(n6586), .A2(n4966), .B1(n4965), .B2(n6521), .ZN(n4961)
         );
  AOI21_X1 U6097 ( .B1(n6560), .B2(n5229), .A(n4961), .ZN(n4962) );
  OAI211_X1 U6098 ( .C1(n6603), .C2(n6592), .A(n4963), .B(n4962), .ZN(U3119)
         );
  NAND2_X1 U6099 ( .A1(n4964), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4969)
         );
  INV_X1 U6100 ( .A(n6520), .ZN(n6026) );
  OAI22_X1 U6101 ( .A1(n6515), .A2(n4966), .B1(n4965), .B2(n6514), .ZN(n4967)
         );
  AOI21_X1 U6102 ( .B1(n6026), .B2(n5229), .A(n4967), .ZN(n4968) );
  OAI211_X1 U6103 ( .C1(n6603), .C2(n6029), .A(n4969), .B(n4968), .ZN(U3118)
         );
  INV_X1 U6104 ( .A(n4782), .ZN(n4970) );
  NAND4_X1 U6105 ( .A1(n4970), .A2(n5316), .A3(n4747), .A4(n3772), .ZN(n5053)
         );
  AOI21_X1 U6106 ( .B1(n4972), .B2(n5187), .A(n4971), .ZN(n4973) );
  OAI21_X1 U6107 ( .B1(n6499), .B2(n5053), .A(n4973), .ZN(n4977) );
  OR2_X1 U6108 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4974), .ZN(n5003)
         );
  NOR2_X1 U6109 ( .A1(n6488), .A2(n4975), .ZN(n5978) );
  OAI21_X1 U6110 ( .B1(n5978), .B2(n4510), .A(n5263), .ZN(n5975) );
  AOI211_X1 U6111 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5003), .A(n5979), .B(
        n5975), .ZN(n4976) );
  NAND2_X1 U6112 ( .A1(n4977), .A2(n4976), .ZN(n5001) );
  NAND2_X1 U6113 ( .A1(n5001), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4982) );
  INV_X1 U6114 ( .A(n5187), .ZN(n4978) );
  NOR3_X1 U6115 ( .A1(n4712), .A2(n4978), .A3(n6496), .ZN(n4979) );
  AOI21_X1 U6116 ( .B1(n5978), .B2(n6489), .A(n4979), .ZN(n5002) );
  OAI22_X1 U6117 ( .A1(n6515), .A2(n5003), .B1(n5002), .B2(n6514), .ZN(n4980)
         );
  AOI21_X1 U6118 ( .B1(n5005), .B2(n6026), .A(n4980), .ZN(n4981) );
  OAI211_X1 U6119 ( .C1(n5053), .C2(n6029), .A(n4982), .B(n4981), .ZN(U3054)
         );
  NAND2_X1 U6120 ( .A1(n5001), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4985) );
  OAI22_X1 U6121 ( .A1(n6601), .A2(n5003), .B1(n5002), .B2(n6543), .ZN(n4983)
         );
  AOI21_X1 U6122 ( .B1(n5005), .B2(n6579), .A(n4983), .ZN(n4984) );
  OAI211_X1 U6123 ( .C1(n5053), .C2(n6611), .A(n4985), .B(n4984), .ZN(U3059)
         );
  NAND2_X1 U6124 ( .A1(n5001), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4988) );
  OAI22_X1 U6125 ( .A1(n6552), .A2(n5003), .B1(n5002), .B2(n6508), .ZN(n4986)
         );
  AOI21_X1 U6126 ( .B1(n5005), .B2(n6554), .A(n4986), .ZN(n4987) );
  OAI211_X1 U6127 ( .C1(n5053), .C2(n6558), .A(n4988), .B(n4987), .ZN(U3053)
         );
  NAND2_X1 U6128 ( .A1(n5001), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4991) );
  OAI22_X1 U6129 ( .A1(n6493), .A2(n5003), .B1(n5002), .B2(n6492), .ZN(n4989)
         );
  AOI21_X1 U6130 ( .B1(n5005), .B2(n6018), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6131 ( .C1(n5053), .C2(n6021), .A(n4991), .B(n4990), .ZN(U3052)
         );
  NAND2_X1 U6132 ( .A1(n5001), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4994) );
  OAI22_X1 U6133 ( .A1(n6570), .A2(n5003), .B1(n5002), .B2(n6537), .ZN(n4992)
         );
  AOI21_X1 U6134 ( .B1(n5005), .B2(n6572), .A(n4992), .ZN(n4993) );
  OAI211_X1 U6135 ( .C1(n5053), .C2(n6576), .A(n4994), .B(n4993), .ZN(U3058)
         );
  NAND2_X1 U6136 ( .A1(n5001), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4997) );
  OAI22_X1 U6137 ( .A1(n6593), .A2(n5003), .B1(n5002), .B2(n6532), .ZN(n4995)
         );
  AOI21_X1 U6138 ( .B1(n5005), .B2(n6037), .A(n4995), .ZN(n4996) );
  OAI211_X1 U6139 ( .C1(n5053), .C2(n6599), .A(n4997), .B(n4996), .ZN(U3057)
         );
  NAND2_X1 U6140 ( .A1(n5001), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5000) );
  OAI22_X1 U6141 ( .A1(n6563), .A2(n5003), .B1(n5002), .B2(n6526), .ZN(n4998)
         );
  AOI21_X1 U6142 ( .B1(n5005), .B2(n6565), .A(n4998), .ZN(n4999) );
  OAI211_X1 U6143 ( .C1(n5053), .C2(n6569), .A(n5000), .B(n4999), .ZN(U3056)
         );
  NAND2_X1 U6144 ( .A1(n5001), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6145 ( .A1(n6586), .A2(n5003), .B1(n5002), .B2(n6521), .ZN(n5004)
         );
  AOI21_X1 U6146 ( .B1(n5005), .B2(n6560), .A(n5004), .ZN(n5006) );
  OAI211_X1 U6147 ( .C1(n5053), .C2(n6592), .A(n5007), .B(n5006), .ZN(U3055)
         );
  OR2_X1 U6148 ( .A1(n5009), .A2(n5008), .ZN(n6265) );
  INV_X1 U6149 ( .A(n6265), .ZN(n6287) );
  AOI22_X1 U6150 ( .A1(n5010), .A2(n6287), .B1(n6288), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5016) );
  INV_X1 U6151 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U6152 ( .A1(n6258), .A2(n5012), .B1(n5621), .B2(n5011), .ZN(n5014)
         );
  OAI22_X1 U6153 ( .A1(n4642), .A2(n6274), .B1(n6272), .B2(REIP_REG_1__SCAN_IN), .ZN(n5013) );
  AOI211_X1 U6154 ( .C1(n6294), .C2(n5012), .A(n5014), .B(n5013), .ZN(n5015)
         );
  OAI211_X1 U6155 ( .C1(n5017), .C2(n5305), .A(n5016), .B(n5015), .ZN(U2826)
         );
  INV_X1 U6156 ( .A(n3772), .ZN(n5139) );
  NOR3_X1 U6157 ( .A1(n5019), .A2(n5139), .A3(n5018), .ZN(n5020) );
  NOR2_X1 U6158 ( .A1(n5020), .A2(n6496), .ZN(n5029) );
  INV_X1 U6159 ( .A(n4712), .ZN(n6485) );
  NOR2_X1 U6160 ( .A1(n5022), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5026)
         );
  AOI21_X1 U6161 ( .B1(n5380), .B2(n5495), .A(n5026), .ZN(n5028) );
  INV_X1 U6162 ( .A(n5028), .ZN(n5023) );
  NAND3_X1 U6163 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6487), .A3(n6623), .ZN(n5371) );
  INV_X1 U6164 ( .A(n5371), .ZN(n5031) );
  NOR4_X1 U6165 ( .A1(n4782), .A2(n5139), .A3(n5024), .A4(n5316), .ZN(n5025)
         );
  INV_X1 U6166 ( .A(n5026), .ZN(n5052) );
  OAI22_X1 U6167 ( .A1(n5053), .A2(n6602), .B1(n6601), .B2(n5052), .ZN(n5027)
         );
  AOI21_X1 U6168 ( .B1(n6548), .B2(n5406), .A(n5027), .ZN(n5033) );
  NAND2_X1 U6169 ( .A1(n5029), .A2(n5028), .ZN(n5030) );
  NAND2_X1 U6170 ( .A1(n5055), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5032) );
  OAI211_X1 U6171 ( .C1(n5058), .C2(n6543), .A(n5033), .B(n5032), .ZN(U3051)
         );
  OAI22_X1 U6172 ( .A1(n5053), .A2(n6513), .B1(n6552), .B2(n5052), .ZN(n5034)
         );
  AOI21_X1 U6173 ( .B1(n6510), .B2(n5406), .A(n5034), .ZN(n5036) );
  NAND2_X1 U6174 ( .A1(n5055), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n5035) );
  OAI211_X1 U6175 ( .C1(n5058), .C2(n6508), .A(n5036), .B(n5035), .ZN(U3045)
         );
  OAI22_X1 U6176 ( .A1(n5053), .A2(n6531), .B1(n6563), .B2(n5052), .ZN(n5037)
         );
  AOI21_X1 U6177 ( .B1(n6528), .B2(n5406), .A(n5037), .ZN(n5039) );
  NAND2_X1 U6178 ( .A1(n5055), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5038) );
  OAI211_X1 U6179 ( .C1(n5058), .C2(n6526), .A(n5039), .B(n5038), .ZN(U3048)
         );
  OAI22_X1 U6180 ( .A1(n5053), .A2(n6594), .B1(n6593), .B2(n5052), .ZN(n5040)
         );
  AOI21_X1 U6181 ( .B1(n6534), .B2(n5406), .A(n5040), .ZN(n5042) );
  NAND2_X1 U6182 ( .A1(n5055), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5041) );
  OAI211_X1 U6183 ( .C1(n5058), .C2(n6532), .A(n5042), .B(n5041), .ZN(U3049)
         );
  OAI22_X1 U6184 ( .A1(n5053), .A2(n6507), .B1(n6493), .B2(n5052), .ZN(n5043)
         );
  AOI21_X1 U6185 ( .B1(n6504), .B2(n5406), .A(n5043), .ZN(n5045) );
  NAND2_X1 U6186 ( .A1(n5055), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n5044) );
  OAI211_X1 U6187 ( .C1(n5058), .C2(n6492), .A(n5045), .B(n5044), .ZN(U3044)
         );
  OAI22_X1 U6188 ( .A1(n5053), .A2(n6542), .B1(n6570), .B2(n5052), .ZN(n5046)
         );
  AOI21_X1 U6189 ( .B1(n6539), .B2(n5406), .A(n5046), .ZN(n5048) );
  NAND2_X1 U6190 ( .A1(n5055), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5047) );
  OAI211_X1 U6191 ( .C1(n5058), .C2(n6537), .A(n5048), .B(n5047), .ZN(U3050)
         );
  OAI22_X1 U6192 ( .A1(n5053), .A2(n6520), .B1(n6515), .B2(n5052), .ZN(n5049)
         );
  AOI21_X1 U6193 ( .B1(n6517), .B2(n5406), .A(n5049), .ZN(n5051) );
  NAND2_X1 U6194 ( .A1(n5055), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5050) );
  OAI211_X1 U6195 ( .C1(n5058), .C2(n6514), .A(n5051), .B(n5050), .ZN(U3046)
         );
  OAI22_X1 U6196 ( .A1(n5053), .A2(n6587), .B1(n6586), .B2(n5052), .ZN(n5054)
         );
  AOI21_X1 U6197 ( .B1(n6523), .B2(n5406), .A(n5054), .ZN(n5057) );
  NAND2_X1 U6198 ( .A1(n5055), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5056) );
  OAI211_X1 U6199 ( .C1(n5058), .C2(n6521), .A(n5057), .B(n5056), .ZN(U3047)
         );
  OR2_X1 U6200 ( .A1(n5066), .A2(n6177), .ZN(n5060) );
  NAND2_X1 U6201 ( .A1(n4712), .A2(n5495), .ZN(n6010) );
  INV_X1 U6202 ( .A(n6010), .ZN(n5188) );
  NAND2_X1 U6203 ( .A1(n4608), .A2(n4577), .ZN(n5138) );
  INV_X1 U6204 ( .A(n5138), .ZN(n5061) );
  NAND3_X1 U6205 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6623), .A3(n6618), .ZN(n5097) );
  NOR2_X1 U6206 ( .A1(n6613), .A2(n5097), .ZN(n5067) );
  AOI21_X1 U6207 ( .B1(n5188), .B2(n5061), .A(n5067), .ZN(n5065) );
  AOI22_X1 U6208 ( .A1(n5063), .A2(n5065), .B1(n6496), .B2(n5097), .ZN(n5062)
         );
  NAND2_X1 U6209 ( .A1(n6012), .A2(n5062), .ZN(n5090) );
  INV_X1 U6210 ( .A(n5063), .ZN(n5064) );
  OAI22_X1 U6211 ( .A1(n5065), .A2(n5064), .B1(n4510), .B2(n5097), .ZN(n5089)
         );
  AOI22_X1 U6212 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5090), .B1(n5212), 
        .B2(n5089), .ZN(n5070) );
  INV_X1 U6213 ( .A(n5067), .ZN(n5091) );
  OAI22_X1 U6214 ( .A1(n5269), .A2(n6520), .B1(n6515), .B2(n5091), .ZN(n5068)
         );
  AOI21_X1 U6215 ( .B1(n6517), .B2(n5095), .A(n5068), .ZN(n5069) );
  NAND2_X1 U6216 ( .A1(n5070), .A2(n5069), .ZN(U3094) );
  AOI22_X1 U6217 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5090), .B1(n5231), 
        .B2(n5089), .ZN(n5073) );
  OAI22_X1 U6218 ( .A1(n5269), .A2(n6507), .B1(n6493), .B2(n5091), .ZN(n5071)
         );
  AOI21_X1 U6219 ( .B1(n6504), .B2(n5095), .A(n5071), .ZN(n5072) );
  NAND2_X1 U6220 ( .A1(n5073), .A2(n5072), .ZN(U3092) );
  AOI22_X1 U6221 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5090), .B1(n6566), 
        .B2(n5089), .ZN(n5076) );
  OAI22_X1 U6222 ( .A1(n5269), .A2(n6531), .B1(n6563), .B2(n5091), .ZN(n5074)
         );
  AOI21_X1 U6223 ( .B1(n6528), .B2(n5095), .A(n5074), .ZN(n5075) );
  NAND2_X1 U6224 ( .A1(n5076), .A2(n5075), .ZN(U3096) );
  AOI22_X1 U6225 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5090), .B1(n6573), 
        .B2(n5089), .ZN(n5079) );
  OAI22_X1 U6226 ( .A1(n5269), .A2(n6542), .B1(n6570), .B2(n5091), .ZN(n5077)
         );
  AOI21_X1 U6227 ( .B1(n6539), .B2(n5095), .A(n5077), .ZN(n5078) );
  NAND2_X1 U6228 ( .A1(n5079), .A2(n5078), .ZN(U3098) );
  AOI22_X1 U6229 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5090), .B1(n6555), 
        .B2(n5089), .ZN(n5082) );
  OAI22_X1 U6230 ( .A1(n5269), .A2(n6513), .B1(n6552), .B2(n5091), .ZN(n5080)
         );
  AOI21_X1 U6231 ( .B1(n6510), .B2(n5095), .A(n5080), .ZN(n5081) );
  NAND2_X1 U6232 ( .A1(n5082), .A2(n5081), .ZN(U3093) );
  AOI22_X1 U6233 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5090), .B1(n6596), 
        .B2(n5089), .ZN(n5085) );
  OAI22_X1 U6234 ( .A1(n5269), .A2(n6594), .B1(n6593), .B2(n5091), .ZN(n5083)
         );
  AOI21_X1 U6235 ( .B1(n6534), .B2(n5095), .A(n5083), .ZN(n5084) );
  NAND2_X1 U6236 ( .A1(n5085), .A2(n5084), .ZN(U3097) );
  AOI22_X1 U6237 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5090), .B1(n6589), 
        .B2(n5089), .ZN(n5088) );
  OAI22_X1 U6238 ( .A1(n5269), .A2(n6587), .B1(n6586), .B2(n5091), .ZN(n5086)
         );
  AOI21_X1 U6239 ( .B1(n6523), .B2(n5095), .A(n5086), .ZN(n5087) );
  NAND2_X1 U6240 ( .A1(n5088), .A2(n5087), .ZN(U3095) );
  AOI22_X1 U6241 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5090), .B1(n6606), 
        .B2(n5089), .ZN(n5094) );
  OAI22_X1 U6242 ( .A1(n5269), .A2(n6602), .B1(n6601), .B2(n5091), .ZN(n5092)
         );
  AOI21_X1 U6243 ( .B1(n6548), .B2(n5095), .A(n5092), .ZN(n5093) );
  NAND2_X1 U6244 ( .A1(n5094), .A2(n5093), .ZN(U3099) );
  NOR3_X1 U6245 ( .A1(n5095), .A2(n6580), .A3(n6496), .ZN(n5096) );
  NOR2_X1 U6246 ( .A1(n5096), .A2(n6499), .ZN(n5100) );
  NOR2_X1 U6247 ( .A1(n6485), .A2(n5138), .ZN(n5102) );
  OR2_X1 U6248 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5097), .ZN(n5126)
         );
  AOI211_X1 U6249 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5126), .A(n6489), .B(
        n5098), .ZN(n5099) );
  NAND2_X1 U6250 ( .A1(n5124), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5105) );
  AOI22_X1 U6251 ( .A1(n5102), .A2(n6015), .B1(n5979), .B2(n5101), .ZN(n5125)
         );
  OAI22_X1 U6252 ( .A1(n6586), .A2(n5126), .B1(n5125), .B2(n6521), .ZN(n5103)
         );
  AOI21_X1 U6253 ( .B1(n6580), .B2(n6523), .A(n5103), .ZN(n5104) );
  OAI211_X1 U6254 ( .C1(n5130), .C2(n6587), .A(n5105), .B(n5104), .ZN(U3087)
         );
  NAND2_X1 U6255 ( .A1(n5124), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n5108) );
  OAI22_X1 U6256 ( .A1(n6552), .A2(n5126), .B1(n5125), .B2(n6508), .ZN(n5106)
         );
  AOI21_X1 U6257 ( .B1(n6580), .B2(n6510), .A(n5106), .ZN(n5107) );
  OAI211_X1 U6258 ( .C1(n5130), .C2(n6513), .A(n5108), .B(n5107), .ZN(U3085)
         );
  NAND2_X1 U6259 ( .A1(n5124), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5111) );
  OAI22_X1 U6260 ( .A1(n6563), .A2(n5126), .B1(n5125), .B2(n6526), .ZN(n5109)
         );
  AOI21_X1 U6261 ( .B1(n6580), .B2(n6528), .A(n5109), .ZN(n5110) );
  OAI211_X1 U6262 ( .C1(n5130), .C2(n6531), .A(n5111), .B(n5110), .ZN(U3088)
         );
  NAND2_X1 U6263 ( .A1(n5124), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5114) );
  OAI22_X1 U6264 ( .A1(n6601), .A2(n5126), .B1(n5125), .B2(n6543), .ZN(n5112)
         );
  AOI21_X1 U6265 ( .B1(n6580), .B2(n6548), .A(n5112), .ZN(n5113) );
  OAI211_X1 U6266 ( .C1(n5130), .C2(n6602), .A(n5114), .B(n5113), .ZN(U3091)
         );
  NAND2_X1 U6267 ( .A1(n5124), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U6268 ( .A1(n6515), .A2(n5126), .B1(n5125), .B2(n6514), .ZN(n5115)
         );
  AOI21_X1 U6269 ( .B1(n6580), .B2(n6517), .A(n5115), .ZN(n5116) );
  OAI211_X1 U6270 ( .C1(n5130), .C2(n6520), .A(n5117), .B(n5116), .ZN(U3086)
         );
  NAND2_X1 U6271 ( .A1(n5124), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5120) );
  OAI22_X1 U6272 ( .A1(n6570), .A2(n5126), .B1(n5125), .B2(n6537), .ZN(n5118)
         );
  AOI21_X1 U6273 ( .B1(n6580), .B2(n6539), .A(n5118), .ZN(n5119) );
  OAI211_X1 U6274 ( .C1(n5130), .C2(n6542), .A(n5120), .B(n5119), .ZN(U3090)
         );
  NAND2_X1 U6275 ( .A1(n5124), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5123) );
  OAI22_X1 U6276 ( .A1(n6493), .A2(n5126), .B1(n5125), .B2(n6492), .ZN(n5121)
         );
  AOI21_X1 U6277 ( .B1(n6580), .B2(n6504), .A(n5121), .ZN(n5122) );
  OAI211_X1 U6278 ( .C1(n5130), .C2(n6507), .A(n5123), .B(n5122), .ZN(U3084)
         );
  NAND2_X1 U6279 ( .A1(n5124), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5129) );
  OAI22_X1 U6280 ( .A1(n6593), .A2(n5126), .B1(n5125), .B2(n6532), .ZN(n5127)
         );
  AOI21_X1 U6281 ( .B1(n6580), .B2(n6534), .A(n5127), .ZN(n5128) );
  OAI211_X1 U6282 ( .C1(n5130), .C2(n6594), .A(n5129), .B(n5128), .ZN(U3089)
         );
  XOR2_X1 U6283 ( .A(n4856), .B(n5131), .Z(n6366) );
  OAI22_X1 U6284 ( .A1(n5709), .A2(n6256), .B1(n6307), .B2(n6252), .ZN(n5132)
         );
  AOI21_X1 U6285 ( .B1(n6366), .B2(n6304), .A(n5132), .ZN(n5133) );
  INV_X1 U6286 ( .A(n5133), .ZN(U2853) );
  XOR2_X1 U6287 ( .A(n5135), .B(n5134), .Z(n5244) );
  INV_X1 U6288 ( .A(n5244), .ZN(n5184) );
  AOI21_X1 U6289 ( .B1(n5136), .B2(n4899), .A(n5252), .ZN(n6424) );
  AOI22_X1 U6290 ( .A1(n6303), .A2(n6424), .B1(EBX_REG_7__SCAN_IN), .B2(n4391), 
        .ZN(n5137) );
  OAI21_X1 U6291 ( .B1(n5184), .B2(n5704), .A(n5137), .ZN(U2852) );
  NOR2_X1 U6292 ( .A1(n4712), .A2(n5138), .ZN(n5980) );
  NAND3_X1 U6293 ( .A1(n6487), .A2(n6623), .A3(n6618), .ZN(n5974) );
  NOR2_X1 U6294 ( .A1(n6613), .A2(n5974), .ZN(n5146) );
  AOI21_X1 U6295 ( .B1(n5980), .B2(n5495), .A(n5146), .ZN(n5143) );
  OR2_X1 U6296 ( .A1(n5145), .A2(n6177), .ZN(n5140) );
  NAND2_X1 U6297 ( .A1(n5140), .A2(n6015), .ZN(n5144) );
  INV_X1 U6298 ( .A(n5144), .ZN(n5141) );
  AOI22_X1 U6299 ( .A1(n5143), .A2(n5141), .B1(n6496), .B2(n5974), .ZN(n5142)
         );
  NAND2_X1 U6300 ( .A1(n6012), .A2(n5142), .ZN(n5169) );
  OAI22_X1 U6301 ( .A1(n5144), .A2(n5143), .B1(n4510), .B2(n5974), .ZN(n5168)
         );
  AOI22_X1 U6302 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5169), .B1(n6589), 
        .B2(n5168), .ZN(n5149) );
  INV_X1 U6303 ( .A(n5146), .ZN(n5170) );
  OAI22_X1 U6304 ( .A1(n5409), .A2(n6587), .B1(n6586), .B2(n5170), .ZN(n5147)
         );
  AOI21_X1 U6305 ( .B1(n6523), .B2(n5972), .A(n5147), .ZN(n5148) );
  NAND2_X1 U6306 ( .A1(n5149), .A2(n5148), .ZN(U3031) );
  AOI22_X1 U6307 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5169), .B1(n6555), 
        .B2(n5168), .ZN(n5152) );
  OAI22_X1 U6308 ( .A1(n5409), .A2(n6513), .B1(n6552), .B2(n5170), .ZN(n5150)
         );
  AOI21_X1 U6309 ( .B1(n6510), .B2(n5972), .A(n5150), .ZN(n5151) );
  NAND2_X1 U6310 ( .A1(n5152), .A2(n5151), .ZN(U3029) );
  AOI22_X1 U6311 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5169), .B1(n5231), 
        .B2(n5168), .ZN(n5155) );
  OAI22_X1 U6312 ( .A1(n5409), .A2(n6507), .B1(n6493), .B2(n5170), .ZN(n5153)
         );
  AOI21_X1 U6313 ( .B1(n6504), .B2(n5972), .A(n5153), .ZN(n5154) );
  NAND2_X1 U6314 ( .A1(n5155), .A2(n5154), .ZN(U3028) );
  AOI22_X1 U6315 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5169), .B1(n6596), 
        .B2(n5168), .ZN(n5158) );
  OAI22_X1 U6316 ( .A1(n5409), .A2(n6594), .B1(n6593), .B2(n5170), .ZN(n5156)
         );
  AOI21_X1 U6317 ( .B1(n6534), .B2(n5972), .A(n5156), .ZN(n5157) );
  NAND2_X1 U6318 ( .A1(n5158), .A2(n5157), .ZN(U3033) );
  AOI22_X1 U6319 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5169), .B1(n6566), 
        .B2(n5168), .ZN(n5161) );
  OAI22_X1 U6320 ( .A1(n5409), .A2(n6531), .B1(n6563), .B2(n5170), .ZN(n5159)
         );
  AOI21_X1 U6321 ( .B1(n6528), .B2(n5972), .A(n5159), .ZN(n5160) );
  NAND2_X1 U6322 ( .A1(n5161), .A2(n5160), .ZN(U3032) );
  AOI22_X1 U6323 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5169), .B1(n6606), 
        .B2(n5168), .ZN(n5164) );
  OAI22_X1 U6324 ( .A1(n5409), .A2(n6602), .B1(n6601), .B2(n5170), .ZN(n5162)
         );
  AOI21_X1 U6325 ( .B1(n6548), .B2(n5972), .A(n5162), .ZN(n5163) );
  NAND2_X1 U6326 ( .A1(n5164), .A2(n5163), .ZN(U3035) );
  AOI22_X1 U6327 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5169), .B1(n6573), 
        .B2(n5168), .ZN(n5167) );
  OAI22_X1 U6328 ( .A1(n5409), .A2(n6542), .B1(n6570), .B2(n5170), .ZN(n5165)
         );
  AOI21_X1 U6329 ( .B1(n6539), .B2(n5972), .A(n5165), .ZN(n5166) );
  NAND2_X1 U6330 ( .A1(n5167), .A2(n5166), .ZN(U3034) );
  AOI22_X1 U6331 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5169), .B1(n5212), 
        .B2(n5168), .ZN(n5173) );
  OAI22_X1 U6332 ( .A1(n5409), .A2(n6520), .B1(n6515), .B2(n5170), .ZN(n5171)
         );
  AOI21_X1 U6333 ( .B1(n6517), .B2(n5972), .A(n5171), .ZN(n5172) );
  NAND2_X1 U6334 ( .A1(n5173), .A2(n5172), .ZN(U3030) );
  INV_X1 U6335 ( .A(n6366), .ZN(n5174) );
  OAI222_X1 U6336 ( .A1(n6086), .A2(n5174), .B1(n5738), .B2(n3814), .C1(n7103), 
        .C2(n5739), .ZN(U2885) );
  INV_X1 U6337 ( .A(n5242), .ZN(n5180) );
  INV_X1 U6338 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5176) );
  AOI22_X1 U6339 ( .A1(n6286), .A2(n6424), .B1(n6288), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5175) );
  OAI211_X1 U6340 ( .C1(n6258), .C2(n5176), .A(n5175), .B(n6257), .ZN(n5179)
         );
  INV_X1 U6341 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6686) );
  AND3_X1 U6342 ( .A1(n6247), .A2(n6686), .A3(n5177), .ZN(n5178) );
  AOI211_X1 U6343 ( .C1(n6294), .C2(n5180), .A(n5179), .B(n5178), .ZN(n5183)
         );
  NOR3_X1 U6344 ( .A1(n6272), .A2(REIP_REG_6__SCAN_IN), .A3(n5181), .ZN(n6254)
         );
  OAI21_X1 U6345 ( .B1(n6254), .B2(n6255), .A(REIP_REG_7__SCAN_IN), .ZN(n5182)
         );
  OAI211_X1 U6346 ( .C1(n5184), .C2(n6212), .A(n5183), .B(n5182), .ZN(U2820)
         );
  OAI222_X1 U6347 ( .A1(n6086), .A2(n5184), .B1(n5738), .B2(n3820), .C1(n7065), 
        .C2(n5739), .ZN(U2884) );
  NOR2_X2 U6348 ( .A1(n5185), .A2(n5969), .ZN(n5350) );
  AND2_X1 U6349 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5196), .ZN(n5186)
         );
  INV_X1 U6350 ( .A(n5186), .ZN(n5235) );
  NAND2_X1 U6351 ( .A1(n5229), .A2(n6510), .ZN(n5201) );
  AOI21_X1 U6352 ( .B1(n5188), .B2(n5187), .A(n5186), .ZN(n5195) );
  OR2_X1 U6353 ( .A1(n5195), .A2(n6496), .ZN(n5193) );
  INV_X1 U6354 ( .A(n5189), .ZN(n5191) );
  AND2_X1 U6355 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6356 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  NAND2_X1 U6357 ( .A1(n5193), .A2(n5192), .ZN(n5232) );
  NAND2_X1 U6358 ( .A1(n5195), .A2(n5194), .ZN(n5199) );
  INV_X1 U6359 ( .A(n5196), .ZN(n5197) );
  NAND2_X1 U6360 ( .A1(n6496), .A2(n5197), .ZN(n5198) );
  OAI211_X1 U6361 ( .C1(n6496), .C2(n5199), .A(n6012), .B(n5198), .ZN(n5230)
         );
  AOI22_X1 U6362 ( .A1(n5232), .A2(n6555), .B1(INSTQUEUE_REG_13__1__SCAN_IN), 
        .B2(n5230), .ZN(n5200) );
  OAI211_X1 U6363 ( .C1(n5235), .C2(n6552), .A(n5201), .B(n5200), .ZN(n5202)
         );
  AOI21_X1 U6364 ( .B1(n6554), .B2(n5350), .A(n5202), .ZN(n5203) );
  INV_X1 U6365 ( .A(n5203), .ZN(U3125) );
  NAND2_X1 U6366 ( .A1(n5229), .A2(n6523), .ZN(n5205) );
  AOI22_X1 U6367 ( .A1(n5232), .A2(n6589), .B1(INSTQUEUE_REG_13__3__SCAN_IN), 
        .B2(n5230), .ZN(n5204) );
  OAI211_X1 U6368 ( .C1(n5235), .C2(n6586), .A(n5205), .B(n5204), .ZN(n5206)
         );
  AOI21_X1 U6369 ( .B1(n6560), .B2(n5350), .A(n5206), .ZN(n5207) );
  INV_X1 U6370 ( .A(n5207), .ZN(U3127) );
  NAND2_X1 U6371 ( .A1(n5229), .A2(n6528), .ZN(n5209) );
  AOI22_X1 U6372 ( .A1(n5232), .A2(n6566), .B1(INSTQUEUE_REG_13__4__SCAN_IN), 
        .B2(n5230), .ZN(n5208) );
  OAI211_X1 U6373 ( .C1(n5235), .C2(n6563), .A(n5209), .B(n5208), .ZN(n5210)
         );
  AOI21_X1 U6374 ( .B1(n6565), .B2(n5350), .A(n5210), .ZN(n5211) );
  INV_X1 U6375 ( .A(n5211), .ZN(U3128) );
  NAND2_X1 U6376 ( .A1(n5229), .A2(n6517), .ZN(n5214) );
  AOI22_X1 U6377 ( .A1(n5232), .A2(n5212), .B1(INSTQUEUE_REG_13__2__SCAN_IN), 
        .B2(n5230), .ZN(n5213) );
  OAI211_X1 U6378 ( .C1(n5235), .C2(n6515), .A(n5214), .B(n5213), .ZN(n5215)
         );
  AOI21_X1 U6379 ( .B1(n6026), .B2(n5350), .A(n5215), .ZN(n5216) );
  INV_X1 U6380 ( .A(n5216), .ZN(U3126) );
  NAND2_X1 U6381 ( .A1(n5229), .A2(n6534), .ZN(n5218) );
  AOI22_X1 U6382 ( .A1(n5232), .A2(n6596), .B1(INSTQUEUE_REG_13__5__SCAN_IN), 
        .B2(n5230), .ZN(n5217) );
  OAI211_X1 U6383 ( .C1(n5235), .C2(n6593), .A(n5218), .B(n5217), .ZN(n5219)
         );
  AOI21_X1 U6384 ( .B1(n6037), .B2(n5350), .A(n5219), .ZN(n5220) );
  INV_X1 U6385 ( .A(n5220), .ZN(U3129) );
  NAND2_X1 U6386 ( .A1(n5229), .A2(n6548), .ZN(n5222) );
  AOI22_X1 U6387 ( .A1(n5232), .A2(n6606), .B1(INSTQUEUE_REG_13__7__SCAN_IN), 
        .B2(n5230), .ZN(n5221) );
  OAI211_X1 U6388 ( .C1(n5235), .C2(n6601), .A(n5222), .B(n5221), .ZN(n5223)
         );
  AOI21_X1 U6389 ( .B1(n6579), .B2(n5350), .A(n5223), .ZN(n5224) );
  INV_X1 U6390 ( .A(n5224), .ZN(U3131) );
  NAND2_X1 U6391 ( .A1(n5229), .A2(n6539), .ZN(n5226) );
  AOI22_X1 U6392 ( .A1(n5232), .A2(n6573), .B1(INSTQUEUE_REG_13__6__SCAN_IN), 
        .B2(n5230), .ZN(n5225) );
  OAI211_X1 U6393 ( .C1(n5235), .C2(n6570), .A(n5226), .B(n5225), .ZN(n5227)
         );
  AOI21_X1 U6394 ( .B1(n6572), .B2(n5350), .A(n5227), .ZN(n5228) );
  INV_X1 U6395 ( .A(n5228), .ZN(U3130) );
  NAND2_X1 U6396 ( .A1(n5229), .A2(n6504), .ZN(n5234) );
  AOI22_X1 U6397 ( .A1(n5232), .A2(n5231), .B1(INSTQUEUE_REG_13__0__SCAN_IN), 
        .B2(n5230), .ZN(n5233) );
  OAI211_X1 U6398 ( .C1(n6493), .C2(n5235), .A(n5234), .B(n5233), .ZN(n5236)
         );
  AOI21_X1 U6399 ( .B1(n6018), .B2(n5350), .A(n5236), .ZN(n5237) );
  INV_X1 U6400 ( .A(n5237), .ZN(U3124) );
  OAI21_X1 U6401 ( .B1(n5238), .B2(n5240), .A(n5239), .ZN(n6425) );
  NAND2_X1 U6402 ( .A1(n6476), .A2(REIP_REG_7__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U6403 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5241)
         );
  OAI211_X1 U6404 ( .C1(n6390), .C2(n5242), .A(n6422), .B(n5241), .ZN(n5243)
         );
  AOI21_X1 U6405 ( .B1(n5244), .B2(n6385), .A(n5243), .ZN(n5245) );
  OAI21_X1 U6406 ( .B1(n6425), .B2(n6364), .A(n5245), .ZN(U2979) );
  OAI21_X1 U6407 ( .B1(n5246), .B2(n5249), .A(n5248), .ZN(n5354) );
  NOR2_X1 U6408 ( .A1(n6246), .A2(n5250), .ZN(n5259) );
  OAI21_X1 U6409 ( .B1(n5253), .B2(n5252), .A(n5251), .ZN(n6416) );
  INV_X1 U6410 ( .A(n5367), .ZN(n5254) );
  NAND2_X1 U6411 ( .A1(n6294), .A2(n5254), .ZN(n5255) );
  OAI21_X1 U6412 ( .B1(n6274), .B2(n6416), .A(n5255), .ZN(n5258) );
  OAI21_X1 U6413 ( .B1(n6272), .B2(n6246), .A(n5621), .ZN(n6242) );
  AOI22_X1 U6414 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6285), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6242), .ZN(n5256) );
  OAI211_X1 U6415 ( .C1(n6270), .C2(n5355), .A(n5256), .B(n6257), .ZN(n5257)
         );
  AOI211_X1 U6416 ( .C1(n6247), .C2(n5259), .A(n5258), .B(n5257), .ZN(n5260)
         );
  OAI21_X1 U6417 ( .B1(n6212), .B2(n5354), .A(n5260), .ZN(U2819) );
  NAND2_X1 U6418 ( .A1(n5269), .A2(n6610), .ZN(n5261) );
  AOI21_X1 U6419 ( .B1(n5261), .B2(STATEBS16_REG_SCAN_IN), .A(n6496), .ZN(
        n5267) );
  INV_X1 U6420 ( .A(n5979), .ZN(n5378) );
  NOR2_X1 U6421 ( .A1(n5378), .A2(n6487), .ZN(n5262) );
  OAI21_X1 U6422 ( .B1(n6488), .B2(n4510), .A(n5263), .ZN(n5319) );
  NOR2_X1 U6423 ( .A1(n6489), .A2(n5319), .ZN(n5375) );
  INV_X1 U6424 ( .A(n5264), .ZN(n5266) );
  OR2_X1 U6425 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5265), .ZN(n5292)
         );
  AOI22_X1 U6426 ( .A1(n5267), .A2(n5266), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5292), .ZN(n5268) );
  NAND2_X1 U6427 ( .A1(n5291), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5272)
         );
  OAI22_X1 U6428 ( .A1(n6610), .A2(n6531), .B1(n5292), .B2(n6563), .ZN(n5270)
         );
  AOI21_X1 U6429 ( .B1(n5294), .B2(n6528), .A(n5270), .ZN(n5271) );
  OAI211_X1 U6430 ( .C1(n5297), .C2(n6526), .A(n5272), .B(n5271), .ZN(U3104)
         );
  NAND2_X1 U6431 ( .A1(n5291), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5275)
         );
  OAI22_X1 U6432 ( .A1(n6610), .A2(n6594), .B1(n5292), .B2(n6593), .ZN(n5273)
         );
  AOI21_X1 U6433 ( .B1(n5294), .B2(n6534), .A(n5273), .ZN(n5274) );
  OAI211_X1 U6434 ( .C1(n5297), .C2(n6532), .A(n5275), .B(n5274), .ZN(U3105)
         );
  NAND2_X1 U6435 ( .A1(n5291), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5278)
         );
  OAI22_X1 U6436 ( .A1(n6610), .A2(n6542), .B1(n5292), .B2(n6570), .ZN(n5276)
         );
  AOI21_X1 U6437 ( .B1(n5294), .B2(n6539), .A(n5276), .ZN(n5277) );
  OAI211_X1 U6438 ( .C1(n5297), .C2(n6537), .A(n5278), .B(n5277), .ZN(U3106)
         );
  NAND2_X1 U6439 ( .A1(n5291), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5281)
         );
  OAI22_X1 U6440 ( .A1(n6610), .A2(n6602), .B1(n5292), .B2(n6601), .ZN(n5279)
         );
  AOI21_X1 U6441 ( .B1(n5294), .B2(n6548), .A(n5279), .ZN(n5280) );
  OAI211_X1 U6442 ( .C1(n5297), .C2(n6543), .A(n5281), .B(n5280), .ZN(U3107)
         );
  NAND2_X1 U6443 ( .A1(n5291), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5284)
         );
  OAI22_X1 U6444 ( .A1(n6610), .A2(n6513), .B1(n5292), .B2(n6552), .ZN(n5282)
         );
  AOI21_X1 U6445 ( .B1(n5294), .B2(n6510), .A(n5282), .ZN(n5283) );
  OAI211_X1 U6446 ( .C1(n5297), .C2(n6508), .A(n5284), .B(n5283), .ZN(U3101)
         );
  NAND2_X1 U6447 ( .A1(n5291), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5287)
         );
  OAI22_X1 U6448 ( .A1(n6610), .A2(n6520), .B1(n5292), .B2(n6515), .ZN(n5285)
         );
  AOI21_X1 U6449 ( .B1(n5294), .B2(n6517), .A(n5285), .ZN(n5286) );
  OAI211_X1 U6450 ( .C1(n5297), .C2(n6514), .A(n5287), .B(n5286), .ZN(U3102)
         );
  NAND2_X1 U6451 ( .A1(n5291), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5290)
         );
  OAI22_X1 U6452 ( .A1(n6610), .A2(n6587), .B1(n5292), .B2(n6586), .ZN(n5288)
         );
  AOI21_X1 U6453 ( .B1(n5294), .B2(n6523), .A(n5288), .ZN(n5289) );
  OAI211_X1 U6454 ( .C1(n5297), .C2(n6521), .A(n5290), .B(n5289), .ZN(U3103)
         );
  NAND2_X1 U6455 ( .A1(n5291), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5296)
         );
  OAI22_X1 U6456 ( .A1(n6610), .A2(n6507), .B1(n6493), .B2(n5292), .ZN(n5293)
         );
  AOI21_X1 U6457 ( .B1(n5294), .B2(n6504), .A(n5293), .ZN(n5295) );
  OAI211_X1 U6458 ( .C1(n5297), .C2(n6492), .A(n5296), .B(n5295), .ZN(U3100)
         );
  OAI22_X1 U6459 ( .A1(n5298), .A2(n6270), .B1(n6265), .B2(n4752), .ZN(n5302)
         );
  OAI21_X1 U6460 ( .B1(n6285), .B2(n6294), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5299) );
  OAI21_X1 U6461 ( .B1(n5300), .B2(n6274), .A(n5299), .ZN(n5301) );
  AOI211_X1 U6462 ( .C1(REIP_REG_0__SCAN_IN), .C2(n6263), .A(n5302), .B(n5301), 
        .ZN(n5303) );
  OAI21_X1 U6463 ( .B1(n5305), .B2(n5304), .A(n5303), .ZN(U2827) );
  INV_X1 U6464 ( .A(n5305), .ZN(n6283) );
  NAND2_X1 U6465 ( .A1(n6384), .A2(n6283), .ZN(n5313) );
  OAI21_X1 U6466 ( .B1(n6272), .B2(REIP_REG_1__SCAN_IN), .A(n5621), .ZN(n6281)
         );
  OAI22_X1 U6467 ( .A1(n4608), .A2(n6265), .B1(n6270), .B2(n5306), .ZN(n5311)
         );
  INV_X1 U6468 ( .A(n6389), .ZN(n5307) );
  AOI22_X1 U6469 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6285), .B1(n6294), 
        .B2(n5307), .ZN(n5309) );
  INV_X1 U6470 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6280) );
  NAND3_X1 U6471 ( .A1(n6247), .A2(REIP_REG_1__SCAN_IN), .A3(n6280), .ZN(n5308) );
  NAND2_X1 U6472 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  AOI211_X1 U6473 ( .C1(REIP_REG_2__SCAN_IN), .C2(n6281), .A(n5311), .B(n5310), 
        .ZN(n5312) );
  OAI211_X1 U6474 ( .C1(n6465), .C2(n6274), .A(n5313), .B(n5312), .ZN(U2825)
         );
  INV_X1 U6475 ( .A(n5971), .ZN(n5315) );
  NAND2_X1 U6476 ( .A1(n5315), .A2(n5314), .ZN(n6009) );
  NOR3_X1 U6477 ( .A1(n5317), .A2(n5350), .A3(n6496), .ZN(n5318) );
  OAI21_X1 U6478 ( .B1(n5318), .B2(n6499), .A(n6498), .ZN(n5322) );
  NOR2_X1 U6479 ( .A1(n5979), .A2(n5319), .ZN(n6502) );
  OR2_X1 U6480 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5320), .ZN(n5348)
         );
  AOI21_X1 U6481 ( .B1(n5348), .B2(STATE2_REG_3__SCAN_IN), .A(n6487), .ZN(
        n5321) );
  NAND3_X1 U6482 ( .A1(n5322), .A2(n6502), .A3(n5321), .ZN(n5346) );
  NAND2_X1 U6483 ( .A1(n5346), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5327)
         );
  NOR2_X1 U6484 ( .A1(n6498), .A2(n6496), .ZN(n6486) );
  INV_X1 U6485 ( .A(n6489), .ZN(n5323) );
  NOR2_X1 U6486 ( .A1(n5323), .A2(n6487), .ZN(n5324) );
  AOI22_X1 U6487 ( .A1(n6486), .A2(n4712), .B1(n6488), .B2(n5324), .ZN(n5347)
         );
  OAI22_X1 U6488 ( .A1(n6515), .A2(n5348), .B1(n5347), .B2(n6514), .ZN(n5325)
         );
  AOI21_X1 U6489 ( .B1(n6517), .B2(n5350), .A(n5325), .ZN(n5326) );
  OAI211_X1 U6490 ( .C1(n6050), .C2(n6520), .A(n5327), .B(n5326), .ZN(U3134)
         );
  NAND2_X1 U6491 ( .A1(n5346), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5330)
         );
  OAI22_X1 U6492 ( .A1(n6593), .A2(n5348), .B1(n5347), .B2(n6532), .ZN(n5328)
         );
  AOI21_X1 U6493 ( .B1(n6534), .B2(n5350), .A(n5328), .ZN(n5329) );
  OAI211_X1 U6494 ( .C1(n6050), .C2(n6594), .A(n5330), .B(n5329), .ZN(U3137)
         );
  NAND2_X1 U6495 ( .A1(n5346), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5333)
         );
  OAI22_X1 U6496 ( .A1(n6586), .A2(n5348), .B1(n5347), .B2(n6521), .ZN(n5331)
         );
  AOI21_X1 U6497 ( .B1(n6523), .B2(n5350), .A(n5331), .ZN(n5332) );
  OAI211_X1 U6498 ( .C1(n6050), .C2(n6587), .A(n5333), .B(n5332), .ZN(U3135)
         );
  NAND2_X1 U6499 ( .A1(n5346), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5336)
         );
  OAI22_X1 U6500 ( .A1(n6563), .A2(n5348), .B1(n5347), .B2(n6526), .ZN(n5334)
         );
  AOI21_X1 U6501 ( .B1(n6528), .B2(n5350), .A(n5334), .ZN(n5335) );
  OAI211_X1 U6502 ( .C1(n6050), .C2(n6531), .A(n5336), .B(n5335), .ZN(U3136)
         );
  NAND2_X1 U6503 ( .A1(n5346), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5339)
         );
  OAI22_X1 U6504 ( .A1(n6601), .A2(n5348), .B1(n5347), .B2(n6543), .ZN(n5337)
         );
  AOI21_X1 U6505 ( .B1(n6548), .B2(n5350), .A(n5337), .ZN(n5338) );
  OAI211_X1 U6506 ( .C1(n6050), .C2(n6602), .A(n5339), .B(n5338), .ZN(U3139)
         );
  NAND2_X1 U6507 ( .A1(n5346), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5342)
         );
  OAI22_X1 U6508 ( .A1(n6493), .A2(n5348), .B1(n5347), .B2(n6492), .ZN(n5340)
         );
  AOI21_X1 U6509 ( .B1(n6504), .B2(n5350), .A(n5340), .ZN(n5341) );
  OAI211_X1 U6510 ( .C1(n6050), .C2(n6507), .A(n5342), .B(n5341), .ZN(U3132)
         );
  NAND2_X1 U6511 ( .A1(n5346), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5345)
         );
  OAI22_X1 U6512 ( .A1(n6552), .A2(n5348), .B1(n5347), .B2(n6508), .ZN(n5343)
         );
  AOI21_X1 U6513 ( .B1(n6510), .B2(n5350), .A(n5343), .ZN(n5344) );
  OAI211_X1 U6514 ( .C1(n6050), .C2(n6513), .A(n5345), .B(n5344), .ZN(U3133)
         );
  NAND2_X1 U6515 ( .A1(n5346), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5352)
         );
  OAI22_X1 U6516 ( .A1(n6570), .A2(n5348), .B1(n5347), .B2(n6537), .ZN(n5349)
         );
  AOI21_X1 U6517 ( .B1(n6539), .B2(n5350), .A(n5349), .ZN(n5351) );
  OAI211_X1 U6518 ( .C1(n6050), .C2(n6542), .A(n5352), .B(n5351), .ZN(U3138)
         );
  INV_X1 U6519 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6336) );
  OAI222_X1 U6520 ( .A1(n5354), .A2(n6086), .B1(n5739), .B2(n5353), .C1(n5738), 
        .C2(n6336), .ZN(U2883) );
  INV_X1 U6521 ( .A(n5354), .ZN(n5369) );
  OAI22_X1 U6522 ( .A1(n5709), .A2(n6416), .B1(n6307), .B2(n5355), .ZN(n5356)
         );
  AOI21_X1 U6523 ( .B1(n5369), .B2(n6304), .A(n5356), .ZN(n5357) );
  INV_X1 U6524 ( .A(n5357), .ZN(U2851) );
  NAND2_X1 U6525 ( .A1(n5248), .A2(n5359), .ZN(n5360) );
  NAND2_X1 U6526 ( .A1(n5358), .A2(n5360), .ZN(n6243) );
  AOI21_X1 U6527 ( .B1(n5361), .B2(n5251), .A(n3182), .ZN(n6409) );
  AOI22_X1 U6528 ( .A1(n6303), .A2(n6409), .B1(EBX_REG_9__SCAN_IN), .B2(n4391), 
        .ZN(n5362) );
  OAI21_X1 U6529 ( .B1(n6243), .B2(n5704), .A(n5362), .ZN(U2850) );
  OAI21_X1 U6530 ( .B1(n5365), .B2(n5364), .A(n5363), .ZN(n6415) );
  AOI22_X1 U6531 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6476), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5366) );
  OAI21_X1 U6532 ( .B1(n5367), .B2(n6390), .A(n5366), .ZN(n5368) );
  AOI21_X1 U6533 ( .B1(n5369), .B2(n6385), .A(n5368), .ZN(n5370) );
  OAI21_X1 U6534 ( .B1(n6415), .B2(n6364), .A(n5370), .ZN(U2978) );
  NOR2_X1 U6535 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5371), .ZN(n5377)
         );
  INV_X1 U6536 ( .A(n5409), .ZN(n5372) );
  NOR2_X1 U6537 ( .A1(n5406), .A2(n5372), .ZN(n5374) );
  INV_X1 U6538 ( .A(n5380), .ZN(n5373) );
  OAI21_X1 U6539 ( .B1(n5374), .B2(n6499), .A(n5373), .ZN(n5376) );
  NAND2_X1 U6540 ( .A1(n5402), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5383) );
  INV_X1 U6541 ( .A(n5377), .ZN(n5404) );
  NOR2_X1 U6542 ( .A1(n5378), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5379)
         );
  AOI22_X1 U6543 ( .A1(n5380), .A2(n6015), .B1(n6488), .B2(n5379), .ZN(n5403)
         );
  OAI22_X1 U6544 ( .A1(n6493), .A2(n5404), .B1(n5403), .B2(n6492), .ZN(n5381)
         );
  AOI21_X1 U6545 ( .B1(n5406), .B2(n6018), .A(n5381), .ZN(n5382) );
  OAI211_X1 U6546 ( .C1(n5409), .C2(n6021), .A(n5383), .B(n5382), .ZN(U3036)
         );
  NAND2_X1 U6547 ( .A1(n5402), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5386) );
  OAI22_X1 U6548 ( .A1(n6552), .A2(n5404), .B1(n5403), .B2(n6508), .ZN(n5384)
         );
  AOI21_X1 U6549 ( .B1(n5406), .B2(n6554), .A(n5384), .ZN(n5385) );
  OAI211_X1 U6550 ( .C1(n6558), .C2(n5409), .A(n5386), .B(n5385), .ZN(U3037)
         );
  NAND2_X1 U6551 ( .A1(n5402), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5389) );
  OAI22_X1 U6552 ( .A1(n6570), .A2(n5404), .B1(n5403), .B2(n6537), .ZN(n5387)
         );
  AOI21_X1 U6553 ( .B1(n5406), .B2(n6572), .A(n5387), .ZN(n5388) );
  OAI211_X1 U6554 ( .C1(n5409), .C2(n6576), .A(n5389), .B(n5388), .ZN(U3042)
         );
  NAND2_X1 U6555 ( .A1(n5402), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5392) );
  OAI22_X1 U6556 ( .A1(n6563), .A2(n5404), .B1(n5403), .B2(n6526), .ZN(n5390)
         );
  AOI21_X1 U6557 ( .B1(n5406), .B2(n6565), .A(n5390), .ZN(n5391) );
  OAI211_X1 U6558 ( .C1(n5409), .C2(n6569), .A(n5392), .B(n5391), .ZN(U3040)
         );
  NAND2_X1 U6559 ( .A1(n5402), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5395) );
  OAI22_X1 U6560 ( .A1(n6586), .A2(n5404), .B1(n5403), .B2(n6521), .ZN(n5393)
         );
  AOI21_X1 U6561 ( .B1(n5406), .B2(n6560), .A(n5393), .ZN(n5394) );
  OAI211_X1 U6562 ( .C1(n5409), .C2(n6592), .A(n5395), .B(n5394), .ZN(U3039)
         );
  NAND2_X1 U6563 ( .A1(n5402), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5398) );
  OAI22_X1 U6564 ( .A1(n6515), .A2(n5404), .B1(n5403), .B2(n6514), .ZN(n5396)
         );
  AOI21_X1 U6565 ( .B1(n5406), .B2(n6026), .A(n5396), .ZN(n5397) );
  OAI211_X1 U6566 ( .C1(n5409), .C2(n6029), .A(n5398), .B(n5397), .ZN(U3038)
         );
  NAND2_X1 U6567 ( .A1(n5402), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5401) );
  OAI22_X1 U6568 ( .A1(n6601), .A2(n5404), .B1(n5403), .B2(n6543), .ZN(n5399)
         );
  AOI21_X1 U6569 ( .B1(n5406), .B2(n6579), .A(n5399), .ZN(n5400) );
  OAI211_X1 U6570 ( .C1(n5409), .C2(n6611), .A(n5401), .B(n5400), .ZN(U3043)
         );
  NAND2_X1 U6571 ( .A1(n5402), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5408) );
  OAI22_X1 U6572 ( .A1(n6593), .A2(n5404), .B1(n5403), .B2(n6532), .ZN(n5405)
         );
  AOI21_X1 U6573 ( .B1(n5406), .B2(n6037), .A(n5405), .ZN(n5407) );
  OAI211_X1 U6574 ( .C1(n5409), .C2(n6599), .A(n5408), .B(n5407), .ZN(U3041)
         );
  INV_X1 U6575 ( .A(DATAI_9_), .ZN(n6978) );
  INV_X1 U6576 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6334) );
  OAI222_X1 U6577 ( .A1(n6243), .A2(n6086), .B1(n5739), .B2(n6978), .C1(n5738), 
        .C2(n6334), .ZN(U2882) );
  NAND2_X1 U6578 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  XNOR2_X1 U6579 ( .A(n5410), .B(n5413), .ZN(n6411) );
  NAND2_X1 U6580 ( .A1(n6411), .A2(n6386), .ZN(n5417) );
  INV_X1 U6581 ( .A(REIP_REG_9__SCAN_IN), .ZN(n5414) );
  NOR2_X1 U6582 ( .A1(n6454), .A2(n5414), .ZN(n6408) );
  AND2_X1 U6583 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5415)
         );
  AOI211_X1 U6584 ( .C1(n6244), .C2(n6360), .A(n6408), .B(n5415), .ZN(n5416)
         );
  OAI211_X1 U6585 ( .C1(n5839), .C2(n6243), .A(n5417), .B(n5416), .ZN(U2977)
         );
  AOI21_X1 U6586 ( .B1(n5420), .B2(n5358), .A(n5419), .ZN(n5643) );
  INV_X1 U6587 ( .A(n5643), .ZN(n5423) );
  INV_X1 U6588 ( .A(DATAI_10_), .ZN(n6897) );
  INV_X1 U6589 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6332) );
  OAI222_X1 U6590 ( .A1(n5423), .A2(n6086), .B1(n5739), .B2(n6897), .C1(n5738), 
        .C2(n6332), .ZN(U2881) );
  INV_X1 U6591 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5422) );
  XNOR2_X1 U6592 ( .A(n3182), .B(n5421), .ZN(n5645) );
  OAI222_X1 U6593 ( .A1(n5704), .A2(n5423), .B1(n5422), .B2(n6307), .C1(n5709), 
        .C2(n5645), .ZN(U2849) );
  NAND2_X1 U6594 ( .A1(n6354), .A2(n5425), .ZN(n5426) );
  XNOR2_X1 U6595 ( .A(n5424), .B(n5426), .ZN(n6404) );
  INV_X1 U6596 ( .A(n6404), .ZN(n5430) );
  NAND2_X1 U6597 ( .A1(n6476), .A2(REIP_REG_10__SCAN_IN), .ZN(n6399) );
  NAND2_X1 U6598 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5427)
         );
  OAI211_X1 U6599 ( .C1(n6390), .C2(n5644), .A(n6399), .B(n5427), .ZN(n5428)
         );
  AOI21_X1 U6600 ( .B1(n5643), .B2(n6385), .A(n5428), .ZN(n5429) );
  OAI21_X1 U6601 ( .B1(n5430), .B2(n6364), .A(n5429), .ZN(U2976) );
  INV_X1 U6602 ( .A(n5431), .ZN(n5434) );
  INV_X1 U6603 ( .A(n5419), .ZN(n5433) );
  AOI21_X1 U6604 ( .B1(n5434), .B2(n5433), .A(n5432), .ZN(n6361) );
  INV_X1 U6605 ( .A(n6361), .ZN(n5435) );
  INV_X1 U6606 ( .A(DATAI_11_), .ZN(n6757) );
  INV_X1 U6607 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6330) );
  OAI222_X1 U6608 ( .A1(n5435), .A2(n6086), .B1(n5739), .B2(n6757), .C1(n5738), 
        .C2(n6330), .ZN(U2880) );
  XOR2_X1 U6609 ( .A(n5436), .B(n5432), .Z(n5454) );
  INV_X1 U6610 ( .A(n5440), .ZN(n5437) );
  NOR2_X1 U6611 ( .A1(n6272), .A2(n5437), .ZN(n6221) );
  INV_X1 U6612 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5450) );
  OAI21_X1 U6613 ( .B1(n5439), .B2(n6229), .A(n5438), .ZN(n5474) );
  OAI22_X1 U6614 ( .A1(n6279), .A2(n5452), .B1(n6274), .B2(n5474), .ZN(n5444)
         );
  INV_X1 U6615 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5442) );
  OAI21_X1 U6616 ( .B1(n6272), .B2(n5440), .A(n5621), .ZN(n6228) );
  AOI22_X1 U6617 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6288), .B1(
        REIP_REG_12__SCAN_IN), .B2(n6228), .ZN(n5441) );
  OAI211_X1 U6618 ( .C1(n6258), .C2(n5442), .A(n5441), .B(n6257), .ZN(n5443)
         );
  AOI211_X1 U6619 ( .C1(n6221), .C2(n5450), .A(n5444), .B(n5443), .ZN(n5445)
         );
  OAI21_X1 U6620 ( .B1(n5473), .B2(n6212), .A(n5445), .ZN(U2815) );
  INV_X1 U6621 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6328) );
  OAI222_X1 U6622 ( .A1(n6086), .A2(n5473), .B1(n5738), .B2(n6328), .C1(n5446), 
        .C2(n5739), .ZN(U2879) );
  NOR2_X1 U6623 ( .A1(n5448), .A2(n3198), .ZN(n5449) );
  XNOR2_X1 U6624 ( .A(n5447), .B(n5449), .ZN(n5472) );
  NOR2_X1 U6625 ( .A1(n6454), .A2(n5450), .ZN(n5468) );
  AOI21_X1 U6626 ( .B1(n6380), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n5468), 
        .ZN(n5451) );
  OAI21_X1 U6627 ( .B1(n5452), .B2(n6390), .A(n5451), .ZN(n5453) );
  AOI21_X1 U6628 ( .B1(n5454), .B2(n6385), .A(n5453), .ZN(n5455) );
  OAI21_X1 U6629 ( .B1(n5472), .B2(n6364), .A(n5455), .ZN(U2974) );
  NOR2_X1 U6630 ( .A1(n6433), .A2(n5456), .ZN(n5465) );
  INV_X1 U6631 ( .A(n5457), .ZN(n6397) );
  OAI21_X1 U6632 ( .B1(n5459), .B2(n5458), .A(n5462), .ZN(n5460) );
  AOI21_X1 U6633 ( .B1(n6433), .B2(n6397), .A(n5460), .ZN(n6431) );
  AOI22_X1 U6634 ( .A1(n5462), .A2(n6403), .B1(n5461), .B2(n6431), .ZN(n6393)
         );
  INV_X1 U6635 ( .A(n6393), .ZN(n5463) );
  OAI221_X1 U6636 ( .B1(n6146), .B2(n5465), .C1(n6146), .C2(n5464), .A(n5463), 
        .ZN(n5470) );
  INV_X1 U6637 ( .A(n6392), .ZN(n6163) );
  OAI21_X1 U6638 ( .B1(n6163), .B2(n3686), .A(n5466), .ZN(n5469) );
  NOR2_X1 U6639 ( .A1(n6448), .A2(n5474), .ZN(n5467) );
  AOI211_X1 U6640 ( .C1(n5470), .C2(n5469), .A(n5468), .B(n5467), .ZN(n5471)
         );
  OAI21_X1 U6641 ( .B1(n5472), .B2(n6455), .A(n5471), .ZN(U3006) );
  OAI222_X1 U6642 ( .A1(n5709), .A2(n5474), .B1(n6307), .B2(n4327), .C1(n5704), 
        .C2(n5473), .ZN(U2847) );
  NOR2_X1 U6643 ( .A1(n6454), .A2(n6861), .ZN(n5861) );
  NOR2_X1 U6644 ( .A1(n6390), .A2(n5486), .ZN(n5475) );
  AOI211_X1 U6645 ( .C1(PHYADDRPOINTER_REG_30__SCAN_IN), .C2(n6380), .A(n5861), 
        .B(n5475), .ZN(n5480) );
  XNOR2_X1 U6646 ( .A(n5478), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5856)
         );
  NAND2_X1 U6647 ( .A1(n5856), .A2(n6386), .ZN(n5479) );
  OAI211_X1 U6648 ( .C1(n5492), .C2(n5839), .A(n5480), .B(n5479), .ZN(U2956)
         );
  AOI22_X1 U6649 ( .A1(n6314), .A2(DATAI_30_), .B1(n6317), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6650 ( .A1(n6318), .A2(DATAI_14_), .ZN(n5481) );
  OAI211_X1 U6651 ( .C1(n5492), .C2(n6086), .A(n5482), .B(n5481), .ZN(U2861)
         );
  NOR2_X1 U6652 ( .A1(n5483), .A2(n6861), .ZN(n5490) );
  NAND2_X1 U6653 ( .A1(n6861), .A2(REIP_REG_29__SCAN_IN), .ZN(n5484) );
  NOR2_X1 U6654 ( .A1(n5514), .A2(n5484), .ZN(n5489) );
  AOI22_X1 U6655 ( .A1(EBX_REG_30__SCAN_IN), .A2(n6288), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6285), .ZN(n5485) );
  OAI21_X1 U6656 ( .B1(n5486), .B2(n6279), .A(n5485), .ZN(n5488) );
  NOR2_X1 U6657 ( .A1(n5857), .A2(n6274), .ZN(n5487) );
  NOR4_X1 U6658 ( .A1(n5490), .A2(n5489), .A3(n5488), .A4(n5487), .ZN(n5491)
         );
  OAI21_X1 U6659 ( .B1(n5492), .B2(n6212), .A(n5491), .ZN(U2797) );
  AOI22_X1 U6660 ( .A1(n5495), .A2(n5494), .B1(n5493), .B2(n3169), .ZN(n6612)
         );
  AOI22_X1 U6661 ( .A1(n5496), .A2(n3169), .B1(n4903), .B2(
        STATE2_REG_1__SCAN_IN), .ZN(n5497) );
  OAI21_X1 U6662 ( .B1(n6612), .B2(n5965), .A(n5497), .ZN(n5500) );
  NOR2_X1 U6663 ( .A1(n5498), .A2(n3169), .ZN(n6614) );
  AOI22_X1 U6664 ( .A1(n6170), .A2(n5500), .B1(n5499), .B2(n6614), .ZN(n5501)
         );
  OAI21_X1 U6665 ( .B1(n3169), .B2(n6170), .A(n5501), .ZN(U3461) );
  OAI22_X1 U6666 ( .A1(n5851), .A2(n5709), .B1(n6307), .B2(n5502), .ZN(U2828)
         );
  INV_X1 U6667 ( .A(n5504), .ZN(n5510) );
  INV_X1 U6668 ( .A(n4383), .ZN(n5508) );
  AOI21_X1 U6669 ( .B1(n5506), .B2(n4324), .A(n5505), .ZN(n5507) );
  NAND2_X1 U6670 ( .A1(n5508), .A2(n5507), .ZN(n5509) );
  NAND2_X1 U6671 ( .A1(n5510), .A2(n5509), .ZN(n5867) );
  AOI22_X1 U6672 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6285), .B1(n6294), 
        .B2(n5511), .ZN(n5513) );
  NAND2_X1 U6673 ( .A1(n6288), .A2(EBX_REG_29__SCAN_IN), .ZN(n5512) );
  OAI211_X1 U6674 ( .C1(n5867), .C2(n6274), .A(n5513), .B(n5512), .ZN(n5516)
         );
  NOR2_X1 U6675 ( .A1(n5514), .A2(REIP_REG_29__SCAN_IN), .ZN(n5515) );
  AOI211_X1 U6676 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5528), .A(n5516), .B(n5515), .ZN(n5517) );
  OAI21_X1 U6677 ( .B1(n5503), .B2(n6212), .A(n5517), .ZN(U2798) );
  AOI21_X1 U6678 ( .B1(n5520), .B2(n5518), .A(n5519), .ZN(n5748) );
  INV_X1 U6679 ( .A(n5748), .ZN(n5719) );
  INV_X1 U6680 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U6681 ( .A1(n5521), .A2(n6871), .ZN(n5526) );
  AOI21_X1 U6682 ( .B1(n5522), .B2(n5535), .A(n4383), .ZN(n5876) );
  INV_X1 U6683 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5523) );
  OAI22_X1 U6684 ( .A1(n5523), .A2(n6258), .B1(n6279), .B2(n5746), .ZN(n5524)
         );
  AOI21_X1 U6685 ( .B1(n5876), .B2(n6286), .A(n5524), .ZN(n5525) );
  OAI211_X1 U6686 ( .C1(n4377), .C2(n6270), .A(n5526), .B(n5525), .ZN(n5527)
         );
  AOI21_X1 U6687 ( .B1(n5528), .B2(REIP_REG_28__SCAN_IN), .A(n5527), .ZN(n5529) );
  OAI21_X1 U6688 ( .B1(n5719), .B2(n6212), .A(n5529), .ZN(U2799) );
  OAI21_X1 U6689 ( .B1(n5530), .B2(n5531), .A(n5518), .ZN(n5758) );
  INV_X1 U6690 ( .A(REIP_REG_27__SCAN_IN), .ZN(n7087) );
  AOI22_X1 U6691 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6288), .B1(n5752), .B2(n6294), .ZN(n5532) );
  OAI21_X1 U6692 ( .B1(n5750), .B2(n6258), .A(n5532), .ZN(n5537) );
  NAND2_X1 U6693 ( .A1(n5665), .A2(n5533), .ZN(n5534) );
  NAND2_X1 U6694 ( .A1(n5535), .A2(n5534), .ZN(n5886) );
  NOR2_X1 U6695 ( .A1(n5886), .A2(n6274), .ZN(n5536) );
  NOR2_X1 U6696 ( .A1(n5537), .A2(n5536), .ZN(n5541) );
  INV_X1 U6697 ( .A(n6051), .ZN(n5539) );
  NAND3_X1 U6698 ( .A1(n5539), .A2(n7087), .A3(n5538), .ZN(n5540) );
  OAI211_X1 U6699 ( .C1(n6053), .C2(n7087), .A(n5541), .B(n5540), .ZN(n5542)
         );
  INV_X1 U6700 ( .A(n5542), .ZN(n5543) );
  OAI21_X1 U6701 ( .B1(n5758), .B2(n6212), .A(n5543), .ZN(U2800) );
  OAI21_X1 U6702 ( .B1(n5546), .B2(n5545), .A(n5670), .ZN(n5781) );
  INV_X1 U6703 ( .A(n5784), .ZN(n5548) );
  NOR2_X1 U6704 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6051), .ZN(n6064) );
  AOI21_X1 U6705 ( .B1(n6285), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6064), 
        .ZN(n5547) );
  OAI21_X1 U6706 ( .B1(n6279), .B2(n5548), .A(n5547), .ZN(n5554) );
  INV_X1 U6707 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5552) );
  INV_X1 U6708 ( .A(n5549), .ZN(n5550) );
  OAI21_X1 U6709 ( .B1(n4464), .B2(n5551), .A(n5550), .ZN(n5906) );
  OAI22_X1 U6710 ( .A1(n5552), .A2(n6270), .B1(n6274), .B2(n5906), .ZN(n5553)
         );
  AOI211_X1 U6711 ( .C1(n6075), .C2(REIP_REG_24__SCAN_IN), .A(n5554), .B(n5553), .ZN(n5555) );
  OAI21_X1 U6712 ( .B1(n5781), .B2(n6212), .A(n5555), .ZN(U2803) );
  AND2_X1 U6713 ( .A1(n5557), .A2(n5556), .ZN(n5558) );
  NOR2_X1 U6714 ( .A1(n3179), .A2(n5558), .ZN(n6087) );
  INV_X1 U6715 ( .A(n6087), .ZN(n5677) );
  AOI21_X1 U6716 ( .B1(n5560), .B2(n5574), .A(n4360), .ZN(n5914) );
  INV_X1 U6717 ( .A(n5914), .ZN(n5561) );
  OAI22_X1 U6718 ( .A1(n6279), .A2(n5790), .B1(n6274), .B2(n5561), .ZN(n5564)
         );
  NAND2_X1 U6719 ( .A1(n5562), .A2(n6868), .ZN(n5572) );
  AOI21_X1 U6720 ( .B1(n6084), .B2(n5572), .A(n7068), .ZN(n5563) );
  AOI211_X1 U6721 ( .C1(EBX_REG_22__SCAN_IN), .C2(n6288), .A(n5564), .B(n5563), 
        .ZN(n5569) );
  INV_X1 U6722 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5565) );
  OAI22_X1 U6723 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5566), .B1(n5565), .B2(
        n6258), .ZN(n5567) );
  INV_X1 U6724 ( .A(n5567), .ZN(n5568) );
  OAI211_X1 U6725 ( .C1(n5677), .C2(n6212), .A(n5569), .B(n5568), .ZN(U2805)
         );
  XOR2_X1 U6726 ( .A(n5571), .B(n5570), .Z(n6090) );
  INV_X1 U6727 ( .A(n6090), .ZN(n5679) );
  INV_X1 U6728 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5796) );
  OAI22_X1 U6729 ( .A1(n5796), .A2(n6258), .B1(n6868), .B2(n6084), .ZN(n5582)
         );
  INV_X1 U6730 ( .A(n5572), .ZN(n5581) );
  INV_X1 U6731 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5579) );
  INV_X1 U6732 ( .A(n5573), .ZN(n5577) );
  INV_X1 U6733 ( .A(n5574), .ZN(n5575) );
  AOI21_X1 U6734 ( .B1(n5577), .B2(n5576), .A(n5575), .ZN(n5923) );
  AOI22_X1 U6735 ( .A1(n6286), .A2(n5923), .B1(n6294), .B2(n5798), .ZN(n5578)
         );
  OAI21_X1 U6736 ( .B1(n6270), .B2(n5579), .A(n5578), .ZN(n5580) );
  NOR3_X1 U6737 ( .A1(n5582), .A2(n5581), .A3(n5580), .ZN(n5583) );
  OAI21_X1 U6738 ( .B1(n5679), .B2(n6212), .A(n5583), .ZN(U2806) );
  AOI21_X1 U6739 ( .B1(n5587), .B2(n5584), .A(n5586), .ZN(n5814) );
  INV_X1 U6740 ( .A(n5814), .ZN(n5732) );
  INV_X1 U6741 ( .A(n5588), .ZN(n5812) );
  INV_X1 U6742 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U6743 ( .A1(n5590), .A2(n4295), .ZN(n5591) );
  OAI21_X1 U6744 ( .B1(n5681), .B2(n4295), .A(n5591), .ZN(n5689) );
  INV_X1 U6745 ( .A(n5610), .ZN(n5690) );
  NAND2_X1 U6746 ( .A1(n5689), .A2(n5690), .ZN(n5692) );
  XOR2_X1 U6747 ( .A(n5592), .B(n5692), .Z(n6119) );
  INV_X1 U6748 ( .A(n6119), .ZN(n5593) );
  OAI22_X1 U6749 ( .A1(n6279), .A2(n5812), .B1(n6274), .B2(n5593), .ZN(n5601)
         );
  INV_X1 U6750 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6899) );
  NOR2_X1 U6751 ( .A1(n5595), .A2(n6899), .ZN(n6079) );
  INV_X1 U6752 ( .A(n6079), .ZN(n5597) );
  AND2_X1 U6753 ( .A1(n6263), .A2(n5594), .ZN(n6195) );
  NOR2_X1 U6754 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5595), .ZN(n6196) );
  NOR2_X1 U6755 ( .A1(n6195), .A2(n6196), .ZN(n5596) );
  MUX2_X1 U6756 ( .A(n5597), .B(n5596), .S(REIP_REG_19__SCAN_IN), .Z(n5598) );
  OAI211_X1 U6757 ( .C1(n6258), .C2(n5599), .A(n5598), .B(n6257), .ZN(n5600)
         );
  AOI211_X1 U6758 ( .C1(n6288), .C2(EBX_REG_19__SCAN_IN), .A(n5601), .B(n5600), 
        .ZN(n5602) );
  OAI21_X1 U6759 ( .B1(n5732), .B2(n6212), .A(n5602), .ZN(U2808) );
  XOR2_X1 U6760 ( .A(n5604), .B(n5603), .Z(n6311) );
  INV_X1 U6761 ( .A(n6311), .ZN(n5700) );
  OAI21_X1 U6762 ( .B1(n6272), .B2(n5605), .A(n6755), .ZN(n5614) );
  INV_X1 U6763 ( .A(EBX_REG_17__SCAN_IN), .ZN(n5607) );
  OAI22_X1 U6764 ( .A1(n5607), .A2(n6270), .B1(n5606), .B2(n6258), .ZN(n5613)
         );
  NAND2_X1 U6765 ( .A1(n5608), .A2(n5619), .ZN(n5609) );
  NAND2_X1 U6766 ( .A1(n5610), .A2(n5609), .ZN(n5698) );
  INV_X1 U6767 ( .A(n6257), .ZN(n6268) );
  AOI21_X1 U6768 ( .B1(n6294), .B2(n6103), .A(n6268), .ZN(n5611) );
  OAI21_X1 U6769 ( .B1(n6274), .B2(n5698), .A(n5611), .ZN(n5612) );
  AOI211_X1 U6770 ( .C1(n6195), .C2(n5614), .A(n5613), .B(n5612), .ZN(n5615)
         );
  OAI21_X1 U6771 ( .B1(n5700), .B2(n6212), .A(n5615), .ZN(U2810) );
  OR2_X1 U6772 ( .A1(n5616), .A2(n5617), .ZN(n5618) );
  AND2_X1 U6773 ( .A1(n5603), .A2(n5618), .ZN(n6316) );
  INV_X1 U6774 ( .A(n6316), .ZN(n5701) );
  OAI21_X1 U6775 ( .B1(n5620), .B2(n5636), .A(n5619), .ZN(n5954) );
  INV_X1 U6776 ( .A(n5621), .ZN(n6264) );
  OAI21_X1 U6777 ( .B1(n6264), .B2(n5622), .A(n6263), .ZN(n6217) );
  OR3_X1 U6778 ( .A1(n6272), .A2(REIP_REG_15__SCAN_IN), .A3(n5622), .ZN(n5634)
         );
  INV_X1 U6779 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6985) );
  AOI21_X1 U6780 ( .B1(n6217), .B2(n5634), .A(n6985), .ZN(n5623) );
  AOI21_X1 U6781 ( .B1(n6294), .B2(n5819), .A(n5623), .ZN(n5624) );
  OAI21_X1 U6782 ( .B1(n6274), .B2(n5954), .A(n5624), .ZN(n5629) );
  NAND3_X1 U6783 ( .A1(n6247), .A2(n6985), .A3(n5625), .ZN(n5626) );
  OAI211_X1 U6784 ( .C1(n6258), .C2(n5627), .A(n6257), .B(n5626), .ZN(n5628)
         );
  AOI211_X1 U6785 ( .C1(EBX_REG_16__SCAN_IN), .C2(n6288), .A(n5629), .B(n5628), 
        .ZN(n5630) );
  OAI21_X1 U6786 ( .B1(n5701), .B2(n6212), .A(n5630), .ZN(U2811) );
  AOI21_X1 U6787 ( .B1(n5632), .B2(n5631), .A(n5616), .ZN(n5829) );
  INV_X1 U6788 ( .A(n5829), .ZN(n5733) );
  OAI22_X1 U6789 ( .A1(n5633), .A2(n6270), .B1(n6691), .B2(n6217), .ZN(n5641)
         );
  OAI211_X1 U6790 ( .C1(n6258), .C2(n5635), .A(n6257), .B(n5634), .ZN(n5640)
         );
  AOI21_X1 U6791 ( .B1(n5637), .B2(n5707), .A(n5636), .ZN(n6136) );
  INV_X1 U6792 ( .A(n6136), .ZN(n5638) );
  OAI22_X1 U6793 ( .A1(n6279), .A2(n5827), .B1(n6274), .B2(n5638), .ZN(n5639)
         );
  NOR3_X1 U6794 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n5642) );
  OAI21_X1 U6795 ( .B1(n5733), .B2(n6212), .A(n5642), .ZN(U2812) );
  NAND2_X1 U6796 ( .A1(n5643), .A2(n4408), .ZN(n5655) );
  INV_X1 U6797 ( .A(n5644), .ZN(n5649) );
  INV_X1 U6798 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5647) );
  INV_X1 U6799 ( .A(n5645), .ZN(n6401) );
  AOI22_X1 U6800 ( .A1(n6286), .A2(n6401), .B1(n6288), .B2(EBX_REG_10__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U6801 ( .C1(n6258), .C2(n5647), .A(n5646), .B(n6257), .ZN(n5648)
         );
  AOI21_X1 U6802 ( .B1(n6294), .B2(n5649), .A(n5648), .ZN(n5654) );
  NOR2_X1 U6803 ( .A1(n6272), .A2(REIP_REG_9__SCAN_IN), .ZN(n5650) );
  OAI21_X1 U6804 ( .B1(n6242), .B2(n5650), .A(REIP_REG_10__SCAN_IN), .ZN(n5653) );
  NOR2_X1 U6805 ( .A1(n6272), .A2(n5651), .ZN(n6227) );
  NAND2_X1 U6806 ( .A1(n6227), .A2(n6688), .ZN(n5652) );
  NAND4_X1 U6807 ( .A1(n5655), .A2(n5654), .A3(n5653), .A4(n5652), .ZN(U2817)
         );
  INV_X1 U6808 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5656) );
  OAI222_X1 U6809 ( .A1(n5704), .A2(n5503), .B1(n5656), .B2(n6307), .C1(n5867), 
        .C2(n5709), .ZN(U2830) );
  INV_X1 U6810 ( .A(n5876), .ZN(n5657) );
  OAI222_X1 U6811 ( .A1(n5704), .A2(n5719), .B1(n6307), .B2(n4377), .C1(n5657), 
        .C2(n5709), .ZN(U2831) );
  INV_X1 U6812 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5658) );
  OAI222_X1 U6813 ( .A1(n5704), .A2(n5758), .B1(n5658), .B2(n6307), .C1(n5886), 
        .C2(n5709), .ZN(U2832) );
  AND2_X1 U6814 ( .A1(n5659), .A2(n5660), .ZN(n5661) );
  OR2_X1 U6815 ( .A1(n5661), .A2(n5530), .ZN(n5761) );
  NAND2_X1 U6816 ( .A1(n5662), .A2(n5663), .ZN(n5664) );
  NAND2_X1 U6817 ( .A1(n5665), .A2(n5664), .ZN(n6052) );
  OAI22_X1 U6818 ( .A1(n6052), .A2(n5709), .B1(n5666), .B2(n6307), .ZN(n5667)
         );
  INV_X1 U6819 ( .A(n5667), .ZN(n5668) );
  OAI21_X1 U6820 ( .B1(n5761), .B2(n5704), .A(n5668), .ZN(U2833) );
  NAND2_X1 U6821 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  AND2_X1 U6822 ( .A1(n5659), .A2(n5671), .ZN(n6063) );
  INV_X1 U6823 ( .A(n6063), .ZN(n5771) );
  INV_X1 U6824 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5674) );
  OR2_X1 U6825 ( .A1(n5549), .A2(n5672), .ZN(n5673) );
  NAND2_X1 U6826 ( .A1(n5662), .A2(n5673), .ZN(n6111) );
  OAI222_X1 U6827 ( .A1(n5771), .A2(n5704), .B1(n5674), .B2(n6307), .C1(n5709), 
        .C2(n6111), .ZN(U2834) );
  OAI222_X1 U6828 ( .A1(n5704), .A2(n5781), .B1(n6307), .B2(n5552), .C1(n5906), 
        .C2(n5709), .ZN(U2835) );
  AOI22_X1 U6829 ( .A1(n6303), .A2(n6070), .B1(EBX_REG_23__SCAN_IN), .B2(n4391), .ZN(n5675) );
  OAI21_X1 U6830 ( .B1(n6072), .B2(n5704), .A(n5675), .ZN(U2836) );
  AOI22_X1 U6831 ( .A1(n6303), .A2(n5914), .B1(EBX_REG_22__SCAN_IN), .B2(n4391), .ZN(n5676) );
  OAI21_X1 U6832 ( .B1(n5677), .B2(n5704), .A(n5676), .ZN(U2837) );
  AOI22_X1 U6833 ( .A1(n6303), .A2(n5923), .B1(EBX_REG_21__SCAN_IN), .B2(n4391), .ZN(n5678) );
  OAI21_X1 U6834 ( .B1(n5679), .B2(n5704), .A(n5678), .ZN(U2838) );
  OAI21_X1 U6835 ( .B1(n5586), .B2(n5680), .A(n5570), .ZN(n5803) );
  INV_X1 U6836 ( .A(n5681), .ZN(n5682) );
  NAND2_X1 U6837 ( .A1(n3196), .A2(n5682), .ZN(n5683) );
  OAI21_X1 U6838 ( .B1(n3196), .B2(n4324), .A(n5683), .ZN(n5686) );
  INV_X1 U6839 ( .A(n5684), .ZN(n5685) );
  XNOR2_X1 U6840 ( .A(n5686), .B(n5685), .ZN(n6081) );
  AOI22_X1 U6841 ( .A1(n6303), .A2(n6081), .B1(EBX_REG_20__SCAN_IN), .B2(n4391), .ZN(n5687) );
  OAI21_X1 U6842 ( .B1(n5803), .B2(n5704), .A(n5687), .ZN(U2839) );
  AOI22_X1 U6843 ( .A1(n6303), .A2(n6119), .B1(EBX_REG_19__SCAN_IN), .B2(n4391), .ZN(n5688) );
  OAI21_X1 U6844 ( .B1(n5732), .B2(n5704), .A(n5688), .ZN(U2840) );
  OR2_X1 U6845 ( .A1(n5690), .A2(n5689), .ZN(n5691) );
  NAND2_X1 U6846 ( .A1(n5692), .A2(n5691), .ZN(n6199) );
  NAND2_X1 U6847 ( .A1(n5693), .A2(n5694), .ZN(n5695) );
  AND2_X1 U6848 ( .A1(n5584), .A2(n5695), .ZN(n6308) );
  INV_X1 U6849 ( .A(n6308), .ZN(n5696) );
  OAI222_X1 U6850 ( .A1(n6199), .A2(n5709), .B1(n5697), .B2(n6307), .C1(n5696), 
        .C2(n5704), .ZN(U2841) );
  INV_X1 U6851 ( .A(n5698), .ZN(n6130) );
  AOI22_X1 U6852 ( .A1(n6303), .A2(n6130), .B1(EBX_REG_17__SCAN_IN), .B2(n4391), .ZN(n5699) );
  OAI21_X1 U6853 ( .B1(n5700), .B2(n5704), .A(n5699), .ZN(U2842) );
  OAI222_X1 U6854 ( .A1(n5954), .A2(n5709), .B1(n5702), .B2(n6307), .C1(n5701), 
        .C2(n5704), .ZN(U2843) );
  AOI22_X1 U6855 ( .A1(n6303), .A2(n6136), .B1(n4391), .B2(EBX_REG_15__SCAN_IN), .ZN(n5703) );
  OAI21_X1 U6856 ( .B1(n5733), .B2(n5704), .A(n5703), .ZN(U2844) );
  OAI21_X1 U6857 ( .B1(n5705), .B2(n5706), .A(n5631), .ZN(n6213) );
  OAI21_X1 U6858 ( .B1(n5708), .B2(n6155), .A(n5707), .ZN(n6208) );
  OAI222_X1 U6859 ( .A1(n6213), .A2(n5704), .B1(n5710), .B2(n6307), .C1(n6208), 
        .C2(n5709), .ZN(U2845) );
  AND2_X1 U6860 ( .A1(n5738), .A2(n4390), .ZN(n5711) );
  NAND2_X1 U6861 ( .A1(n5712), .A2(n5711), .ZN(n5714) );
  AOI22_X1 U6862 ( .A1(n6314), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6317), .ZN(n5713) );
  NAND2_X1 U6863 ( .A1(n5714), .A2(n5713), .ZN(U2860) );
  AOI22_X1 U6864 ( .A1(n6314), .A2(DATAI_29_), .B1(n6317), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U6865 ( .A1(n6318), .A2(DATAI_13_), .ZN(n5715) );
  OAI211_X1 U6866 ( .C1(n5503), .C2(n6086), .A(n5716), .B(n5715), .ZN(U2862)
         );
  AOI22_X1 U6867 ( .A1(n6314), .A2(DATAI_28_), .B1(n6317), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U6868 ( .A1(n6318), .A2(DATAI_12_), .ZN(n5717) );
  OAI211_X1 U6869 ( .C1(n5719), .C2(n6086), .A(n5718), .B(n5717), .ZN(U2863)
         );
  AOI22_X1 U6870 ( .A1(n6314), .A2(DATAI_27_), .B1(n6317), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5721) );
  NAND2_X1 U6871 ( .A1(n6318), .A2(DATAI_11_), .ZN(n5720) );
  OAI211_X1 U6872 ( .C1(n5758), .C2(n6086), .A(n5721), .B(n5720), .ZN(U2864)
         );
  AOI22_X1 U6873 ( .A1(n6318), .A2(DATAI_10_), .B1(n6317), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6874 ( .A1(n6314), .A2(DATAI_26_), .ZN(n5722) );
  OAI211_X1 U6875 ( .C1(n5761), .C2(n6086), .A(n5723), .B(n5722), .ZN(U2865)
         );
  AOI22_X1 U6876 ( .A1(n6318), .A2(DATAI_9_), .B1(n6317), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6877 ( .A1(n6314), .A2(DATAI_25_), .ZN(n5724) );
  OAI211_X1 U6878 ( .C1(n5771), .C2(n6086), .A(n5725), .B(n5724), .ZN(U2866)
         );
  AOI22_X1 U6879 ( .A1(n6314), .A2(DATAI_24_), .B1(n6317), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U6880 ( .A1(n6318), .A2(DATAI_8_), .ZN(n5726) );
  OAI211_X1 U6881 ( .C1(n5781), .C2(n6086), .A(n5727), .B(n5726), .ZN(U2867)
         );
  AOI22_X1 U6882 ( .A1(n6318), .A2(DATAI_7_), .B1(n6317), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5729) );
  NAND2_X1 U6883 ( .A1(n6314), .A2(DATAI_23_), .ZN(n5728) );
  OAI211_X1 U6884 ( .C1(n6072), .C2(n6086), .A(n5729), .B(n5728), .ZN(U2868)
         );
  AOI22_X1 U6885 ( .A1(n6314), .A2(DATAI_19_), .B1(n6317), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5731) );
  NAND2_X1 U6886 ( .A1(n6318), .A2(DATAI_3_), .ZN(n5730) );
  OAI211_X1 U6887 ( .C1(n5732), .C2(n6086), .A(n5731), .B(n5730), .ZN(U2872)
         );
  OAI222_X1 U6888 ( .A1(n5733), .A2(n6086), .B1(n6829), .B2(n5739), .C1(n5738), 
        .C2(n4535), .ZN(U2876) );
  INV_X1 U6889 ( .A(DATAI_14_), .ZN(n6972) );
  INV_X1 U6890 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U6891 ( .A1(n6213), .A2(n6086), .B1(n5739), .B2(n6972), .C1(n5738), 
        .C2(n6324), .ZN(U2877) );
  NAND2_X1 U6892 ( .A1(n5735), .A2(n5736), .ZN(n5737) );
  INV_X1 U6893 ( .A(n6300), .ZN(n5740) );
  INV_X1 U6894 ( .A(DATAI_13_), .ZN(n6841) );
  INV_X1 U6895 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6326) );
  OAI222_X1 U6896 ( .A1(n5740), .A2(n6086), .B1(n5739), .B2(n6841), .C1(n5738), 
        .C2(n6326), .ZN(U2878) );
  NAND3_X1 U6897 ( .A1(n3706), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n6356), .ZN(n5743) );
  NOR2_X1 U6898 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5895) );
  NAND3_X1 U6899 ( .A1(n5742), .A2(n5944), .A3(n5895), .ZN(n5753) );
  AOI22_X1 U6900 ( .A1(n5743), .A2(n5753), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5759), .ZN(n5744) );
  XNOR2_X1 U6901 ( .A(n5744), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5882)
         );
  NAND2_X1 U6902 ( .A1(n6476), .A2(REIP_REG_28__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6903 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5745)
         );
  OAI211_X1 U6904 ( .C1(n6390), .C2(n5746), .A(n5878), .B(n5745), .ZN(n5747)
         );
  AOI21_X1 U6905 ( .B1(n5748), .B2(n6385), .A(n5747), .ZN(n5749) );
  OAI21_X1 U6906 ( .B1(n6364), .B2(n5882), .A(n5749), .ZN(U2958) );
  NOR2_X1 U6907 ( .A1(n6454), .A2(n7087), .ZN(n5887) );
  NOR2_X1 U6908 ( .A1(n5836), .A2(n5750), .ZN(n5751) );
  AOI211_X1 U6909 ( .C1(n6360), .C2(n5752), .A(n5887), .B(n5751), .ZN(n5757)
         );
  NAND2_X1 U6910 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  XNOR2_X1 U6911 ( .A(n5755), .B(n5892), .ZN(n5884) );
  NAND2_X1 U6912 ( .A1(n5884), .A2(n6386), .ZN(n5756) );
  OAI211_X1 U6913 ( .C1(n5758), .C2(n5839), .A(n5757), .B(n5756), .ZN(U2959)
         );
  XNOR2_X1 U6914 ( .A(n6356), .B(n5759), .ZN(n5760) );
  XNOR2_X1 U6915 ( .A(n5741), .B(n5760), .ZN(n5901) );
  INV_X1 U6916 ( .A(n5761), .ZN(n6056) );
  NAND2_X1 U6917 ( .A1(n6476), .A2(REIP_REG_26__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U6918 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5762)
         );
  OAI211_X1 U6919 ( .C1(n6390), .C2(n6059), .A(n5894), .B(n5762), .ZN(n5763)
         );
  AOI21_X1 U6920 ( .B1(n6056), .B2(n6385), .A(n5763), .ZN(n5764) );
  OAI21_X1 U6921 ( .B1(n6364), .B2(n5901), .A(n5764), .ZN(U2960) );
  INV_X1 U6922 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5765) );
  OAI22_X1 U6923 ( .A1(n5836), .A2(n5766), .B1(n6454), .B2(n5765), .ZN(n5767)
         );
  AOI21_X1 U6924 ( .B1(n6360), .B2(n6061), .A(n5767), .ZN(n5770) );
  OAI21_X1 U6925 ( .B1(n5742), .B2(n5768), .A(n4229), .ZN(n6113) );
  NAND2_X1 U6926 ( .A1(n6113), .A2(n6386), .ZN(n5769) );
  OAI211_X1 U6927 ( .C1(n5771), .C2(n5839), .A(n5770), .B(n5769), .ZN(U2961)
         );
  INV_X1 U6928 ( .A(n5772), .ZN(n5773) );
  NAND2_X1 U6929 ( .A1(n5773), .A2(n4495), .ZN(n5778) );
  AND2_X1 U6930 ( .A1(n5774), .A2(n3278), .ZN(n5776) );
  NAND2_X1 U6931 ( .A1(n5787), .A2(n5776), .ZN(n5777) );
  NAND2_X1 U6932 ( .A1(n5778), .A2(n5777), .ZN(n5779) );
  XNOR2_X1 U6933 ( .A(n5779), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5911)
         );
  NAND2_X1 U6934 ( .A1(n6476), .A2(REIP_REG_24__SCAN_IN), .ZN(n5905) );
  OAI21_X1 U6935 ( .B1(n5836), .B2(n5780), .A(n5905), .ZN(n5783) );
  NOR2_X1 U6936 ( .A1(n5781), .A2(n5839), .ZN(n5782) );
  AOI211_X1 U6937 ( .C1(n6360), .C2(n5784), .A(n5783), .B(n5782), .ZN(n5785)
         );
  OAI21_X1 U6938 ( .B1(n5911), .B2(n6364), .A(n5785), .ZN(U2962) );
  AOI21_X1 U6939 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n6356), .A(n5786), 
        .ZN(n5788) );
  XOR2_X1 U6940 ( .A(n5788), .B(n5787), .Z(n5920) );
  NOR2_X1 U6941 ( .A1(n6454), .A2(n7068), .ZN(n5913) );
  AOI21_X1 U6942 ( .B1(n6380), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5913), 
        .ZN(n5789) );
  OAI21_X1 U6943 ( .B1(n5790), .B2(n6390), .A(n5789), .ZN(n5791) );
  AOI21_X1 U6944 ( .B1(n6087), .B2(n6385), .A(n5791), .ZN(n5792) );
  OAI21_X1 U6945 ( .B1(n5920), .B2(n6364), .A(n5792), .ZN(U2964) );
  AOI21_X1 U6946 ( .B1(n5795), .B2(n5794), .A(n5793), .ZN(n5930) );
  NOR2_X1 U6947 ( .A1(n6454), .A2(n6868), .ZN(n5922) );
  NOR2_X1 U6948 ( .A1(n5836), .A2(n5796), .ZN(n5797) );
  AOI211_X1 U6949 ( .C1(n6360), .C2(n5798), .A(n5922), .B(n5797), .ZN(n5800)
         );
  NAND2_X1 U6950 ( .A1(n6090), .A2(n6385), .ZN(n5799) );
  OAI211_X1 U6951 ( .C1(n5930), .C2(n6364), .A(n5800), .B(n5799), .ZN(U2965)
         );
  OAI21_X1 U6952 ( .B1(n5802), .B2(n5801), .A(n4439), .ZN(n5943) );
  INV_X1 U6953 ( .A(n5803), .ZN(n6093) );
  INV_X1 U6954 ( .A(REIP_REG_20__SCAN_IN), .ZN(n5804) );
  NOR2_X1 U6955 ( .A1(n6454), .A2(n5804), .ZN(n5934) );
  AOI21_X1 U6956 ( .B1(n6380), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5934), 
        .ZN(n5805) );
  OAI21_X1 U6957 ( .B1(n5806), .B2(n6390), .A(n5805), .ZN(n5807) );
  AOI21_X1 U6958 ( .B1(n6093), .B2(n6385), .A(n5807), .ZN(n5808) );
  OAI21_X1 U6959 ( .B1(n5943), .B2(n6364), .A(n5808), .ZN(U2966) );
  AOI21_X1 U6960 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5809), .A(n4434), 
        .ZN(n5810) );
  XNOR2_X1 U6961 ( .A(n5810), .B(n6356), .ZN(n6120) );
  INV_X1 U6962 ( .A(n6120), .ZN(n5816) );
  AOI22_X1 U6963 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n6476), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n5811) );
  OAI21_X1 U6964 ( .B1(n5812), .B2(n6390), .A(n5811), .ZN(n5813) );
  AOI21_X1 U6965 ( .B1(n5814), .B2(n6385), .A(n5813), .ZN(n5815) );
  OAI21_X1 U6966 ( .B1(n5816), .B2(n6364), .A(n5815), .ZN(U2967) );
  XNOR2_X1 U6967 ( .A(n6356), .B(n5953), .ZN(n5818) );
  XNOR2_X1 U6968 ( .A(n5817), .B(n5818), .ZN(n5963) );
  INV_X1 U6969 ( .A(n5819), .ZN(n5821) );
  AOI22_X1 U6970 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6476), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5820) );
  OAI21_X1 U6971 ( .B1(n6390), .B2(n5821), .A(n5820), .ZN(n5822) );
  AOI21_X1 U6972 ( .B1(n6316), .B2(n6385), .A(n5822), .ZN(n5823) );
  OAI21_X1 U6973 ( .B1(n5963), .B2(n6364), .A(n5823), .ZN(U2970) );
  XNOR2_X1 U6974 ( .A(n6356), .B(n6140), .ZN(n5825) );
  XNOR2_X1 U6975 ( .A(n5824), .B(n5825), .ZN(n6137) );
  INV_X1 U6976 ( .A(n6137), .ZN(n5831) );
  AOI22_X1 U6977 ( .A1(n6380), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6476), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5826) );
  OAI21_X1 U6978 ( .B1(n5827), .B2(n6390), .A(n5826), .ZN(n5828) );
  AOI21_X1 U6979 ( .B1(n5829), .B2(n6385), .A(n5828), .ZN(n5830) );
  OAI21_X1 U6980 ( .B1(n5831), .B2(n6364), .A(n5830), .ZN(U2971) );
  XNOR2_X1 U6981 ( .A(n6356), .B(n5833), .ZN(n5834) );
  XNOR2_X1 U6982 ( .A(n5832), .B(n5834), .ZN(n6149) );
  INV_X1 U6983 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5835) );
  OAI22_X1 U6984 ( .A1(n5836), .A2(n6209), .B1(n6454), .B2(n5835), .ZN(n5837)
         );
  AOI21_X1 U6985 ( .B1(n6360), .B2(n5838), .A(n5837), .ZN(n5841) );
  OR2_X1 U6986 ( .A1(n6213), .A2(n5839), .ZN(n5840) );
  OAI211_X1 U6987 ( .C1(n6149), .C2(n6364), .A(n5841), .B(n5840), .ZN(U2972)
         );
  AND2_X1 U6988 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5896) );
  OR2_X1 U6989 ( .A1(n6478), .A2(n6433), .ZN(n5931) );
  INV_X1 U6990 ( .A(n5842), .ZN(n5843) );
  NAND2_X1 U6991 ( .A1(n5931), .A2(n5843), .ZN(n5844) );
  OAI21_X1 U6992 ( .B1(n6403), .B2(n5896), .A(n6117), .ZN(n5883) );
  AOI21_X1 U6993 ( .B1(n5846), .B2(n5959), .A(n5883), .ZN(n5863) );
  OAI21_X1 U6994 ( .B1(n6403), .B2(n5847), .A(n5863), .ZN(n5853) );
  NAND2_X1 U6995 ( .A1(n6110), .A2(n5896), .ZN(n5885) );
  NOR2_X1 U6996 ( .A1(n5885), .A2(n5846), .ZN(n5872) );
  NAND3_X1 U6997 ( .A1(n5872), .A2(n5847), .A3(n4233), .ZN(n5850) );
  INV_X1 U6998 ( .A(n5848), .ZN(n5849) );
  OAI211_X1 U6999 ( .C1(n6448), .C2(n5851), .A(n5850), .B(n5849), .ZN(n5852)
         );
  AOI21_X1 U7000 ( .B1(n5853), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5852), 
        .ZN(n5854) );
  OAI21_X1 U7001 ( .B1(n5855), .B2(n6455), .A(n5854), .ZN(U2987) );
  INV_X1 U7002 ( .A(n5856), .ZN(n5866) );
  INV_X1 U7003 ( .A(n5857), .ZN(n5862) );
  INV_X1 U7004 ( .A(n5872), .ZN(n5859) );
  NOR3_X1 U7005 ( .A1(n5859), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5858), 
        .ZN(n5860) );
  AOI211_X1 U7006 ( .C1(n6467), .C2(n5862), .A(n5861), .B(n5860), .ZN(n5865)
         );
  INV_X1 U7007 ( .A(n6117), .ZN(n5909) );
  NAND2_X1 U7008 ( .A1(n5863), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5871) );
  OAI211_X1 U7009 ( .C1(n5959), .C2(n5909), .A(n5871), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5864) );
  OAI211_X1 U7010 ( .C1(n5866), .C2(n6455), .A(n5865), .B(n5864), .ZN(U2988)
         );
  INV_X1 U7011 ( .A(n5867), .ZN(n5870) );
  INV_X1 U7012 ( .A(n5868), .ZN(n5869) );
  AOI21_X1 U7013 ( .B1(n5870), .B2(n6467), .A(n5869), .ZN(n5874) );
  OAI21_X1 U7014 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5872), .A(n5871), 
        .ZN(n5873) );
  OAI211_X1 U7015 ( .C1(n5875), .C2(n6455), .A(n5874), .B(n5873), .ZN(U2989)
         );
  XNOR2_X1 U7016 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7017 ( .A1(n5876), .A2(n6467), .ZN(n5877) );
  OAI211_X1 U7018 ( .C1(n5885), .C2(n5879), .A(n5878), .B(n5877), .ZN(n5880)
         );
  AOI21_X1 U7019 ( .B1(n5883), .B2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5880), 
        .ZN(n5881) );
  OAI21_X1 U7020 ( .B1(n5882), .B2(n6455), .A(n5881), .ZN(U2990) );
  INV_X1 U7021 ( .A(n5883), .ZN(n5893) );
  NAND2_X1 U7022 ( .A1(n5884), .A2(n6474), .ZN(n5891) );
  INV_X1 U7023 ( .A(n5885), .ZN(n5889) );
  NOR2_X1 U7024 ( .A1(n5886), .A2(n6448), .ZN(n5888) );
  AOI211_X1 U7025 ( .C1(n5889), .C2(n5892), .A(n5888), .B(n5887), .ZN(n5890)
         );
  OAI211_X1 U7026 ( .C1(n5893), .C2(n5892), .A(n5891), .B(n5890), .ZN(U2991)
         );
  OAI21_X1 U7027 ( .B1(n6052), .B2(n6448), .A(n5894), .ZN(n5899) );
  INV_X1 U7028 ( .A(n6110), .ZN(n5897) );
  NOR3_X1 U7029 ( .A1(n5897), .A2(n5896), .A3(n5895), .ZN(n5898) );
  AOI211_X1 U7030 ( .C1(n5909), .C2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5899), .B(n5898), .ZN(n5900) );
  OAI21_X1 U7031 ( .B1(n5901), .B2(n6455), .A(n5900), .ZN(U2992) );
  NAND2_X1 U7032 ( .A1(n5902), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U7033 ( .B1(n5921), .B2(n5904), .A(n5903), .ZN(n5908) );
  OAI21_X1 U7034 ( .B1(n5906), .B2(n6448), .A(n5905), .ZN(n5907) );
  AOI21_X1 U7035 ( .B1(n5909), .B2(n5908), .A(n5907), .ZN(n5910) );
  OAI21_X1 U7036 ( .B1(n5911), .B2(n6455), .A(n5910), .ZN(U2994) );
  INV_X1 U7037 ( .A(n5912), .ZN(n5918) );
  AOI21_X1 U7038 ( .B1(n6467), .B2(n5914), .A(n5913), .ZN(n5915) );
  OAI21_X1 U7039 ( .B1(n5916), .B2(n5927), .A(n5915), .ZN(n5917) );
  AOI21_X1 U7040 ( .B1(n5918), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5917), 
        .ZN(n5919) );
  OAI21_X1 U7041 ( .B1(n5920), .B2(n6455), .A(n5919), .ZN(U2996) );
  INV_X1 U7042 ( .A(n5921), .ZN(n5928) );
  AOI21_X1 U7043 ( .B1(n6467), .B2(n5923), .A(n5922), .ZN(n5924) );
  OAI21_X1 U7044 ( .B1(n5925), .B2(n5927), .A(n5924), .ZN(n5926) );
  AOI21_X1 U7045 ( .B1(n5928), .B2(n5927), .A(n5926), .ZN(n5929) );
  OAI21_X1 U7046 ( .B1(n5930), .B2(n6455), .A(n5929), .ZN(U2997) );
  NAND2_X1 U7047 ( .A1(n5931), .A2(n6127), .ZN(n5932) );
  AND2_X1 U7048 ( .A1(n6126), .A2(n5932), .ZN(n5952) );
  NAND2_X1 U7049 ( .A1(n5959), .A2(n5951), .ZN(n5933) );
  AND2_X1 U7050 ( .A1(n5952), .A2(n5933), .ZN(n6124) );
  AOI21_X1 U7051 ( .B1(n6467), .B2(n6081), .A(n5934), .ZN(n5939) );
  INV_X1 U7052 ( .A(n5935), .ZN(n5937) );
  NAND2_X1 U7053 ( .A1(n6123), .A2(n5940), .ZN(n5936) );
  NAND3_X1 U7054 ( .A1(n6118), .A2(n5937), .A3(n5936), .ZN(n5938) );
  OAI211_X1 U7055 ( .C1(n6124), .C2(n5940), .A(n5939), .B(n5938), .ZN(n5941)
         );
  INV_X1 U7056 ( .A(n5941), .ZN(n5942) );
  OAI21_X1 U7057 ( .B1(n5943), .B2(n6455), .A(n5942), .ZN(U2998) );
  NAND3_X1 U7058 ( .A1(n5817), .A2(n5944), .A3(n5953), .ZN(n6099) );
  NOR3_X1 U7059 ( .A1(n5817), .A2(n5944), .A3(n5953), .ZN(n6101) );
  NAND2_X1 U7060 ( .A1(n6101), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5945) );
  OAI21_X1 U7061 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6099), .A(n5945), 
        .ZN(n5946) );
  XNOR2_X1 U7062 ( .A(n5946), .B(n5951), .ZN(n6096) );
  NAND2_X1 U7063 ( .A1(n6096), .A2(n6474), .ZN(n5950) );
  NOR3_X1 U7064 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6127), .A3(n6128), 
        .ZN(n5948) );
  NOR2_X1 U7065 ( .A1(n6448), .A2(n6199), .ZN(n5947) );
  AOI211_X1 U7066 ( .C1(n6476), .C2(REIP_REG_18__SCAN_IN), .A(n5948), .B(n5947), .ZN(n5949) );
  OAI211_X1 U7067 ( .C1(n5952), .C2(n5951), .A(n5950), .B(n5949), .ZN(U3000)
         );
  AOI211_X1 U7068 ( .C1(n6140), .C2(n5953), .A(n6163), .B(n6134), .ZN(n5958)
         );
  NOR2_X1 U7069 ( .A1(n6454), .A2(n6985), .ZN(n5956) );
  NOR2_X1 U7070 ( .A1(n6448), .A2(n5954), .ZN(n5955) );
  AOI211_X1 U7071 ( .C1(n5958), .C2(n5957), .A(n5956), .B(n5955), .ZN(n5962)
         );
  AND2_X1 U7072 ( .A1(n5959), .A2(n6134), .ZN(n5960) );
  OR2_X1 U7073 ( .A1(n6393), .A2(n5960), .ZN(n6133) );
  NAND2_X1 U7074 ( .A1(n6133), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5961) );
  OAI211_X1 U7075 ( .C1(n5963), .C2(n6455), .A(n5962), .B(n5961), .ZN(U3002)
         );
  OAI22_X1 U7076 ( .A1(n5966), .A2(n5965), .B1(n5964), .B2(n6646), .ZN(n5968)
         );
  MUX2_X1 U7077 ( .A(n5968), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n5967), 
        .Z(U3456) );
  NOR3_X4 U7078 ( .A1(n5971), .A2(n5970), .A3(n5969), .ZN(n6047) );
  NOR3_X1 U7079 ( .A1(n6047), .A2(n5972), .A3(n6496), .ZN(n5973) );
  NOR2_X1 U7080 ( .A1(n5973), .A2(n6499), .ZN(n5977) );
  OR2_X1 U7081 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5974), .ZN(n6004)
         );
  AOI211_X1 U7082 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6004), .A(n6489), .B(
        n5975), .ZN(n5976) );
  NAND2_X1 U7083 ( .A1(n6002), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5983) );
  AOI22_X1 U7084 ( .A1(n5980), .A2(n6015), .B1(n5979), .B2(n5978), .ZN(n6003)
         );
  OAI22_X1 U7085 ( .A1(n6493), .A2(n6004), .B1(n6003), .B2(n6492), .ZN(n5981)
         );
  AOI21_X1 U7086 ( .B1(n6047), .B2(n6504), .A(n5981), .ZN(n5982) );
  OAI211_X1 U7087 ( .C1(n6008), .C2(n6507), .A(n5983), .B(n5982), .ZN(U3020)
         );
  NAND2_X1 U7088 ( .A1(n6002), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5986) );
  OAI22_X1 U7089 ( .A1(n6552), .A2(n6004), .B1(n6003), .B2(n6508), .ZN(n5984)
         );
  AOI21_X1 U7090 ( .B1(n6047), .B2(n6510), .A(n5984), .ZN(n5985) );
  OAI211_X1 U7091 ( .C1(n6008), .C2(n6513), .A(n5986), .B(n5985), .ZN(U3021)
         );
  NAND2_X1 U7092 ( .A1(n6002), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5989) );
  OAI22_X1 U7093 ( .A1(n6515), .A2(n6004), .B1(n6003), .B2(n6514), .ZN(n5987)
         );
  AOI21_X1 U7094 ( .B1(n6047), .B2(n6517), .A(n5987), .ZN(n5988) );
  OAI211_X1 U7095 ( .C1(n6008), .C2(n6520), .A(n5989), .B(n5988), .ZN(U3022)
         );
  NAND2_X1 U7096 ( .A1(n6002), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5992) );
  OAI22_X1 U7097 ( .A1(n6586), .A2(n6004), .B1(n6003), .B2(n6521), .ZN(n5990)
         );
  AOI21_X1 U7098 ( .B1(n6047), .B2(n6523), .A(n5990), .ZN(n5991) );
  OAI211_X1 U7099 ( .C1(n6008), .C2(n6587), .A(n5992), .B(n5991), .ZN(U3023)
         );
  NAND2_X1 U7100 ( .A1(n6002), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5995) );
  OAI22_X1 U7101 ( .A1(n6563), .A2(n6004), .B1(n6003), .B2(n6526), .ZN(n5993)
         );
  AOI21_X1 U7102 ( .B1(n6047), .B2(n6528), .A(n5993), .ZN(n5994) );
  OAI211_X1 U7103 ( .C1(n6008), .C2(n6531), .A(n5995), .B(n5994), .ZN(U3024)
         );
  NAND2_X1 U7104 ( .A1(n6002), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5998) );
  OAI22_X1 U7105 ( .A1(n6593), .A2(n6004), .B1(n6003), .B2(n6532), .ZN(n5996)
         );
  AOI21_X1 U7106 ( .B1(n6047), .B2(n6534), .A(n5996), .ZN(n5997) );
  OAI211_X1 U7107 ( .C1(n6008), .C2(n6594), .A(n5998), .B(n5997), .ZN(U3025)
         );
  NAND2_X1 U7108 ( .A1(n6002), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6001) );
  OAI22_X1 U7109 ( .A1(n6570), .A2(n6004), .B1(n6003), .B2(n6537), .ZN(n5999)
         );
  AOI21_X1 U7110 ( .B1(n6047), .B2(n6539), .A(n5999), .ZN(n6000) );
  OAI211_X1 U7111 ( .C1(n6008), .C2(n6542), .A(n6001), .B(n6000), .ZN(U3026)
         );
  NAND2_X1 U7112 ( .A1(n6002), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6007) );
  OAI22_X1 U7113 ( .A1(n6601), .A2(n6004), .B1(n6003), .B2(n6543), .ZN(n6005)
         );
  AOI21_X1 U7114 ( .B1(n6047), .B2(n6548), .A(n6005), .ZN(n6006) );
  OAI211_X1 U7115 ( .C1(n6008), .C2(n6602), .A(n6007), .B(n6006), .ZN(U3027)
         );
  AOI21_X1 U7116 ( .B1(n6009), .B2(n6385), .A(n6499), .ZN(n6011) );
  OAI21_X1 U7117 ( .B1(n6010), .B2(n6498), .A(n6045), .ZN(n6016) );
  OR2_X1 U7118 ( .A1(n6011), .A2(n6016), .ZN(n6013) );
  NAND2_X1 U7119 ( .A1(n6043), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n6020)
         );
  AOI22_X1 U7120 ( .A1(n6016), .A2(n6015), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6014), .ZN(n6044) );
  OAI22_X1 U7121 ( .A1(n6493), .A2(n6045), .B1(n6044), .B2(n6492), .ZN(n6017)
         );
  AOI21_X1 U7122 ( .B1(n6047), .B2(n6018), .A(n6017), .ZN(n6019) );
  OAI211_X1 U7123 ( .C1(n6050), .C2(n6021), .A(n6020), .B(n6019), .ZN(U3140)
         );
  NAND2_X1 U7124 ( .A1(n6043), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6024)
         );
  OAI22_X1 U7125 ( .A1(n6552), .A2(n6045), .B1(n6044), .B2(n6508), .ZN(n6022)
         );
  AOI21_X1 U7126 ( .B1(n6047), .B2(n6554), .A(n6022), .ZN(n6023) );
  OAI211_X1 U7127 ( .C1(n6050), .C2(n6558), .A(n6024), .B(n6023), .ZN(U3141)
         );
  NAND2_X1 U7128 ( .A1(n6043), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6028)
         );
  OAI22_X1 U7129 ( .A1(n6515), .A2(n6045), .B1(n6044), .B2(n6514), .ZN(n6025)
         );
  AOI21_X1 U7130 ( .B1(n6047), .B2(n6026), .A(n6025), .ZN(n6027) );
  OAI211_X1 U7131 ( .C1(n6050), .C2(n6029), .A(n6028), .B(n6027), .ZN(U3142)
         );
  NAND2_X1 U7132 ( .A1(n6043), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6032)
         );
  OAI22_X1 U7133 ( .A1(n6586), .A2(n6045), .B1(n6044), .B2(n6521), .ZN(n6030)
         );
  AOI21_X1 U7134 ( .B1(n6047), .B2(n6560), .A(n6030), .ZN(n6031) );
  OAI211_X1 U7135 ( .C1(n6050), .C2(n6592), .A(n6032), .B(n6031), .ZN(U3143)
         );
  NAND2_X1 U7136 ( .A1(n6043), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6035)
         );
  OAI22_X1 U7137 ( .A1(n6563), .A2(n6045), .B1(n6044), .B2(n6526), .ZN(n6033)
         );
  AOI21_X1 U7138 ( .B1(n6047), .B2(n6565), .A(n6033), .ZN(n6034) );
  OAI211_X1 U7139 ( .C1(n6050), .C2(n6569), .A(n6035), .B(n6034), .ZN(U3144)
         );
  NAND2_X1 U7140 ( .A1(n6043), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6039)
         );
  OAI22_X1 U7141 ( .A1(n6593), .A2(n6045), .B1(n6044), .B2(n6532), .ZN(n6036)
         );
  AOI21_X1 U7142 ( .B1(n6047), .B2(n6037), .A(n6036), .ZN(n6038) );
  OAI211_X1 U7143 ( .C1(n6050), .C2(n6599), .A(n6039), .B(n6038), .ZN(U3145)
         );
  NAND2_X1 U7144 ( .A1(n6043), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6042)
         );
  OAI22_X1 U7145 ( .A1(n6570), .A2(n6045), .B1(n6044), .B2(n6537), .ZN(n6040)
         );
  AOI21_X1 U7146 ( .B1(n6047), .B2(n6572), .A(n6040), .ZN(n6041) );
  OAI211_X1 U7147 ( .C1(n6050), .C2(n6576), .A(n6042), .B(n6041), .ZN(U3146)
         );
  NAND2_X1 U7148 ( .A1(n6043), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6049)
         );
  OAI22_X1 U7149 ( .A1(n6601), .A2(n6045), .B1(n6044), .B2(n6543), .ZN(n6046)
         );
  AOI21_X1 U7150 ( .B1(n6047), .B2(n6579), .A(n6046), .ZN(n6048) );
  OAI211_X1 U7151 ( .C1(n6050), .C2(n6611), .A(n6049), .B(n6048), .ZN(U3147)
         );
  AOI22_X1 U7152 ( .A1(EBX_REG_26__SCAN_IN), .A2(n6288), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6285), .ZN(n6058) );
  INV_X1 U7153 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6697) );
  NOR2_X1 U7154 ( .A1(n6697), .A2(n6051), .ZN(n6060) );
  AOI21_X1 U7155 ( .B1(REIP_REG_25__SCAN_IN), .B2(n6060), .A(
        REIP_REG_26__SCAN_IN), .ZN(n6054) );
  OAI22_X1 U7156 ( .A1(n6054), .A2(n6053), .B1(n6052), .B2(n6274), .ZN(n6055)
         );
  AOI21_X1 U7157 ( .B1(n6056), .B2(n4408), .A(n6055), .ZN(n6057) );
  OAI211_X1 U7158 ( .C1(n6059), .C2(n6279), .A(n6058), .B(n6057), .ZN(U2801)
         );
  AOI22_X1 U7159 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6288), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6285), .ZN(n6068) );
  AOI22_X1 U7160 ( .A1(n6061), .A2(n6294), .B1(n6060), .B2(n5765), .ZN(n6067)
         );
  NOR2_X1 U7161 ( .A1(n6274), .A2(n6111), .ZN(n6062) );
  AOI21_X1 U7162 ( .B1(n6063), .B2(n4408), .A(n6062), .ZN(n6066) );
  OAI21_X1 U7163 ( .B1(n6064), .B2(n6075), .A(REIP_REG_25__SCAN_IN), .ZN(n6065) );
  NAND4_X1 U7164 ( .A1(n6068), .A2(n6067), .A3(n6066), .A4(n6065), .ZN(U2802)
         );
  INV_X1 U7165 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6078) );
  AOI22_X1 U7166 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n6285), .B1(n6069), 
        .B2(n6294), .ZN(n6077) );
  INV_X1 U7167 ( .A(n6070), .ZN(n6071) );
  OAI22_X1 U7168 ( .A1(n6072), .A2(n6212), .B1(n6071), .B2(n6274), .ZN(n6073)
         );
  OAI211_X1 U7169 ( .C1(n6078), .C2(n6270), .A(n6077), .B(n6076), .ZN(U2804)
         );
  AOI21_X1 U7170 ( .B1(REIP_REG_19__SCAN_IN), .B2(n6079), .A(
        REIP_REG_20__SCAN_IN), .ZN(n6085) );
  AOI22_X1 U7171 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6288), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6285), .ZN(n6083) );
  AOI222_X1 U7172 ( .A1(n6081), .A2(n6286), .B1(n4408), .B2(n6093), .C1(n6080), 
        .C2(n6294), .ZN(n6082) );
  OAI211_X1 U7173 ( .C1(n6085), .C2(n6084), .A(n6083), .B(n6082), .ZN(U2807)
         );
  AOI22_X1 U7174 ( .A1(n6087), .A2(n6315), .B1(n6314), .B2(DATAI_22_), .ZN(
        n6089) );
  AOI22_X1 U7175 ( .A1(n6318), .A2(DATAI_6_), .B1(n6317), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7176 ( .A1(n6089), .A2(n6088), .ZN(U2869) );
  AOI22_X1 U7177 ( .A1(n6090), .A2(n6315), .B1(n6314), .B2(DATAI_21_), .ZN(
        n6092) );
  AOI22_X1 U7178 ( .A1(n6318), .A2(DATAI_5_), .B1(n6317), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7179 ( .A1(n6092), .A2(n6091), .ZN(U2870) );
  AOI22_X1 U7180 ( .A1(n6093), .A2(n6315), .B1(n6314), .B2(DATAI_20_), .ZN(
        n6095) );
  AOI22_X1 U7181 ( .A1(n6318), .A2(DATAI_4_), .B1(n6317), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6094) );
  NAND2_X1 U7182 ( .A1(n6095), .A2(n6094), .ZN(U2871) );
  AOI22_X1 U7183 ( .A1(n6476), .A2(REIP_REG_18__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6098) );
  AOI22_X1 U7184 ( .A1(n6096), .A2(n6386), .B1(n6385), .B2(n6308), .ZN(n6097)
         );
  OAI211_X1 U7185 ( .C1(n6390), .C2(n6207), .A(n6098), .B(n6097), .ZN(U2968)
         );
  INV_X1 U7186 ( .A(n6099), .ZN(n6100) );
  NOR2_X1 U7187 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  XNOR2_X1 U7188 ( .A(n6102), .B(n6127), .ZN(n6132) );
  AOI22_X1 U7189 ( .A1(n6476), .A2(REIP_REG_17__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6105) );
  AOI22_X1 U7190 ( .A1(n6311), .A2(n6385), .B1(n6360), .B2(n6103), .ZN(n6104)
         );
  OAI211_X1 U7191 ( .C1(n6132), .C2(n6364), .A(n6105), .B(n6104), .ZN(U2969)
         );
  AOI22_X1 U7192 ( .A1(n6476), .A2(REIP_REG_13__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6109) );
  XNOR2_X1 U7193 ( .A(n6106), .B(n6107), .ZN(n6159) );
  AOI22_X1 U7194 ( .A1(n6159), .A2(n6386), .B1(n6385), .B2(n6300), .ZN(n6108)
         );
  OAI211_X1 U7195 ( .C1(n6390), .C2(n6226), .A(n6109), .B(n6108), .ZN(U2973)
         );
  AOI22_X1 U7196 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6476), .B1(n6110), .B2(
        n6116), .ZN(n6115) );
  INV_X1 U7197 ( .A(n6111), .ZN(n6112) );
  AOI22_X1 U7198 ( .A1(n6113), .A2(n6474), .B1(n6467), .B2(n6112), .ZN(n6114)
         );
  OAI211_X1 U7199 ( .C1(n6117), .C2(n6116), .A(n6115), .B(n6114), .ZN(U2993)
         );
  AOI22_X1 U7200 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6476), .B1(n6118), .B2(
        n6123), .ZN(n6122) );
  AOI22_X1 U7201 ( .A1(n6120), .A2(n6474), .B1(n6467), .B2(n6119), .ZN(n6121)
         );
  OAI211_X1 U7202 ( .C1(n6124), .C2(n6123), .A(n6122), .B(n6121), .ZN(U2999)
         );
  NAND2_X1 U7203 ( .A1(n6476), .A2(REIP_REG_17__SCAN_IN), .ZN(n6125) );
  OAI221_X1 U7204 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n6128), .C1(
        n6127), .C2(n6126), .A(n6125), .ZN(n6129) );
  AOI21_X1 U7205 ( .B1(n6130), .B2(n6467), .A(n6129), .ZN(n6131) );
  OAI21_X1 U7206 ( .B1(n6132), .B2(n6455), .A(n6131), .ZN(U3001) );
  INV_X1 U7207 ( .A(n6133), .ZN(n6141) );
  NOR2_X1 U7208 ( .A1(n6163), .A2(n6134), .ZN(n6135) );
  AOI22_X1 U7209 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6476), .B1(n6135), .B2(
        n6140), .ZN(n6139) );
  AOI22_X1 U7210 ( .A1(n6137), .A2(n6474), .B1(n6467), .B2(n6136), .ZN(n6138)
         );
  OAI211_X1 U7211 ( .C1(n6141), .C2(n6140), .A(n6139), .B(n6138), .ZN(U3003)
         );
  NAND2_X1 U7212 ( .A1(n6144), .A2(n6392), .ZN(n6154) );
  INV_X1 U7213 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7214 ( .A1(n6146), .A2(n6142), .ZN(n6162) );
  OAI22_X1 U7215 ( .A1(n6146), .A2(n6145), .B1(n6144), .B2(n6143), .ZN(n6147)
         );
  NOR2_X1 U7216 ( .A1(n6393), .A2(n6147), .ZN(n6157) );
  OAI21_X1 U7217 ( .B1(n6148), .B2(n6162), .A(n6157), .ZN(n6151) );
  OAI22_X1 U7218 ( .A1(n6149), .A2(n6455), .B1(n6448), .B2(n6208), .ZN(n6150)
         );
  AOI21_X1 U7219 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6151), .A(n6150), 
        .ZN(n6153) );
  NAND2_X1 U7220 ( .A1(n6476), .A2(REIP_REG_14__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7221 ( .C1(INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n6154), .A(n6153), .B(n6152), .ZN(U3004) );
  AOI21_X1 U7222 ( .B1(n6156), .B2(n5438), .A(n6155), .ZN(n6299) );
  AOI22_X1 U7223 ( .A1(n6467), .A2(n6299), .B1(n6476), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n6161) );
  INV_X1 U7224 ( .A(n6157), .ZN(n6158) );
  AOI22_X1 U7225 ( .A1(n6159), .A2(n6474), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6158), .ZN(n6160) );
  OAI211_X1 U7226 ( .C1(n6163), .C2(n6162), .A(n6161), .B(n6160), .ZN(U3005)
         );
  INV_X1 U7227 ( .A(n6164), .ZN(n6167) );
  NAND3_X1 U7228 ( .A1(n6167), .A2(n6166), .A3(n6165), .ZN(n6168) );
  OAI21_X1 U7229 ( .B1(n6170), .B2(n6169), .A(n6168), .ZN(U3455) );
  INV_X1 U7230 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6677) );
  AOI21_X1 U7231 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6814), .A(n6677), .ZN(n6175) );
  INV_X1 U7232 ( .A(ADS_N_REG_SCAN_IN), .ZN(n7083) );
  AOI21_X1 U7233 ( .B1(n6175), .B2(n7083), .A(n7129), .ZN(U2789) );
  OAI21_X1 U7234 ( .B1(n6171), .B2(n6655), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6172) );
  OAI21_X1 U7235 ( .B1(n6173), .B2(n6659), .A(n6172), .ZN(U2790) );
  INV_X1 U7236 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6962) );
  NOR2_X1 U7237 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6176) );
  NOR2_X1 U7238 ( .A1(n7129), .A2(n6176), .ZN(n6174) );
  AOI22_X1 U7239 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7129), .B1(n6962), .B2(
        n6174), .ZN(U2791) );
  NOR2_X2 U7240 ( .A1(n7129), .A2(n6175), .ZN(n6707) );
  OAI21_X1 U7241 ( .B1(BS16_N), .B2(n6176), .A(n6707), .ZN(n6705) );
  OAI21_X1 U7242 ( .B1(n6707), .B2(n6177), .A(n6705), .ZN(U2792) );
  INV_X1 U7243 ( .A(n6178), .ZN(n6180) );
  OAI21_X1 U7244 ( .B1(n6180), .B2(n6179), .A(n6364), .ZN(U2793) );
  NOR4_X1 U7245 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_9__SCAN_IN), .A4(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6184) );
  NOR4_X1 U7246 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_13__SCAN_IN), .A4(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6183)
         );
  NOR4_X1 U7247 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6182) );
  NOR4_X1 U7248 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6181) );
  NAND4_X1 U7249 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n6190)
         );
  NOR4_X1 U7250 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), .A3(DATAWIDTH_REG_18__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6188) );
  AOI211_X1 U7251 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_20__SCAN_IN), .B(
        DATAWIDTH_REG_12__SCAN_IN), .ZN(n6187) );
  NOR4_X1 U7252 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6186) );
  NOR4_X1 U7253 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6185) );
  NAND4_X1 U7254 ( .A1(n6188), .A2(n6187), .A3(n6186), .A4(n6185), .ZN(n6189)
         );
  NOR2_X1 U7255 ( .A1(n6190), .A2(n6189), .ZN(n6716) );
  INV_X1 U7256 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n7067) );
  NOR3_X1 U7257 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6192) );
  OAI21_X1 U7258 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6192), .A(n6716), .ZN(n6191)
         );
  OAI21_X1 U7259 ( .B1(n6716), .B2(n7067), .A(n6191), .ZN(U2794) );
  INV_X1 U7260 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6706) );
  AOI21_X1 U7261 ( .B1(n5011), .B2(n6706), .A(n6192), .ZN(n6194) );
  INV_X1 U7262 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6193) );
  INV_X1 U7263 ( .A(n6716), .ZN(n6714) );
  AOI22_X1 U7264 ( .A1(n6716), .A2(n6194), .B1(n6193), .B2(n6714), .ZN(U2795)
         );
  NAND2_X1 U7265 ( .A1(n6195), .A2(REIP_REG_18__SCAN_IN), .ZN(n6204) );
  INV_X1 U7266 ( .A(n6196), .ZN(n6197) );
  NAND2_X1 U7267 ( .A1(n6257), .A2(n6197), .ZN(n6198) );
  AOI21_X1 U7268 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6285), .A(n6198), 
        .ZN(n6203) );
  NAND2_X1 U7269 ( .A1(n6288), .A2(EBX_REG_18__SCAN_IN), .ZN(n6202) );
  INV_X1 U7270 ( .A(n6199), .ZN(n6200) );
  NAND2_X1 U7271 ( .A1(n6286), .A2(n6200), .ZN(n6201) );
  NAND4_X1 U7272 ( .A1(n6204), .A2(n6203), .A3(n6202), .A4(n6201), .ZN(n6205)
         );
  AOI21_X1 U7273 ( .B1(n6308), .B2(n4408), .A(n6205), .ZN(n6206) );
  OAI21_X1 U7274 ( .B1(n6207), .B2(n6279), .A(n6206), .ZN(U2809) );
  INV_X1 U7275 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6690) );
  NOR2_X1 U7276 ( .A1(n6690), .A2(n5450), .ZN(n6219) );
  AOI21_X1 U7277 ( .B1(n6219), .B2(n6221), .A(REIP_REG_14__SCAN_IN), .ZN(n6218) );
  OAI22_X1 U7278 ( .A1(n6258), .A2(n6209), .B1(n6274), .B2(n6208), .ZN(n6210)
         );
  AOI211_X1 U7279 ( .C1(n6288), .C2(EBX_REG_14__SCAN_IN), .A(n6268), .B(n6210), 
        .ZN(n6216) );
  OAI22_X1 U7280 ( .A1(n6213), .A2(n6212), .B1(n6279), .B2(n6211), .ZN(n6214)
         );
  INV_X1 U7281 ( .A(n6214), .ZN(n6215) );
  OAI211_X1 U7282 ( .C1(n6218), .C2(n6217), .A(n6216), .B(n6215), .ZN(U2813)
         );
  AOI22_X1 U7283 ( .A1(n6228), .A2(REIP_REG_13__SCAN_IN), .B1(n6286), .B2(
        n6299), .ZN(n6225) );
  INV_X1 U7284 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6302) );
  AOI21_X1 U7285 ( .B1(n6690), .B2(n5450), .A(n6219), .ZN(n6220) );
  AOI22_X1 U7286 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6285), .B1(n6221), 
        .B2(n6220), .ZN(n6222) );
  OAI211_X1 U7287 ( .C1(n6302), .C2(n6270), .A(n6222), .B(n6257), .ZN(n6223)
         );
  AOI21_X1 U7288 ( .B1(n6300), .B2(n4408), .A(n6223), .ZN(n6224) );
  OAI211_X1 U7289 ( .C1(n6226), .C2(n6279), .A(n6225), .B(n6224), .ZN(U2814)
         );
  AOI21_X1 U7290 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6227), .A(
        REIP_REG_11__SCAN_IN), .ZN(n6238) );
  INV_X1 U7291 ( .A(n6228), .ZN(n6237) );
  AOI21_X1 U7292 ( .B1(n6231), .B2(n6230), .A(n6229), .ZN(n6391) );
  INV_X1 U7293 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6306) );
  NOR2_X1 U7294 ( .A1(n6270), .A2(n6306), .ZN(n6234) );
  OAI21_X1 U7295 ( .B1(n6258), .B2(n6232), .A(n6257), .ZN(n6233) );
  AOI211_X1 U7296 ( .C1(n6391), .C2(n6286), .A(n6234), .B(n6233), .ZN(n6236)
         );
  AOI22_X1 U7297 ( .A1(n6361), .A2(n4408), .B1(n6294), .B2(n6359), .ZN(n6235)
         );
  OAI211_X1 U7298 ( .C1(n6238), .C2(n6237), .A(n6236), .B(n6235), .ZN(U2816)
         );
  INV_X1 U7299 ( .A(n6409), .ZN(n6240) );
  NAND2_X1 U7300 ( .A1(n6285), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6239)
         );
  OAI211_X1 U7301 ( .C1(n6274), .C2(n6240), .A(n6257), .B(n6239), .ZN(n6241)
         );
  INV_X1 U7302 ( .A(n6241), .ZN(n6251) );
  AOI22_X1 U7303 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6288), .B1(
        REIP_REG_9__SCAN_IN), .B2(n6242), .ZN(n6250) );
  INV_X1 U7304 ( .A(n6243), .ZN(n6245) );
  AOI22_X1 U7305 ( .A1(n6245), .A2(n4408), .B1(n6294), .B2(n6244), .ZN(n6249)
         );
  NAND3_X1 U7306 ( .A1(n6247), .A2(n6246), .A3(n5414), .ZN(n6248) );
  NAND4_X1 U7307 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(U2818)
         );
  NOR2_X1 U7308 ( .A1(n6252), .A2(n6270), .ZN(n6253) );
  AOI211_X1 U7309 ( .C1(n6255), .C2(REIP_REG_6__SCAN_IN), .A(n6254), .B(n6253), 
        .ZN(n6262) );
  NOR2_X1 U7310 ( .A1(n6274), .A2(n6256), .ZN(n6260) );
  OAI21_X1 U7311 ( .B1(n6258), .B2(n3813), .A(n6257), .ZN(n6259) );
  AOI211_X1 U7312 ( .C1(n6366), .C2(n4408), .A(n6260), .B(n6259), .ZN(n6261)
         );
  OAI211_X1 U7313 ( .C1(n6370), .C2(n6279), .A(n6262), .B(n6261), .ZN(U2821)
         );
  OAI21_X1 U7314 ( .B1(n6264), .B2(n6271), .A(n6263), .ZN(n6298) );
  OAI22_X1 U7315 ( .A1(n6298), .A2(n6684), .B1(n6266), .B2(n6265), .ZN(n6267)
         );
  AOI211_X1 U7316 ( .C1(n6285), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6268), 
        .B(n6267), .ZN(n6278) );
  NOR2_X1 U7317 ( .A1(n6270), .A2(n6269), .ZN(n6276) );
  OR3_X1 U7318 ( .A1(n6272), .A2(REIP_REG_4__SCAN_IN), .A3(n6271), .ZN(n6273)
         );
  OAI21_X1 U7319 ( .B1(n6274), .B2(n6447), .A(n6273), .ZN(n6275) );
  AOI211_X1 U7320 ( .C1(n6375), .C2(n6283), .A(n6276), .B(n6275), .ZN(n6277)
         );
  OAI211_X1 U7321 ( .C1(n6379), .C2(n6279), .A(n6278), .B(n6277), .ZN(U2823)
         );
  OR2_X1 U7322 ( .A1(n6281), .A2(n6280), .ZN(n6297) );
  INV_X1 U7323 ( .A(n6282), .ZN(n6284) );
  NAND2_X1 U7324 ( .A1(n6284), .A2(n6283), .ZN(n6292) );
  AOI22_X1 U7325 ( .A1(n6286), .A2(n6460), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .B2(n6285), .ZN(n6291) );
  NAND2_X1 U7326 ( .A1(n6287), .A2(n4712), .ZN(n6290) );
  NAND2_X1 U7327 ( .A1(n6288), .A2(EBX_REG_3__SCAN_IN), .ZN(n6289) );
  NAND4_X1 U7328 ( .A1(n6292), .A2(n6291), .A3(n6290), .A4(n6289), .ZN(n6293)
         );
  AOI21_X1 U7329 ( .B1(n6295), .B2(n6294), .A(n6293), .ZN(n6296) );
  OAI221_X1 U7330 ( .B1(n6298), .B2(n4775), .C1(n6298), .C2(n6297), .A(n6296), 
        .ZN(U2824) );
  AOI22_X1 U7331 ( .A1(n6300), .A2(n6304), .B1(n6303), .B2(n6299), .ZN(n6301)
         );
  OAI21_X1 U7332 ( .B1(n6307), .B2(n6302), .A(n6301), .ZN(U2846) );
  AOI22_X1 U7333 ( .A1(n6361), .A2(n6304), .B1(n6303), .B2(n6391), .ZN(n6305)
         );
  OAI21_X1 U7334 ( .B1(n6307), .B2(n6306), .A(n6305), .ZN(U2848) );
  AOI22_X1 U7335 ( .A1(n6308), .A2(n6315), .B1(n6314), .B2(DATAI_18_), .ZN(
        n6310) );
  AOI22_X1 U7336 ( .A1(n6318), .A2(DATAI_2_), .B1(n6317), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U7337 ( .A1(n6310), .A2(n6309), .ZN(U2873) );
  AOI22_X1 U7338 ( .A1(n6311), .A2(n6315), .B1(n6314), .B2(DATAI_17_), .ZN(
        n6313) );
  AOI22_X1 U7339 ( .A1(n6318), .A2(DATAI_1_), .B1(n6317), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7340 ( .A1(n6313), .A2(n6312), .ZN(U2874) );
  AOI22_X1 U7341 ( .A1(n6316), .A2(n6315), .B1(n6314), .B2(DATAI_16_), .ZN(
        n6320) );
  AOI22_X1 U7342 ( .A1(n6318), .A2(DATAI_0_), .B1(n6317), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7343 ( .A1(n6320), .A2(n6319), .ZN(U2875) );
  AOI22_X1 U7344 ( .A1(n6720), .A2(LWORD_REG_15__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6322) );
  OAI21_X1 U7345 ( .B1(n4535), .B2(n6352), .A(n6322), .ZN(U2908) );
  AOI22_X1 U7346 ( .A1(n6720), .A2(LWORD_REG_14__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6323) );
  OAI21_X1 U7347 ( .B1(n6324), .B2(n6352), .A(n6323), .ZN(U2909) );
  AOI22_X1 U7348 ( .A1(n6720), .A2(LWORD_REG_13__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6325) );
  OAI21_X1 U7349 ( .B1(n6326), .B2(n6352), .A(n6325), .ZN(U2910) );
  AOI22_X1 U7350 ( .A1(n6720), .A2(LWORD_REG_12__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6327) );
  OAI21_X1 U7351 ( .B1(n6328), .B2(n6352), .A(n6327), .ZN(U2911) );
  AOI22_X1 U7352 ( .A1(n6720), .A2(LWORD_REG_11__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6329) );
  OAI21_X1 U7353 ( .B1(n6330), .B2(n6352), .A(n6329), .ZN(U2912) );
  AOI22_X1 U7354 ( .A1(n6720), .A2(LWORD_REG_10__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6331) );
  OAI21_X1 U7355 ( .B1(n6332), .B2(n6352), .A(n6331), .ZN(U2913) );
  AOI22_X1 U7356 ( .A1(n6720), .A2(LWORD_REG_9__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6333) );
  OAI21_X1 U7357 ( .B1(n6334), .B2(n6352), .A(n6333), .ZN(U2914) );
  AOI22_X1 U7358 ( .A1(n6720), .A2(LWORD_REG_8__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6335) );
  OAI21_X1 U7359 ( .B1(n6336), .B2(n6352), .A(n6335), .ZN(U2915) );
  AOI22_X1 U7360 ( .A1(n6720), .A2(LWORD_REG_7__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6337) );
  OAI21_X1 U7361 ( .B1(n3820), .B2(n6352), .A(n6337), .ZN(U2916) );
  AOI22_X1 U7362 ( .A1(n6720), .A2(LWORD_REG_6__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7363 ( .B1(n3814), .B2(n6352), .A(n6338), .ZN(U2917) );
  AOI22_X1 U7364 ( .A1(n6720), .A2(LWORD_REG_5__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U7365 ( .B1(n6340), .B2(n6352), .A(n6339), .ZN(U2918) );
  AOI22_X1 U7366 ( .A1(n6720), .A2(LWORD_REG_4__SCAN_IN), .B1(n6341), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6342) );
  OAI21_X1 U7367 ( .B1(n6343), .B2(n6352), .A(n6342), .ZN(U2919) );
  AOI22_X1 U7368 ( .A1(n6720), .A2(LWORD_REG_3__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6344) );
  OAI21_X1 U7369 ( .B1(n6345), .B2(n6352), .A(n6344), .ZN(U2920) );
  AOI22_X1 U7370 ( .A1(n6720), .A2(LWORD_REG_2__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6346) );
  OAI21_X1 U7371 ( .B1(n6347), .B2(n6352), .A(n6346), .ZN(U2921) );
  AOI22_X1 U7372 ( .A1(n6720), .A2(LWORD_REG_1__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7373 ( .B1(n6349), .B2(n6352), .A(n6348), .ZN(U2922) );
  AOI22_X1 U7374 ( .A1(n6720), .A2(LWORD_REG_0__SCAN_IN), .B1(n6350), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6351) );
  OAI21_X1 U7375 ( .B1(n6353), .B2(n6352), .A(n6351), .ZN(U2923) );
  NAND2_X1 U7376 ( .A1(n6355), .A2(n6354), .ZN(n6358) );
  XNOR2_X1 U7377 ( .A(n6356), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6357)
         );
  XNOR2_X1 U7378 ( .A(n6358), .B(n6357), .ZN(n6396) );
  AOI22_X1 U7379 ( .A1(n6476), .A2(REIP_REG_11__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6363) );
  AOI22_X1 U7380 ( .A1(n6361), .A2(n6385), .B1(n6360), .B2(n6359), .ZN(n6362)
         );
  OAI211_X1 U7381 ( .C1(n6396), .C2(n6364), .A(n6363), .B(n6362), .ZN(U2975)
         );
  AOI22_X1 U7382 ( .A1(n6476), .A2(REIP_REG_6__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6369) );
  INV_X1 U7383 ( .A(n6365), .ZN(n6367) );
  AOI22_X1 U7384 ( .A1(n6367), .A2(n6386), .B1(n6385), .B2(n6366), .ZN(n6368)
         );
  OAI211_X1 U7385 ( .C1(n6390), .C2(n6370), .A(n6369), .B(n6368), .ZN(U2980)
         );
  AOI22_X1 U7386 ( .A1(n6476), .A2(REIP_REG_4__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6378) );
  OR2_X1 U7387 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  NAND2_X1 U7388 ( .A1(n6374), .A2(n6373), .ZN(n6446) );
  INV_X1 U7389 ( .A(n6446), .ZN(n6376) );
  AOI22_X1 U7390 ( .A1(n6376), .A2(n6386), .B1(n6385), .B2(n6375), .ZN(n6377)
         );
  OAI211_X1 U7391 ( .C1(n6390), .C2(n6379), .A(n6378), .B(n6377), .ZN(U2982)
         );
  AOI22_X1 U7392 ( .A1(n6476), .A2(REIP_REG_2__SCAN_IN), .B1(n6380), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6388) );
  XNOR2_X1 U7393 ( .A(n6381), .B(n6477), .ZN(n6383) );
  XNOR2_X1 U7394 ( .A(n6383), .B(n6382), .ZN(n6473) );
  AOI22_X1 U7395 ( .A1(n6473), .A2(n6386), .B1(n6385), .B2(n6384), .ZN(n6387)
         );
  OAI211_X1 U7396 ( .C1(n6390), .C2(n6389), .A(n6388), .B(n6387), .ZN(U2984)
         );
  AOI22_X1 U7397 ( .A1(n6467), .A2(n6391), .B1(n6476), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n6395) );
  AOI22_X1 U7398 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6393), .B1(n6392), .B2(n3686), .ZN(n6394) );
  OAI211_X1 U7399 ( .C1(n6396), .C2(n6455), .A(n6395), .B(n6394), .ZN(U3007)
         );
  NOR2_X1 U7400 ( .A1(n6397), .A2(n6443), .ZN(n6426) );
  NAND2_X1 U7401 ( .A1(n6402), .A2(n6426), .ZN(n6414) );
  AOI22_X1 U7402 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n3685), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6398), .ZN(n6407) );
  INV_X1 U7403 ( .A(n6399), .ZN(n6400) );
  AOI21_X1 U7404 ( .B1(n6467), .B2(n6401), .A(n6400), .ZN(n6406) );
  OAI21_X1 U7405 ( .B1(n6403), .B2(n6402), .A(n6431), .ZN(n6410) );
  AOI22_X1 U7406 ( .A1(n6404), .A2(n6474), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6410), .ZN(n6405) );
  OAI211_X1 U7407 ( .C1(n6414), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3008)
         );
  AOI21_X1 U7408 ( .B1(n6467), .B2(n6409), .A(n6408), .ZN(n6413) );
  AOI22_X1 U7409 ( .A1(n6411), .A2(n6474), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6410), .ZN(n6412) );
  OAI211_X1 U7410 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6414), .A(n6413), 
        .B(n6412), .ZN(U3009) );
  OAI222_X1 U7411 ( .A1(n6416), .A2(n6448), .B1(n6454), .B2(n6687), .C1(n6455), 
        .C2(n6415), .ZN(n6417) );
  INV_X1 U7412 ( .A(n6417), .ZN(n6420) );
  OAI211_X1 U7413 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6426), .B(n6418), .ZN(n6419) );
  OAI211_X1 U7414 ( .C1(n6431), .C2(n6421), .A(n6420), .B(n6419), .ZN(U3010)
         );
  INV_X1 U7415 ( .A(n6422), .ZN(n6423) );
  AOI21_X1 U7416 ( .B1(n6467), .B2(n6424), .A(n6423), .ZN(n6429) );
  INV_X1 U7417 ( .A(n6425), .ZN(n6427) );
  AOI22_X1 U7418 ( .A1(n6427), .A2(n6474), .B1(n6426), .B2(n6430), .ZN(n6428)
         );
  OAI211_X1 U7419 ( .C1(n6431), .C2(n6430), .A(n6429), .B(n6428), .ZN(U3011)
         );
  AOI21_X1 U7420 ( .B1(n6433), .B2(n6432), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6441) );
  AOI21_X1 U7421 ( .B1(n6467), .B2(n6435), .A(n6434), .ZN(n6440) );
  NOR2_X1 U7422 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6436), .ZN(n6437)
         );
  AOI22_X1 U7423 ( .A1(n6438), .A2(n6474), .B1(n6437), .B2(n6478), .ZN(n6439)
         );
  OAI211_X1 U7424 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n6439), .ZN(U3013)
         );
  NOR2_X1 U7425 ( .A1(n6471), .A2(n6444), .ZN(n6466) );
  NOR2_X1 U7426 ( .A1(n6466), .A2(n6469), .ZN(n6462) );
  INV_X1 U7427 ( .A(n6443), .ZN(n6445) );
  NAND2_X1 U7428 ( .A1(n6445), .A2(n6444), .ZN(n6464) );
  AOI221_X1 U7429 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n6463), .C2(n6453), .A(n6464), 
        .ZN(n6451) );
  NOR2_X1 U7430 ( .A1(n6446), .A2(n6455), .ZN(n6450) );
  OAI22_X1 U7431 ( .A1(n6448), .A2(n6447), .B1(n6684), .B2(n6454), .ZN(n6449)
         );
  NOR3_X1 U7432 ( .A1(n6451), .A2(n6450), .A3(n6449), .ZN(n6452) );
  OAI21_X1 U7433 ( .B1(n6462), .B2(n6453), .A(n6452), .ZN(U3014) );
  NOR2_X1 U7434 ( .A1(n6454), .A2(n4775), .ZN(n6459) );
  NOR3_X1 U7435 ( .A1(n6457), .A2(n6456), .A3(n6455), .ZN(n6458) );
  AOI211_X1 U7436 ( .C1(n6467), .C2(n6460), .A(n6459), .B(n6458), .ZN(n6461)
         );
  OAI221_X1 U7437 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6464), .C1(n6463), .C2(n6462), .A(n6461), .ZN(U3015) );
  INV_X1 U7438 ( .A(n6465), .ZN(n6468) );
  AOI21_X1 U7439 ( .B1(n6468), .B2(n6467), .A(n6466), .ZN(n6482) );
  INV_X1 U7440 ( .A(n6469), .ZN(n6470) );
  OAI21_X1 U7441 ( .B1(n6472), .B2(n6471), .A(n6470), .ZN(n6475) );
  AOI22_X1 U7442 ( .A1(n6475), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6474), 
        .B2(n6473), .ZN(n6481) );
  NAND2_X1 U7443 ( .A1(n6476), .A2(REIP_REG_2__SCAN_IN), .ZN(n6480) );
  NAND3_X1 U7444 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6478), .A3(n6477), 
        .ZN(n6479) );
  NAND4_X1 U7445 ( .A1(n6482), .A2(n6481), .A3(n6480), .A4(n6479), .ZN(U3016)
         );
  INV_X1 U7446 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U7447 ( .A1(n6628), .A2(n6483), .ZN(U3019) );
  OR2_X1 U7448 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6484), .ZN(n6545)
         );
  NAND2_X1 U7449 ( .A1(n6486), .A2(n6485), .ZN(n6491) );
  NAND3_X1 U7450 ( .A1(n6489), .A2(n6488), .A3(n6487), .ZN(n6490) );
  OAI22_X1 U7451 ( .A1(n6493), .A2(n6545), .B1(n6544), .B2(n6492), .ZN(n6494)
         );
  INV_X1 U7452 ( .A(n6494), .ZN(n6506) );
  NOR3_X1 U7453 ( .A1(n6547), .A2(n6497), .A3(n6496), .ZN(n6500) );
  OAI21_X1 U7454 ( .B1(n6500), .B2(n6499), .A(n6498), .ZN(n6503) );
  AOI21_X1 U7455 ( .B1(n6545), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6501) );
  NAND3_X1 U7456 ( .A1(n6503), .A2(n6502), .A3(n6501), .ZN(n6549) );
  AOI22_X1 U7457 ( .A1(n6549), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6504), 
        .B2(n6547), .ZN(n6505) );
  OAI211_X1 U7458 ( .C1(n6507), .C2(n6585), .A(n6506), .B(n6505), .ZN(U3068)
         );
  OAI22_X1 U7459 ( .A1(n6552), .A2(n6545), .B1(n6544), .B2(n6508), .ZN(n6509)
         );
  INV_X1 U7460 ( .A(n6509), .ZN(n6512) );
  AOI22_X1 U7461 ( .A1(n6549), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6510), 
        .B2(n6547), .ZN(n6511) );
  OAI211_X1 U7462 ( .C1(n6513), .C2(n6585), .A(n6512), .B(n6511), .ZN(U3069)
         );
  OAI22_X1 U7463 ( .A1(n6515), .A2(n6545), .B1(n6544), .B2(n6514), .ZN(n6516)
         );
  INV_X1 U7464 ( .A(n6516), .ZN(n6519) );
  AOI22_X1 U7465 ( .A1(n6549), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6517), 
        .B2(n6547), .ZN(n6518) );
  OAI211_X1 U7466 ( .C1(n6520), .C2(n6585), .A(n6519), .B(n6518), .ZN(U3070)
         );
  OAI22_X1 U7467 ( .A1(n6586), .A2(n6545), .B1(n6544), .B2(n6521), .ZN(n6522)
         );
  INV_X1 U7468 ( .A(n6522), .ZN(n6525) );
  AOI22_X1 U7469 ( .A1(n6549), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6523), 
        .B2(n6547), .ZN(n6524) );
  OAI211_X1 U7470 ( .C1(n6587), .C2(n6585), .A(n6525), .B(n6524), .ZN(U3071)
         );
  OAI22_X1 U7471 ( .A1(n6563), .A2(n6545), .B1(n6544), .B2(n6526), .ZN(n6527)
         );
  INV_X1 U7472 ( .A(n6527), .ZN(n6530) );
  AOI22_X1 U7473 ( .A1(n6549), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6528), 
        .B2(n6547), .ZN(n6529) );
  OAI211_X1 U7474 ( .C1(n6531), .C2(n6585), .A(n6530), .B(n6529), .ZN(U3072)
         );
  OAI22_X1 U7475 ( .A1(n6593), .A2(n6545), .B1(n6544), .B2(n6532), .ZN(n6533)
         );
  INV_X1 U7476 ( .A(n6533), .ZN(n6536) );
  AOI22_X1 U7477 ( .A1(n6549), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6534), 
        .B2(n6547), .ZN(n6535) );
  OAI211_X1 U7478 ( .C1(n6594), .C2(n6585), .A(n6536), .B(n6535), .ZN(U3073)
         );
  OAI22_X1 U7479 ( .A1(n6570), .A2(n6545), .B1(n6544), .B2(n6537), .ZN(n6538)
         );
  INV_X1 U7480 ( .A(n6538), .ZN(n6541) );
  AOI22_X1 U7481 ( .A1(n6549), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6539), 
        .B2(n6547), .ZN(n6540) );
  OAI211_X1 U7482 ( .C1(n6542), .C2(n6585), .A(n6541), .B(n6540), .ZN(U3074)
         );
  OAI22_X1 U7483 ( .A1(n6601), .A2(n6545), .B1(n6544), .B2(n6543), .ZN(n6546)
         );
  INV_X1 U7484 ( .A(n6546), .ZN(n6551) );
  AOI22_X1 U7485 ( .A1(n6549), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6548), 
        .B2(n6547), .ZN(n6550) );
  OAI211_X1 U7486 ( .C1(n6602), .C2(n6585), .A(n6551), .B(n6550), .ZN(U3075)
         );
  NOR2_X1 U7487 ( .A1(n6552), .A2(n6577), .ZN(n6553) );
  AOI21_X1 U7488 ( .B1(n6580), .B2(n6554), .A(n6553), .ZN(n6557) );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6582), .B1(n6555), 
        .B2(n6581), .ZN(n6556) );
  OAI211_X1 U7490 ( .C1(n6558), .C2(n6585), .A(n6557), .B(n6556), .ZN(U3077)
         );
  NOR2_X1 U7491 ( .A1(n6586), .A2(n6577), .ZN(n6559) );
  AOI21_X1 U7492 ( .B1(n6580), .B2(n6560), .A(n6559), .ZN(n6562) );
  AOI22_X1 U7493 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6582), .B1(n6589), 
        .B2(n6581), .ZN(n6561) );
  OAI211_X1 U7494 ( .C1(n6592), .C2(n6585), .A(n6562), .B(n6561), .ZN(U3079)
         );
  NOR2_X1 U7495 ( .A1(n6563), .A2(n6577), .ZN(n6564) );
  AOI21_X1 U7496 ( .B1(n6580), .B2(n6565), .A(n6564), .ZN(n6568) );
  AOI22_X1 U7497 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6582), .B1(n6566), 
        .B2(n6581), .ZN(n6567) );
  OAI211_X1 U7498 ( .C1(n6569), .C2(n6585), .A(n6568), .B(n6567), .ZN(U3080)
         );
  NOR2_X1 U7499 ( .A1(n6570), .A2(n6577), .ZN(n6571) );
  AOI21_X1 U7500 ( .B1(n6580), .B2(n6572), .A(n6571), .ZN(n6575) );
  AOI22_X1 U7501 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6582), .B1(n6573), 
        .B2(n6581), .ZN(n6574) );
  OAI211_X1 U7502 ( .C1(n6576), .C2(n6585), .A(n6575), .B(n6574), .ZN(U3082)
         );
  NOR2_X1 U7503 ( .A1(n6601), .A2(n6577), .ZN(n6578) );
  AOI21_X1 U7504 ( .B1(n6580), .B2(n6579), .A(n6578), .ZN(n6584) );
  AOI22_X1 U7505 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6582), .B1(n6606), 
        .B2(n6581), .ZN(n6583) );
  OAI211_X1 U7506 ( .C1(n6611), .C2(n6585), .A(n6584), .B(n6583), .ZN(U3083)
         );
  OAI22_X1 U7507 ( .A1(n6603), .A2(n6587), .B1(n6586), .B2(n6600), .ZN(n6588)
         );
  INV_X1 U7508 ( .A(n6588), .ZN(n6591) );
  AOI22_X1 U7509 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6607), .B1(n6589), 
        .B2(n6605), .ZN(n6590) );
  OAI211_X1 U7510 ( .C1(n6592), .C2(n6610), .A(n6591), .B(n6590), .ZN(U3111)
         );
  OAI22_X1 U7511 ( .A1(n6603), .A2(n6594), .B1(n6593), .B2(n6600), .ZN(n6595)
         );
  INV_X1 U7512 ( .A(n6595), .ZN(n6598) );
  AOI22_X1 U7513 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6607), .B1(n6596), 
        .B2(n6605), .ZN(n6597) );
  OAI211_X1 U7514 ( .C1(n6599), .C2(n6610), .A(n6598), .B(n6597), .ZN(U3113)
         );
  OAI22_X1 U7515 ( .A1(n6603), .A2(n6602), .B1(n6601), .B2(n6600), .ZN(n6604)
         );
  INV_X1 U7516 ( .A(n6604), .ZN(n6609) );
  AOI22_X1 U7517 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6607), .B1(n6606), 
        .B2(n6605), .ZN(n6608) );
  OAI211_X1 U7518 ( .C1(n6611), .C2(n6610), .A(n6609), .B(n6608), .ZN(U3115)
         );
  INV_X1 U7519 ( .A(n6612), .ZN(n6615) );
  NOR3_X1 U7520 ( .A1(n6615), .A2(n6614), .A3(n6613), .ZN(n6621) );
  INV_X1 U7521 ( .A(n6621), .ZN(n6619) );
  OAI211_X1 U7522 ( .C1(n6619), .C2(n6618), .A(n6617), .B(n6616), .ZN(n6620)
         );
  OAI21_X1 U7523 ( .B1(n6621), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6620), 
        .ZN(n6622) );
  AOI222_X1 U7524 ( .A1(n6624), .A2(n6623), .B1(n6624), .B2(n6622), .C1(n6623), 
        .C2(n6622), .ZN(n6627) );
  OR2_X1 U7525 ( .A1(n6627), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6626)
         );
  NAND2_X1 U7526 ( .A1(n6626), .A2(n6625), .ZN(n6630) );
  NAND2_X1 U7527 ( .A1(n6627), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6629) );
  NAND3_X1 U7528 ( .A1(n6630), .A2(n6629), .A3(n6628), .ZN(n6639) );
  OAI21_X1 U7529 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6631), 
        .ZN(n6632) );
  NAND4_X1 U7530 ( .A1(n6635), .A2(n6634), .A3(n6633), .A4(n6632), .ZN(n6636)
         );
  NOR2_X1 U7531 ( .A1(n6637), .A2(n6636), .ZN(n6638) );
  NOR2_X1 U7532 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6719), .ZN(n6667) );
  NAND2_X1 U7533 ( .A1(n6656), .A2(n6657), .ZN(n6641) );
  NAND2_X1 U7534 ( .A1(READY_N), .A2(n6720), .ZN(n6640) );
  NAND2_X1 U7535 ( .A1(n6641), .A2(n6640), .ZN(n6645) );
  OR2_X1 U7536 ( .A1(n6643), .A2(n6642), .ZN(n6644) );
  NOR2_X1 U7537 ( .A1(n6667), .A2(n6710), .ZN(n6652) );
  OAI21_X1 U7538 ( .B1(n6663), .B2(n6646), .A(n6659), .ZN(n6647) );
  OR2_X1 U7539 ( .A1(n6710), .A2(n6647), .ZN(n6651) );
  INV_X1 U7540 ( .A(n6662), .ZN(n6708) );
  AOI21_X1 U7541 ( .B1(n6649), .B2(n6708), .A(n6648), .ZN(n6650) );
  OAI211_X1 U7542 ( .C1(n6652), .C2(n6659), .A(n6651), .B(n6650), .ZN(n6653)
         );
  INV_X1 U7543 ( .A(n6653), .ZN(n6654) );
  OAI21_X1 U7544 ( .B1(n6656), .B2(n6655), .A(n6654), .ZN(U3148) );
  AOI21_X1 U7545 ( .B1(n6658), .B2(n6719), .A(n6657), .ZN(n6661) );
  NAND2_X1 U7546 ( .A1(n6659), .A2(n4510), .ZN(n6664) );
  OAI211_X1 U7547 ( .C1(n6710), .C2(n6667), .A(STATE2_REG_1__SCAN_IN), .B(
        n6664), .ZN(n6660) );
  OAI211_X1 U7548 ( .C1(n6710), .C2(n6661), .A(n3197), .B(n6660), .ZN(U3149)
         );
  NAND3_X1 U7549 ( .A1(n6664), .A2(n6663), .A3(n6662), .ZN(n6666) );
  OAI21_X1 U7550 ( .B1(n6667), .B2(n6666), .A(n6665), .ZN(U3150) );
  AND2_X1 U7551 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6703), .ZN(U3151) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6703), .ZN(U3152) );
  AND2_X1 U7553 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6703), .ZN(U3153) );
  AND2_X1 U7554 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6703), .ZN(U3154) );
  AND2_X1 U7555 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6703), .ZN(U3155) );
  AND2_X1 U7556 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6703), .ZN(U3156) );
  AND2_X1 U7557 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6703), .ZN(U3157) );
  AND2_X1 U7558 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6703), .ZN(U3158) );
  INV_X1 U7559 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6971) );
  NOR2_X1 U7560 ( .A1(n6707), .A2(n6971), .ZN(U3159) );
  INV_X1 U7561 ( .A(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6942) );
  NOR2_X1 U7562 ( .A1(n6707), .A2(n6942), .ZN(U3160) );
  AND2_X1 U7563 ( .A1(n6703), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  INV_X1 U7564 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6805) );
  NOR2_X1 U7565 ( .A1(n6707), .A2(n6805), .ZN(U3162) );
  INV_X1 U7566 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6827) );
  NOR2_X1 U7567 ( .A1(n6707), .A2(n6827), .ZN(U3163) );
  AND2_X1 U7568 ( .A1(n6703), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  INV_X1 U7569 ( .A(DATAWIDTH_REG_17__SCAN_IN), .ZN(n7081) );
  NOR2_X1 U7570 ( .A1(n6707), .A2(n7081), .ZN(U3165) );
  INV_X1 U7571 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6802) );
  NOR2_X1 U7572 ( .A1(n6707), .A2(n6802), .ZN(U3166) );
  INV_X1 U7573 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6875) );
  NOR2_X1 U7574 ( .A1(n6707), .A2(n6875), .ZN(U3167) );
  INV_X1 U7575 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6825) );
  NOR2_X1 U7576 ( .A1(n6707), .A2(n6825), .ZN(U3168) );
  INV_X1 U7577 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6816) );
  NOR2_X1 U7578 ( .A1(n6707), .A2(n6816), .ZN(U3169) );
  AND2_X1 U7579 ( .A1(n6703), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U7580 ( .A1(n6703), .A2(DATAWIDTH_REG_11__SCAN_IN), .ZN(U3171) );
  AND2_X1 U7581 ( .A1(n6703), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  INV_X1 U7582 ( .A(DATAWIDTH_REG_9__SCAN_IN), .ZN(n6845) );
  NOR2_X1 U7583 ( .A1(n6707), .A2(n6845), .ZN(U3173) );
  INV_X1 U7584 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6994) );
  NOR2_X1 U7585 ( .A1(n6707), .A2(n6994), .ZN(U3174) );
  INV_X1 U7586 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6858) );
  NOR2_X1 U7587 ( .A1(n6707), .A2(n6858), .ZN(U3175) );
  AND2_X1 U7588 ( .A1(n6703), .A2(DATAWIDTH_REG_6__SCAN_IN), .ZN(U3176) );
  AND2_X1 U7589 ( .A1(n6703), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  AND2_X1 U7590 ( .A1(n6703), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  INV_X1 U7591 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6807) );
  NOR2_X1 U7592 ( .A1(n6707), .A2(n6807), .ZN(U3179) );
  INV_X1 U7593 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6840) );
  NOR2_X1 U7594 ( .A1(n6707), .A2(n6840), .ZN(U3180) );
  INV_X1 U7595 ( .A(n6681), .ZN(n6669) );
  AOI22_X1 U7596 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6682) );
  INV_X1 U7597 ( .A(HOLD), .ZN(n6877) );
  NOR2_X1 U7598 ( .A1(n7000), .A2(n6877), .ZN(n6670) );
  INV_X1 U7599 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6955) );
  OAI21_X1 U7600 ( .B1(n6670), .B2(n6955), .A(n7128), .ZN(n6668) );
  OAI221_X1 U7601 ( .B1(n6814), .B2(NA_N), .C1(n6814), .C2(n7000), .A(n6677), 
        .ZN(n6675) );
  OAI211_X1 U7602 ( .C1(n6669), .C2(n6682), .A(n6668), .B(n6675), .ZN(U3181)
         );
  NOR2_X1 U7603 ( .A1(n6677), .A2(n6955), .ZN(n6671) );
  OAI22_X1 U7604 ( .A1(n6671), .A2(n6670), .B1(n6814), .B2(n6877), .ZN(n6672)
         );
  OAI211_X1 U7605 ( .C1(n7000), .C2(n6719), .A(n6673), .B(n6672), .ZN(U3182)
         );
  NOR2_X1 U7606 ( .A1(n6719), .A2(NA_N), .ZN(n6678) );
  INV_X1 U7607 ( .A(n6678), .ZN(n6674) );
  OAI221_X1 U7608 ( .B1(REQUESTPENDING_REG_SCAN_IN), .B2(STATE_REG_1__SCAN_IN), 
        .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6674), .A(n6814), .ZN(n6676) );
  OAI211_X1 U7609 ( .C1(n6677), .C2(HOLD), .A(n6676), .B(n6675), .ZN(n6680) );
  NAND4_X1 U7610 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .A3(
        REQUESTPENDING_REG_SCAN_IN), .A4(n6678), .ZN(n6679) );
  OAI211_X1 U7611 ( .C1(n6682), .C2(n6681), .A(n6680), .B(n6679), .ZN(U3183)
         );
  INV_X1 U7612 ( .A(ADDRESS_REG_0__SCAN_IN), .ZN(n6683) );
  INV_X2 U7613 ( .A(n7128), .ZN(n7129) );
  OAI222_X1 U7614 ( .A1(n6694), .A2(n6280), .B1(n6683), .B2(n7129), .C1(n5011), 
        .C2(n6696), .ZN(U3184) );
  INV_X1 U7615 ( .A(ADDRESS_REG_1__SCAN_IN), .ZN(n6984) );
  OAI222_X1 U7616 ( .A1(n6696), .A2(n6280), .B1(n6984), .B2(n7129), .C1(n4775), 
        .C2(n6694), .ZN(U3185) );
  INV_X1 U7617 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6974) );
  OAI222_X1 U7618 ( .A1(n6696), .A2(n4775), .B1(n6974), .B2(n7129), .C1(n6684), 
        .C2(n6694), .ZN(U3186) );
  INV_X1 U7619 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U7620 ( .A1(n6696), .A2(n6684), .B1(n6831), .B2(n7129), .C1(n4892), 
        .C2(n6694), .ZN(U3187) );
  INV_X1 U7621 ( .A(ADDRESS_REG_4__SCAN_IN), .ZN(n6889) );
  OAI222_X1 U7622 ( .A1(n6696), .A2(n4892), .B1(n6889), .B2(n7129), .C1(n6685), 
        .C2(n6694), .ZN(U3188) );
  INV_X1 U7623 ( .A(ADDRESS_REG_5__SCAN_IN), .ZN(n6846) );
  OAI222_X1 U7624 ( .A1(n6696), .A2(n6685), .B1(n6846), .B2(n7129), .C1(n6686), 
        .C2(n6694), .ZN(U3189) );
  INV_X1 U7625 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n7003) );
  OAI222_X1 U7626 ( .A1(n6696), .A2(n6686), .B1(n7003), .B2(n7129), .C1(n6687), 
        .C2(n6694), .ZN(U3190) );
  INV_X1 U7627 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n7057) );
  OAI222_X1 U7628 ( .A1(n6696), .A2(n6687), .B1(n7057), .B2(n7129), .C1(n5414), 
        .C2(n6694), .ZN(U3191) );
  INV_X1 U7629 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n7124) );
  OAI222_X1 U7630 ( .A1(n6696), .A2(n5414), .B1(n7124), .B2(n7129), .C1(n6688), 
        .C2(n6694), .ZN(U3192) );
  INV_X1 U7631 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n7052) );
  OAI222_X1 U7632 ( .A1(n6696), .A2(n6688), .B1(n7052), .B2(n6700), .C1(n6689), 
        .C2(n6694), .ZN(U3193) );
  INV_X1 U7633 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6874) );
  OAI222_X1 U7634 ( .A1(n6694), .A2(n5450), .B1(n6874), .B2(n7129), .C1(n6689), 
        .C2(n6696), .ZN(U3194) );
  INV_X1 U7635 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6818) );
  OAI222_X1 U7636 ( .A1(n6696), .A2(n5450), .B1(n6818), .B2(n6700), .C1(n6690), 
        .C2(n6694), .ZN(U3195) );
  INV_X1 U7637 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n7093) );
  OAI222_X1 U7638 ( .A1(n6696), .A2(n6690), .B1(n7093), .B2(n7129), .C1(n5835), 
        .C2(n6694), .ZN(U3196) );
  INV_X1 U7639 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6959) );
  OAI222_X1 U7640 ( .A1(n6696), .A2(n5835), .B1(n6959), .B2(n7129), .C1(n6691), 
        .C2(n6694), .ZN(U3197) );
  INV_X1 U7641 ( .A(ADDRESS_REG_14__SCAN_IN), .ZN(n6895) );
  OAI222_X1 U7642 ( .A1(n6696), .A2(n6691), .B1(n6895), .B2(n6700), .C1(n6985), 
        .C2(n6694), .ZN(U3198) );
  INV_X1 U7643 ( .A(ADDRESS_REG_15__SCAN_IN), .ZN(n6692) );
  OAI222_X1 U7644 ( .A1(n6696), .A2(n6985), .B1(n6692), .B2(n6700), .C1(n6755), 
        .C2(n6694), .ZN(U3199) );
  INV_X1 U7645 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6968) );
  OAI222_X1 U7646 ( .A1(n6694), .A2(n6899), .B1(n6968), .B2(n6700), .C1(n6755), 
        .C2(n6696), .ZN(U3200) );
  INV_X1 U7647 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6991) );
  INV_X1 U7648 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6693) );
  OAI222_X1 U7649 ( .A1(n6694), .A2(n6991), .B1(n6693), .B2(n6700), .C1(n6899), 
        .C2(n6696), .ZN(U3201) );
  INV_X1 U7650 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6975) );
  OAI222_X1 U7651 ( .A1(n6696), .A2(n6991), .B1(n6975), .B2(n6700), .C1(n5804), 
        .C2(n6694), .ZN(U3202) );
  INV_X1 U7652 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6813) );
  OAI222_X1 U7653 ( .A1(n6696), .A2(n5804), .B1(n6813), .B2(n7129), .C1(n6868), 
        .C2(n6694), .ZN(U3203) );
  INV_X1 U7654 ( .A(ADDRESS_REG_20__SCAN_IN), .ZN(n7054) );
  OAI222_X1 U7655 ( .A1(n6696), .A2(n6868), .B1(n7054), .B2(n6700), .C1(n7068), 
        .C2(n6694), .ZN(U3204) );
  INV_X1 U7656 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6869) );
  OAI222_X1 U7657 ( .A1(n6696), .A2(n7068), .B1(n6869), .B2(n7129), .C1(n6695), 
        .C2(n6694), .ZN(U3205) );
  INV_X1 U7658 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n7102) );
  OAI222_X1 U7659 ( .A1(n6696), .A2(n6695), .B1(n7102), .B2(n6700), .C1(n6697), 
        .C2(n6694), .ZN(U3206) );
  INV_X1 U7660 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n7070) );
  OAI222_X1 U7661 ( .A1(n6694), .A2(n5765), .B1(n7070), .B2(n7129), .C1(n6697), 
        .C2(n6696), .ZN(U3207) );
  INV_X1 U7662 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n7094) );
  INV_X1 U7663 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6886) );
  OAI222_X1 U7664 ( .A1(n6696), .A2(n5765), .B1(n7094), .B2(n7129), .C1(n6886), 
        .C2(n6694), .ZN(U3208) );
  INV_X1 U7665 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6698) );
  OAI222_X1 U7666 ( .A1(n6696), .A2(n6886), .B1(n6698), .B2(n7129), .C1(n7087), 
        .C2(n6694), .ZN(U3209) );
  INV_X1 U7667 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6699) );
  OAI222_X1 U7668 ( .A1(n6696), .A2(n7087), .B1(n6699), .B2(n7129), .C1(n6871), 
        .C2(n6694), .ZN(U3210) );
  INV_X1 U7669 ( .A(ADDRESS_REG_27__SCAN_IN), .ZN(n7080) );
  OAI222_X1 U7670 ( .A1(n6696), .A2(n6871), .B1(n7080), .B2(n7129), .C1(n6860), 
        .C2(n6694), .ZN(U3211) );
  INV_X1 U7671 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6952) );
  OAI222_X1 U7672 ( .A1(n6696), .A2(n6860), .B1(n6952), .B2(n6700), .C1(n6861), 
        .C2(n6694), .ZN(U3212) );
  INV_X1 U7673 ( .A(ADDRESS_REG_29__SCAN_IN), .ZN(n6701) );
  OAI222_X1 U7674 ( .A1(n6694), .A2(n6872), .B1(n6701), .B2(n7129), .C1(n6861), 
        .C2(n6696), .ZN(U3213) );
  INV_X1 U7675 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n7099) );
  INV_X1 U7676 ( .A(BE_N_REG_2__SCAN_IN), .ZN(n7004) );
  AOI22_X1 U7677 ( .A1(n7129), .A2(n7099), .B1(n7004), .B2(n7128), .ZN(U3446)
         );
  INV_X1 U7678 ( .A(BE_N_REG_1__SCAN_IN), .ZN(n7097) );
  AOI22_X1 U7679 ( .A1(n7129), .A2(n7067), .B1(n7097), .B2(n7128), .ZN(U3447)
         );
  INV_X1 U7680 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n7001) );
  INV_X1 U7681 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U7682 ( .A1(n7129), .A2(n7001), .B1(n6838), .B2(n7128), .ZN(U3448)
         );
  INV_X1 U7683 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6704) );
  INV_X1 U7684 ( .A(n6705), .ZN(n6702) );
  AOI21_X1 U7685 ( .B1(n6704), .B2(n6703), .A(n6702), .ZN(U3451) );
  OAI21_X1 U7686 ( .B1(n6707), .B2(n6706), .A(n6705), .ZN(U3452) );
  AOI211_X1 U7687 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6710), .A(n6709), .B(
        n6708), .ZN(n6711) );
  INV_X1 U7688 ( .A(n6711), .ZN(U3453) );
  AOI211_X1 U7689 ( .C1(REIP_REG_0__SCAN_IN), .C2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(REIP_REG_1__SCAN_IN), .B(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6712) );
  AOI21_X1 U7690 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6712), .ZN(n6713) );
  AOI22_X1 U7691 ( .A1(n6716), .A2(n6713), .B1(n7099), .B2(n6714), .ZN(U3468)
         );
  NOR2_X1 U7692 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6715) );
  AOI22_X1 U7693 ( .A1(n6716), .A2(n6715), .B1(n7001), .B2(n6714), .ZN(U3469)
         );
  INV_X1 U7694 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6953) );
  AOI22_X1 U7695 ( .A1(n7129), .A2(READREQUEST_REG_SCAN_IN), .B1(n6953), .B2(
        n7128), .ZN(U3470) );
  AOI211_X1 U7696 ( .C1(n6720), .C2(n6719), .A(n6718), .B(n6717), .ZN(n6727)
         );
  OAI211_X1 U7697 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6722), .A(n6721), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6724) );
  AOI21_X1 U7698 ( .B1(n6724), .B2(STATE2_REG_0__SCAN_IN), .A(n6723), .ZN(
        n6726) );
  NAND2_X1 U7699 ( .A1(n6727), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6725) );
  OAI21_X1 U7700 ( .B1(n6727), .B2(n6726), .A(n6725), .ZN(U3472) );
  INV_X1 U7701 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7055) );
  AOI22_X1 U7702 ( .A1(n7129), .A2(n6832), .B1(n7055), .B2(n7128), .ZN(U3473)
         );
  OAI22_X1 U7703 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(keyinput_g100), .ZN(n6728) );
  AOI221_X1 U7704 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(keyinput_g100), .C2(
        ADDRESS_REG_0__SCAN_IN), .A(n6728), .ZN(n6735) );
  OAI22_X1 U7705 ( .A1(REIP_REG_23__SCAN_IN), .A2(keyinput_g59), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_g39), .ZN(n6729) );
  AOI221_X1 U7706 ( .B1(REIP_REG_23__SCAN_IN), .B2(keyinput_g59), .C1(
        keyinput_g39), .C2(CODEFETCH_REG_SCAN_IN), .A(n6729), .ZN(n6734) );
  OAI22_X1 U7707 ( .A1(ADDRESS_REG_13__SCAN_IN), .A2(keyinput_g87), .B1(
        keyinput_g49), .B2(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6730) );
  AOI221_X1 U7708 ( .B1(ADDRESS_REG_13__SCAN_IN), .B2(keyinput_g87), .C1(
        BYTEENABLE_REG_2__SCAN_IN), .C2(keyinput_g49), .A(n6730), .ZN(n6733)
         );
  OAI22_X1 U7709 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(keyinput_g11), .B2(
        DATAI_20_), .ZN(n6731) );
  AOI221_X1 U7710 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(DATAI_20_), .C2(
        keyinput_g11), .A(n6731), .ZN(n6732) );
  NAND4_X1 U7711 ( .A1(n6735), .A2(n6734), .A3(n6733), .A4(n6732), .ZN(n6765)
         );
  OAI22_X1 U7712 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(keyinput_g122), .B1(
        keyinput_g50), .B2(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6736) );
  AOI221_X1 U7713 ( .B1(DATAWIDTH_REG_18__SCAN_IN), .B2(keyinput_g122), .C1(
        BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_g50), .A(n6736), .ZN(n6743)
         );
  OAI22_X1 U7714 ( .A1(ADDRESS_REG_15__SCAN_IN), .A2(keyinput_g85), .B1(
        keyinput_g105), .B2(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6737) );
  AOI221_X1 U7715 ( .B1(ADDRESS_REG_15__SCAN_IN), .B2(keyinput_g85), .C1(
        DATAWIDTH_REG_1__SCAN_IN), .C2(keyinput_g105), .A(n6737), .ZN(n6742)
         );
  OAI22_X1 U7716 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(keyinput_g33), .B2(
        NA_N), .ZN(n6738) );
  AOI221_X1 U7717 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(NA_N), .C2(
        keyinput_g33), .A(n6738), .ZN(n6741) );
  OAI22_X1 U7718 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(keyinput_g110), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(keyinput_g80), .ZN(n6739) );
  AOI221_X1 U7719 ( .B1(DATAWIDTH_REG_6__SCAN_IN), .B2(keyinput_g110), .C1(
        keyinput_g80), .C2(ADDRESS_REG_20__SCAN_IN), .A(n6739), .ZN(n6740) );
  NAND4_X1 U7720 ( .A1(n6743), .A2(n6742), .A3(n6741), .A4(n6740), .ZN(n6764)
         );
  OAI22_X1 U7721 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_g45), .B1(keyinput_g69), .B2(BE_N_REG_1__SCAN_IN), .ZN(n6744) );
  AOI221_X1 U7722 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        BE_N_REG_1__SCAN_IN), .C2(keyinput_g69), .A(n6744), .ZN(n6751) );
  OAI22_X1 U7723 ( .A1(ADDRESS_REG_26__SCAN_IN), .A2(keyinput_g74), .B1(
        keyinput_g99), .B2(ADDRESS_REG_1__SCAN_IN), .ZN(n6745) );
  AOI221_X1 U7724 ( .B1(ADDRESS_REG_26__SCAN_IN), .B2(keyinput_g74), .C1(
        ADDRESS_REG_1__SCAN_IN), .C2(keyinput_g99), .A(n6745), .ZN(n6750) );
  OAI22_X1 U7725 ( .A1(STATE_REG_0__SCAN_IN), .A2(keyinput_g103), .B1(
        DATAI_14_), .B2(keyinput_g17), .ZN(n6746) );
  AOI221_X1 U7726 ( .B1(STATE_REG_0__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g17), .C2(DATAI_14_), .A(n6746), .ZN(n6749) );
  OAI22_X1 U7727 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(keyinput_g114), .B1(
        keyinput_g121), .B2(DATAWIDTH_REG_17__SCAN_IN), .ZN(n6747) );
  AOI221_X1 U7728 ( .B1(DATAWIDTH_REG_10__SCAN_IN), .B2(keyinput_g114), .C1(
        DATAWIDTH_REG_17__SCAN_IN), .C2(keyinput_g121), .A(n6747), .ZN(n6748)
         );
  NAND4_X1 U7729 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6763)
         );
  AOI22_X1 U7730 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput_g94), .B1(
        DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput_g108), .ZN(n6752) );
  OAI221_X1 U7731 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput_g94), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput_g108), .A(n6752), .ZN(n6761)
         );
  INV_X1 U7732 ( .A(DATAI_31_), .ZN(n7071) );
  AOI22_X1 U7733 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(keyinput_g115), .B1(
        n7071), .B2(keyinput_g0), .ZN(n6753) );
  OAI221_X1 U7734 ( .B1(DATAWIDTH_REG_11__SCAN_IN), .B2(keyinput_g115), .C1(
        n7071), .C2(keyinput_g0), .A(n6753), .ZN(n6760) );
  AOI22_X1 U7735 ( .A1(n7093), .A2(keyinput_g88), .B1(n6755), .B2(keyinput_g65), .ZN(n6754) );
  OAI221_X1 U7736 ( .B1(n7093), .B2(keyinput_g88), .C1(n6755), .C2(
        keyinput_g65), .A(n6754), .ZN(n6759) );
  AOI22_X1 U7737 ( .A1(n6757), .A2(keyinput_g20), .B1(n6985), .B2(keyinput_g66), .ZN(n6756) );
  OAI221_X1 U7738 ( .B1(n6757), .B2(keyinput_g20), .C1(n6985), .C2(
        keyinput_g66), .A(n6756), .ZN(n6758) );
  OR4_X1 U7739 ( .A1(n6761), .A2(n6760), .A3(n6759), .A4(n6758), .ZN(n6762) );
  NOR4_X1 U7740 ( .A1(n6765), .A2(n6764), .A3(n6763), .A4(n6762), .ZN(n7127)
         );
  OAI22_X1 U7741 ( .A1(ADDRESS_REG_29__SCAN_IN), .A2(keyinput_g71), .B1(
        keyinput_g126), .B2(DATAWIDTH_REG_22__SCAN_IN), .ZN(n6766) );
  AOI221_X1 U7742 ( .B1(ADDRESS_REG_29__SCAN_IN), .B2(keyinput_g71), .C1(
        DATAWIDTH_REG_22__SCAN_IN), .C2(keyinput_g126), .A(n6766), .ZN(n6773)
         );
  OAI22_X1 U7743 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(keyinput_g44), .B2(
        MORE_REG_SCAN_IN), .ZN(n6767) );
  AOI221_X1 U7744 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(MORE_REG_SCAN_IN), 
        .C2(keyinput_g44), .A(n6767), .ZN(n6772) );
  OAI22_X1 U7745 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_g60), .B1(
        DATAWIDTH_REG_12__SCAN_IN), .B2(keyinput_g116), .ZN(n6768) );
  AOI221_X1 U7746 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_g60), .C1(
        keyinput_g116), .C2(DATAWIDTH_REG_12__SCAN_IN), .A(n6768), .ZN(n6771)
         );
  OAI22_X1 U7747 ( .A1(REIP_REG_27__SCAN_IN), .A2(keyinput_g55), .B1(
        DATAWIDTH_REG_8__SCAN_IN), .B2(keyinput_g112), .ZN(n6769) );
  AOI221_X1 U7748 ( .B1(REIP_REG_27__SCAN_IN), .B2(keyinput_g55), .C1(
        keyinput_g112), .C2(DATAWIDTH_REG_8__SCAN_IN), .A(n6769), .ZN(n6770)
         );
  NAND4_X1 U7749 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6913)
         );
  OAI22_X1 U7750 ( .A1(DATAI_12_), .A2(keyinput_g19), .B1(keyinput_g15), .B2(
        DATAI_16_), .ZN(n6774) );
  AOI221_X1 U7751 ( .B1(DATAI_12_), .B2(keyinput_g19), .C1(DATAI_16_), .C2(
        keyinput_g15), .A(n6774), .ZN(n6800) );
  OAI22_X1 U7752 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_g58), .B1(
        keyinput_g29), .B2(DATAI_2_), .ZN(n6775) );
  AOI221_X1 U7753 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_g58), .C1(DATAI_2_), .C2(keyinput_g29), .A(n6775), .ZN(n6778) );
  OAI22_X1 U7754 ( .A1(READY_N), .A2(keyinput_g35), .B1(keyinput_g125), .B2(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6776) );
  AOI221_X1 U7755 ( .B1(READY_N), .B2(keyinput_g35), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(keyinput_g125), .A(n6776), .ZN(n6777)
         );
  OAI211_X1 U7756 ( .C1(n6780), .C2(keyinput_g27), .A(n6778), .B(n6777), .ZN(
        n6779) );
  AOI21_X1 U7757 ( .B1(n6780), .B2(keyinput_g27), .A(n6779), .ZN(n6799) );
  AOI22_X1 U7758 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput_g83), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_g42), .ZN(n6781) );
  OAI221_X1 U7759 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput_g83), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_g42), .A(n6781), .ZN(n6788)
         );
  AOI22_X1 U7760 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(DATAI_30_), .B2(
        keyinput_g1), .ZN(n6782) );
  OAI221_X1 U7761 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_30_), .C2(
        keyinput_g1), .A(n6782), .ZN(n6787) );
  AOI22_X1 U7762 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput_g127), .B1(
        DATAI_25_), .B2(keyinput_g6), .ZN(n6783) );
  OAI221_X1 U7763 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput_g127), .C1(
        DATAI_25_), .C2(keyinput_g6), .A(n6783), .ZN(n6786) );
  AOI22_X1 U7764 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput_g104), .B1(
        DATAI_29_), .B2(keyinput_g2), .ZN(n6784) );
  OAI221_X1 U7765 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput_g104), .C1(
        DATAI_29_), .C2(keyinput_g2), .A(n6784), .ZN(n6785) );
  NOR4_X1 U7766 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6798)
         );
  AOI22_X1 U7767 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_21_), .B2(
        keyinput_g10), .ZN(n6789) );
  OAI221_X1 U7768 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_21_), .C2(
        keyinput_g10), .A(n6789), .ZN(n6796) );
  AOI22_X1 U7769 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_g40), .B1(
        BE_N_REG_2__SCAN_IN), .B2(keyinput_g68), .ZN(n6790) );
  OAI221_X1 U7770 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_g40), .C1(
        BE_N_REG_2__SCAN_IN), .C2(keyinput_g68), .A(n6790), .ZN(n6795) );
  AOI22_X1 U7771 ( .A1(ADDRESS_REG_25__SCAN_IN), .A2(keyinput_g75), .B1(
        DATAI_24_), .B2(keyinput_g7), .ZN(n6791) );
  OAI221_X1 U7772 ( .B1(ADDRESS_REG_25__SCAN_IN), .B2(keyinput_g75), .C1(
        DATAI_24_), .C2(keyinput_g7), .A(n6791), .ZN(n6794) );
  AOI22_X1 U7773 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(keyinput_g109), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_g43), .ZN(n6792) );
  OAI221_X1 U7774 ( .B1(DATAWIDTH_REG_5__SCAN_IN), .B2(keyinput_g109), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_g43), .A(n6792), .ZN(n6793) );
  NOR4_X1 U7775 ( .A1(n6796), .A2(n6795), .A3(n6794), .A4(n6793), .ZN(n6797)
         );
  NAND4_X1 U7776 ( .A1(n6800), .A2(n6799), .A3(n6798), .A4(n6797), .ZN(n6912)
         );
  AOI22_X1 U7777 ( .A1(n6802), .A2(keyinput_g120), .B1(n7000), .B2(
        keyinput_g102), .ZN(n6801) );
  OAI221_X1 U7778 ( .B1(n6802), .B2(keyinput_g120), .C1(n7000), .C2(
        keyinput_g102), .A(n6801), .ZN(n6811) );
  AOI22_X1 U7779 ( .A1(n7080), .A2(keyinput_g73), .B1(n7067), .B2(keyinput_g48), .ZN(n6803) );
  OAI221_X1 U7780 ( .B1(n7080), .B2(keyinput_g73), .C1(n7067), .C2(
        keyinput_g48), .A(n6803), .ZN(n6810) );
  INV_X1 U7781 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n6988) );
  AOI22_X1 U7782 ( .A1(n6805), .A2(keyinput_g124), .B1(n6988), .B2(
        keyinput_g37), .ZN(n6804) );
  OAI221_X1 U7783 ( .B1(n6805), .B2(keyinput_g124), .C1(n6988), .C2(
        keyinput_g37), .A(n6804), .ZN(n6809) );
  INV_X1 U7784 ( .A(DATAI_27_), .ZN(n6961) );
  AOI22_X1 U7785 ( .A1(n6961), .A2(keyinput_g4), .B1(keyinput_g107), .B2(n6807), .ZN(n6806) );
  OAI221_X1 U7786 ( .B1(n6961), .B2(keyinput_g4), .C1(n6807), .C2(
        keyinput_g107), .A(n6806), .ZN(n6808) );
  NOR4_X1 U7787 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6854)
         );
  AOI22_X1 U7788 ( .A1(n6814), .A2(keyinput_g101), .B1(keyinput_g81), .B2(
        n6813), .ZN(n6812) );
  OAI221_X1 U7789 ( .B1(n6814), .B2(keyinput_g101), .C1(n6813), .C2(
        keyinput_g81), .A(n6812), .ZN(n6823) );
  AOI22_X1 U7790 ( .A1(n7103), .A2(keyinput_g25), .B1(keyinput_g117), .B2(
        n6816), .ZN(n6815) );
  OAI221_X1 U7791 ( .B1(n7103), .B2(keyinput_g25), .C1(n6816), .C2(
        keyinput_g117), .A(n6815), .ZN(n6822) );
  AOI22_X1 U7792 ( .A1(n6975), .A2(keyinput_g82), .B1(n6818), .B2(keyinput_g89), .ZN(n6817) );
  OAI221_X1 U7793 ( .B1(n6975), .B2(keyinput_g82), .C1(n6818), .C2(
        keyinput_g89), .A(n6817), .ZN(n6821) );
  AOI22_X1 U7794 ( .A1(n6991), .A2(keyinput_g63), .B1(keyinput_g76), .B2(n7094), .ZN(n6819) );
  OAI221_X1 U7795 ( .B1(n6991), .B2(keyinput_g63), .C1(n7094), .C2(
        keyinput_g76), .A(n6819), .ZN(n6820) );
  NOR4_X1 U7796 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6853)
         );
  INV_X1 U7797 ( .A(DATAI_23_), .ZN(n7086) );
  AOI22_X1 U7798 ( .A1(n7086), .A2(keyinput_g8), .B1(keyinput_g118), .B2(n6825), .ZN(n6824) );
  OAI221_X1 U7799 ( .B1(n7086), .B2(keyinput_g8), .C1(n6825), .C2(
        keyinput_g118), .A(n6824), .ZN(n6836) );
  AOI22_X1 U7800 ( .A1(n7084), .A2(keyinput_g31), .B1(keyinput_g123), .B2(
        n6827), .ZN(n6826) );
  OAI221_X1 U7801 ( .B1(n7084), .B2(keyinput_g31), .C1(n6827), .C2(
        keyinput_g123), .A(n6826), .ZN(n6835) );
  AOI22_X1 U7802 ( .A1(n7065), .A2(keyinput_g24), .B1(keyinput_g16), .B2(n6829), .ZN(n6828) );
  OAI221_X1 U7803 ( .B1(n7065), .B2(keyinput_g24), .C1(n6829), .C2(
        keyinput_g16), .A(n6828), .ZN(n6834) );
  AOI22_X1 U7804 ( .A1(n6832), .A2(keyinput_g32), .B1(keyinput_g97), .B2(n6831), .ZN(n6830) );
  OAI221_X1 U7805 ( .B1(n6832), .B2(keyinput_g32), .C1(n6831), .C2(
        keyinput_g97), .A(n6830), .ZN(n6833) );
  NOR4_X1 U7806 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6852)
         );
  INV_X1 U7807 ( .A(DATAI_17_), .ZN(n6956) );
  AOI22_X1 U7808 ( .A1(n6838), .A2(keyinput_g70), .B1(n6956), .B2(keyinput_g14), .ZN(n6837) );
  OAI221_X1 U7809 ( .B1(n6838), .B2(keyinput_g70), .C1(n6956), .C2(
        keyinput_g14), .A(n6837), .ZN(n6850) );
  AOI22_X1 U7810 ( .A1(n6841), .A2(keyinput_g18), .B1(keyinput_g106), .B2(
        n6840), .ZN(n6839) );
  OAI221_X1 U7811 ( .B1(n6841), .B2(keyinput_g18), .C1(n6840), .C2(
        keyinput_g106), .A(n6839), .ZN(n6849) );
  AOI22_X1 U7812 ( .A1(n6843), .A2(keyinput_g30), .B1(keyinput_g78), .B2(n7102), .ZN(n6842) );
  OAI221_X1 U7813 ( .B1(n6843), .B2(keyinput_g30), .C1(n7102), .C2(
        keyinput_g78), .A(n6842), .ZN(n6848) );
  AOI22_X1 U7814 ( .A1(n6846), .A2(keyinput_g95), .B1(keyinput_g113), .B2(
        n6845), .ZN(n6844) );
  OAI221_X1 U7815 ( .B1(n6846), .B2(keyinput_g95), .C1(n6845), .C2(
        keyinput_g113), .A(n6844), .ZN(n6847) );
  NOR4_X1 U7816 ( .A1(n6850), .A2(n6849), .A3(n6848), .A4(n6847), .ZN(n6851)
         );
  NAND4_X1 U7817 ( .A1(n6854), .A2(n6853), .A3(n6852), .A4(n6851), .ZN(n6911)
         );
  INV_X1 U7818 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7819 ( .A1(n7001), .A2(keyinput_g47), .B1(n6856), .B2(keyinput_g67), .ZN(n6855) );
  OAI221_X1 U7820 ( .B1(n7001), .B2(keyinput_g47), .C1(n6856), .C2(
        keyinput_g67), .A(n6855), .ZN(n6866) );
  AOI22_X1 U7821 ( .A1(n6858), .A2(keyinput_g111), .B1(n5804), .B2(
        keyinput_g62), .ZN(n6857) );
  OAI221_X1 U7822 ( .B1(n6858), .B2(keyinput_g111), .C1(n5804), .C2(
        keyinput_g62), .A(n6857), .ZN(n6865) );
  AOI22_X1 U7823 ( .A1(n6861), .A2(keyinput_g52), .B1(keyinput_g53), .B2(n6860), .ZN(n6859) );
  OAI221_X1 U7824 ( .B1(n6861), .B2(keyinput_g52), .C1(n6860), .C2(
        keyinput_g53), .A(n6859), .ZN(n6864) );
  INV_X1 U7825 ( .A(DATAI_26_), .ZN(n7100) );
  AOI22_X1 U7826 ( .A1(n6974), .A2(keyinput_g98), .B1(n7100), .B2(keyinput_g5), 
        .ZN(n6862) );
  OAI221_X1 U7827 ( .B1(n6974), .B2(keyinput_g98), .C1(n7100), .C2(keyinput_g5), .A(n6862), .ZN(n6863) );
  NOR4_X1 U7828 ( .A1(n6866), .A2(n6865), .A3(n6864), .A4(n6863), .ZN(n6909)
         );
  AOI22_X1 U7829 ( .A1(n6869), .A2(keyinput_g79), .B1(n6868), .B2(keyinput_g61), .ZN(n6867) );
  OAI221_X1 U7830 ( .B1(n6869), .B2(keyinput_g79), .C1(n6868), .C2(
        keyinput_g61), .A(n6867), .ZN(n6881) );
  AOI22_X1 U7831 ( .A1(n6872), .A2(keyinput_g51), .B1(keyinput_g54), .B2(n6871), .ZN(n6870) );
  OAI221_X1 U7832 ( .B1(n6872), .B2(keyinput_g51), .C1(n6871), .C2(
        keyinput_g54), .A(n6870), .ZN(n6880) );
  AOI22_X1 U7833 ( .A1(n6875), .A2(keyinput_g119), .B1(n6874), .B2(
        keyinput_g90), .ZN(n6873) );
  OAI221_X1 U7834 ( .B1(n6875), .B2(keyinput_g119), .C1(n6874), .C2(
        keyinput_g90), .A(n6873), .ZN(n6879) );
  AOI22_X1 U7835 ( .A1(n6877), .A2(keyinput_g36), .B1(keyinput_g93), .B2(n7057), .ZN(n6876) );
  OAI221_X1 U7836 ( .B1(n6877), .B2(keyinput_g36), .C1(n7057), .C2(
        keyinput_g93), .A(n6876), .ZN(n6878) );
  NOR4_X1 U7837 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n6908)
         );
  INV_X1 U7838 ( .A(BS16_N), .ZN(n6883) );
  AOI22_X1 U7839 ( .A1(n7052), .A2(keyinput_g91), .B1(n6883), .B2(keyinput_g34), .ZN(n6882) );
  OAI221_X1 U7840 ( .B1(n7052), .B2(keyinput_g91), .C1(n6883), .C2(
        keyinput_g34), .A(n6882), .ZN(n6893) );
  AOI22_X1 U7841 ( .A1(n6962), .A2(keyinput_g41), .B1(n6952), .B2(keyinput_g72), .ZN(n6884) );
  OAI221_X1 U7842 ( .B1(n6962), .B2(keyinput_g41), .C1(n6952), .C2(
        keyinput_g72), .A(n6884), .ZN(n6892) );
  INV_X1 U7843 ( .A(DATAI_19_), .ZN(n6887) );
  AOI22_X1 U7844 ( .A1(n6887), .A2(keyinput_g12), .B1(n6886), .B2(keyinput_g56), .ZN(n6885) );
  OAI221_X1 U7845 ( .B1(n6887), .B2(keyinput_g12), .C1(n6886), .C2(
        keyinput_g56), .A(n6885), .ZN(n6891) );
  AOI22_X1 U7846 ( .A1(n6889), .A2(keyinput_g96), .B1(keyinput_g38), .B2(n7083), .ZN(n6888) );
  OAI221_X1 U7847 ( .B1(n6889), .B2(keyinput_g96), .C1(n7083), .C2(
        keyinput_g38), .A(n6888), .ZN(n6890) );
  NOR4_X1 U7848 ( .A1(n6893), .A2(n6892), .A3(n6891), .A4(n6890), .ZN(n6907)
         );
  AOI22_X1 U7849 ( .A1(n5765), .A2(keyinput_g57), .B1(keyinput_g86), .B2(n6895), .ZN(n6894) );
  OAI221_X1 U7850 ( .B1(n5765), .B2(keyinput_g57), .C1(n6895), .C2(
        keyinput_g86), .A(n6894), .ZN(n6905) );
  AOI22_X1 U7851 ( .A1(n6897), .A2(keyinput_g21), .B1(keyinput_g84), .B2(n6968), .ZN(n6896) );
  OAI221_X1 U7852 ( .B1(n6897), .B2(keyinput_g21), .C1(n6968), .C2(
        keyinput_g84), .A(n6896), .ZN(n6904) );
  INV_X1 U7853 ( .A(DATAI_22_), .ZN(n6900) );
  AOI22_X1 U7854 ( .A1(n6900), .A2(keyinput_g9), .B1(n6899), .B2(keyinput_g64), 
        .ZN(n6898) );
  OAI221_X1 U7855 ( .B1(n6900), .B2(keyinput_g9), .C1(n6899), .C2(keyinput_g64), .A(n6898), .ZN(n6903) );
  AOI22_X1 U7856 ( .A1(n7070), .A2(keyinput_g77), .B1(n6953), .B2(keyinput_g46), .ZN(n6901) );
  OAI221_X1 U7857 ( .B1(n7070), .B2(keyinput_g77), .C1(n6953), .C2(
        keyinput_g46), .A(n6901), .ZN(n6902) );
  NOR4_X1 U7858 ( .A1(n6905), .A2(n6904), .A3(n6903), .A4(n6902), .ZN(n6906)
         );
  NAND4_X1 U7859 ( .A1(n6909), .A2(n6908), .A3(n6907), .A4(n6906), .ZN(n6910)
         );
  NOR4_X1 U7860 ( .A1(n6913), .A2(n6912), .A3(n6911), .A4(n6910), .ZN(n7126)
         );
  OAI22_X1 U7861 ( .A1(REIP_REG_28__SCAN_IN), .A2(keyinput_f54), .B1(DATAI_12_), .B2(keyinput_f19), .ZN(n6914) );
  AOI221_X1 U7862 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_f54), .C1(
        keyinput_f19), .C2(DATAI_12_), .A(n6914), .ZN(n6921) );
  OAI22_X1 U7863 ( .A1(REIP_REG_20__SCAN_IN), .A2(keyinput_f62), .B1(DATAI_24_), .B2(keyinput_f7), .ZN(n6915) );
  AOI221_X1 U7864 ( .B1(REIP_REG_20__SCAN_IN), .B2(keyinput_f62), .C1(
        keyinput_f7), .C2(DATAI_24_), .A(n6915), .ZN(n6920) );
  OAI22_X1 U7865 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_f39), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(keyinput_f85), .ZN(n6916) );
  AOI221_X1 U7866 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f85), .C2(ADDRESS_REG_15__SCAN_IN), .A(n6916), .ZN(n6919) );
  OAI22_X1 U7867 ( .A1(REIP_REG_18__SCAN_IN), .A2(keyinput_f64), .B1(
        keyinput_f96), .B2(ADDRESS_REG_4__SCAN_IN), .ZN(n6917) );
  AOI221_X1 U7868 ( .B1(REIP_REG_18__SCAN_IN), .B2(keyinput_f64), .C1(
        ADDRESS_REG_4__SCAN_IN), .C2(keyinput_f96), .A(n6917), .ZN(n6918) );
  NAND4_X1 U7869 ( .A1(n6921), .A2(n6920), .A3(n6919), .A4(n6918), .ZN(n6950)
         );
  OAI22_X1 U7870 ( .A1(keyinput_f90), .A2(ADDRESS_REG_10__SCAN_IN), .B1(
        keyinput_f122), .B2(DATAWIDTH_REG_18__SCAN_IN), .ZN(n6922) );
  AOI221_X1 U7871 ( .B1(keyinput_f90), .B2(ADDRESS_REG_10__SCAN_IN), .C1(
        DATAWIDTH_REG_18__SCAN_IN), .C2(keyinput_f122), .A(n6922), .ZN(n6929)
         );
  OAI22_X1 U7872 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(DATAI_21_), .B2(
        keyinput_f10), .ZN(n6923) );
  AOI221_X1 U7873 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(keyinput_f10), .C2(
        DATAI_21_), .A(n6923), .ZN(n6928) );
  OAI22_X1 U7874 ( .A1(keyinput_f111), .A2(DATAWIDTH_REG_7__SCAN_IN), .B1(
        keyinput_f83), .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n6924) );
  AOI221_X1 U7875 ( .B1(keyinput_f111), .B2(DATAWIDTH_REG_7__SCAN_IN), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput_f83), .A(n6924), .ZN(n6927) );
  OAI22_X1 U7876 ( .A1(REIP_REG_17__SCAN_IN), .A2(keyinput_f65), .B1(DATAI_19_), .B2(keyinput_f12), .ZN(n6925) );
  AOI221_X1 U7877 ( .B1(REIP_REG_17__SCAN_IN), .B2(keyinput_f65), .C1(
        keyinput_f12), .C2(DATAI_19_), .A(n6925), .ZN(n6926) );
  NAND4_X1 U7878 ( .A1(n6929), .A2(n6928), .A3(n6927), .A4(n6926), .ZN(n6949)
         );
  OAI22_X1 U7879 ( .A1(REIP_REG_21__SCAN_IN), .A2(keyinput_f61), .B1(NA_N), 
        .B2(keyinput_f33), .ZN(n6930) );
  AOI221_X1 U7880 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f33), .C2(NA_N), .A(n6930), .ZN(n6937) );
  OAI22_X1 U7881 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f32), .ZN(n6931) );
  AOI221_X1 U7882 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f32), .C2(MEMORYFETCH_REG_SCAN_IN), .A(n6931), .ZN(n6936) );
  OAI22_X1 U7883 ( .A1(REIP_REG_31__SCAN_IN), .A2(keyinput_f51), .B1(
        REIP_REG_23__SCAN_IN), .B2(keyinput_f59), .ZN(n6932) );
  AOI221_X1 U7884 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f59), .C2(REIP_REG_23__SCAN_IN), .A(n6932), .ZN(n6935) );
  OAI22_X1 U7885 ( .A1(REIP_REG_26__SCAN_IN), .A2(keyinput_f56), .B1(
        keyinput_f108), .B2(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6933) );
  AOI221_X1 U7886 ( .B1(REIP_REG_26__SCAN_IN), .B2(keyinput_f56), .C1(
        DATAWIDTH_REG_4__SCAN_IN), .C2(keyinput_f108), .A(n6933), .ZN(n6934)
         );
  NAND4_X1 U7887 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6948)
         );
  OAI22_X1 U7888 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput_f58), .B1(
        keyinput_f123), .B2(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6938) );
  AOI221_X1 U7889 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput_f58), .C1(
        DATAWIDTH_REG_19__SCAN_IN), .C2(keyinput_f123), .A(n6938), .ZN(n6946)
         );
  OAI22_X1 U7890 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput_f120), .ZN(n6939) );
  AOI221_X1 U7891 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(keyinput_f120), .C2(
        DATAWIDTH_REG_16__SCAN_IN), .A(n6939), .ZN(n6945) );
  OAI22_X1 U7892 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(keyinput_f109), .B2(
        DATAWIDTH_REG_5__SCAN_IN), .ZN(n6940) );
  AOI221_X1 U7893 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(
        DATAWIDTH_REG_5__SCAN_IN), .C2(keyinput_f109), .A(n6940), .ZN(n6944)
         );
  OAI22_X1 U7894 ( .A1(keyinput_f126), .A2(n6942), .B1(keyinput_f104), .B2(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n6941) );
  AOI221_X1 U7895 ( .B1(n6942), .B2(keyinput_f126), .C1(keyinput_f104), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(n6941), .ZN(n6943) );
  NAND4_X1 U7896 ( .A1(n6946), .A2(n6945), .A3(n6944), .A4(n6943), .ZN(n6947)
         );
  NOR4_X1 U7897 ( .A1(n6950), .A2(n6949), .A3(n6948), .A4(n6947), .ZN(n7119)
         );
  AOI22_X1 U7898 ( .A1(n6953), .A2(keyinput_f46), .B1(keyinput_f72), .B2(n6952), .ZN(n6951) );
  OAI221_X1 U7899 ( .B1(n6953), .B2(keyinput_f46), .C1(n6952), .C2(
        keyinput_f72), .A(n6951), .ZN(n6966) );
  AOI22_X1 U7900 ( .A1(n6956), .A2(keyinput_f14), .B1(keyinput_f42), .B2(n6955), .ZN(n6954) );
  OAI221_X1 U7901 ( .B1(n6956), .B2(keyinput_f14), .C1(n6955), .C2(
        keyinput_f42), .A(n6954), .ZN(n6965) );
  INV_X1 U7902 ( .A(keyinput_f105), .ZN(n6958) );
  AOI22_X1 U7903 ( .A1(n6959), .A2(keyinput_f87), .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6958), .ZN(n6957) );
  OAI221_X1 U7904 ( .B1(n6959), .B2(keyinput_f87), .C1(n6958), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(n6957), .ZN(n6964) );
  AOI22_X1 U7905 ( .A1(n6962), .A2(keyinput_f41), .B1(n6961), .B2(keyinput_f4), 
        .ZN(n6960) );
  OAI221_X1 U7906 ( .B1(n6962), .B2(keyinput_f41), .C1(n6961), .C2(keyinput_f4), .A(n6960), .ZN(n6963) );
  NOR4_X1 U7907 ( .A1(n6966), .A2(n6965), .A3(n6964), .A4(n6963), .ZN(n7118)
         );
  INV_X1 U7908 ( .A(DATAI_25_), .ZN(n6969) );
  OAI22_X1 U7909 ( .A1(n6969), .A2(keyinput_f6), .B1(n6968), .B2(keyinput_f84), 
        .ZN(n6967) );
  AOI221_X1 U7910 ( .B1(n6969), .B2(keyinput_f6), .C1(keyinput_f84), .C2(n6968), .A(n6967), .ZN(n6982) );
  OAI22_X1 U7911 ( .A1(n6972), .A2(keyinput_f17), .B1(n6971), .B2(
        keyinput_f127), .ZN(n6970) );
  AOI221_X1 U7912 ( .B1(n6972), .B2(keyinput_f17), .C1(keyinput_f127), .C2(
        n6971), .A(n6970), .ZN(n6981) );
  OAI22_X1 U7913 ( .A1(n6975), .A2(keyinput_f82), .B1(n6974), .B2(keyinput_f98), .ZN(n6973) );
  AOI221_X1 U7914 ( .B1(n6975), .B2(keyinput_f82), .C1(keyinput_f98), .C2(
        n6974), .A(n6973), .ZN(n6980) );
  INV_X1 U7915 ( .A(keyinput_f106), .ZN(n6977) );
  OAI22_X1 U7916 ( .A1(n6978), .A2(keyinput_f22), .B1(n6977), .B2(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n6976) );
  AOI221_X1 U7917 ( .B1(n6978), .B2(keyinput_f22), .C1(
        DATAWIDTH_REG_2__SCAN_IN), .C2(n6977), .A(n6976), .ZN(n6979) );
  NAND4_X1 U7918 ( .A1(n6982), .A2(n6981), .A3(n6980), .A4(n6979), .ZN(n7014)
         );
  OAI22_X1 U7919 ( .A1(n6985), .A2(keyinput_f66), .B1(n6984), .B2(keyinput_f99), .ZN(n6983) );
  AOI221_X1 U7920 ( .B1(n6985), .B2(keyinput_f66), .C1(keyinput_f99), .C2(
        n6984), .A(n6983), .ZN(n6998) );
  INV_X1 U7921 ( .A(keyinput_f36), .ZN(n6987) );
  OAI22_X1 U7922 ( .A1(n6988), .A2(keyinput_f37), .B1(n6987), .B2(HOLD), .ZN(
        n6986) );
  AOI221_X1 U7923 ( .B1(n6988), .B2(keyinput_f37), .C1(HOLD), .C2(n6987), .A(
        n6986), .ZN(n6997) );
  INV_X1 U7924 ( .A(keyinput_f125), .ZN(n6990) );
  OAI22_X1 U7925 ( .A1(n6991), .A2(keyinput_f63), .B1(n6990), .B2(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6989) );
  AOI221_X1 U7926 ( .B1(n6991), .B2(keyinput_f63), .C1(
        DATAWIDTH_REG_21__SCAN_IN), .C2(n6990), .A(n6989), .ZN(n6996) );
  INV_X1 U7927 ( .A(keyinput_f115), .ZN(n6993) );
  OAI22_X1 U7928 ( .A1(keyinput_f112), .A2(n6994), .B1(n6993), .B2(
        DATAWIDTH_REG_11__SCAN_IN), .ZN(n6992) );
  AOI221_X1 U7929 ( .B1(n6994), .B2(keyinput_f112), .C1(n6993), .C2(
        DATAWIDTH_REG_11__SCAN_IN), .A(n6992), .ZN(n6995) );
  NAND4_X1 U7930 ( .A1(n6998), .A2(n6997), .A3(n6996), .A4(n6995), .ZN(n7013)
         );
  AOI22_X1 U7931 ( .A1(n7001), .A2(keyinput_f47), .B1(n7000), .B2(
        keyinput_f102), .ZN(n6999) );
  OAI221_X1 U7932 ( .B1(n7001), .B2(keyinput_f47), .C1(n7000), .C2(
        keyinput_f102), .A(n6999), .ZN(n7012) );
  OAI22_X1 U7933 ( .A1(n7004), .A2(keyinput_f68), .B1(n7003), .B2(keyinput_f94), .ZN(n7002) );
  AOI221_X1 U7934 ( .B1(n7004), .B2(keyinput_f68), .C1(keyinput_f94), .C2(
        n7003), .A(n7002), .ZN(n7010) );
  INV_X1 U7935 ( .A(keyinput_f119), .ZN(n7006) );
  OAI22_X1 U7936 ( .A1(n5765), .A2(keyinput_f57), .B1(n7006), .B2(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n7005) );
  AOI221_X1 U7937 ( .B1(n5765), .B2(keyinput_f57), .C1(
        DATAWIDTH_REG_15__SCAN_IN), .C2(n7006), .A(n7005), .ZN(n7009) );
  XNOR2_X1 U7938 ( .A(keyinput_f117), .B(DATAWIDTH_REG_13__SCAN_IN), .ZN(n7008) );
  XNOR2_X1 U7939 ( .A(ADDRESS_REG_21__SCAN_IN), .B(keyinput_f79), .ZN(n7007)
         );
  NAND4_X1 U7940 ( .A1(n7010), .A2(n7009), .A3(n7008), .A4(n7007), .ZN(n7011)
         );
  NOR4_X1 U7941 ( .A1(n7014), .A2(n7013), .A3(n7012), .A4(n7011), .ZN(n7117)
         );
  XOR2_X1 U7942 ( .A(ADDRESS_REG_0__SCAN_IN), .B(keyinput_f100), .Z(n7021) );
  AOI22_X1 U7943 ( .A1(keyinput_f124), .A2(DATAWIDTH_REG_20__SCAN_IN), .B1(
        STATE_REG_0__SCAN_IN), .B2(keyinput_f103), .ZN(n7015) );
  OAI221_X1 U7944 ( .B1(keyinput_f124), .B2(DATAWIDTH_REG_20__SCAN_IN), .C1(
        STATE_REG_0__SCAN_IN), .C2(keyinput_f103), .A(n7015), .ZN(n7020) );
  AOI22_X1 U7945 ( .A1(keyinput_f116), .A2(DATAWIDTH_REG_12__SCAN_IN), .B1(
        DATAI_22_), .B2(keyinput_f9), .ZN(n7016) );
  OAI221_X1 U7946 ( .B1(keyinput_f116), .B2(DATAWIDTH_REG_12__SCAN_IN), .C1(
        DATAI_22_), .C2(keyinput_f9), .A(n7016), .ZN(n7019) );
  AOI22_X1 U7947 ( .A1(DATAI_28_), .A2(keyinput_f3), .B1(REIP_REG_30__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n7017) );
  OAI221_X1 U7948 ( .B1(DATAI_28_), .B2(keyinput_f3), .C1(REIP_REG_30__SCAN_IN), .C2(keyinput_f52), .A(n7017), .ZN(n7018) );
  NOR4_X1 U7949 ( .A1(n7021), .A2(n7020), .A3(n7019), .A4(n7018), .ZN(n7049)
         );
  AOI22_X1 U7950 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput_f89), .B1(
        DATAI_4_), .B2(keyinput_f27), .ZN(n7022) );
  OAI221_X1 U7951 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput_f89), .C1(
        DATAI_4_), .C2(keyinput_f27), .A(n7022), .ZN(n7029) );
  AOI22_X1 U7952 ( .A1(keyinput_f75), .A2(ADDRESS_REG_25__SCAN_IN), .B1(
        DATAI_13_), .B2(keyinput_f18), .ZN(n7023) );
  OAI221_X1 U7953 ( .B1(keyinput_f75), .B2(ADDRESS_REG_25__SCAN_IN), .C1(
        DATAI_13_), .C2(keyinput_f18), .A(n7023), .ZN(n7028) );
  AOI22_X1 U7954 ( .A1(keyinput_f34), .A2(BS16_N), .B1(READY_N), .B2(
        keyinput_f35), .ZN(n7024) );
  OAI221_X1 U7955 ( .B1(keyinput_f34), .B2(BS16_N), .C1(READY_N), .C2(
        keyinput_f35), .A(n7024), .ZN(n7027) );
  AOI22_X1 U7956 ( .A1(keyinput_f114), .A2(DATAWIDTH_REG_10__SCAN_IN), .B1(
        BE_N_REG_0__SCAN_IN), .B2(keyinput_f70), .ZN(n7025) );
  OAI221_X1 U7957 ( .B1(keyinput_f114), .B2(DATAWIDTH_REG_10__SCAN_IN), .C1(
        BE_N_REG_0__SCAN_IN), .C2(keyinput_f70), .A(n7025), .ZN(n7026) );
  NOR4_X1 U7958 ( .A1(n7029), .A2(n7028), .A3(n7027), .A4(n7026), .ZN(n7048)
         );
  AOI22_X1 U7959 ( .A1(keyinput_f71), .A2(ADDRESS_REG_29__SCAN_IN), .B1(
        DATAI_11_), .B2(keyinput_f20), .ZN(n7030) );
  OAI221_X1 U7960 ( .B1(keyinput_f71), .B2(ADDRESS_REG_29__SCAN_IN), .C1(
        DATAI_11_), .C2(keyinput_f20), .A(n7030), .ZN(n7037) );
  AOI22_X1 U7961 ( .A1(REIP_REG_29__SCAN_IN), .A2(keyinput_f53), .B1(
        STATEBS16_REG_SCAN_IN), .B2(keyinput_f43), .ZN(n7031) );
  OAI221_X1 U7962 ( .B1(REIP_REG_29__SCAN_IN), .B2(keyinput_f53), .C1(
        STATEBS16_REG_SCAN_IN), .C2(keyinput_f43), .A(n7031), .ZN(n7036) );
  AOI22_X1 U7963 ( .A1(ADDRESS_REG_5__SCAN_IN), .A2(keyinput_f95), .B1(
        DATAI_2_), .B2(keyinput_f29), .ZN(n7032) );
  OAI221_X1 U7964 ( .B1(ADDRESS_REG_5__SCAN_IN), .B2(keyinput_f95), .C1(
        DATAI_2_), .C2(keyinput_f29), .A(n7032), .ZN(n7035) );
  AOI22_X1 U7965 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(STATE_REG_2__SCAN_IN), .B2(keyinput_f101), .ZN(n7033) );
  OAI221_X1 U7966 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput_f101), .A(n7033), .ZN(n7034) );
  NOR4_X1 U7967 ( .A1(n7037), .A2(n7036), .A3(n7035), .A4(n7034), .ZN(n7047)
         );
  AOI22_X1 U7968 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_10_), .B2(
        keyinput_f21), .ZN(n7038) );
  OAI221_X1 U7969 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(DATAI_10_), .C2(
        keyinput_f21), .A(n7038), .ZN(n7045) );
  AOI22_X1 U7970 ( .A1(keyinput_f81), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        DATAI_18_), .B2(keyinput_f13), .ZN(n7039) );
  OAI221_X1 U7971 ( .B1(keyinput_f81), .B2(ADDRESS_REG_19__SCAN_IN), .C1(
        DATAI_18_), .C2(keyinput_f13), .A(n7039), .ZN(n7044) );
  AOI22_X1 U7972 ( .A1(keyinput_f74), .A2(ADDRESS_REG_26__SCAN_IN), .B1(
        DATAI_15_), .B2(keyinput_f16), .ZN(n7040) );
  OAI221_X1 U7973 ( .B1(keyinput_f74), .B2(ADDRESS_REG_26__SCAN_IN), .C1(
        DATAI_15_), .C2(keyinput_f16), .A(n7040), .ZN(n7043) );
  AOI22_X1 U7974 ( .A1(keyinput_f67), .A2(BE_N_REG_3__SCAN_IN), .B1(
        keyinput_f110), .B2(DATAWIDTH_REG_6__SCAN_IN), .ZN(n7041) );
  OAI221_X1 U7975 ( .B1(keyinput_f67), .B2(BE_N_REG_3__SCAN_IN), .C1(
        keyinput_f110), .C2(DATAWIDTH_REG_6__SCAN_IN), .A(n7041), .ZN(n7042)
         );
  NOR4_X1 U7976 ( .A1(n7045), .A2(n7044), .A3(n7043), .A4(n7042), .ZN(n7046)
         );
  NAND4_X1 U7977 ( .A1(n7049), .A2(n7048), .A3(n7047), .A4(n7046), .ZN(n7115)
         );
  INV_X1 U7978 ( .A(keyinput_f107), .ZN(n7051) );
  AOI22_X1 U7979 ( .A1(n7052), .A2(keyinput_f91), .B1(DATAWIDTH_REG_3__SCAN_IN), .B2(n7051), .ZN(n7050) );
  OAI221_X1 U7980 ( .B1(n7052), .B2(keyinput_f91), .C1(n7051), .C2(
        DATAWIDTH_REG_3__SCAN_IN), .A(n7050), .ZN(n7114) );
  OAI22_X1 U7981 ( .A1(n7055), .A2(keyinput_f40), .B1(n7054), .B2(keyinput_f80), .ZN(n7053) );
  AOI221_X1 U7982 ( .B1(n7055), .B2(keyinput_f40), .C1(keyinput_f80), .C2(
        n7054), .A(n7053), .ZN(n7062) );
  INV_X1 U7983 ( .A(DATAI_29_), .ZN(n7058) );
  OAI22_X1 U7984 ( .A1(n7058), .A2(keyinput_f2), .B1(n7057), .B2(keyinput_f93), 
        .ZN(n7056) );
  AOI221_X1 U7985 ( .B1(n7058), .B2(keyinput_f2), .C1(keyinput_f93), .C2(n7057), .A(n7056), .ZN(n7061) );
  XNOR2_X1 U7986 ( .A(ADDRESS_REG_14__SCAN_IN), .B(keyinput_f86), .ZN(n7060)
         );
  XNOR2_X1 U7987 ( .A(keyinput_f118), .B(DATAWIDTH_REG_14__SCAN_IN), .ZN(n7059) );
  NAND4_X1 U7988 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n7113)
         );
  INV_X1 U7989 ( .A(DATAI_20_), .ZN(n7064) );
  AOI22_X1 U7990 ( .A1(n7065), .A2(keyinput_f24), .B1(keyinput_f11), .B2(n7064), .ZN(n7063) );
  OAI221_X1 U7991 ( .B1(n7065), .B2(keyinput_f24), .C1(n7064), .C2(
        keyinput_f11), .A(n7063), .ZN(n7078) );
  AOI22_X1 U7992 ( .A1(n7068), .A2(keyinput_f60), .B1(keyinput_f48), .B2(n7067), .ZN(n7066) );
  OAI221_X1 U7993 ( .B1(n7068), .B2(keyinput_f60), .C1(n7067), .C2(
        keyinput_f48), .A(n7066), .ZN(n7077) );
  AOI22_X1 U7994 ( .A1(n7071), .A2(keyinput_f0), .B1(keyinput_f77), .B2(n7070), 
        .ZN(n7069) );
  OAI221_X1 U7995 ( .B1(n7071), .B2(keyinput_f0), .C1(n7070), .C2(keyinput_f77), .A(n7069), .ZN(n7076) );
  INV_X1 U7996 ( .A(keyinput_f113), .ZN(n7073) );
  AOI22_X1 U7997 ( .A1(n7074), .A2(keyinput_f28), .B1(DATAWIDTH_REG_9__SCAN_IN), .B2(n7073), .ZN(n7072) );
  OAI221_X1 U7998 ( .B1(n7074), .B2(keyinput_f28), .C1(n7073), .C2(
        DATAWIDTH_REG_9__SCAN_IN), .A(n7072), .ZN(n7075) );
  NOR4_X1 U7999 ( .A1(n7078), .A2(n7077), .A3(n7076), .A4(n7075), .ZN(n7111)
         );
  OAI22_X1 U8000 ( .A1(keyinput_f121), .A2(n7081), .B1(n7080), .B2(
        keyinput_f73), .ZN(n7079) );
  AOI221_X1 U8001 ( .B1(n7081), .B2(keyinput_f121), .C1(n7080), .C2(
        keyinput_f73), .A(n7079), .ZN(n7110) );
  XOR2_X1 U8002 ( .A(ADDRESS_REG_3__SCAN_IN), .B(keyinput_f97), .Z(n7091) );
  XOR2_X1 U8003 ( .A(keyinput_f50), .B(BYTEENABLE_REG_3__SCAN_IN), .Z(n7090)
         );
  AOI22_X1 U8004 ( .A1(n7084), .A2(keyinput_f31), .B1(keyinput_f38), .B2(n7083), .ZN(n7082) );
  OAI221_X1 U8005 ( .B1(n7084), .B2(keyinput_f31), .C1(n7083), .C2(
        keyinput_f38), .A(n7082), .ZN(n7089) );
  AOI22_X1 U8006 ( .A1(n7087), .A2(keyinput_f55), .B1(keyinput_f8), .B2(n7086), 
        .ZN(n7085) );
  OAI221_X1 U8007 ( .B1(n7087), .B2(keyinput_f55), .C1(n7086), .C2(keyinput_f8), .A(n7085), .ZN(n7088) );
  NOR4_X1 U8008 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .ZN(n7109)
         );
  AOI22_X1 U8009 ( .A1(n7094), .A2(keyinput_f76), .B1(keyinput_f88), .B2(n7093), .ZN(n7092) );
  OAI221_X1 U8010 ( .B1(n7094), .B2(keyinput_f76), .C1(n7093), .C2(
        keyinput_f88), .A(n7092), .ZN(n7107) );
  INV_X1 U8011 ( .A(MORE_REG_SCAN_IN), .ZN(n7096) );
  AOI22_X1 U8012 ( .A1(n7097), .A2(keyinput_f69), .B1(n7096), .B2(keyinput_f44), .ZN(n7095) );
  OAI221_X1 U8013 ( .B1(n7097), .B2(keyinput_f69), .C1(n7096), .C2(
        keyinput_f44), .A(n7095), .ZN(n7106) );
  AOI22_X1 U8014 ( .A1(n7100), .A2(keyinput_f5), .B1(keyinput_f49), .B2(n7099), 
        .ZN(n7098) );
  OAI221_X1 U8015 ( .B1(n7100), .B2(keyinput_f5), .C1(n7099), .C2(keyinput_f49), .A(n7098), .ZN(n7105) );
  AOI22_X1 U8016 ( .A1(n7103), .A2(keyinput_f25), .B1(keyinput_f78), .B2(n7102), .ZN(n7101) );
  OAI221_X1 U8017 ( .B1(n7103), .B2(keyinput_f25), .C1(n7102), .C2(
        keyinput_f78), .A(n7101), .ZN(n7104) );
  NOR4_X1 U8018 ( .A1(n7107), .A2(n7106), .A3(n7105), .A4(n7104), .ZN(n7108)
         );
  NAND4_X1 U8019 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7112)
         );
  NOR4_X1 U8020 ( .A1(n7115), .A2(n7114), .A3(n7113), .A4(n7112), .ZN(n7116)
         );
  NAND4_X1 U8021 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7121)
         );
  AOI21_X1 U8022 ( .B1(keyinput_f92), .B2(n7121), .A(keyinput_g92), .ZN(n7123)
         );
  INV_X1 U8023 ( .A(keyinput_f92), .ZN(n7120) );
  AOI21_X1 U8024 ( .B1(n7121), .B2(n7120), .A(n7124), .ZN(n7122) );
  AOI22_X1 U8025 ( .A1(n7124), .A2(n7123), .B1(keyinput_g92), .B2(n7122), .ZN(
        n7125) );
  AOI21_X1 U8026 ( .B1(n7127), .B2(n7126), .A(n7125), .ZN(n7131) );
  AOI22_X1 U8027 ( .A1(n7129), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n7128), .ZN(n7130) );
  XNOR2_X1 U8028 ( .A(n7131), .B(n7130), .ZN(U3445) );
  NAND2_X2 U3783 ( .A1(n3306), .A2(n3305), .ZN(n3373) );
  BUF_X1 U3604 ( .A(n4293), .Z(n3157) );
  INV_X2 U3603 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3791) );
  INV_X1 U3654 ( .A(n5774), .ZN(n5944) );
  CLKBUF_X1 U3664 ( .A(n3439), .Z(n4446) );
  AND2_X1 U3763 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4733) );
  CLKBUF_X1 U3893 ( .A(n4228), .Z(n4229) );
  CLKBUF_X2 U5163 ( .A(n3385), .Z(n3357) );
endmodule

