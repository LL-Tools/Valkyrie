

module b15_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD, 
        READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN, 
        M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN, 
        STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN, 
        W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N,
         BS16_N, READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
         CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
         REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
         FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846,
         n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
         n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
         n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
         n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886,
         n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896,
         n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906,
         n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916,
         n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926,
         n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936,
         n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946,
         n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956,
         n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
         n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
         n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
         n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996,
         n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006,
         n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
         n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
         n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
         n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
         n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
         n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
         n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
         n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
         n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
         n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126,
         n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136,
         n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146,
         n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156,
         n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166,
         n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176,
         n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186,
         n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
         n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
         n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216,
         n7217, n7218;

  OR2_X1 U3458 ( .A1(n5938), .A2(n5920), .ZN(n5922) );
  NAND2_X1 U34590 ( .A1(n5491), .A2(n5490), .ZN(n5628) );
  NAND2_X1 U34600 ( .A1(n3897), .A2(n3896), .ZN(n5189) );
  NAND2_X1 U34610 ( .A1(n3452), .A2(n3703), .ZN(n4777) );
  NOR2_X1 U34620 ( .A1(n3460), .A2(n7072), .ZN(n4247) );
  AND2_X1 U34630 ( .A1(n3460), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4239) );
  CLKBUF_X2 U34640 ( .A(n3572), .Z(n4604) );
  CLKBUF_X2 U34650 ( .A(n3682), .Z(n4612) );
  NAND2_X1 U3466 ( .A1(n3451), .A2(n3536), .ZN(n3602) );
  NAND2_X1 U3467 ( .A1(n3504), .A2(n3503), .ZN(n3622) );
  AND4_X1 U34680 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3525)
         );
  AND2_X2 U34690 ( .A1(n4842), .A2(n3468), .ZN(n3756) );
  INV_X1 U34710 ( .A(n7218), .ZN(n3425) );
  CLKBUF_X2 U34720 ( .A(n3636), .Z(n4602) );
  AND2_X2 U34730 ( .A1(n5139), .A2(n5164), .ZN(n3751) );
  INV_X1 U34740 ( .A(n3587), .ZN(n3527) );
  NAND2_X1 U3475 ( .A1(n3623), .A2(n3584), .ZN(n3595) );
  INV_X1 U3476 ( .A(n3602), .ZN(n4944) );
  OR2_X1 U3477 ( .A1(n5956), .A2(n4325), .ZN(n5995) );
  NOR2_X1 U3478 ( .A1(n3431), .A2(n5628), .ZN(n5706) );
  INV_X1 U3480 ( .A(n6981), .ZN(n7010) );
  OR2_X1 U3481 ( .A1(n5854), .A2(n4475), .ZN(n6696) );
  NOR2_X1 U3482 ( .A1(n4733), .A2(n4751), .ZN(n5349) );
  NOR2_X1 U3483 ( .A1(n3602), .A2(n4733), .ZN(n3630) );
  AND2_X2 U3484 ( .A1(n4733), .A2(n4751), .ZN(n4767) );
  XNOR2_X2 U3486 ( .A(n3847), .B(n3848), .ZN(n4412) );
  AND2_X2 U3488 ( .A1(n5167), .A2(n3468), .ZN(n3750) );
  OAI21_X2 U3489 ( .B1(n4408), .B2(n4446), .A(n4407), .ZN(n4411) );
  NOR2_X1 U3490 ( .A1(n5189), .A2(n5418), .ZN(n5452) );
  AOI21_X2 U3491 ( .B1(n5638), .B2(n5637), .A(n3454), .ZN(n4459) );
  NOR2_X2 U3492 ( .A1(n5562), .A2(n4455), .ZN(n5638) );
  AOI211_X2 U3493 ( .C1(n6693), .C2(n5890), .A(n5782), .B(n5781), .ZN(n5783)
         );
  AND2_X1 U3494 ( .A1(n4733), .A2(n4751), .ZN(n3426) );
  NAND2_X1 U3496 ( .A1(n4418), .A2(n4417), .ZN(n4428) );
  AOI21_X2 U3497 ( .B1(n4396), .B2(n4435), .A(n4395), .ZN(n6664) );
  OAI21_X2 U3498 ( .B1(n4386), .B2(n4446), .A(n4385), .ZN(n4861) );
  NAND2_X4 U3500 ( .A1(n3710), .A2(n3709), .ZN(n4386) );
  AND2_X1 U3501 ( .A1(n5917), .A2(n5916), .ZN(n5931) );
  NAND2_X1 U3502 ( .A1(n6062), .A2(n6061), .ZN(n6060) );
  NAND2_X1 U3503 ( .A1(n4777), .A2(n4776), .ZN(n4775) );
  AND2_X1 U3504 ( .A1(n5981), .A2(n4354), .ZN(n5936) );
  NOR2_X1 U3505 ( .A1(n3801), .A2(n3800), .ZN(n3815) );
  OAI21_X1 U3507 ( .B1(n4914), .B2(STATE2_REG_0__SCAN_IN), .A(n3764), .ZN(
        n3765) );
  OR2_X1 U3508 ( .A1(n5194), .A2(n5193), .ZN(n5419) );
  CLKBUF_X1 U3509 ( .A(n3736), .Z(n3737) );
  OAI21_X1 U3510 ( .B1(n3736), .B2(n5818), .A(n3615), .ZN(n3668) );
  AOI22_X1 U3511 ( .A1(n4649), .A2(n5856), .B1(n4474), .B2(n4268), .ZN(n3634)
         );
  NAND2_X1 U3512 ( .A1(n3586), .A2(n3602), .ZN(n3627) );
  AND2_X1 U3513 ( .A1(n3587), .A2(n4733), .ZN(n3460) );
  CLKBUF_X2 U3514 ( .A(n3622), .Z(n4378) );
  INV_X2 U3515 ( .A(n4733), .ZN(n4939) );
  AND4_X1 U3516 ( .A1(n3478), .A2(n3477), .A3(n3476), .A4(n3475), .ZN(n3484)
         );
  CLKBUF_X2 U3517 ( .A(n3676), .Z(n4613) );
  NOR2_X1 U3518 ( .A1(n4634), .A2(n4633), .ZN(n4635) );
  AND2_X1 U3519 ( .A1(n5977), .A2(n5976), .ZN(n7115) );
  OR2_X1 U3520 ( .A1(n5975), .A2(n5974), .ZN(n5977) );
  NAND2_X1 U3521 ( .A1(n4188), .A2(n5932), .ZN(n6073) );
  AOI21_X1 U3522 ( .B1(n5907), .B2(n5918), .A(n5906), .ZN(n6049) );
  OAI21_X1 U3523 ( .B1(n5931), .B2(n5919), .A(n5918), .ZN(n6054) );
  NAND2_X1 U3524 ( .A1(n6060), .A2(n3456), .ZN(n6053) );
  AOI21_X1 U3525 ( .B1(n6060), .B2(n4490), .A(n4639), .ZN(n6031) );
  OAI21_X1 U3526 ( .B1(n4464), .B2(n4463), .A(n4460), .ZN(n4465) );
  OAI22_X1 U3527 ( .A1(n5437), .A2(n5438), .B1(n4453), .B2(n5445), .ZN(n5581)
         );
  AND2_X1 U3528 ( .A1(n4426), .A2(n4425), .ZN(n5509) );
  XNOR2_X1 U3529 ( .A(n4449), .B(n3873), .ZN(n4436) );
  NAND2_X1 U3530 ( .A1(n3827), .A2(n3826), .ZN(n4789) );
  NAND2_X1 U3531 ( .A1(n3846), .A2(n3845), .ZN(n4852) );
  NAND2_X1 U3532 ( .A1(n4775), .A2(n3768), .ZN(n4763) );
  NAND2_X1 U3533 ( .A1(n3798), .A2(n3797), .ZN(n4798) );
  OAI21_X1 U3534 ( .B1(n5575), .B2(n4388), .A(n4387), .ZN(n6666) );
  OR2_X1 U3535 ( .A1(n3766), .A2(n3765), .ZN(n3440) );
  NAND2_X1 U3536 ( .A1(n3731), .A2(n3730), .ZN(n3766) );
  NAND2_X1 U3537 ( .A1(n4861), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4860)
         );
  CLKBUF_X1 U3538 ( .A(n4914), .Z(n5344) );
  NAND2_X1 U3539 ( .A1(n5171), .A2(n3748), .ZN(n4914) );
  NAND2_X1 U3540 ( .A1(n3745), .A2(n3744), .ZN(n5171) );
  AND2_X2 U3541 ( .A1(n4253), .A2(n4252), .ZN(n5854) );
  INV_X1 U3542 ( .A(n3747), .ZN(n3744) );
  AND2_X1 U3543 ( .A1(n3743), .A2(n3742), .ZN(n3747) );
  NOR2_X1 U3544 ( .A1(n4857), .A2(n4807), .ZN(n5025) );
  OR2_X1 U3545 ( .A1(n4692), .A2(n3635), .ZN(n3450) );
  OR2_X1 U3546 ( .A1(n3428), .A2(n4802), .ZN(n4857) );
  OAI21_X1 U3547 ( .B1(n5137), .B2(n3613), .A(n3439), .ZN(n3614) );
  AND2_X1 U3548 ( .A1(n4772), .A2(n4771), .ZN(n4800) );
  AOI21_X1 U3549 ( .B1(n5362), .B2(n4767), .A(n4276), .ZN(n4772) );
  NAND2_X1 U3550 ( .A1(n3616), .A2(n3589), .ZN(n4698) );
  OR2_X1 U3551 ( .A1(n5626), .A2(n5627), .ZN(n4311) );
  NAND2_X1 U3552 ( .A1(n3581), .A2(n4939), .ZN(n3616) );
  INV_X1 U3553 ( .A(n3628), .ZN(n4016) );
  NAND2_X1 U3554 ( .A1(n3695), .A2(n3694), .ZN(n3707) );
  MUX2_X1 U3555 ( .A(n3691), .B(n4447), .S(n3690), .Z(n3706) );
  AND3_X1 U3556 ( .A1(n3667), .A2(n3666), .A3(n3691), .ZN(n3728) );
  AND2_X1 U3557 ( .A1(n3599), .A2(n4944), .ZN(n4768) );
  AND3_X1 U3558 ( .A1(n3693), .A2(n3692), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3694) );
  INV_X1 U3559 ( .A(n3623), .ZN(n3711) );
  INV_X2 U3560 ( .A(n4268), .ZN(n5859) );
  AND2_X2 U3561 ( .A1(n3602), .A2(n4751), .ZN(n4268) );
  OR2_X1 U3562 ( .A1(n3664), .A2(n3663), .ZN(n4445) );
  OR2_X1 U3563 ( .A1(n3651), .A2(n3650), .ZN(n4375) );
  INV_X1 U3564 ( .A(n4687), .ZN(n4377) );
  INV_X1 U3565 ( .A(n3622), .ZN(n5734) );
  AND4_X1 U3566 ( .A1(n3531), .A2(n3530), .A3(n3529), .A4(n3528), .ZN(n3451)
         );
  AND4_X1 U3567 ( .A1(n3567), .A2(n3566), .A3(n3565), .A4(n3564), .ZN(n3579)
         );
  AND4_X1 U3568 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3580)
         );
  AND4_X1 U3569 ( .A1(n3571), .A2(n3570), .A3(n3569), .A4(n3568), .ZN(n3578)
         );
  AND4_X1 U3570 ( .A1(n3552), .A2(n3551), .A3(n3550), .A4(n3549), .ZN(n3553)
         );
  AND4_X1 U3571 ( .A1(n3548), .A2(n3547), .A3(n3546), .A4(n3545), .ZN(n3554)
         );
  AND4_X1 U3572 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3555)
         );
  AND4_X1 U3573 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(n3556)
         );
  AND4_X1 U3574 ( .A1(n3502), .A2(n3501), .A3(n3500), .A4(n3499), .ZN(n3503)
         );
  AND4_X1 U3575 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(n3504)
         );
  AND4_X1 U3576 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3483)
         );
  AND4_X1 U3577 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3536)
         );
  AND4_X1 U3578 ( .A1(n3488), .A2(n3487), .A3(n3486), .A4(n3485), .ZN(n3494)
         );
  AOI22_X1 U3579 ( .A1(n3750), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3470) );
  BUF_X2 U3580 ( .A(n3642), .Z(n4110) );
  CLKBUF_X2 U3581 ( .A(n3637), .Z(n4565) );
  CLKBUF_X1 U3582 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n5137) );
  AND2_X1 U3583 ( .A1(n3455), .A2(n3433), .ZN(n3427) );
  AND2_X1 U3584 ( .A1(n3432), .A2(n3433), .ZN(n5699) );
  OR2_X1 U3585 ( .A1(n4854), .A2(n4794), .ZN(n3428) );
  OR2_X1 U3586 ( .A1(n4802), .A2(n4794), .ZN(n4855) );
  INV_X1 U3587 ( .A(n5985), .ZN(n3429) );
  NAND2_X1 U3588 ( .A1(n3430), .A2(n6657), .ZN(n6198) );
  NOR2_X1 U3589 ( .A1(n6195), .A2(n3429), .ZN(n3430) );
  OR2_X1 U3590 ( .A1(n5649), .A2(n4311), .ZN(n3431) );
  OR2_X1 U3591 ( .A1(n5628), .A2(n4311), .ZN(n5650) );
  AND2_X1 U3592 ( .A1(n6655), .A2(n6654), .ZN(n6657) );
  NAND2_X1 U3593 ( .A1(n5648), .A2(n3435), .ZN(n3432) );
  OR2_X1 U3594 ( .A1(n3434), .A2(n3457), .ZN(n3433) );
  INV_X1 U3595 ( .A(n5700), .ZN(n3434) );
  AND2_X1 U3596 ( .A1(n5647), .A2(n5700), .ZN(n3435) );
  NAND2_X1 U3597 ( .A1(n5706), .A2(n5705), .ZN(n5956) );
  NAND2_X1 U3598 ( .A1(n3766), .A2(n3765), .ZN(n3436) );
  NAND2_X1 U3599 ( .A1(n3766), .A2(n3765), .ZN(n3801) );
  NOR2_X1 U3600 ( .A1(n4860), .A2(n6764), .ZN(n4388) );
  AND2_X1 U3601 ( .A1(n4470), .A2(n3588), .ZN(n3589) );
  NAND2_X1 U3602 ( .A1(n3437), .A2(n3438), .ZN(n5487) );
  AND2_X1 U3603 ( .A1(n5489), .A2(n5453), .ZN(n3438) );
  AND2_X1 U3604 ( .A1(n3607), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3439) );
  OAI211_X2 U3605 ( .C1(n4254), .C2(n3606), .A(n4663), .B(n5175), .ZN(n3607)
         );
  NAND2_X2 U3606 ( .A1(n3593), .A2(n3700), .ZN(n3623) );
  NAND2_X1 U3607 ( .A1(n3815), .A2(n3814), .ZN(n3847) );
  OAI22_X2 U3608 ( .A1(n4488), .A2(n4487), .B1(n4460), .B2(n4701), .ZN(n6062)
         );
  INV_X1 U3609 ( .A(n5991), .ZN(n3441) );
  INV_X1 U3610 ( .A(n5991), .ZN(n5992) );
  NAND2_X2 U3611 ( .A1(n3605), .A2(n3604), .ZN(n5175) );
  AND2_X4 U3612 ( .A1(n5146), .A2(n5139), .ZN(n3658) );
  INV_X1 U3613 ( .A(n4765), .ZN(n3442) );
  BUF_X2 U3614 ( .A(n3699), .Z(n4765) );
  NOR3_X2 U3615 ( .A1(n4765), .A2(n4687), .A3(n3587), .ZN(n3596) );
  INV_X1 U3616 ( .A(n3587), .ZN(n3594) );
  AND2_X2 U3617 ( .A1(n3468), .A2(n5139), .ZN(n3643) );
  AND3_X1 U3618 ( .A1(n3491), .A2(n3490), .A3(n3489), .ZN(n3492) );
  INV_X1 U3619 ( .A(n3586), .ZN(n3443) );
  INV_X1 U3620 ( .A(n3443), .ZN(n3444) );
  NAND2_X1 U3621 ( .A1(n3593), .A2(n3622), .ZN(n3586) );
  NOR2_X2 U3622 ( .A1(n6198), .A2(n4348), .ZN(n5981) );
  NAND2_X1 U3623 ( .A1(n3981), .A2(n3980), .ZN(n5677) );
  AND2_X1 U3624 ( .A1(n3734), .A2(n3614), .ZN(n3445) );
  AOI22_X1 U3625 ( .A1(n3636), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3448), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3469) );
  NAND4_X4 U3626 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3587)
         );
  AND2_X4 U3627 ( .A1(n4843), .A2(n5164), .ZN(n3563) );
  AND2_X1 U3628 ( .A1(n5146), .A2(n5139), .ZN(n3446) );
  AND2_X1 U3629 ( .A1(n5146), .A2(n5139), .ZN(n3447) );
  BUF_X4 U3630 ( .A(n4396), .Z(n5210) );
  AOI22_X1 U3631 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n3683), .B1(n3563), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3465) );
  AND2_X4 U3632 ( .A1(n3738), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5140)
         );
  AND2_X2 U3633 ( .A1(n3699), .A2(n3700), .ZN(n3600) );
  INV_X2 U3634 ( .A(n3699), .ZN(n3593) );
  AND2_X4 U3635 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5164) );
  NOR2_X4 U3636 ( .A1(n5779), .A2(n5801), .ZN(n5868) );
  AND2_X1 U3637 ( .A1(n5139), .A2(n5164), .ZN(n3448) );
  AND2_X2 U3638 ( .A1(n5139), .A2(n5164), .ZN(n3449) );
  NAND2_X2 U3639 ( .A1(n3668), .A2(n3450), .ZN(n3733) );
  OAI21_X2 U3640 ( .B1(n4837), .B2(STATE2_REG_0__SCAN_IN), .A(n3652), .ZN(
        n3727) );
  CLKBUF_X1 U3641 ( .A(n3683), .Z(n4582) );
  CLKBUF_X2 U3642 ( .A(n3563), .Z(n4603) );
  INV_X1 U3643 ( .A(n3799), .ZN(n3800) );
  CLKBUF_X1 U3644 ( .A(n3751), .Z(n4614) );
  CLKBUF_X1 U3645 ( .A(n3674), .Z(n4611) );
  XNOR2_X1 U3646 ( .A(n5171), .B(n5172), .ZN(n4912) );
  OR2_X1 U3647 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  AND2_X1 U3648 ( .A1(n6122), .A2(n4721), .ZN(n6145) );
  NAND2_X1 U3649 ( .A1(n3583), .A2(n3602), .ZN(n3621) );
  AND2_X1 U3650 ( .A1(n3627), .A2(n3604), .ZN(n3557) );
  CLKBUF_X1 U3651 ( .A(n3674), .Z(n4560) );
  CLKBUF_X1 U3652 ( .A(n3683), .Z(n3749) );
  OR2_X1 U3653 ( .A1(n3763), .A2(n3762), .ZN(n4389) );
  AOI22_X1 U3654 ( .A1(n3642), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3475) );
  INV_X1 U3655 ( .A(n3874), .ZN(n3880) );
  OAI21_X1 U3656 ( .B1(n6080), .B2(n4466), .A(n4465), .ZN(n4488) );
  AND2_X1 U3657 ( .A1(n6106), .A2(n4454), .ZN(n4455) );
  NAND2_X1 U3658 ( .A1(n3870), .A2(n3869), .ZN(n4449) );
  INV_X1 U3659 ( .A(n3868), .ZN(n3869) );
  OR2_X1 U3660 ( .A1(n4836), .A2(n4835), .ZN(n5169) );
  NAND2_X1 U3661 ( .A1(n3791), .A2(n3790), .ZN(n3799) );
  OAI21_X1 U3662 ( .B1(n7070), .B2(n7058), .A(n5767), .ZN(n4923) );
  OR2_X1 U3663 ( .A1(n6739), .A2(n4266), .ZN(n5826) );
  INV_X1 U3664 ( .A(n4767), .ZN(n5861) );
  INV_X1 U3665 ( .A(n4179), .ZN(n5865) );
  NAND2_X1 U3666 ( .A1(n5917), .A2(n4371), .ZN(n5973) );
  INV_X1 U3667 ( .A(n5715), .ZN(n4013) );
  AND2_X1 U3668 ( .A1(n3914), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3938)
         );
  INV_X1 U3669 ( .A(n5190), .ZN(n3896) );
  OR2_X1 U3670 ( .A1(n3840), .A2(n3843), .ZN(n3875) );
  NOR2_X1 U3671 ( .A1(n6790), .A2(n5631), .ZN(n5668) );
  AND2_X1 U3672 ( .A1(n5567), .A2(n6798), .ZN(n6754) );
  INV_X1 U3673 ( .A(n4374), .ZN(n4917) );
  NAND2_X1 U3674 ( .A1(n7072), .A2(n4923), .ZN(n5253) );
  INV_X1 U3675 ( .A(n5185), .ZN(n6229) );
  AND2_X1 U3676 ( .A1(n7062), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4255) );
  INV_X1 U3677 ( .A(n6663), .ZN(n5970) );
  NAND2_X1 U3678 ( .A1(n6663), .A2(n6006), .ZN(n6658) );
  NAND2_X1 U3679 ( .A1(n4911), .A2(n4817), .ZN(n6026) );
  AOI21_X1 U3680 ( .B1(n6693), .B2(n5822), .A(n4631), .ZN(n4632) );
  AOI21_X1 U3681 ( .B1(n6693), .B2(n5757), .A(n4482), .ZN(n4483) );
  NAND2_X1 U3682 ( .A1(n5973), .A2(n4372), .ZN(n5759) );
  OR2_X1 U3683 ( .A1(n4371), .A2(n5917), .ZN(n4372) );
  NAND2_X1 U3684 ( .A1(n6101), .A2(n4862), .ZN(n6717) );
  INV_X1 U3685 ( .A(n6707), .ZN(n6101) );
  INV_X1 U3686 ( .A(n6717), .ZN(n6693) );
  AND2_X2 U3687 ( .A1(n6696), .A2(n4477), .ZN(n6707) );
  XNOR2_X1 U3688 ( .A(n4493), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6141)
         );
  NAND2_X1 U3689 ( .A1(n4492), .A2(n4491), .ZN(n4493) );
  OR2_X1 U3690 ( .A1(n6031), .A2(n4460), .ZN(n4492) );
  NOR2_X1 U3691 ( .A1(n6179), .A2(n4719), .ZN(n6169) );
  NAND2_X1 U3692 ( .A1(n4706), .A2(n4667), .ZN(n6793) );
  INV_X1 U3693 ( .A(n6793), .ZN(n6860) );
  NAND2_X1 U3694 ( .A1(n3708), .A2(n3707), .ZN(n3709) );
  NAND2_X1 U3695 ( .A1(n3705), .A2(n3706), .ZN(n3710) );
  INV_X1 U3696 ( .A(n3706), .ZN(n3708) );
  INV_X1 U3697 ( .A(n4917), .ZN(n5415) );
  INV_X1 U3698 ( .A(n6327), .ZN(n5797) );
  OR2_X1 U3699 ( .A1(n6327), .A2(n7132), .ZN(n5794) );
  NOR2_X1 U3700 ( .A1(n4687), .A2(n3527), .ZN(n3526) );
  NOR2_X1 U3701 ( .A1(n3585), .A2(n3621), .ZN(n4470) );
  OR2_X1 U3702 ( .A1(n4213), .A2(n5349), .ZN(n4229) );
  NAND3_X1 U3703 ( .A1(n4474), .A2(n3600), .A3(n4687), .ZN(n3601) );
  CLKBUF_X1 U3704 ( .A(n3750), .Z(n3657) );
  CLKBUF_X1 U3705 ( .A(n3756), .Z(n3644) );
  AND2_X1 U3706 ( .A1(n6106), .A2(n6105), .ZN(n4461) );
  OR2_X1 U3707 ( .A1(n3811), .A2(n3810), .ZN(n4413) );
  CLKBUF_X1 U3708 ( .A(n4470), .Z(n4471) );
  NAND2_X1 U3709 ( .A1(n4204), .A2(n4203), .ZN(n4264) );
  NAND2_X1 U3710 ( .A1(n3505), .A2(n5734), .ZN(n3598) );
  AOI22_X1 U3711 ( .A1(n3676), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3683), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3479) );
  AND2_X1 U3712 ( .A1(n4556), .A2(n5905), .ZN(n5778) );
  AND2_X2 U3713 ( .A1(n3527), .A2(n3622), .ZN(n4474) );
  OR2_X1 U3714 ( .A1(n3859), .A2(n3858), .ZN(n4438) );
  OR2_X1 U3715 ( .A1(n3789), .A2(n3788), .ZN(n4400) );
  OR2_X1 U3716 ( .A1(n3689), .A2(n3688), .ZN(n4383) );
  NAND2_X1 U3717 ( .A1(n3734), .A2(n3614), .ZN(n3732) );
  INV_X1 U3718 ( .A(n6230), .ZN(n5104) );
  AND2_X1 U3719 ( .A1(n5160), .A2(n5159), .ZN(n7030) );
  NAND2_X1 U3720 ( .A1(n4239), .A2(n4435), .ZN(n4251) );
  CLKBUF_X1 U3721 ( .A(n4257), .Z(n4258) );
  AND2_X1 U3722 ( .A1(n4317), .A2(n4316), .ZN(n5705) );
  AND2_X1 U3723 ( .A1(n4293), .A2(n4292), .ZN(n5024) );
  NOR2_X1 U3724 ( .A1(n4750), .A2(READY_N), .ZN(n4754) );
  OR2_X1 U3725 ( .A1(n4547), .A2(n4548), .ZN(n4495) );
  OR2_X1 U3726 ( .A1(n4495), .A2(n4494), .ZN(n4557) );
  NOR2_X1 U3727 ( .A1(n4190), .A2(n4189), .ZN(n4535) );
  NOR2_X1 U3728 ( .A1(n4104), .A2(n4117), .ZN(n4151) );
  NOR2_X1 U3729 ( .A1(n4067), .A2(n4066), .ZN(n4068) );
  AND2_X1 U3730 ( .A1(n4068), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4103)
         );
  INV_X1 U3731 ( .A(n6652), .ZN(n4086) );
  AND2_X1 U3732 ( .A1(n4043), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4044)
         );
  NAND2_X1 U3733 ( .A1(n4044), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4067)
         );
  CLKBUF_X1 U3734 ( .A(n5946), .Z(n5947) );
  NOR2_X1 U3735 ( .A1(n4015), .A2(n5725), .ZN(n4043) );
  NAND2_X1 U3736 ( .A1(n3996), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4015)
         );
  NOR2_X1 U3737 ( .A1(n3992), .A2(n6946), .ZN(n3996) );
  NAND2_X1 U3738 ( .A1(n5608), .A2(n3979), .ZN(n3980) );
  NOR2_X1 U3739 ( .A1(n3943), .A2(n3939), .ZN(n3974) );
  NAND2_X1 U3740 ( .A1(n3938), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3943)
         );
  CLKBUF_X1 U3741 ( .A(n5487), .Z(n5488) );
  NOR2_X1 U3742 ( .A1(n3899), .A2(n3898), .ZN(n3914) );
  AND3_X1 U3743 ( .A1(n3895), .A2(n3894), .A3(n3893), .ZN(n5190) );
  NAND2_X1 U3744 ( .A1(n3882), .A2(n3881), .ZN(n5022) );
  NOR2_X1 U3745 ( .A1(n3880), .A2(n3879), .ZN(n3881) );
  NOR2_X1 U3746 ( .A1(n3878), .A2(n4623), .ZN(n3879) );
  INV_X1 U3747 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3843) );
  INV_X1 U3748 ( .A(n3821), .ZN(n3820) );
  INV_X1 U3750 ( .A(n3792), .ZN(n3793) );
  NAND2_X1 U3751 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3793), .ZN(n3821)
         );
  NAND2_X1 U3752 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3792) );
  NOR2_X1 U3753 ( .A1(n6106), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6029)
         );
  AND2_X1 U3754 ( .A1(n6106), .A2(n6051), .ZN(n4636) );
  AND2_X1 U3755 ( .A1(n6106), .A2(n4457), .ZN(n4458) );
  AND2_X1 U3756 ( .A1(n4310), .A2(n4309), .ZN(n5627) );
  AND2_X1 U3757 ( .A1(n5456), .A2(n5455), .ZN(n5491) );
  AND2_X1 U3758 ( .A1(n4305), .A2(n4304), .ZN(n5490) );
  AOI22_X1 U3759 ( .A1(n5581), .A2(n5582), .B1(n4460), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5562) );
  NOR2_X2 U3760 ( .A1(n5419), .A2(n5420), .ZN(n5456) );
  AOI21_X1 U3761 ( .B1(n5586), .B2(n5588), .A(n4444), .ZN(n5437) );
  AND2_X1 U3762 ( .A1(n4443), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4444)
         );
  AND2_X1 U3763 ( .A1(n4291), .A2(n4290), .ZN(n4807) );
  NAND2_X1 U3764 ( .A1(n4706), .A2(n5843), .ZN(n6798) );
  AND2_X1 U3765 ( .A1(n5859), .A2(n4679), .ZN(n4823) );
  CLKBUF_X1 U3766 ( .A(n4912), .Z(n4913) );
  CLKBUF_X1 U3767 ( .A(n3591), .Z(n3592) );
  INV_X1 U3768 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3463) );
  NAND2_X1 U3769 ( .A1(n3779), .A2(n3778), .ZN(n5172) );
  AND2_X1 U3770 ( .A1(n5263), .A2(n5030), .ZN(n5090) );
  INV_X1 U3771 ( .A(n5527), .ZN(n5217) );
  NAND2_X1 U3772 ( .A1(n5210), .A2(n4917), .ZN(n6230) );
  AND2_X1 U3773 ( .A1(n4952), .A2(n5209), .ZN(n5255) );
  NAND2_X1 U3774 ( .A1(n7063), .A2(n4923), .ZN(n5252) );
  AOI21_X1 U3775 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7020), .A(n5253), .ZN(
        n7143) );
  NAND2_X1 U3776 ( .A1(n4750), .A2(n4731), .ZN(n6739) );
  NAND2_X1 U3777 ( .A1(n5872), .A2(n4360), .ZN(n6986) );
  INV_X1 U3778 ( .A(n6978), .ZN(n7007) );
  AND2_X1 U3779 ( .A1(n6038), .A2(n4363), .ZN(n6981) );
  INV_X1 U3780 ( .A(n6999), .ZN(n6968) );
  INV_X1 U3781 ( .A(n6001), .ZN(n6660) );
  INV_X1 U3782 ( .A(n6658), .ZN(n6649) );
  NAND2_X1 U3783 ( .A1(n4770), .A2(n4769), .ZN(n6663) );
  OR2_X1 U3784 ( .A1(n4834), .A2(n7077), .ZN(n4770) );
  INV_X1 U3785 ( .A(n6026), .ZN(n7116) );
  AND2_X1 U3786 ( .A1(n6026), .A2(n5735), .ZN(n7117) );
  NAND2_X1 U3787 ( .A1(n6026), .A2(n4819), .ZN(n6027) );
  INV_X1 U3788 ( .A(n5973), .ZN(n5975) );
  OR2_X1 U3789 ( .A1(n4697), .A2(n5567), .ZN(n6790) );
  AND2_X1 U3790 ( .A1(n4706), .A2(n5814), .ZN(n6858) );
  CLKBUF_X1 U3791 ( .A(n3712), .Z(n5800) );
  INV_X1 U3792 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5523) );
  INV_X1 U3794 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5181) );
  AND2_X1 U3795 ( .A1(n5180), .A2(n5253), .ZN(n6327) );
  INV_X1 U3796 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5818) );
  CLKBUF_X1 U3797 ( .A(n3738), .Z(n3739) );
  NOR2_X1 U3799 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n7055) );
  INV_X1 U3800 ( .A(n5255), .ZN(n5321) );
  AND2_X1 U3801 ( .A1(n5090), .A2(n4386), .ZN(n5304) );
  INV_X1 U3802 ( .A(n5220), .ZN(n5472) );
  NOR2_X1 U3803 ( .A1(n5184), .A2(n4998), .ZN(n7207) );
  INV_X1 U3804 ( .A(n7147), .ZN(n7211) );
  INV_X1 U3805 ( .A(n6279), .ZN(n7159) );
  INV_X1 U3806 ( .A(n6291), .ZN(n7175) );
  INV_X1 U3807 ( .A(n6297), .ZN(n7183) );
  INV_X1 U3808 ( .A(n6303), .ZN(n7191) );
  INV_X1 U3809 ( .A(n6309), .ZN(n7199) );
  AND2_X1 U3810 ( .A1(n7046), .A2(n7045), .ZN(n7078) );
  NOR2_X1 U3811 ( .A1(n5854), .A2(n7066), .ZN(n7069) );
  INV_X1 U3812 ( .A(n7068), .ZN(n7067) );
  INV_X1 U3813 ( .A(n4632), .ZN(n4633) );
  INV_X1 U3814 ( .A(n6073), .ZN(n6078) );
  OAI21_X1 U3815 ( .B1(n6194), .B2(n6696), .A(n4483), .ZN(n4484) );
  AND2_X1 U3816 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  INV_X2 U3817 ( .A(n4640), .ZN(n4460) );
  INV_X2 U3818 ( .A(n4460), .ZN(n6106) );
  INV_X1 U3819 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6226) );
  OR2_X1 U3820 ( .A1(n4917), .A2(n4010), .ZN(n3452) );
  NAND2_X1 U3821 ( .A1(n5992), .A2(n4086), .ZN(n5987) );
  INV_X1 U3822 ( .A(n6696), .ZN(n6714) );
  NOR2_X1 U3823 ( .A1(n4765), .A2(n6226), .ZN(n3973) );
  INV_X1 U3824 ( .A(n3973), .ZN(n4010) );
  XNOR2_X1 U3825 ( .A(n3732), .B(n3733), .ZN(n4837) );
  OR2_X1 U3826 ( .A1(n3700), .A2(n6226), .ZN(n3453) );
  INV_X1 U3827 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n7072) );
  OR2_X1 U3828 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4623) );
  NOR2_X4 U3829 ( .A1(n5350), .A2(n4366), .ZN(n7003) );
  NAND2_X1 U3830 ( .A1(n5826), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5350) );
  NOR3_X2 U3831 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n5266), .ZN(n5323) );
  NAND2_X1 U3832 ( .A1(n5648), .A2(n5647), .ZN(n5646) );
  INV_X1 U3833 ( .A(n3978), .ZN(n5608) );
  NAND2_X1 U3834 ( .A1(n4449), .A2(n4448), .ZN(n4640) );
  BUF_X1 U3835 ( .A(n4087), .Z(n4497) );
  AND2_X1 U3836 ( .A1(n4460), .A2(n4456), .ZN(n3454) );
  OR2_X1 U3837 ( .A1(n4460), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3455)
         );
  OR2_X1 U3838 ( .A1(n4460), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3456)
         );
  OR2_X1 U3839 ( .A1(n4460), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3457)
         );
  XOR2_X1 U3840 ( .A(n6106), .B(n5776), .Z(n3458) );
  OR2_X1 U3841 ( .A1(n6914), .A2(n4349), .ZN(n3459) );
  AND2_X1 U3842 ( .A1(n3660), .A2(n3659), .ZN(n3461) );
  OR2_X1 U3843 ( .A1(n5759), .A2(n6121), .ZN(n3462) );
  INV_X1 U3844 ( .A(n4257), .ZN(n3605) );
  INV_X1 U3845 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4200) );
  INV_X1 U3846 ( .A(n4751), .ZN(n4212) );
  NOR2_X1 U3847 ( .A1(n5854), .A2(READY_N), .ZN(n4826) );
  INV_X1 U3848 ( .A(n5993), .ZN(n4064) );
  OR2_X1 U3849 ( .A1(n3815), .A2(n3814), .ZN(n3816) );
  INV_X1 U3850 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4462) );
  OR2_X1 U3851 ( .A1(n3837), .A2(n3836), .ZN(n4422) );
  AOI22_X1 U3852 ( .A1(n3676), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3683), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3487) );
  INV_X1 U3853 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4243) );
  INV_X1 U3854 ( .A(n5509), .ZN(n4432) );
  AND2_X2 U3855 ( .A1(n3591), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4843)
         );
  AOI22_X1 U3856 ( .A1(n4247), .A2(n4400), .B1(n4239), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U3857 ( .A1(n3676), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3683), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3501) );
  OR2_X1 U3858 ( .A1(n4244), .A2(n4243), .ZN(n4242) );
  AND2_X2 U3859 ( .A1(n4843), .A2(n5140), .ZN(n3682) );
  OR2_X1 U3860 ( .A1(n4841), .A2(n7072), .ZN(n4596) );
  INV_X1 U3861 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3898) );
  OR2_X1 U3862 ( .A1(n4408), .A2(n4010), .ZN(n3827) );
  XNOR2_X1 U3863 ( .A(n3727), .B(n3728), .ZN(n3726) );
  INV_X1 U3864 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4637) );
  NAND2_X1 U3865 ( .A1(n4654), .A2(n4733), .ZN(n4254) );
  INV_X1 U3866 ( .A(n4242), .ZN(n4204) );
  INV_X1 U3867 ( .A(n5350), .ZN(n5872) );
  NAND2_X1 U3868 ( .A1(n5859), .A2(n4767), .ZN(n4675) );
  AND2_X1 U3869 ( .A1(n5778), .A2(n5780), .ZN(n4576) );
  OR2_X1 U3870 ( .A1(n4578), .A2(n5880), .ZN(n4599) );
  NAND2_X1 U3871 ( .A1(n4535), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4547)
         );
  AND2_X1 U3872 ( .A1(n4378), .A2(n4751), .ZN(n4435) );
  INV_X1 U3873 ( .A(n4751), .ZN(n3604) );
  AND2_X1 U3874 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5264) );
  AND2_X1 U3875 ( .A1(n4913), .A2(n7146), .ZN(n5031) );
  OAI21_X1 U3876 ( .B1(n5553), .B2(n7066), .A(n5530), .ZN(n5552) );
  AND2_X1 U3877 ( .A1(n4913), .A2(n5811), .ZN(n7122) );
  NAND2_X1 U3878 ( .A1(n4103), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4104)
         );
  NOR2_X1 U3879 ( .A1(n3875), .A2(n3860), .ZN(n3876) );
  INV_X1 U3880 ( .A(n7003), .ZN(n6914) );
  AND4_X1 U3881 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3577)
         );
  NAND2_X1 U3882 ( .A1(n6031), .A2(n6029), .ZN(n4491) );
  NOR2_X1 U3883 ( .A1(n6042), .A2(n5774), .ZN(n5775) );
  AND2_X1 U3884 ( .A1(n5632), .A2(n5622), .ZN(n5567) );
  INV_X1 U3885 ( .A(n7069), .ZN(n5767) );
  INV_X1 U3886 ( .A(n4403), .ZN(n5263) );
  INV_X1 U3887 ( .A(n5253), .ZN(n4974) );
  AND2_X1 U3888 ( .A1(n4984), .A2(n4983), .ZN(n5334) );
  AND2_X2 U3889 ( .A1(n4212), .A2(n4733), .ZN(n5856) );
  OR2_X1 U3890 ( .A1(n4123), .A2(n4145), .ZN(n4190) );
  NOR2_X2 U3891 ( .A1(n5995), .A2(n5994), .ZN(n6655) );
  AND2_X1 U3892 ( .A1(n5685), .A2(REIP_REG_11__SCAN_IN), .ZN(n6953) );
  INV_X1 U3893 ( .A(n6986), .ZN(n6998) );
  NAND2_X1 U3894 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3899)
         );
  NOR2_X1 U3895 ( .A1(n5197), .A2(n6724), .ZN(n6967) );
  NAND2_X1 U3896 ( .A1(n5936), .A2(n5935), .ZN(n5938) );
  NAND2_X1 U3897 ( .A1(n6657), .A2(n5985), .ZN(n6196) );
  NOR2_X1 U3898 ( .A1(n4754), .A2(n4909), .ZN(n4867) );
  INV_X1 U3899 ( .A(n4911), .ZN(n4876) );
  AND2_X1 U3900 ( .A1(n5987), .A2(n6653), .ZN(n7107) );
  CLKBUF_X1 U3901 ( .A(n5021), .Z(n5191) );
  NAND2_X1 U3902 ( .A1(n3820), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3840)
         );
  NOR2_X1 U3903 ( .A1(n5668), .A2(n5618), .ZN(n6842) );
  CLKBUF_X1 U3904 ( .A(n5437), .Z(n5439) );
  AND2_X1 U3905 ( .A1(n4661), .A2(n7047), .ZN(n4706) );
  OR2_X1 U3906 ( .A1(n6858), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6755)
         );
  INV_X1 U3907 ( .A(n6800), .ZN(n6854) );
  OR2_X1 U3908 ( .A1(n5035), .A2(n5034), .ZN(n5319) );
  OAI211_X1 U3909 ( .C1(n5219), .C2(n5221), .A(n5218), .B(n5217), .ZN(n5468)
         );
  AND2_X1 U3910 ( .A1(n5054), .A2(n5263), .ZN(n5378) );
  INV_X1 U3911 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n7020) );
  OR2_X1 U3912 ( .A1(n4980), .A2(n4979), .ZN(n5333) );
  INV_X1 U3913 ( .A(n4386), .ZN(n5209) );
  INV_X1 U3914 ( .A(n7124), .ZN(n7202) );
  OR3_X1 U3915 ( .A1(n6260), .A2(n4922), .A3(n4921), .ZN(n5435) );
  AND2_X1 U3916 ( .A1(n7054), .A2(n7053), .ZN(n7068) );
  OR2_X1 U3917 ( .A1(n5854), .A2(n4256), .ZN(n4750) );
  INV_X1 U3918 ( .A(n6993), .ZN(n7004) );
  OR2_X1 U3919 ( .A1(n6038), .A2(n4362), .ZN(n6978) );
  INV_X1 U3920 ( .A(n6660), .ZN(n6005) );
  INV_X1 U3921 ( .A(n5504), .ZN(n5262) );
  OR2_X1 U3922 ( .A1(n5854), .A2(n4729), .ZN(n6572) );
  INV_X1 U3923 ( .A(n4484), .ZN(n4485) );
  OR2_X1 U3924 ( .A1(n6842), .A2(n4709), .ZN(n6753) );
  NAND2_X1 U3925 ( .A1(n4706), .A2(n4666), .ZN(n6800) );
  INV_X1 U3926 ( .A(n4913), .ZN(n5214) );
  INV_X1 U3927 ( .A(n5304), .ZN(n5326) );
  NAND2_X1 U3928 ( .A1(n5090), .A2(n5209), .ZN(n5475) );
  OR2_X1 U3929 ( .A1(n5087), .A2(n5209), .ZN(n5339) );
  INV_X1 U3930 ( .A(n6273), .ZN(n7151) );
  INV_X1 U3931 ( .A(n6285), .ZN(n7167) );
  INV_X1 U3932 ( .A(n6316), .ZN(n7216) );
  AND2_X1 U3933 ( .A1(n6268), .A2(n6267), .ZN(n6325) );
  AND2_X1 U3934 ( .A1(n7143), .A2(n4951), .ZN(n5261) );
  INV_X1 U3935 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n7062) );
  AND2_X1 U3936 ( .A1(STATE_REG_1__SCAN_IN), .A2(n4357), .ZN(n7099) );
  OR2_X1 U3937 ( .A1(n4370), .A2(n4369), .ZN(U2803) );
  NAND2_X1 U3938 ( .A1(n3462), .A2(n4485), .ZN(U2964) );
  AND2_X4 U3939 ( .A1(n3463), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4842)
         );
  INV_X1 U3940 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3738) );
  AND2_X4 U3941 ( .A1(n4842), .A2(n5140), .ZN(n4087) );
  INV_X1 U3942 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3773) );
  AND2_X2 U3943 ( .A1(n3773), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3468)
         );
  AND2_X4 U3944 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5139) );
  AOI22_X1 U3945 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n4087), .B1(n3643), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3467) );
  AND2_X2 U3946 ( .A1(n4842), .A2(n5164), .ZN(n3642) );
  INV_X1 U3947 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3591) );
  AND2_X4 U3948 ( .A1(n3468), .A2(n4843), .ZN(n3674) );
  AOI22_X2 U3949 ( .A1(n3642), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3466) );
  AND2_X4 U3950 ( .A1(n5140), .A2(n5139), .ZN(n3683) );
  NOR2_X4 U3951 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5167) );
  AND2_X2 U3952 ( .A1(n5167), .A2(n5164), .ZN(n3645) );
  AOI22_X1 U3953 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n3682), .B1(n3645), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3464) );
  NAND4_X1 U3954 ( .A1(n3467), .A2(n3466), .A3(n3465), .A4(n3464), .ZN(n3474)
         );
  AND2_X4 U3955 ( .A1(n5140), .A2(n5167), .ZN(n3676) );
  AOI22_X2 U3956 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n3756), .B1(n3676), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3472) );
  NOR2_X4 U3957 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5146) );
  AND2_X2 U3958 ( .A1(n4843), .A2(n5146), .ZN(n3572) );
  AND2_X2 U3959 ( .A1(n5167), .A2(n5146), .ZN(n3637) );
  AOI22_X1 U3960 ( .A1(n3572), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3471) );
  AND2_X2 U3961 ( .A1(n4842), .A2(n5146), .ZN(n3636) );
  NAND4_X1 U3962 ( .A1(n3472), .A2(n3471), .A3(n3470), .A4(n3469), .ZN(n3473)
         );
  OR2_X2 U3963 ( .A1(n3474), .A2(n3473), .ZN(n3699) );
  AOI22_X1 U3964 ( .A1(n4087), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3478) );
  AOI22_X1 U3965 ( .A1(n3572), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U3966 ( .A1(n3750), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U3967 ( .A1(n3682), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3563), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U3968 ( .A1(n3636), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U3969 ( .A1(n3756), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3480) );
  NAND2_X4 U3970 ( .A1(n3484), .A2(n3483), .ZN(n3700) );
  INV_X1 U3971 ( .A(n3600), .ZN(n5733) );
  AOI22_X1 U3972 ( .A1(n3642), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3682), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U3973 ( .A1(n3756), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U3974 ( .A1(n3637), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U3975 ( .A1(n4087), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U3976 ( .A1(n3674), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3491) );
  AOI22_X1 U3977 ( .A1(n3750), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3572), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3490) );
  AOI22_X1 U3978 ( .A1(n3636), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3563), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3489) );
  NAND3_X2 U3979 ( .A1(n3494), .A2(n3493), .A3(n3492), .ZN(n4687) );
  INV_X1 U3980 ( .A(n4687), .ZN(n3505) );
  AOI22_X1 U3981 ( .A1(n3642), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3756), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U3982 ( .A1(n4087), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U3983 ( .A1(n3636), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U3984 ( .A1(n3750), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U3985 ( .A1(n3682), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3563), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3502) );
  AOI22_X1 U3986 ( .A1(n3674), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3500) );
  AOI22_X1 U3987 ( .A1(n3572), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3499) );
  NAND2_X1 U3988 ( .A1(n4087), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3509)
         );
  NAND2_X1 U3989 ( .A1(n3643), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U3990 ( .A1(n3642), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3507)
         );
  NAND2_X1 U3991 ( .A1(n3674), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U3992 ( .A1(n3756), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3513) );
  NAND2_X1 U3993 ( .A1(n3636), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U3994 ( .A1(n3676), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U3995 ( .A1(n3449), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3510)
         );
  AND4_X2 U3996 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3524)
         );
  NAND2_X1 U3997 ( .A1(n3682), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U3998 ( .A1(n3683), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3516)
         );
  NAND2_X1 U3999 ( .A1(n3563), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3515)
         );
  NAND2_X1 U4000 ( .A1(n3645), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3514)
         );
  AND4_X2 U4001 ( .A1(n3517), .A2(n3516), .A3(n3515), .A4(n3514), .ZN(n3523)
         );
  NAND2_X1 U4002 ( .A1(n3750), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3521) );
  NAND2_X1 U4003 ( .A1(n3572), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3520) );
  NAND2_X1 U4004 ( .A1(n3637), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3519) );
  NAND2_X1 U4005 ( .A1(n3446), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3518) );
  AND4_X2 U4006 ( .A1(n3521), .A2(n3520), .A3(n3519), .A4(n3518), .ZN(n3522)
         );
  NAND2_X1 U4007 ( .A1(n3711), .A2(n3526), .ZN(n3628) );
  OAI211_X1 U4008 ( .C1(n5733), .C2(n3598), .A(n3628), .B(n3601), .ZN(n3558)
         );
  AOI22_X1 U4009 ( .A1(n4087), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3643), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3531) );
  AOI22_X1 U4010 ( .A1(n3642), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3674), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3530) );
  AOI22_X1 U4011 ( .A1(n3563), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3683), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4012 ( .A1(n3682), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3645), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4013 ( .A1(n3572), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3637), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3535) );
  AOI22_X1 U4014 ( .A1(n3756), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3534) );
  AOI22_X1 U4015 ( .A1(n3750), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3533) );
  AOI22_X1 U4016 ( .A1(n3636), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3532) );
  NAND2_X1 U4017 ( .A1(n3682), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U4018 ( .A1(n3643), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3539) );
  NAND2_X1 U4019 ( .A1(n3683), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3538)
         );
  NAND2_X1 U4020 ( .A1(n3563), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3537)
         );
  NAND2_X1 U4021 ( .A1(n4087), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3544)
         );
  NAND2_X1 U4022 ( .A1(n3642), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3543)
         );
  NAND2_X1 U4023 ( .A1(n3674), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3542) );
  NAND2_X1 U4024 ( .A1(n3645), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3541)
         );
  NAND2_X1 U4025 ( .A1(n3750), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4026 ( .A1(n3756), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3547) );
  NAND2_X1 U4027 ( .A1(n3572), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3546) );
  NAND2_X1 U4028 ( .A1(n3637), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3545) );
  NAND2_X1 U4029 ( .A1(n3636), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3552) );
  NAND2_X1 U4030 ( .A1(n3676), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3551) );
  NAND2_X1 U4031 ( .A1(n3449), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3550)
         );
  NAND2_X1 U4032 ( .A1(n3658), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3549) );
  NAND4_X4 U4033 ( .A1(n3556), .A2(n3555), .A3(n3554), .A4(n3553), .ZN(n4751)
         );
  NAND2_X1 U4034 ( .A1(n3558), .A2(n3557), .ZN(n3581) );
  NAND2_X1 U4035 ( .A1(n4087), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3562)
         );
  NAND2_X1 U4036 ( .A1(n3643), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3561) );
  NAND2_X1 U4037 ( .A1(n3642), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3560)
         );
  NAND2_X1 U4038 ( .A1(n3674), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4039 ( .A1(n3682), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3567) );
  NAND2_X1 U4040 ( .A1(n3683), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3566)
         );
  NAND2_X1 U4041 ( .A1(n3563), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3565)
         );
  NAND2_X1 U4042 ( .A1(n3645), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3564)
         );
  NAND2_X1 U4043 ( .A1(n3636), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3571) );
  NAND2_X1 U4044 ( .A1(n3756), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3570) );
  NAND2_X1 U4045 ( .A1(n3676), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3569) );
  NAND2_X1 U4046 ( .A1(n3751), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3568)
         );
  NAND2_X1 U4047 ( .A1(n3750), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U4048 ( .A1(n3572), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4049 ( .A1(n3637), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3574) );
  NAND2_X1 U4050 ( .A1(n3658), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3573) );
  NAND4_X4 U4051 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n4733)
         );
  INV_X1 U4052 ( .A(n3586), .ZN(n3582) );
  NAND2_X1 U4053 ( .A1(n3582), .A2(n3594), .ZN(n3583) );
  NAND2_X1 U4054 ( .A1(n3700), .A2(n3622), .ZN(n3584) );
  NAND2_X1 U4055 ( .A1(n3595), .A2(n4377), .ZN(n3585) );
  NAND2_X1 U4056 ( .A1(n3444), .A2(n3460), .ZN(n3588) );
  INV_X1 U4057 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6731) );
  XNOR2_X1 U4058 ( .A(n6731), .B(STATE_REG_2__SCAN_IN), .ZN(n4358) );
  NOR2_X1 U4059 ( .A1(n4751), .A2(n4358), .ZN(n3606) );
  NAND2_X1 U4060 ( .A1(n3595), .A2(n3594), .ZN(n4649) );
  OAI21_X1 U4061 ( .B1(n3606), .B2(n4378), .A(n3634), .ZN(n3590) );
  OAI21_X2 U4062 ( .B1(n4698), .B2(n3590), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3736) );
  OR2_X2 U4063 ( .A1(n3736), .A2(n3592), .ZN(n3610) );
  INV_X1 U4064 ( .A(n3627), .ZN(n3597) );
  AND3_X2 U4065 ( .A1(n3597), .A2(n3596), .A3(n3595), .ZN(n4654) );
  INV_X1 U4066 ( .A(n3598), .ZN(n3599) );
  AND2_X2 U4067 ( .A1(n4768), .A2(n5349), .ZN(n4693) );
  NAND2_X1 U4068 ( .A1(n4693), .A2(n3600), .ZN(n4663) );
  INV_X1 U4069 ( .A(n3601), .ZN(n3603) );
  NAND2_X1 U4070 ( .A1(n3603), .A2(n3630), .ZN(n4257) );
  NAND2_X1 U4071 ( .A1(n3607), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3612) );
  NOR2_X1 U4072 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3608) );
  NOR2_X1 U4073 ( .A1(n5264), .A2(n3608), .ZN(n5521) );
  NAND2_X1 U4074 ( .A1(n7055), .A2(n7072), .ZN(n4476) );
  INV_X1 U4075 ( .A(n4476), .ZN(n3777) );
  INV_X1 U4076 ( .A(n4255), .ZN(n3776) );
  AOI22_X1 U4077 ( .A1(n5521), .A2(n3777), .B1(n3776), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3611) );
  AND2_X2 U4078 ( .A1(n3612), .A2(n3611), .ZN(n3609) );
  NAND2_X2 U4079 ( .A1(n3610), .A2(n3609), .ZN(n3734) );
  INV_X1 U4080 ( .A(n3611), .ZN(n3613) );
  MUX2_X1 U4081 ( .A(n4476), .B(n4255), .S(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), 
        .Z(n3615) );
  INV_X1 U4082 ( .A(n3616), .ZN(n3618) );
  NAND2_X1 U4083 ( .A1(n4435), .A2(n3594), .ZN(n3617) );
  NAND2_X1 U4084 ( .A1(n3618), .A2(n3617), .ZN(n3620) );
  NAND2_X1 U4085 ( .A1(n4687), .A2(n4733), .ZN(n3619) );
  NAND2_X1 U4086 ( .A1(n3620), .A2(n3619), .ZN(n4692) );
  INV_X1 U4087 ( .A(n3621), .ZN(n3625) );
  OR2_X1 U4088 ( .A1(n3623), .A2(n5734), .ZN(n4472) );
  NAND2_X1 U4089 ( .A1(n4649), .A2(n4472), .ZN(n3624) );
  NAND2_X1 U4090 ( .A1(n3625), .A2(n3624), .ZN(n3626) );
  NAND2_X1 U4091 ( .A1(n3626), .A2(n4751), .ZN(n3633) );
  NAND2_X1 U4092 ( .A1(n7055), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6721) );
  AOI21_X1 U4093 ( .B1(n3627), .B2(n5856), .A(n6721), .ZN(n3632) );
  NAND2_X1 U4095 ( .A1(n4016), .A2(n3630), .ZN(n3631) );
  NAND4_X1 U4096 ( .A1(n3634), .A2(n3633), .A3(n3632), .A4(n3631), .ZN(n3635)
         );
  NOR2_X1 U4097 ( .A1(n3587), .A2(n7072), .ZN(n3673) );
  AOI22_X1 U4098 ( .A1(n4497), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4099 ( .A1(n4602), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4100 ( .A1(n3563), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3639) );
  BUF_X1 U4101 ( .A(n3658), .Z(n4583) );
  AOI22_X1 U4102 ( .A1(n4565), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4103 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3651)
         );
  INV_X1 U4104 ( .A(n3643), .ZN(n5142) );
  AOI22_X1 U4105 ( .A1(n4110), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4106 ( .A1(n3644), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3648) );
  BUF_X1 U4107 ( .A(n3645), .Z(n3757) );
  AOI22_X1 U4109 ( .A1(n4612), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3647) );
  AOI22_X1 U4110 ( .A1(n4604), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3646) );
  NAND4_X1 U4111 ( .A1(n3649), .A2(n3648), .A3(n3647), .A4(n3646), .ZN(n3650)
         );
  NAND2_X1 U4112 ( .A1(n3673), .A2(n4375), .ZN(n3652) );
  NAND2_X1 U4113 ( .A1(n4239), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3667) );
  NAND3_X1 U4114 ( .A1(n4939), .A2(STATE2_REG_0__SCAN_IN), .A3(n4375), .ZN(
        n3666) );
  AOI22_X1 U4115 ( .A1(n4497), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4116 ( .A1(n4110), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4117 ( .A1(n3563), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3683), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4118 ( .A1(n4612), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4119 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3664)
         );
  AOI22_X1 U4120 ( .A1(n4602), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4121 ( .A1(n4604), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3661) );
  CLKBUF_X1 U4122 ( .A(n3756), .Z(n3675) );
  AOI22_X1 U4123 ( .A1(n3644), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3676), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3660) );
  AOI22_X1 U4124 ( .A1(n3657), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3659) );
  NAND3_X1 U4125 ( .A1(n3662), .A2(n3661), .A3(n3461), .ZN(n3663) );
  INV_X1 U4126 ( .A(n4445), .ZN(n3665) );
  NAND2_X1 U4127 ( .A1(n3673), .A2(n3665), .ZN(n3691) );
  INV_X1 U4128 ( .A(n3668), .ZN(n3670) );
  INV_X1 U4129 ( .A(n3450), .ZN(n3669) );
  NAND2_X1 U4130 ( .A1(n3670), .A2(n3669), .ZN(n3671) );
  NAND2_X1 U4131 ( .A1(n3671), .A2(n3733), .ZN(n3712) );
  INV_X1 U4132 ( .A(n3712), .ZN(n3672) );
  NAND2_X1 U4133 ( .A1(n3672), .A2(n7072), .ZN(n3704) );
  NAND2_X1 U4134 ( .A1(n3673), .A2(n4445), .ZN(n4447) );
  AOI22_X1 U4135 ( .A1(n4560), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4136 ( .A1(n3675), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4602), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4137 ( .A1(n3676), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3563), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3679) );
  CLKBUF_X1 U4138 ( .A(n3750), .Z(n3677) );
  AOI22_X1 U4139 ( .A1(n3677), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3678) );
  NAND4_X1 U4140 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3689)
         );
  AOI22_X1 U4141 ( .A1(n4110), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4142 ( .A1(n4612), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4143 ( .A1(n4565), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4144 ( .A1(n3749), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4145 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3688)
         );
  INV_X1 U4146 ( .A(n4383), .ZN(n3690) );
  NAND2_X1 U4147 ( .A1(n3704), .A2(n3706), .ZN(n3696) );
  NAND2_X1 U4148 ( .A1(n4239), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4149 ( .A1(n4939), .A2(n4383), .ZN(n3693) );
  NAND2_X1 U4150 ( .A1(n3594), .A2(n4445), .ZN(n3692) );
  NAND2_X1 U4151 ( .A1(n3696), .A2(n3707), .ZN(n3697) );
  NAND2_X1 U4152 ( .A1(n3697), .A2(n4447), .ZN(n3725) );
  INV_X1 U4153 ( .A(n3725), .ZN(n3698) );
  XNOR2_X1 U4154 ( .A(n3726), .B(n3698), .ZN(n4374) );
  INV_X2 U4155 ( .A(n3453), .ZN(n5866) );
  AOI22_X1 U4156 ( .A1(n5866), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6226), .ZN(n3702) );
  NAND2_X1 U4157 ( .A1(n3600), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3819) );
  INV_X1 U4158 ( .A(n3819), .ZN(n3719) );
  NAND2_X1 U4159 ( .A1(n3719), .A2(n5137), .ZN(n3701) );
  AND2_X1 U4160 ( .A1(n3702), .A2(n3701), .ZN(n3703) );
  NAND2_X1 U4161 ( .A1(n3704), .A2(n3707), .ZN(n3705) );
  AOI21_X1 U4162 ( .B1(n4386), .B2(n3711), .A(n6226), .ZN(n4813) );
  OR2_X1 U4163 ( .A1(n5800), .A2(n4010), .ZN(n3716) );
  AOI22_X1 U4164 ( .A1(n5866), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6226), .ZN(n3714) );
  NAND2_X1 U4165 ( .A1(n3719), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3713) );
  AND2_X1 U4166 ( .A1(n3714), .A2(n3713), .ZN(n3715) );
  NAND2_X1 U4167 ( .A1(n3716), .A2(n3715), .ZN(n4812) );
  NAND2_X1 U4168 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  INV_X1 U4169 ( .A(n4812), .ZN(n3717) );
  INV_X1 U4170 ( .A(n4623), .ZN(n4555) );
  NAND2_X1 U4171 ( .A1(n3717), .A2(n4555), .ZN(n3718) );
  NAND2_X1 U4172 ( .A1(n4811), .A2(n3718), .ZN(n4776) );
  NAND2_X1 U4173 ( .A1(n3719), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3724) );
  OAI21_X1 U4174 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3792), .ZN(n6671) );
  NAND2_X1 U4175 ( .A1(n6671), .A2(n4555), .ZN(n3721) );
  NAND2_X1 U4176 ( .A1(n6226), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4179) );
  NAND2_X1 U4177 ( .A1(n5865), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3720)
         );
  NAND2_X1 U4178 ( .A1(n3721), .A2(n3720), .ZN(n3722) );
  AOI21_X1 U4179 ( .B1(n5866), .B2(EAX_REG_2__SCAN_IN), .A(n3722), .ZN(n3723)
         );
  AND2_X1 U4180 ( .A1(n3724), .A2(n3723), .ZN(n3768) );
  NAND2_X1 U4181 ( .A1(n3726), .A2(n3725), .ZN(n3731) );
  INV_X1 U4182 ( .A(n3728), .ZN(n3729) );
  NAND2_X1 U4183 ( .A1(n3727), .A2(n3729), .ZN(n3730) );
  NAND2_X1 U4184 ( .A1(n3445), .A2(n3733), .ZN(n3735) );
  NAND2_X1 U4185 ( .A1(n3735), .A2(n3734), .ZN(n3746) );
  INV_X1 U4186 ( .A(n3746), .ZN(n3745) );
  OR2_X1 U4187 ( .A1(n3737), .A2(n3739), .ZN(n3743) );
  AND2_X1 U4188 ( .A1(n5264), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3774)
         );
  NOR2_X1 U4189 ( .A1(n5264), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3740)
         );
  NOR2_X1 U4190 ( .A1(n3774), .A2(n3740), .ZN(n4924) );
  NOR2_X1 U4191 ( .A1(n4255), .A2(n5181), .ZN(n3741) );
  AOI21_X1 U4192 ( .B1(n4924), .B2(n3777), .A(n3741), .ZN(n3742) );
  NAND2_X1 U4193 ( .A1(n3746), .A2(n3747), .ZN(n3748) );
  AOI22_X1 U4194 ( .A1(n4110), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4195 ( .A1(n4603), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4196 ( .A1(n3677), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4197 ( .A1(n4602), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4198 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3763)
         );
  INV_X2 U4199 ( .A(n5142), .ZN(n4606) );
  AOI22_X1 U4200 ( .A1(n4611), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4201 ( .A1(n3675), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4202 ( .A1(n4612), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3759) );
  AOI22_X1 U4203 ( .A1(n4565), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3758) );
  NAND4_X1 U4204 ( .A1(n3761), .A2(n3760), .A3(n3759), .A4(n3758), .ZN(n3762)
         );
  AOI22_X1 U4205 ( .A1(n4247), .A2(n4389), .B1(n4239), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3764) );
  AND2_X2 U4206 ( .A1(n3440), .A2(n3436), .ZN(n4396) );
  INV_X1 U4207 ( .A(n5210), .ZN(n3767) );
  OAI21_X2 U4208 ( .B1(n3767), .B2(n4010), .A(n4179), .ZN(n4762) );
  NAND2_X1 U4209 ( .A1(n4763), .A2(n4762), .ZN(n3772) );
  INV_X1 U4210 ( .A(n4775), .ZN(n3770) );
  INV_X1 U4211 ( .A(n3768), .ZN(n3769) );
  NAND2_X1 U4212 ( .A1(n3770), .A2(n3769), .ZN(n3771) );
  NAND2_X2 U4213 ( .A1(n3772), .A2(n3771), .ZN(n4761) );
  OR2_X1 U4214 ( .A1(n3737), .A2(n5762), .ZN(n3779) );
  NAND2_X1 U4215 ( .A1(n3774), .A2(n4200), .ZN(n7137) );
  INV_X1 U4216 ( .A(n3774), .ZN(n4949) );
  NAND2_X1 U4217 ( .A1(n4949), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4218 ( .A1(n7137), .A2(n3775), .ZN(n5063) );
  AOI22_X1 U4219 ( .A1(n5063), .A2(n3777), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n3776), .ZN(n3778) );
  NAND2_X1 U4220 ( .A1(n4912), .A2(n7072), .ZN(n3791) );
  AOI22_X1 U4221 ( .A1(n4497), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4222 ( .A1(n4110), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4223 ( .A1(n4603), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3781) );
  AOI22_X1 U4224 ( .A1(n4612), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3780) );
  NAND4_X1 U4225 ( .A1(n3783), .A2(n3782), .A3(n3781), .A4(n3780), .ZN(n3789)
         );
  AOI22_X1 U4226 ( .A1(n3675), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4227 ( .A1(n4604), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4228 ( .A1(n3677), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3785) );
  AOI22_X1 U4229 ( .A1(n4602), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3784) );
  NAND4_X1 U4230 ( .A1(n3787), .A2(n3786), .A3(n3785), .A4(n3784), .ZN(n3788)
         );
  XNOR2_X2 U4231 ( .A(n3436), .B(n5185), .ZN(n4403) );
  NAND2_X1 U4232 ( .A1(n4403), .A2(n3973), .ZN(n3798) );
  OAI21_X1 U4233 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3793), .A(n3821), 
        .ZN(n6679) );
  AOI22_X1 U4234 ( .A1(n4555), .A2(n6679), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U4235 ( .A1(n5866), .A2(EAX_REG_3__SCAN_IN), .ZN(n3794) );
  OAI211_X1 U4236 ( .C1(n3819), .C2(n5762), .A(n3795), .B(n3794), .ZN(n3796)
         );
  INV_X1 U4237 ( .A(n3796), .ZN(n3797) );
  AOI22_X1 U4238 ( .A1(n4611), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4239 ( .A1(n3675), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4240 ( .A1(n4612), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4241 ( .A1(n3677), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3802) );
  NAND4_X1 U4242 ( .A1(n3805), .A2(n3804), .A3(n3803), .A4(n3802), .ZN(n3811)
         );
  AOI22_X1 U4243 ( .A1(n4110), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4244 ( .A1(n4613), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4245 ( .A1(n4604), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4246 ( .A1(n4602), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3447), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4247 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3810)
         );
  NAND2_X1 U4248 ( .A1(n4247), .A2(n4413), .ZN(n3813) );
  NAND2_X1 U4249 ( .A1(n4239), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3812) );
  NAND2_X1 U4250 ( .A1(n3813), .A2(n3812), .ZN(n3814) );
  NAND2_X1 U4251 ( .A1(n3816), .A2(n3847), .ZN(n4408) );
  INV_X1 U4252 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4203) );
  NAND2_X1 U4253 ( .A1(n6226), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3818)
         );
  NAND2_X1 U4254 ( .A1(n5866), .A2(EAX_REG_4__SCAN_IN), .ZN(n3817) );
  OAI211_X1 U4255 ( .C1(n3819), .C2(n4203), .A(n3818), .B(n3817), .ZN(n3825)
         );
  INV_X1 U4256 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3822) );
  NAND2_X1 U4257 ( .A1(n3822), .A2(n3821), .ZN(n3823) );
  NAND2_X1 U4258 ( .A1(n3840), .A2(n3823), .ZN(n6878) );
  AND2_X1 U4259 ( .A1(n6878), .A2(n4555), .ZN(n3824) );
  AOI21_X1 U4260 ( .B1(n3825), .B2(n4623), .A(n3824), .ZN(n3826) );
  NAND3_X1 U4261 ( .A1(n4761), .A2(n4798), .A3(n4789), .ZN(n4792) );
  AOI22_X1 U4262 ( .A1(n4497), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4263 ( .A1(n4110), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4264 ( .A1(n4603), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4265 ( .A1(n4612), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4266 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3837)
         );
  AOI22_X1 U4267 ( .A1(n3675), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4268 ( .A1(n4604), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3834) );
  AOI22_X1 U4269 ( .A1(n3677), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4270 ( .A1(n4602), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3832) );
  NAND4_X1 U4271 ( .A1(n3835), .A2(n3834), .A3(n3833), .A4(n3832), .ZN(n3836)
         );
  NAND2_X1 U4272 ( .A1(n4247), .A2(n4422), .ZN(n3839) );
  NAND2_X1 U4273 ( .A1(n4239), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3838) );
  NAND2_X1 U4274 ( .A1(n3839), .A2(n3838), .ZN(n3848) );
  NAND2_X1 U4275 ( .A1(n4412), .A2(n3973), .ZN(n3846) );
  NAND2_X1 U4276 ( .A1(n3840), .A2(n3843), .ZN(n3841) );
  NAND2_X1 U4277 ( .A1(n3875), .A2(n3841), .ZN(n6889) );
  NAND2_X1 U4278 ( .A1(n6889), .A2(n4555), .ZN(n3842) );
  OAI21_X1 U4279 ( .B1(n3843), .B2(n4179), .A(n3842), .ZN(n3844) );
  AOI21_X1 U4280 ( .B1(n5866), .B2(EAX_REG_5__SCAN_IN), .A(n3844), .ZN(n3845)
         );
  INV_X1 U4281 ( .A(n3847), .ZN(n3849) );
  NAND2_X1 U4282 ( .A1(n3849), .A2(n3848), .ZN(n3867) );
  AOI22_X1 U4283 ( .A1(n4110), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4284 ( .A1(n3675), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4285 ( .A1(n4612), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4286 ( .A1(n4604), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3850) );
  NAND4_X1 U4287 ( .A1(n3853), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(n3859)
         );
  AOI22_X1 U4288 ( .A1(n4497), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4289 ( .A1(n4603), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4290 ( .A1(n4602), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4291 ( .A1(n3749), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4292 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3858)
         );
  AOI22_X1 U4293 ( .A1(n4247), .A2(n4438), .B1(n4239), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3868) );
  NAND2_X1 U4294 ( .A1(n3867), .A2(n3868), .ZN(n4420) );
  NAND2_X1 U4295 ( .A1(n4420), .A2(n3973), .ZN(n3865) );
  INV_X1 U4296 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3860) );
  XNOR2_X1 U4297 ( .A(n3875), .B(n3860), .ZN(n5513) );
  INV_X1 U4298 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3862) );
  INV_X1 U4299 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n7080) );
  OAI21_X1 U4300 ( .B1(n7080), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6226), 
        .ZN(n3861) );
  OAI21_X1 U4301 ( .B1(n3453), .B2(n3862), .A(n3861), .ZN(n3863) );
  OAI21_X1 U4302 ( .B1(n4623), .B2(n5513), .A(n3863), .ZN(n3864) );
  NAND2_X1 U4303 ( .A1(n3865), .A2(n3864), .ZN(n4804) );
  NAND2_X1 U4304 ( .A1(n4852), .A2(n4804), .ZN(n3866) );
  NOR2_X2 U4305 ( .A1(n4792), .A2(n3866), .ZN(n5023) );
  INV_X1 U4306 ( .A(n3867), .ZN(n3870) );
  NAND2_X1 U4307 ( .A1(n4247), .A2(n4445), .ZN(n3872) );
  NAND2_X1 U4308 ( .A1(n4239), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3871) );
  NAND2_X1 U4309 ( .A1(n3872), .A2(n3871), .ZN(n3873) );
  NAND2_X1 U4310 ( .A1(n4436), .A2(n3973), .ZN(n3882) );
  AOI22_X1 U4311 ( .A1(n5866), .A2(EAX_REG_7__SCAN_IN), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3874) );
  OR2_X1 U4312 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3877) );
  NAND2_X1 U4313 ( .A1(n3877), .A2(n3899), .ZN(n6902) );
  INV_X1 U4314 ( .A(n6902), .ZN(n3878) );
  NAND2_X1 U4315 ( .A1(n5023), .A2(n5022), .ZN(n5021) );
  INV_X1 U4316 ( .A(n5021), .ZN(n3897) );
  AOI22_X1 U4317 ( .A1(n4612), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4318 ( .A1(n4110), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4319 ( .A1(n3677), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3446), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4320 ( .A1(n4582), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4321 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  AOI22_X1 U4322 ( .A1(n4497), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4323 ( .A1(n3675), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4602), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4324 ( .A1(n4611), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4325 ( .A1(n4604), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4326 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  OAI21_X1 U4327 ( .B1(n3892), .B2(n3891), .A(n3973), .ZN(n3895) );
  XNOR2_X1 U4328 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3899), .ZN(n5206) );
  INV_X1 U4329 ( .A(n5206), .ZN(n5502) );
  AOI22_X1 U4330 ( .A1(n5865), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n4555), 
        .B2(n5502), .ZN(n3894) );
  NAND2_X1 U4331 ( .A1(n5866), .A2(EAX_REG_8__SCAN_IN), .ZN(n3893) );
  XNOR2_X1 U4332 ( .A(n3914), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6907) );
  AOI22_X1 U4333 ( .A1(n4497), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4334 ( .A1(n4110), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4335 ( .A1(n4603), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4336 ( .A1(n4604), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3900) );
  NAND4_X1 U4337 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3909)
         );
  AOI22_X1 U4338 ( .A1(n4602), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4339 ( .A1(n3675), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4340 ( .A1(n4612), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4341 ( .A1(n4565), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3658), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3904) );
  NAND4_X1 U4342 ( .A1(n3907), .A2(n3906), .A3(n3905), .A4(n3904), .ZN(n3908)
         );
  NOR2_X1 U4343 ( .A1(n3909), .A2(n3908), .ZN(n3912) );
  NAND2_X1 U4344 ( .A1(n5866), .A2(EAX_REG_9__SCAN_IN), .ZN(n3911) );
  NAND2_X1 U4345 ( .A1(n5865), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3910)
         );
  OAI211_X1 U4346 ( .C1(n4010), .C2(n3912), .A(n3911), .B(n3910), .ZN(n3913)
         );
  AOI21_X1 U4347 ( .B1(n6907), .B2(n4555), .A(n3913), .ZN(n5418) );
  XOR2_X1 U4348 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3938), .Z(n6917) );
  AOI22_X1 U4349 ( .A1(n4110), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4350 ( .A1(n3675), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4351 ( .A1(n4603), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4352 ( .A1(n4604), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4353 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3924)
         );
  AOI22_X1 U4354 ( .A1(n4611), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4355 ( .A1(n4612), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4356 ( .A1(n3677), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4357 ( .A1(n4602), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3751), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4358 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3923)
         );
  OR2_X1 U4359 ( .A1(n3924), .A2(n3923), .ZN(n3925) );
  AOI22_X1 U4360 ( .A1(n3973), .A2(n3925), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3927) );
  NAND2_X1 U4361 ( .A1(n5866), .A2(EAX_REG_10__SCAN_IN), .ZN(n3926) );
  OAI211_X1 U4362 ( .C1(n6917), .C2(n4623), .A(n3927), .B(n3926), .ZN(n5453)
         );
  AND2_X1 U4363 ( .A1(n5452), .A2(n5453), .ZN(n5451) );
  AOI22_X1 U4364 ( .A1(n4497), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4365 ( .A1(n4560), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4612), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4366 ( .A1(n3675), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4367 ( .A1(n4604), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4368 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4369 ( .A1(n4613), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4370 ( .A1(n4110), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4371 ( .A1(n3677), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4372 ( .A1(n4602), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4373 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  NOR2_X1 U4374 ( .A1(n3937), .A2(n3936), .ZN(n3942) );
  INV_X1 U4375 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3939) );
  XNOR2_X1 U4376 ( .A(n3943), .B(n3939), .ZN(n5640) );
  NAND2_X1 U4377 ( .A1(n5640), .A2(n4555), .ZN(n3941) );
  AOI22_X1 U4378 ( .A1(n5866), .A2(EAX_REG_11__SCAN_IN), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3940) );
  OAI211_X1 U4379 ( .C1(n3942), .C2(n4010), .A(n3941), .B(n3940), .ZN(n5489)
         );
  INV_X1 U4380 ( .A(n5487), .ZN(n3961) );
  XOR2_X1 U4381 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3974), .Z(n6930) );
  NAND2_X1 U4382 ( .A1(n6930), .A2(n4555), .ZN(n3959) );
  INV_X1 U4383 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3945) );
  OAI21_X1 U4384 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n7080), .A(n6226), 
        .ZN(n3944) );
  OAI21_X1 U4385 ( .B1(n3453), .B2(n3945), .A(n3944), .ZN(n3958) );
  AOI22_X1 U4386 ( .A1(n4497), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4387 ( .A1(n4110), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4388 ( .A1(n4613), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4389 ( .A1(n4604), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3946) );
  NAND4_X1 U4390 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3955)
         );
  AOI22_X1 U4391 ( .A1(n3644), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4392 ( .A1(n4612), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4393 ( .A1(n3657), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4394 ( .A1(n4602), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3449), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4395 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3954)
         );
  NOR2_X1 U4396 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  NOR2_X1 U4397 ( .A1(n4010), .A2(n3956), .ZN(n3957) );
  AOI21_X1 U4398 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n5609) );
  INV_X1 U4399 ( .A(n5609), .ZN(n3960) );
  NAND2_X1 U4400 ( .A1(n3961), .A2(n3960), .ZN(n3978) );
  AOI22_X1 U4401 ( .A1(n4497), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4402 ( .A1(n4110), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4403 ( .A1(n4603), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4404 ( .A1(n4612), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3962) );
  NAND4_X1 U4405 ( .A1(n3965), .A2(n3964), .A3(n3963), .A4(n3962), .ZN(n3971)
         );
  AOI22_X1 U4406 ( .A1(n3644), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4407 ( .A1(n4604), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4408 ( .A1(n3657), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4409 ( .A1(n4602), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3966) );
  NAND4_X1 U4410 ( .A1(n3969), .A2(n3968), .A3(n3967), .A4(n3966), .ZN(n3970)
         );
  OR2_X1 U4411 ( .A1(n3971), .A2(n3970), .ZN(n3972) );
  AND2_X1 U4412 ( .A1(n3973), .A2(n3972), .ZN(n3979) );
  XNOR2_X2 U4413 ( .A(n3978), .B(n3979), .ZN(n5657) );
  NAND2_X1 U4414 ( .A1(n3974), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3992)
         );
  INV_X1 U4415 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6946) );
  XNOR2_X1 U4416 ( .A(n3992), .B(n6946), .ZN(n6936) );
  NAND2_X1 U4417 ( .A1(n6936), .A2(n4555), .ZN(n3977) );
  NOR2_X1 U4418 ( .A1(n4179), .A2(n6946), .ZN(n3975) );
  AOI21_X1 U4419 ( .B1(n5866), .B2(EAX_REG_13__SCAN_IN), .A(n3975), .ZN(n3976)
         );
  NAND2_X1 U4420 ( .A1(n3977), .A2(n3976), .ZN(n5658) );
  NAND2_X1 U4421 ( .A1(n5657), .A2(n5658), .ZN(n3981) );
  AOI22_X1 U4422 ( .A1(n4110), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3985) );
  AOI22_X1 U4423 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n4603), .B1(n4582), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4424 ( .A1(n3644), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4425 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n3677), .B1(n4604), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3982) );
  NAND4_X1 U4426 ( .A1(n3985), .A2(n3984), .A3(n3983), .A4(n3982), .ZN(n3991)
         );
  AOI22_X1 U4427 ( .A1(n4560), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4428 ( .A1(n4612), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4429 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n4565), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4430 ( .A1(n4602), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3986) );
  NAND4_X1 U4431 ( .A1(n3989), .A2(n3988), .A3(n3987), .A4(n3986), .ZN(n3990)
         );
  NOR2_X1 U4432 ( .A1(n3991), .A2(n3990), .ZN(n3995) );
  XNOR2_X1 U4433 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3996), .ZN(n5684)
         );
  AOI22_X1 U4434 ( .A1(n4555), .A2(n5684), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3994) );
  NAND2_X1 U4435 ( .A1(n5866), .A2(EAX_REG_14__SCAN_IN), .ZN(n3993) );
  OAI211_X1 U4436 ( .C1(n4010), .C2(n3995), .A(n3994), .B(n3993), .ZN(n5678)
         );
  NAND2_X1 U4437 ( .A1(n5677), .A2(n5678), .ZN(n5714) );
  INV_X1 U4438 ( .A(n5714), .ZN(n4014) );
  XNOR2_X1 U4439 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n4015), .ZN(n5727)
         );
  INV_X1 U4440 ( .A(n5727), .ZN(n4012) );
  AOI22_X1 U4441 ( .A1(n4611), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4442 ( .A1(n4110), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4443 ( .A1(n3644), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4444 ( .A1(n4565), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3997) );
  NAND4_X1 U4445 ( .A1(n4000), .A2(n3999), .A3(n3998), .A4(n3997), .ZN(n4006)
         );
  AOI22_X1 U4446 ( .A1(n4602), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4447 ( .A1(n4612), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4448 ( .A1(n4497), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4449 ( .A1(n4604), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4001) );
  NAND4_X1 U4450 ( .A1(n4004), .A2(n4003), .A3(n4002), .A4(n4001), .ZN(n4005)
         );
  NOR2_X1 U4451 ( .A1(n4006), .A2(n4005), .ZN(n4009) );
  NAND2_X1 U4452 ( .A1(n5866), .A2(EAX_REG_15__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U4453 ( .A1(n5865), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n4007)
         );
  OAI211_X1 U4454 ( .C1(n4010), .C2(n4009), .A(n4008), .B(n4007), .ZN(n4011)
         );
  AOI21_X1 U4455 ( .B1(n4012), .B2(n4555), .A(n4011), .ZN(n5715) );
  NAND2_X1 U4456 ( .A1(n4014), .A2(n4013), .ZN(n5712) );
  INV_X1 U4457 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U4458 ( .A(n4043), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6116)
         );
  NAND2_X1 U4459 ( .A1(n4016), .A2(n4378), .ZN(n4841) );
  AOI22_X1 U4460 ( .A1(n4110), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4461 ( .A1(n4602), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4462 ( .A1(n4613), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U4463 ( .A1(n4604), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4017) );
  NAND4_X1 U4464 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4026)
         );
  AOI22_X1 U4465 ( .A1(n4497), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U4466 ( .A1(n3644), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4467 ( .A1(n4612), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4468 ( .A1(n4565), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4021) );
  NAND4_X1 U4469 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4025)
         );
  NOR2_X1 U4470 ( .A1(n4026), .A2(n4025), .ZN(n4028) );
  AOI22_X1 U4471 ( .A1(n5866), .A2(EAX_REG_16__SCAN_IN), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4027) );
  OAI21_X1 U4472 ( .B1(n4596), .B2(n4028), .A(n4027), .ZN(n4029) );
  AOI21_X1 U4473 ( .B1(n6116), .B2(n4555), .A(n4029), .ZN(n5729) );
  NOR2_X2 U4474 ( .A1(n5712), .A2(n5729), .ZN(n5730) );
  AOI22_X1 U4475 ( .A1(n4110), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U4476 ( .A1(n3675), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4477 ( .A1(n4612), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4478 ( .A1(n3657), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U4479 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U4480 ( .A1(n4497), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U4481 ( .A1(n4613), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4482 ( .A1(n4604), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4483 ( .A1(n4602), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U4484 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U4485 ( .A1(n4039), .A2(n4038), .ZN(n4040) );
  OR2_X1 U4486 ( .A1(n4596), .A2(n4040), .ZN(n4047) );
  OAI21_X1 U4487 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n7080), .A(n6226), 
        .ZN(n4041) );
  INV_X1 U4488 ( .A(n4041), .ZN(n4042) );
  AOI21_X1 U4489 ( .B1(n5866), .B2(EAX_REG_17__SCAN_IN), .A(n4042), .ZN(n4046)
         );
  OAI21_X1 U4490 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4044), .A(n4067), 
        .ZN(n6706) );
  NOR2_X1 U4491 ( .A1(n6706), .A2(n4623), .ZN(n4045) );
  AOI21_X1 U4492 ( .B1(n4047), .B2(n4046), .A(n4045), .ZN(n5948) );
  NAND2_X1 U4493 ( .A1(n5730), .A2(n5948), .ZN(n5946) );
  INV_X1 U4494 ( .A(n5946), .ZN(n4065) );
  AOI22_X1 U4495 ( .A1(n4497), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4051) );
  AOI22_X1 U4496 ( .A1(n4110), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4612), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4050) );
  AOI22_X1 U4497 ( .A1(n4603), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4049) );
  AOI22_X1 U4498 ( .A1(n4604), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4048) );
  NAND4_X1 U4499 ( .A1(n4051), .A2(n4050), .A3(n4049), .A4(n4048), .ZN(n4057)
         );
  AOI22_X1 U4500 ( .A1(n4602), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U4501 ( .A1(n3675), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U4502 ( .A1(n4606), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U4503 ( .A1(n4565), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4052) );
  NAND4_X1 U4504 ( .A1(n4055), .A2(n4054), .A3(n4053), .A4(n4052), .ZN(n4056)
         );
  NOR2_X1 U4505 ( .A1(n4057), .A2(n4056), .ZN(n4061) );
  NAND2_X1 U4506 ( .A1(n6226), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4058)
         );
  NAND2_X1 U4507 ( .A1(n4623), .A2(n4058), .ZN(n4059) );
  AOI21_X1 U4508 ( .B1(n5866), .B2(EAX_REG_18__SCAN_IN), .A(n4059), .ZN(n4060)
         );
  OAI21_X1 U4509 ( .B1(n4596), .B2(n4061), .A(n4060), .ZN(n4063) );
  XNOR2_X1 U4510 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4067), .ZN(n6957)
         );
  NAND2_X1 U4511 ( .A1(n4555), .A2(n6957), .ZN(n4062) );
  NAND2_X1 U4512 ( .A1(n4063), .A2(n4062), .ZN(n5993) );
  NAND2_X1 U4513 ( .A1(n4065), .A2(n4064), .ZN(n5991) );
  INV_X1 U4514 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4066) );
  INV_X1 U4515 ( .A(n4103), .ZN(n4070) );
  OR2_X1 U4516 ( .A1(n4068), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4069)
         );
  NAND2_X1 U4517 ( .A1(n4070), .A2(n4069), .ZN(n6973) );
  AOI22_X1 U4518 ( .A1(n4612), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4074) );
  AOI22_X1 U4519 ( .A1(n3644), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4602), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4073) );
  AOI22_X1 U4520 ( .A1(n4613), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U4521 ( .A1(n3677), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4071) );
  NAND4_X1 U4522 ( .A1(n4074), .A2(n4073), .A3(n4072), .A4(n4071), .ZN(n4080)
         );
  AOI22_X1 U4523 ( .A1(n4497), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4078) );
  AOI22_X1 U4524 ( .A1(n4110), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U4525 ( .A1(n4604), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U4526 ( .A1(n4582), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4075) );
  NAND4_X1 U4527 ( .A1(n4078), .A2(n4077), .A3(n4076), .A4(n4075), .ZN(n4079)
         );
  NOR2_X1 U4528 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  NOR2_X1 U4529 ( .A1(n4596), .A2(n4081), .ZN(n4085) );
  INV_X1 U4530 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4083) );
  NAND2_X1 U4531 ( .A1(n6226), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4082)
         );
  OAI211_X1 U4532 ( .C1(n3453), .C2(n4083), .A(n4623), .B(n4082), .ZN(n4084)
         );
  OAI22_X1 U4533 ( .A1(n6973), .A2(n4623), .B1(n4085), .B2(n4084), .ZN(n6652)
         );
  INV_X1 U4534 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6985) );
  XNOR2_X1 U4535 ( .A(n4103), .B(n6985), .ZN(n6982) );
  NAND2_X1 U4536 ( .A1(n6982), .A2(n4555), .ZN(n4102) );
  AOI22_X1 U4537 ( .A1(n4087), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U4538 ( .A1(n4612), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U4539 ( .A1(n3675), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U4540 ( .A1(n4602), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U4541 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4097)
         );
  AOI22_X1 U4542 ( .A1(n4110), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U4543 ( .A1(n4613), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U4544 ( .A1(n4604), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4093) );
  AOI22_X1 U4545 ( .A1(n3677), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4092) );
  NAND4_X1 U4546 ( .A1(n4095), .A2(n4094), .A3(n4093), .A4(n4092), .ZN(n4096)
         );
  NOR2_X1 U4547 ( .A1(n4097), .A2(n4096), .ZN(n4100) );
  AOI21_X1 U4548 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6985), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4098) );
  AOI21_X1 U4549 ( .B1(n5866), .B2(EAX_REG_20__SCAN_IN), .A(n4098), .ZN(n4099)
         );
  OAI21_X1 U4550 ( .B1(n4596), .B2(n4100), .A(n4099), .ZN(n4101) );
  NAND2_X1 U4551 ( .A1(n4102), .A2(n4101), .ZN(n5990) );
  NOR2_X2 U4552 ( .A1(n5987), .A2(n5990), .ZN(n5988) );
  INV_X1 U4553 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4117) );
  AND2_X1 U4554 ( .A1(n4104), .A2(n4117), .ZN(n4105) );
  OR2_X1 U4555 ( .A1(n4105), .A2(n4151), .ZN(n6996) );
  AOI22_X1 U4556 ( .A1(n4087), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U4557 ( .A1(n4560), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4612), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U4558 ( .A1(n4613), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4107) );
  AOI22_X1 U4559 ( .A1(n4565), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4106) );
  NAND4_X1 U4560 ( .A1(n4109), .A2(n4108), .A3(n4107), .A4(n4106), .ZN(n4116)
         );
  AOI22_X1 U4561 ( .A1(n3644), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U4562 ( .A1(n3677), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U4563 ( .A1(n4110), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U4564 ( .A1(n4602), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4111) );
  NAND4_X1 U4565 ( .A1(n4114), .A2(n4113), .A3(n4112), .A4(n4111), .ZN(n4115)
         );
  NOR2_X1 U4566 ( .A1(n4116), .A2(n4115), .ZN(n4120) );
  OAI21_X1 U4567 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4117), .A(n4623), .ZN(
        n4118) );
  AOI21_X1 U4568 ( .B1(n5866), .B2(EAX_REG_21__SCAN_IN), .A(n4118), .ZN(n4119)
         );
  OAI21_X1 U4569 ( .B1(n4596), .B2(n4120), .A(n4119), .ZN(n4121) );
  OAI21_X1 U4570 ( .B1(n6996), .B2(n4623), .A(n4121), .ZN(n6092) );
  INV_X1 U4571 ( .A(n6092), .ZN(n4122) );
  AND2_X2 U4572 ( .A1(n5988), .A2(n4122), .ZN(n4577) );
  BUF_X4 U4573 ( .A(n4577), .Z(n5917) );
  NAND2_X1 U4574 ( .A1(n4151), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4123)
         );
  INV_X1 U4575 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U4576 ( .A1(n4123), .A2(n4145), .ZN(n4124) );
  NAND2_X1 U4577 ( .A1(n4190), .A2(n4124), .ZN(n7011) );
  OR2_X1 U4578 ( .A1(n7011), .A2(n4623), .ZN(n4150) );
  AOI22_X1 U4579 ( .A1(n4497), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4128) );
  AOI22_X1 U4580 ( .A1(n4612), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4127) );
  AOI22_X1 U4581 ( .A1(n4602), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U4582 ( .A1(n4560), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4125) );
  NAND4_X1 U4583 ( .A1(n4128), .A2(n4127), .A3(n4126), .A4(n4125), .ZN(n4134)
         );
  AOI22_X1 U4584 ( .A1(n4110), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U4585 ( .A1(n3675), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U4586 ( .A1(n3657), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U4587 ( .A1(n4565), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4129) );
  NAND4_X1 U4588 ( .A1(n4132), .A2(n4131), .A3(n4130), .A4(n4129), .ZN(n4133)
         );
  NOR2_X1 U4589 ( .A1(n4134), .A2(n4133), .ZN(n4167) );
  AOI22_X1 U4590 ( .A1(n4110), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4138) );
  AOI22_X1 U4591 ( .A1(n4613), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U4592 ( .A1(n3644), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4604), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U4593 ( .A1(n4612), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4135) );
  NAND4_X1 U4594 ( .A1(n4138), .A2(n4137), .A3(n4136), .A4(n4135), .ZN(n4144)
         );
  AOI22_X1 U4595 ( .A1(n4497), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U4596 ( .A1(n4602), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3677), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U4597 ( .A1(n4603), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U4598 ( .A1(n4565), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U4599 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4143)
         );
  NOR2_X1 U4600 ( .A1(n4144), .A2(n4143), .ZN(n4168) );
  XNOR2_X1 U4601 ( .A(n4167), .B(n4168), .ZN(n4148) );
  OAI21_X1 U4602 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4145), .A(n4623), .ZN(
        n4146) );
  AOI21_X1 U4603 ( .B1(n5866), .B2(EAX_REG_23__SCAN_IN), .A(n4146), .ZN(n4147)
         );
  OAI21_X1 U4604 ( .B1(n4596), .B2(n4148), .A(n4147), .ZN(n4149) );
  AND2_X1 U4605 ( .A1(n4150), .A2(n4149), .ZN(n5974) );
  INV_X1 U4606 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4481) );
  XNOR2_X1 U4607 ( .A(n4151), .B(n4481), .ZN(n5757) );
  INV_X1 U4608 ( .A(n4596), .ZN(n4627) );
  AOI22_X1 U4609 ( .A1(n4611), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U4610 ( .A1(n4110), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4612), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4154) );
  AOI22_X1 U4611 ( .A1(n4613), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U4612 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n4602), .B1(n4565), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4152) );
  NAND4_X1 U4613 ( .A1(n4155), .A2(n4154), .A3(n4153), .A4(n4152), .ZN(n4161)
         );
  AOI22_X1 U4614 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n3644), .B1(n3657), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U4615 ( .A1(n4603), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U4616 ( .A1(n4497), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U4617 ( .A1(n4604), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U4618 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4160)
         );
  OR2_X1 U4619 ( .A1(n4161), .A2(n4160), .ZN(n4165) );
  INV_X1 U4620 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U4621 ( .A1(n6226), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4162)
         );
  OAI211_X1 U4622 ( .C1(n3453), .C2(n4163), .A(n4623), .B(n4162), .ZN(n4164)
         );
  AOI21_X1 U4623 ( .B1(n4627), .B2(n4165), .A(n4164), .ZN(n4166) );
  AOI21_X1 U4624 ( .B1(n5757), .B2(n4555), .A(n4166), .ZN(n4371) );
  AND2_X1 U4625 ( .A1(n5974), .A2(n4371), .ZN(n4187) );
  NAND2_X1 U4626 ( .A1(n5917), .A2(n4187), .ZN(n5976) );
  XNOR2_X1 U4627 ( .A(n4190), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6074)
         );
  OR2_X1 U4628 ( .A1(n6074), .A2(n4623), .ZN(n4184) );
  OR2_X1 U4629 ( .A1(n4168), .A2(n4167), .ZN(n4520) );
  AOI22_X1 U4630 ( .A1(n4602), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U4631 ( .A1(n4497), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4171) );
  AOI22_X1 U4632 ( .A1(n4613), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4170) );
  AOI22_X1 U4633 ( .A1(n3644), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4169) );
  NAND4_X1 U4634 ( .A1(n4172), .A2(n4171), .A3(n4170), .A4(n4169), .ZN(n4178)
         );
  AOI22_X1 U4635 ( .A1(n4612), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U4636 ( .A1(n3657), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4637 ( .A1(n4604), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U4638 ( .A1(n4110), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U4639 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4177)
         );
  OR2_X1 U4640 ( .A1(n4178), .A2(n4177), .ZN(n4518) );
  XNOR2_X1 U4641 ( .A(n4520), .B(n4518), .ZN(n4182) );
  INV_X1 U4642 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4180) );
  INV_X1 U4643 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4189) );
  OAI22_X1 U4644 ( .A1(n3453), .A2(n4180), .B1(n4189), .B2(n4179), .ZN(n4181)
         );
  AOI21_X1 U4645 ( .B1(n4627), .B2(n4182), .A(n4181), .ZN(n4183) );
  AND2_X1 U4646 ( .A1(n4184), .A2(n4183), .ZN(n4185) );
  NAND2_X1 U4647 ( .A1(n5976), .A2(n4185), .ZN(n4188) );
  INV_X1 U4648 ( .A(n4185), .ZN(n4186) );
  AND2_X1 U4649 ( .A1(n4187), .A2(n4186), .ZN(n4545) );
  NAND2_X1 U4650 ( .A1(n5917), .A2(n4545), .ZN(n5932) );
  INV_X1 U4651 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4548) );
  INV_X1 U4652 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4494) );
  INV_X1 U4653 ( .A(n4557), .ZN(n4191) );
  NAND2_X1 U4654 ( .A1(n4191), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4578)
         );
  INV_X1 U4655 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5880) );
  INV_X1 U4656 ( .A(n4599), .ZN(n4192) );
  NAND2_X1 U4657 ( .A1(n4192), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4194)
         );
  INV_X1 U4658 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4193) );
  XNOR2_X1 U4659 ( .A(n4194), .B(n4193), .ZN(n6038) );
  XNOR2_X1 U4660 ( .A(n5137), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4205)
         );
  NAND2_X1 U4661 ( .A1(n7020), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4207) );
  INV_X1 U4662 ( .A(n4207), .ZN(n4195) );
  NAND2_X1 U4663 ( .A1(n4205), .A2(n4195), .ZN(n4197) );
  NAND2_X1 U4664 ( .A1(n5523), .A2(n5137), .ZN(n4196) );
  NAND2_X1 U4665 ( .A1(n4197), .A2(n4196), .ZN(n4225) );
  XNOR2_X1 U4666 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U4667 ( .A1(n4225), .A2(n4223), .ZN(n4199) );
  NAND2_X1 U4668 ( .A1(n5181), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4198) );
  NAND2_X1 U4669 ( .A1(n4199), .A2(n4198), .ZN(n4235) );
  MUX2_X1 U4670 ( .A(n4200), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4233) );
  NAND2_X1 U4671 ( .A1(n4235), .A2(n4233), .ZN(n4202) );
  NAND2_X1 U4672 ( .A1(n4200), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U4673 ( .A1(n4202), .A2(n4201), .ZN(n4244) );
  INV_X1 U4674 ( .A(n4239), .ZN(n4227) );
  XNOR2_X1 U4675 ( .A(n4205), .B(n4207), .ZN(n4260) );
  OAI21_X1 U4676 ( .B1(n4227), .B2(n4260), .A(n4378), .ZN(n4206) );
  AOI21_X1 U4677 ( .B1(n4247), .B2(n4751), .A(n4206), .ZN(n4217) );
  NAND2_X1 U4678 ( .A1(n4260), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4216) );
  OAI21_X1 U4679 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n7020), .A(n4207), 
        .ZN(n4209) );
  INV_X1 U4680 ( .A(n4247), .ZN(n4208) );
  AOI211_X1 U4681 ( .C1(n4217), .C2(n4216), .A(n4209), .B(n4208), .ZN(n4215)
         );
  INV_X1 U4682 ( .A(n4251), .ZN(n4220) );
  INV_X1 U4683 ( .A(n4474), .ZN(n4211) );
  INV_X1 U4684 ( .A(n4209), .ZN(n4210) );
  AOI21_X1 U4685 ( .B1(n4211), .B2(n4210), .A(n4939), .ZN(n4214) );
  AND2_X1 U4686 ( .A1(n3604), .A2(n4378), .ZN(n4213) );
  OAI22_X1 U4687 ( .A1(n4215), .A2(n4220), .B1(n4214), .B2(n4229), .ZN(n4222)
         );
  INV_X1 U4688 ( .A(n4216), .ZN(n4219) );
  INV_X1 U4689 ( .A(n4217), .ZN(n4218) );
  OAI21_X1 U4690 ( .B1(n4220), .B2(n4219), .A(n4218), .ZN(n4221) );
  NAND2_X1 U4691 ( .A1(n4222), .A2(n4221), .ZN(n4232) );
  INV_X1 U4692 ( .A(n4223), .ZN(n4224) );
  XNOR2_X1 U4693 ( .A(n4225), .B(n4224), .ZN(n4259) );
  NAND2_X1 U4694 ( .A1(n4247), .A2(n4259), .ZN(n4228) );
  INV_X1 U4695 ( .A(n4229), .ZN(n4226) );
  OAI211_X1 U4696 ( .C1(n4227), .C2(n4259), .A(n4228), .B(n4226), .ZN(n4231)
         );
  INV_X1 U4697 ( .A(n4228), .ZN(n4230) );
  AOI22_X1 U4698 ( .A1(n4232), .A2(n4231), .B1(n4230), .B2(n4229), .ZN(n4237)
         );
  INV_X1 U4699 ( .A(n4233), .ZN(n4234) );
  XNOR2_X1 U4700 ( .A(n4235), .B(n4234), .ZN(n4261) );
  NOR2_X1 U4701 ( .A1(n4239), .A2(n4261), .ZN(n4236) );
  OAI22_X1 U4702 ( .A1(n4237), .A2(n4236), .B1(n4261), .B2(n4251), .ZN(n4238)
         );
  OAI21_X1 U4703 ( .B1(n4239), .B2(n4264), .A(n4238), .ZN(n4240) );
  OAI21_X1 U4704 ( .B1(n4264), .B2(n4251), .A(n4240), .ZN(n4241) );
  AOI21_X1 U4705 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n7072), .A(n4241), 
        .ZN(n4249) );
  NAND2_X1 U4706 ( .A1(n4242), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U4707 ( .A1(n4244), .A2(n4243), .ZN(n4245) );
  NAND2_X1 U4708 ( .A1(n4246), .A2(n4245), .ZN(n4263) );
  NAND2_X1 U4709 ( .A1(n4247), .A2(n4263), .ZN(n4248) );
  NAND2_X1 U4710 ( .A1(n4249), .A2(n4248), .ZN(n4253) );
  INV_X1 U4711 ( .A(n4263), .ZN(n4250) );
  NAND2_X1 U4712 ( .A1(n4255), .A2(STATE2_REG_0__SCAN_IN), .ZN(n7077) );
  OR2_X1 U4713 ( .A1(n4254), .A2(n7077), .ZN(n4256) );
  INV_X1 U4714 ( .A(n7077), .ZN(n7047) );
  AND3_X1 U4715 ( .A1(n4261), .A2(n4260), .A3(n4259), .ZN(n4262) );
  OR2_X1 U4716 ( .A1(n4263), .A2(n4262), .ZN(n4265) );
  NAND2_X1 U4717 ( .A1(n4265), .A2(n4264), .ZN(n5849) );
  NAND3_X1 U4718 ( .A1(n3605), .A2(n7047), .A3(n5849), .ZN(n4731) );
  NOR2_X2 U4719 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n7146) );
  NAND2_X1 U4720 ( .A1(n7146), .A2(n7062), .ZN(n6724) );
  OR2_X1 U4721 ( .A1(n6724), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U4722 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n7070) );
  NAND3_X1 U4723 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), 
        .A3(n7070), .ZN(n7075) );
  NOR2_X1 U4724 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7062), .ZN(n4730) );
  NAND2_X1 U4725 ( .A1(n4555), .A2(n4730), .ZN(n7059) );
  NAND3_X1 U4726 ( .A1(n4480), .A2(n7075), .A3(n7059), .ZN(n4266) );
  NAND2_X1 U4727 ( .A1(n5826), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4362) );
  INV_X1 U4728 ( .A(READY_N), .ZN(n7088) );
  NAND2_X1 U4729 ( .A1(n7080), .A2(n7088), .ZN(n4364) );
  NAND3_X1 U4730 ( .A1(n3426), .A2(EBX_REG_31__SCAN_IN), .A3(n4364), .ZN(n4267) );
  NOR2_X2 U4731 ( .A1(n5350), .A2(n4267), .ZN(n6993) );
  AND2_X2 U4732 ( .A1(n4268), .A2(n3426), .ZN(n4678) );
  INV_X1 U4733 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4269) );
  NAND2_X1 U4734 ( .A1(n4678), .A2(n4269), .ZN(n4273) );
  NAND2_X2 U4735 ( .A1(n4944), .A2(n4733), .ZN(n4679) );
  INV_X1 U4736 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U4737 ( .A1(n4679), .A2(n6764), .ZN(n4271) );
  NAND2_X1 U4738 ( .A1(n4767), .A2(n4269), .ZN(n4270) );
  NAND3_X1 U4739 ( .A1(n4271), .A2(n5859), .A3(n4270), .ZN(n4272) );
  NAND2_X1 U4740 ( .A1(n4273), .A2(n4272), .ZN(n4275) );
  NAND2_X1 U4741 ( .A1(n4679), .A2(EBX_REG_0__SCAN_IN), .ZN(n4274) );
  OAI21_X1 U4742 ( .B1(n4268), .B2(EBX_REG_0__SCAN_IN), .A(n4274), .ZN(n4821)
         );
  XNOR2_X1 U4743 ( .A(n4275), .B(n4821), .ZN(n5362) );
  INV_X1 U4744 ( .A(n4275), .ZN(n4276) );
  INV_X1 U4745 ( .A(n4678), .ZN(n4353) );
  INV_X1 U4746 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6806) );
  NAND2_X1 U4747 ( .A1(n4679), .A2(n6806), .ZN(n4278) );
  INV_X1 U4748 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5345) );
  NAND2_X1 U4749 ( .A1(n4767), .A2(n5345), .ZN(n4277) );
  NAND3_X1 U4750 ( .A1(n4278), .A2(n5859), .A3(n4277), .ZN(n4279) );
  OAI21_X1 U4751 ( .B1(n4353), .B2(EBX_REG_2__SCAN_IN), .A(n4279), .ZN(n4771)
         );
  MUX2_X1 U4752 ( .A(n4675), .B(n5859), .S(EBX_REG_3__SCAN_IN), .Z(n4281) );
  INV_X1 U4753 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U4754 ( .A1(n4823), .A2(n6777), .ZN(n4280) );
  AND2_X1 U4755 ( .A1(n4281), .A2(n4280), .ZN(n4799) );
  NAND2_X1 U4756 ( .A1(n4800), .A2(n4799), .ZN(n4802) );
  INV_X1 U4757 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U4758 ( .A1(n4678), .A2(n6872), .ZN(n4285) );
  INV_X1 U4759 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U4760 ( .A1(n4679), .A2(n6770), .ZN(n4283) );
  NAND2_X1 U4761 ( .A1(n4767), .A2(n6872), .ZN(n4282) );
  NAND3_X1 U4762 ( .A1(n4283), .A2(n5859), .A3(n4282), .ZN(n4284) );
  AND2_X1 U4763 ( .A1(n4285), .A2(n4284), .ZN(n4794) );
  INV_X1 U4764 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U4765 ( .A1(n5598), .A2(n4823), .ZN(n4287) );
  MUX2_X1 U4766 ( .A(n4675), .B(n5859), .S(EBX_REG_5__SCAN_IN), .Z(n4286) );
  NAND2_X1 U4767 ( .A1(n4287), .A2(n4286), .ZN(n4854) );
  INV_X1 U4768 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U4769 ( .A1(n4678), .A2(n5479), .ZN(n4291) );
  INV_X1 U4770 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4427) );
  NAND2_X1 U4771 ( .A1(n4679), .A2(n4427), .ZN(n4289) );
  NAND2_X1 U4772 ( .A1(n4767), .A2(n5479), .ZN(n4288) );
  NAND3_X1 U4773 ( .A1(n4289), .A2(n5859), .A3(n4288), .ZN(n4290) );
  MUX2_X1 U4774 ( .A(n4675), .B(n5859), .S(EBX_REG_7__SCAN_IN), .Z(n4293) );
  INV_X1 U4775 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U4776 ( .A1(n6817), .A2(n4823), .ZN(n4292) );
  NAND2_X1 U4777 ( .A1(n5025), .A2(n5024), .ZN(n5194) );
  INV_X1 U4778 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U4779 ( .A1(n4678), .A2(n5199), .ZN(n4297) );
  INV_X1 U4780 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5445) );
  NAND2_X1 U4781 ( .A1(n4679), .A2(n5445), .ZN(n4295) );
  NAND2_X1 U4782 ( .A1(n4767), .A2(n5199), .ZN(n4294) );
  NAND3_X1 U4783 ( .A1(n4295), .A2(n5859), .A3(n4294), .ZN(n4296) );
  AND2_X1 U4784 ( .A1(n4297), .A2(n4296), .ZN(n5193) );
  INV_X1 U4785 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U4786 ( .A1(n4298), .A2(n4823), .ZN(n4300) );
  MUX2_X1 U4787 ( .A(n4675), .B(n5859), .S(EBX_REG_9__SCAN_IN), .Z(n4299) );
  NAND2_X1 U4788 ( .A1(n4300), .A2(n4299), .ZN(n5420) );
  INV_X1 U4789 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4454) );
  NAND2_X1 U4790 ( .A1(n4679), .A2(n4454), .ZN(n4302) );
  INV_X1 U4791 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6915) );
  NAND2_X1 U4792 ( .A1(n4767), .A2(n6915), .ZN(n4301) );
  NAND3_X1 U4793 ( .A1(n4302), .A2(n5859), .A3(n4301), .ZN(n4303) );
  OAI21_X1 U4794 ( .B1(n4353), .B2(EBX_REG_10__SCAN_IN), .A(n4303), .ZN(n5455)
         );
  MUX2_X1 U4795 ( .A(n4675), .B(n5859), .S(EBX_REG_11__SCAN_IN), .Z(n4305) );
  INV_X1 U4796 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6830) );
  NAND2_X1 U4797 ( .A1(n6830), .A2(n4823), .ZN(n4304) );
  INV_X1 U4798 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5616) );
  NAND2_X1 U4799 ( .A1(n5616), .A2(n4823), .ZN(n4307) );
  MUX2_X1 U4800 ( .A(n4675), .B(n5859), .S(EBX_REG_13__SCAN_IN), .Z(n4306) );
  NAND2_X1 U4801 ( .A1(n4307), .A2(n4306), .ZN(n5626) );
  INV_X1 U4802 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4457) );
  OAI21_X1 U4803 ( .B1(n4268), .B2(n4457), .A(n4679), .ZN(n4308) );
  OAI21_X1 U4804 ( .B1(EBX_REG_12__SCAN_IN), .B2(n5861), .A(n4308), .ZN(n4310)
         );
  INV_X1 U4805 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U4806 ( .A1(n4678), .A2(n5611), .ZN(n4309) );
  INV_X1 U4807 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U4808 ( .A1(n4678), .A2(n5688), .ZN(n4315) );
  INV_X1 U4809 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U4810 ( .A1(n4679), .A2(n5703), .ZN(n4313) );
  NAND2_X1 U4811 ( .A1(n4767), .A2(n5688), .ZN(n4312) );
  NAND3_X1 U4812 ( .A1(n4313), .A2(n5859), .A3(n4312), .ZN(n4314) );
  AND2_X1 U4813 ( .A1(n4315), .A2(n4314), .ZN(n5649) );
  MUX2_X1 U4814 ( .A(n4675), .B(n5859), .S(EBX_REG_15__SCAN_IN), .Z(n4317) );
  INV_X1 U4815 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U4816 ( .A1(n6837), .A2(n4823), .ZN(n4316) );
  INV_X1 U4817 ( .A(n4675), .ZN(n4668) );
  MUX2_X1 U4818 ( .A(n4668), .B(n4268), .S(EBX_REG_17__SCAN_IN), .Z(n4319) );
  INV_X1 U4819 ( .A(n4823), .ZN(n5862) );
  NOR2_X1 U4820 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4318)
         );
  NOR2_X1 U4821 ( .A1(n4319), .A2(n4318), .ZN(n5953) );
  INV_X1 U4822 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4320) );
  NAND2_X1 U4823 ( .A1(n4678), .A2(n4320), .ZN(n4324) );
  INV_X1 U4824 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U4825 ( .A1(n4679), .A2(n6105), .ZN(n4322) );
  NAND2_X1 U4826 ( .A1(n4767), .A2(n4320), .ZN(n4321) );
  NAND3_X1 U4827 ( .A1(n4322), .A2(n5859), .A3(n4321), .ZN(n4323) );
  NAND2_X1 U4828 ( .A1(n4324), .A2(n4323), .ZN(n5952) );
  NAND2_X1 U4829 ( .A1(n5953), .A2(n5952), .ZN(n4325) );
  INV_X1 U4830 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U4831 ( .A1(n4678), .A2(n5997), .ZN(n4329) );
  INV_X1 U4832 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U4833 ( .A1(n4679), .A2(n6108), .ZN(n4327) );
  NAND2_X1 U4834 ( .A1(n4767), .A2(n5997), .ZN(n4326) );
  NAND3_X1 U4835 ( .A1(n4327), .A2(n5859), .A3(n4326), .ZN(n4328) );
  AND2_X1 U4836 ( .A1(n4329), .A2(n4328), .ZN(n5994) );
  INV_X1 U4837 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U4838 ( .A1(n4668), .A2(n6662), .ZN(n4332) );
  INV_X1 U4839 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U4840 ( .A1(n3426), .A2(n6662), .ZN(n4330) );
  OAI211_X1 U4841 ( .C1(n4268), .C2(n6096), .A(n4330), .B(n4679), .ZN(n4331)
         );
  AND2_X1 U4842 ( .A1(n4332), .A2(n4331), .ZN(n6654) );
  INV_X1 U4843 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6069) );
  OAI21_X1 U4844 ( .B1(n4268), .B2(n6069), .A(n4679), .ZN(n4335) );
  INV_X1 U4845 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4333) );
  NAND2_X1 U4846 ( .A1(n4767), .A2(n4333), .ZN(n4334) );
  NAND2_X1 U4847 ( .A1(n4335), .A2(n4334), .ZN(n4336) );
  OAI21_X1 U4848 ( .B1(EBX_REG_20__SCAN_IN), .B2(n4353), .A(n4336), .ZN(n5985)
         );
  INV_X1 U4849 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6651) );
  NAND2_X1 U4850 ( .A1(n4668), .A2(n6651), .ZN(n4340) );
  INV_X1 U4851 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4338) );
  NAND2_X1 U4852 ( .A1(n3426), .A2(n6651), .ZN(n4337) );
  OAI211_X1 U4853 ( .C1(n4268), .C2(n4338), .A(n4337), .B(n4679), .ZN(n4339)
         );
  NAND2_X1 U4854 ( .A1(n4340), .A2(n4339), .ZN(n6195) );
  MUX2_X1 U4855 ( .A(n4675), .B(n5859), .S(EBX_REG_23__SCAN_IN), .Z(n4342) );
  INV_X1 U4856 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U4857 ( .A1(n4823), .A2(n6180), .ZN(n4341) );
  AND2_X1 U4858 ( .A1(n4342), .A2(n4341), .ZN(n5978) );
  INV_X1 U4859 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U4860 ( .A1(n4678), .A2(n5753), .ZN(n4347) );
  INV_X1 U4861 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U4862 ( .A1(n4679), .A2(n4343), .ZN(n4345) );
  NAND2_X1 U4863 ( .A1(n4767), .A2(n5753), .ZN(n4344) );
  NAND3_X1 U4864 ( .A1(n4345), .A2(n5859), .A3(n4344), .ZN(n4346) );
  NAND2_X1 U4865 ( .A1(n4347), .A2(n4346), .ZN(n5979) );
  NAND2_X1 U4866 ( .A1(n5978), .A2(n5979), .ZN(n4348) );
  INV_X1 U4867 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6171) );
  OAI21_X1 U4868 ( .B1(n4268), .B2(n6171), .A(n4679), .ZN(n4351) );
  INV_X1 U4869 ( .A(EBX_REG_24__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U4870 ( .A1(n3426), .A2(n4349), .ZN(n4350) );
  NAND2_X1 U4871 ( .A1(n4351), .A2(n4350), .ZN(n4352) );
  OAI21_X1 U4872 ( .B1(EBX_REG_24__SCAN_IN), .B2(n4353), .A(n4352), .ZN(n4354)
         );
  NOR2_X1 U4873 ( .A1(n5981), .A2(n4354), .ZN(n4355) );
  OR2_X1 U4874 ( .A1(n5936), .A2(n4355), .ZN(n6168) );
  OAI22_X1 U4875 ( .A1(n6073), .A2(n6978), .B1(n7004), .B2(n6168), .ZN(n4370)
         );
  NAND2_X1 U4876 ( .A1(n5826), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6999) );
  INV_X1 U4877 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6608) );
  INV_X1 U4878 ( .A(n5826), .ZN(n5197) );
  INV_X1 U4879 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6604) );
  INV_X1 U4880 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6974) );
  NAND2_X1 U4881 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .ZN(
        n5354) );
  INV_X1 U4882 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U4883 ( .A1(n5354), .A2(n6577), .ZN(n6870) );
  NAND2_X1 U4884 ( .A1(n6870), .A2(REIP_REG_4__SCAN_IN), .ZN(n6883) );
  INV_X1 U4885 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6882) );
  NOR2_X1 U4886 ( .A1(n6883), .A2(n6882), .ZN(n5481) );
  NAND2_X1 U4887 ( .A1(n5481), .A2(REIP_REG_6__SCAN_IN), .ZN(n6891) );
  INV_X1 U4888 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6582) );
  NOR2_X1 U4889 ( .A1(n6891), .A2(n6582), .ZN(n5201) );
  NAND2_X1 U4890 ( .A1(n5201), .A2(REIP_REG_8__SCAN_IN), .ZN(n6904) );
  INV_X1 U4891 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4356) );
  NOR2_X1 U4892 ( .A1(n6904), .A2(n4356), .ZN(n6923) );
  NAND2_X1 U4893 ( .A1(n6923), .A2(REIP_REG_10__SCAN_IN), .ZN(n5497) );
  INV_X1 U4894 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6588) );
  NOR2_X1 U4895 ( .A1(n5497), .A2(n6588), .ZN(n5498) );
  INV_X1 U4896 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6939) );
  INV_X1 U4897 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6592) );
  INV_X1 U4898 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6949) );
  NOR3_X1 U4899 ( .A1(n6939), .A2(n6592), .A3(n6949), .ZN(n5721) );
  NAND2_X1 U4900 ( .A1(n5721), .A2(REIP_REG_15__SCAN_IN), .ZN(n5738) );
  INV_X1 U4901 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6843) );
  INV_X1 U4902 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6594) );
  NOR3_X1 U4903 ( .A1(n5738), .A2(n6843), .A3(n6594), .ZN(n6954) );
  NAND4_X1 U4904 ( .A1(n5498), .A2(n6954), .A3(REIP_REG_18__SCAN_IN), .A4(
        REIP_REG_19__SCAN_IN), .ZN(n6975) );
  NOR2_X1 U4905 ( .A1(n6974), .A2(n6975), .ZN(n6988) );
  NAND2_X1 U4906 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6988), .ZN(n5750) );
  NOR2_X1 U4907 ( .A1(n6604), .A2(n5750), .ZN(n6997) );
  NAND2_X1 U4908 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6997), .ZN(n5823) );
  INV_X1 U4909 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4357) );
  NAND2_X1 U4910 ( .A1(n4358), .A2(n4357), .ZN(n6733) );
  INV_X1 U4911 ( .A(n6733), .ZN(n4727) );
  NAND2_X1 U4912 ( .A1(n4733), .A2(n4727), .ZN(n4359) );
  AOI21_X1 U4913 ( .B1(n5861), .B2(n4359), .A(n4364), .ZN(n4360) );
  AND2_X1 U4914 ( .A1(n6986), .A2(n5826), .ZN(n6941) );
  INV_X1 U4915 ( .A(n6941), .ZN(n5396) );
  OAI21_X1 U4916 ( .B1(n5197), .B2(n5823), .A(n5396), .ZN(n7000) );
  NAND2_X1 U4917 ( .A1(n6998), .A2(n6608), .ZN(n5939) );
  OAI22_X1 U4918 ( .A1(n6608), .A2(n7000), .B1(n5823), .B2(n5939), .ZN(n4361)
         );
  AOI21_X1 U4919 ( .B1(PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6968), .A(n4361), 
        .ZN(n4368) );
  INV_X1 U4920 ( .A(n4362), .ZN(n4363) );
  NAND2_X1 U4921 ( .A1(n6981), .A2(n6074), .ZN(n4367) );
  OR2_X1 U4922 ( .A1(n6733), .A2(n4364), .ZN(n7051) );
  AND2_X1 U4923 ( .A1(n5856), .A2(n7051), .ZN(n5871) );
  INV_X1 U4924 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5963) );
  AND3_X1 U4925 ( .A1(n4733), .A2(n5963), .A3(n4364), .ZN(n4365) );
  NOR2_X1 U4926 ( .A1(n5871), .A2(n4365), .ZN(n4366) );
  NAND3_X1 U4927 ( .A1(n4368), .A2(n4367), .A3(n3459), .ZN(n4369) );
  NAND2_X1 U4928 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n4730), .ZN(n6736) );
  INV_X1 U4929 ( .A(n6736), .ZN(n4373) );
  NAND2_X1 U4930 ( .A1(n7146), .A2(n4373), .ZN(n6121) );
  NAND2_X1 U4931 ( .A1(n4374), .A2(n4435), .ZN(n4382) );
  NAND2_X1 U4932 ( .A1(n4383), .A2(n4375), .ZN(n4390) );
  OAI21_X1 U4933 ( .B1(n4383), .B2(n4375), .A(n4390), .ZN(n4376) );
  INV_X1 U4934 ( .A(n4376), .ZN(n4380) );
  NAND3_X1 U4935 ( .A1(n4377), .A2(n4378), .A3(n3602), .ZN(n4379) );
  AOI21_X1 U4936 ( .B1(n4380), .B2(n5856), .A(n4379), .ZN(n4381) );
  NAND2_X1 U4937 ( .A1(n4382), .A2(n4381), .ZN(n5575) );
  INV_X1 U4938 ( .A(n4435), .ZN(n4446) );
  INV_X1 U4939 ( .A(n5856), .ZN(n6741) );
  NAND2_X1 U4940 ( .A1(n4939), .A2(n3602), .ZN(n4393) );
  OAI21_X1 U4941 ( .B1(n6741), .B2(n4383), .A(n4393), .ZN(n4384) );
  INV_X1 U4942 ( .A(n4384), .ZN(n4385) );
  NAND2_X1 U4943 ( .A1(n4860), .A2(n6764), .ZN(n4387) );
  INV_X1 U4944 ( .A(n4389), .ZN(n4391) );
  NAND2_X1 U4945 ( .A1(n4390), .A2(n4391), .ZN(n4399) );
  OAI21_X1 U4946 ( .B1(n4391), .B2(n4390), .A(n4399), .ZN(n4392) );
  NAND2_X1 U4947 ( .A1(n4392), .A2(n5856), .ZN(n4394) );
  NAND2_X1 U4948 ( .A1(n4394), .A2(n4393), .ZN(n4395) );
  OAI21_X1 U4949 ( .B1(n6666), .B2(n6806), .A(n6664), .ZN(n4398) );
  NAND2_X1 U4950 ( .A1(n6666), .A2(n6806), .ZN(n4397) );
  NAND2_X1 U4951 ( .A1(n4398), .A2(n4397), .ZN(n6674) );
  NAND2_X1 U4952 ( .A1(n4399), .A2(n4400), .ZN(n4415) );
  OAI211_X1 U4953 ( .C1(n4400), .C2(n4399), .A(n4415), .B(n5856), .ZN(n4401)
         );
  INV_X1 U4954 ( .A(n4401), .ZN(n4402) );
  AOI21_X1 U4955 ( .B1(n4403), .B2(n4435), .A(n4402), .ZN(n6672) );
  OAI21_X1 U4956 ( .B1(n6674), .B2(n6777), .A(n6672), .ZN(n4405) );
  NAND2_X1 U4957 ( .A1(n6674), .A2(n6777), .ZN(n4404) );
  NAND2_X1 U4958 ( .A1(n4405), .A2(n4404), .ZN(n6681) );
  INV_X1 U4959 ( .A(n6681), .ZN(n4410) );
  XNOR2_X1 U4960 ( .A(n4415), .B(n4413), .ZN(n4406) );
  NAND2_X1 U4961 ( .A1(n4406), .A2(n5856), .ZN(n4407) );
  XNOR2_X1 U4962 ( .A(n4411), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6682)
         );
  INV_X1 U4963 ( .A(n6682), .ZN(n4409) );
  NAND2_X1 U4964 ( .A1(n4410), .A2(n4409), .ZN(n6680) );
  NAND2_X1 U4965 ( .A1(n4411), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6686)
         );
  NAND2_X1 U4966 ( .A1(n4412), .A2(n4435), .ZN(n4418) );
  INV_X1 U4967 ( .A(n4413), .ZN(n4414) );
  OR2_X1 U4968 ( .A1(n4415), .A2(n4414), .ZN(n4421) );
  XNOR2_X1 U4969 ( .A(n4421), .B(n4422), .ZN(n4416) );
  NAND2_X1 U4970 ( .A1(n4416), .A2(n5856), .ZN(n4417) );
  NAND2_X1 U4971 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4429)
         );
  AND2_X1 U4972 ( .A1(n6686), .A2(n4429), .ZN(n4419) );
  NAND2_X1 U4973 ( .A1(n6680), .A2(n4419), .ZN(n5508) );
  NAND3_X1 U4974 ( .A1(n4449), .A2(n4420), .A3(n4435), .ZN(n4426) );
  INV_X1 U4975 ( .A(n4421), .ZN(n4423) );
  NAND2_X1 U4976 ( .A1(n4423), .A2(n4422), .ZN(n4437) );
  XNOR2_X1 U4977 ( .A(n4437), .B(n4438), .ZN(n4424) );
  NAND2_X1 U4978 ( .A1(n4424), .A2(n5856), .ZN(n4425) );
  NAND2_X1 U4979 ( .A1(n5509), .A2(n4427), .ZN(n4431) );
  INV_X1 U4980 ( .A(n6687), .ZN(n4430) );
  NAND2_X1 U4981 ( .A1(n4430), .A2(n4429), .ZN(n5507) );
  NAND3_X1 U4982 ( .A1(n5508), .A2(n4431), .A3(n5507), .ZN(n4434) );
  NAND2_X1 U4983 ( .A1(n4432), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4433)
         );
  NAND2_X1 U4984 ( .A1(n4434), .A2(n4433), .ZN(n5586) );
  NAND2_X1 U4985 ( .A1(n4436), .A2(n4435), .ZN(n4442) );
  INV_X1 U4986 ( .A(n4437), .ZN(n4439) );
  NAND2_X1 U4987 ( .A1(n4439), .A2(n4438), .ZN(n4451) );
  XNOR2_X1 U4988 ( .A(n4451), .B(n4445), .ZN(n4440) );
  NAND2_X1 U4989 ( .A1(n4440), .A2(n5856), .ZN(n4441) );
  NAND2_X1 U4990 ( .A1(n4442), .A2(n4441), .ZN(n4443) );
  XNOR2_X1 U4991 ( .A(n4443), .B(n6817), .ZN(n5588) );
  NAND2_X1 U4992 ( .A1(n5856), .A2(n4445), .ZN(n4450) );
  NOR2_X1 U4993 ( .A1(n4447), .A2(n4446), .ZN(n4448) );
  OAI21_X1 U4994 ( .B1(n4451), .B2(n4450), .A(n4640), .ZN(n4452) );
  XNOR2_X1 U4995 ( .A(n4452), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5438)
         );
  INV_X1 U4996 ( .A(n4452), .ZN(n4453) );
  XNOR2_X1 U4997 ( .A(n4640), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5582)
         );
  NAND2_X1 U4998 ( .A1(n6106), .A2(n6830), .ZN(n5637) );
  OR3_X1 U4999 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n4456) );
  NOR2_X2 U5000 ( .A1(n4459), .A2(n4458), .ZN(n5614) );
  XNOR2_X1 U5001 ( .A(n6106), .B(n5616), .ZN(n5615) );
  OAI22_X1 U5002 ( .A1(n5614), .A2(n5615), .B1(n4460), .B2(
        INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5648) );
  XNOR2_X1 U5003 ( .A(n6106), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5647)
         );
  NAND2_X1 U5004 ( .A1(n5646), .A2(n3457), .ZN(n5698) );
  XNOR2_X1 U5005 ( .A(n6106), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5700)
         );
  NAND2_X1 U5006 ( .A1(n3427), .A2(n3432), .ZN(n6115) );
  NOR2_X2 U5007 ( .A1(n6115), .A2(n4461), .ZN(n4464) );
  INV_X1 U5008 ( .A(n4464), .ZN(n6080) );
  NAND2_X1 U5009 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4466) );
  NAND3_X1 U5010 ( .A1(n6108), .A2(n6105), .A3(n4462), .ZN(n4463) );
  XNOR2_X1 U5012 ( .A(n4460), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6709)
         );
  NOR2_X2 U5013 ( .A1(n6708), .A2(n6709), .ZN(n6097) );
  XNOR2_X1 U5014 ( .A(n4460), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6089)
         );
  NOR2_X1 U5015 ( .A1(n6106), .A2(n6069), .ZN(n6088) );
  NOR2_X1 U5016 ( .A1(n6089), .A2(n6088), .ZN(n4468) );
  AND2_X1 U5017 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6207) );
  AOI21_X1 U5018 ( .B1(n6207), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n4460), 
        .ZN(n4467) );
  AOI21_X1 U5019 ( .B1(n6097), .B2(n4468), .A(n4467), .ZN(n6070) );
  XNOR2_X1 U5020 ( .A(n6106), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4469)
         );
  XNOR2_X1 U5021 ( .A(n6070), .B(n4469), .ZN(n6194) );
  NAND2_X1 U5022 ( .A1(n4472), .A2(n4939), .ZN(n4473) );
  AND2_X1 U5023 ( .A1(n4471), .A2(n4473), .ZN(n4662) );
  AND2_X1 U5024 ( .A1(n4474), .A2(n4662), .ZN(n7034) );
  NAND2_X1 U5025 ( .A1(n7034), .A2(n7047), .ZN(n4475) );
  INV_X1 U5026 ( .A(n7146), .ZN(n7132) );
  NAND2_X1 U5027 ( .A1(n7132), .A2(n4476), .ZN(n6740) );
  NAND2_X1 U5028 ( .A1(n6740), .A2(n7072), .ZN(n4477) );
  NAND2_X1 U5029 ( .A1(n7072), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4479) );
  NAND2_X1 U5030 ( .A1(n7080), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4478) );
  NAND2_X1 U5031 ( .A1(n4479), .A2(n4478), .ZN(n4862) );
  INV_X1 U5032 ( .A(n4480), .ZN(n6771) );
  NAND2_X1 U5033 ( .A1(n6771), .A2(REIP_REG_22__SCAN_IN), .ZN(n6186) );
  OAI21_X1 U5034 ( .B1(n6101), .B2(n4481), .A(n6186), .ZN(n4482) );
  NOR2_X1 U5035 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6190) );
  NOR2_X1 U5036 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6208) );
  NAND4_X1 U5037 ( .A1(n6190), .A2(n6208), .A3(n6171), .A4(n6180), .ZN(n4486)
         );
  AND2_X1 U5038 ( .A1(n4460), .A2(n4486), .ZN(n4487) );
  AND2_X1 U5039 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U5040 ( .A1(n6207), .A2(n6189), .ZN(n6081) );
  NAND2_X1 U5041 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4717) );
  NOR2_X1 U5042 ( .A1(n6081), .A2(n4717), .ZN(n4701) );
  XNOR2_X1 U5043 ( .A(n6106), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6061)
         );
  NAND2_X1 U5044 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4702) );
  AND2_X1 U5045 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U5046 ( .A1(n4722), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n6133) );
  OAI21_X1 U5047 ( .B1(n4702), .B2(n6133), .A(n6106), .ZN(n4490) );
  NOR3_X1 U5048 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n4489) );
  NOR2_X1 U5049 ( .A1(n6106), .A2(n4489), .ZN(n4639) );
  NAND2_X1 U5050 ( .A1(n4495), .A2(n4494), .ZN(n4496) );
  NAND2_X1 U5051 ( .A1(n4557), .A2(n4496), .ZN(n6047) );
  AOI22_X1 U5052 ( .A1(n4110), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4497), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4501) );
  AOI22_X1 U5053 ( .A1(n4612), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4500) );
  AOI22_X1 U5054 ( .A1(n4602), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4499) );
  AOI22_X1 U5055 ( .A1(n3675), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4498) );
  NAND4_X1 U5056 ( .A1(n4501), .A2(n4500), .A3(n4499), .A4(n4498), .ZN(n4507)
         );
  AOI22_X1 U5057 ( .A1(n4611), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4505) );
  AOI22_X1 U5058 ( .A1(n3657), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4504) );
  AOI22_X1 U5059 ( .A1(n4603), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5060 ( .A1(n4604), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4502) );
  NAND4_X1 U5061 ( .A1(n4505), .A2(n4504), .A3(n4503), .A4(n4502), .ZN(n4506)
         );
  NOR2_X1 U5062 ( .A1(n4507), .A2(n4506), .ZN(n4559) );
  AOI22_X1 U5063 ( .A1(n4497), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4511) );
  AOI22_X1 U5064 ( .A1(n4603), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4510) );
  AOI22_X1 U5065 ( .A1(n3677), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5066 ( .A1(n4602), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4508) );
  NAND4_X1 U5067 ( .A1(n4511), .A2(n4510), .A3(n4509), .A4(n4508), .ZN(n4517)
         );
  AOI22_X1 U5068 ( .A1(n4110), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5069 ( .A1(n3675), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4514) );
  AOI22_X1 U5070 ( .A1(n4612), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4513) );
  AOI22_X1 U5071 ( .A1(n4604), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4512) );
  NAND4_X1 U5072 ( .A1(n4515), .A2(n4514), .A3(n4513), .A4(n4512), .ZN(n4516)
         );
  NOR2_X1 U5073 ( .A1(n4517), .A2(n4516), .ZN(n4539) );
  INV_X1 U5074 ( .A(n4518), .ZN(n4519) );
  OR2_X1 U5075 ( .A1(n4520), .A2(n4519), .ZN(n4540) );
  NOR2_X1 U5076 ( .A1(n4539), .A2(n4540), .ZN(n4550) );
  AOI22_X1 U5077 ( .A1(n4497), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4524) );
  AOI22_X1 U5078 ( .A1(n4110), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4523) );
  AOI22_X1 U5079 ( .A1(n4603), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5080 ( .A1(n4612), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3757), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4521) );
  NAND4_X1 U5081 ( .A1(n4524), .A2(n4523), .A3(n4522), .A4(n4521), .ZN(n4530)
         );
  AOI22_X1 U5082 ( .A1(n3675), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5083 ( .A1(n4604), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4527) );
  AOI22_X1 U5084 ( .A1(n3677), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4526) );
  AOI22_X1 U5085 ( .A1(n4602), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4525) );
  NAND4_X1 U5086 ( .A1(n4528), .A2(n4527), .A3(n4526), .A4(n4525), .ZN(n4529)
         );
  OR2_X1 U5087 ( .A1(n4530), .A2(n4529), .ZN(n4551) );
  NAND2_X1 U5088 ( .A1(n4550), .A2(n4551), .ZN(n4558) );
  XNOR2_X1 U5089 ( .A(n4559), .B(n4558), .ZN(n4533) );
  AOI21_X1 U5090 ( .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6226), .A(n4555), 
        .ZN(n4532) );
  NAND2_X1 U5091 ( .A1(n5866), .A2(EAX_REG_27__SCAN_IN), .ZN(n4531) );
  OAI211_X1 U5092 ( .C1(n4533), .C2(n4596), .A(n4532), .B(n4531), .ZN(n4534)
         );
  OAI21_X1 U5093 ( .B1(n6047), .B2(n4623), .A(n4534), .ZN(n5907) );
  INV_X1 U5094 ( .A(n5907), .ZN(n4556) );
  INV_X1 U5095 ( .A(n4535), .ZN(n4537) );
  INV_X1 U5096 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4536) );
  NAND2_X1 U5097 ( .A1(n4537), .A2(n4536), .ZN(n4538) );
  NAND2_X1 U5098 ( .A1(n4547), .A2(n4538), .ZN(n6065) );
  XNOR2_X1 U5099 ( .A(n4540), .B(n4539), .ZN(n4543) );
  AOI21_X1 U5100 ( .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6226), .A(n4555), 
        .ZN(n4542) );
  NAND2_X1 U5101 ( .A1(n5866), .A2(EAX_REG_25__SCAN_IN), .ZN(n4541) );
  OAI211_X1 U5102 ( .C1(n4543), .C2(n4596), .A(n4542), .B(n4541), .ZN(n4544)
         );
  OAI21_X1 U5103 ( .B1(n6065), .B2(n4623), .A(n4544), .ZN(n5933) );
  INV_X1 U5104 ( .A(n5933), .ZN(n4546) );
  AND2_X1 U5105 ( .A1(n4546), .A2(n4545), .ZN(n5916) );
  XNOR2_X1 U5106 ( .A(n4547), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5923)
         );
  NOR2_X1 U5107 ( .A1(n4548), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4549) );
  AOI211_X1 U5108 ( .C1(n5866), .C2(EAX_REG_26__SCAN_IN), .A(n4555), .B(n4549), 
        .ZN(n4554) );
  XOR2_X1 U5109 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND2_X1 U5110 ( .A1(n4552), .A2(n4627), .ZN(n4553) );
  AOI22_X1 U5111 ( .A1(n5923), .A2(n4555), .B1(n4554), .B2(n4553), .ZN(n5919)
         );
  AND2_X1 U5112 ( .A1(n5916), .A2(n5919), .ZN(n5905) );
  XNOR2_X1 U5113 ( .A(n4557), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5890)
         );
  INV_X1 U5114 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5891) );
  AOI21_X1 U5115 ( .B1(n5891), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4574) );
  NOR2_X1 U5116 ( .A1(n4559), .A2(n4558), .ZN(n4581) );
  AOI22_X1 U5117 ( .A1(n4497), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4564) );
  AOI22_X1 U5118 ( .A1(n4110), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4560), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5119 ( .A1(n4603), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4582), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4562) );
  AOI22_X1 U5120 ( .A1(n4612), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4561) );
  NAND4_X1 U5121 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4571)
         );
  AOI22_X1 U5122 ( .A1(n3644), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5123 ( .A1(n4604), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5124 ( .A1(n3677), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4567) );
  AOI22_X1 U5125 ( .A1(n4602), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4566) );
  NAND4_X1 U5126 ( .A1(n4569), .A2(n4568), .A3(n4567), .A4(n4566), .ZN(n4570)
         );
  OR2_X1 U5127 ( .A1(n4571), .A2(n4570), .ZN(n4580) );
  XNOR2_X1 U5128 ( .A(n4581), .B(n4580), .ZN(n4572) );
  NOR2_X1 U5129 ( .A1(n4572), .A2(n4596), .ZN(n4573) );
  AOI211_X1 U5130 ( .C1(n5866), .C2(EAX_REG_28__SCAN_IN), .A(n4574), .B(n4573), 
        .ZN(n4575) );
  AOI21_X1 U5131 ( .B1(n5890), .B2(n4555), .A(n4575), .ZN(n5780) );
  NAND2_X2 U5132 ( .A1(n4577), .A2(n4576), .ZN(n5779) );
  NAND2_X1 U5133 ( .A1(n4578), .A2(n5880), .ZN(n4579) );
  NAND2_X1 U5134 ( .A1(n4599), .A2(n4579), .ZN(n5884) );
  NAND2_X1 U5135 ( .A1(n4581), .A2(n4580), .ZN(n4600) );
  AOI22_X1 U5136 ( .A1(n4087), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4587) );
  AOI22_X1 U5137 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n4582), .B1(n3757), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4586) );
  AOI22_X1 U5138 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n4604), .B1(n4583), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5139 ( .A1(n3675), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4584) );
  NAND4_X1 U5140 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4593)
         );
  AOI22_X1 U5141 ( .A1(n4110), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4606), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4591) );
  AOI22_X1 U5142 ( .A1(n4612), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4603), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4590) );
  AOI22_X1 U5143 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n4602), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5144 ( .A1(n3657), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4588) );
  NAND4_X1 U5145 ( .A1(n4591), .A2(n4590), .A3(n4589), .A4(n4588), .ZN(n4592)
         );
  NOR2_X1 U5146 ( .A1(n4593), .A2(n4592), .ZN(n4601) );
  XNOR2_X1 U5147 ( .A(n4600), .B(n4601), .ZN(n4597) );
  AOI21_X1 U5148 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6226), .A(n4555), 
        .ZN(n4595) );
  NAND2_X1 U5149 ( .A1(n5866), .A2(EAX_REG_29__SCAN_IN), .ZN(n4594) );
  OAI211_X1 U5150 ( .C1(n4597), .C2(n4596), .A(n4595), .B(n4594), .ZN(n4598)
         );
  OAI21_X1 U5151 ( .B1(n5884), .B2(n4623), .A(n4598), .ZN(n5801) );
  XNOR2_X1 U5152 ( .A(n4599), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5822)
         );
  NOR2_X1 U5153 ( .A1(n4601), .A2(n4600), .ZN(n4622) );
  AOI22_X1 U5154 ( .A1(n4602), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3657), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4610) );
  AOI22_X1 U5155 ( .A1(n4603), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3749), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4609) );
  AOI22_X1 U5156 ( .A1(n4604), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4565), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4608) );
  AOI22_X1 U5157 ( .A1(n4606), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4605), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4607) );
  NAND4_X1 U5158 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4620)
         );
  AOI22_X1 U5159 ( .A1(n4087), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4611), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4618) );
  AOI22_X1 U5160 ( .A1(n4110), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4612), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4617) );
  AOI22_X1 U5161 ( .A1(n3675), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4613), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U5162 ( .A1(n4583), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4614), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4615) );
  NAND4_X1 U5163 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4619)
         );
  NOR2_X1 U5164 ( .A1(n4620), .A2(n4619), .ZN(n4621) );
  XNOR2_X1 U5165 ( .A(n4622), .B(n4621), .ZN(n4628) );
  INV_X1 U5166 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4625) );
  NAND2_X1 U5167 ( .A1(n6226), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4624)
         );
  OAI211_X1 U5168 ( .C1(n3453), .C2(n4625), .A(n4624), .B(n4623), .ZN(n4626)
         );
  AOI21_X1 U5169 ( .B1(n4628), .B2(n4627), .A(n4626), .ZN(n4629) );
  AOI21_X1 U5170 ( .B1(n5822), .B2(n4555), .A(n4629), .ZN(n5867) );
  XNOR2_X1 U5171 ( .A(n5868), .B(n5867), .ZN(n5841) );
  NOR2_X1 U5172 ( .A1(n5841), .A2(n6121), .ZN(n4634) );
  INV_X1 U5173 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4630) );
  NAND2_X1 U5174 ( .A1(n6771), .A2(REIP_REG_30__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U5175 ( .B1(n6101), .B2(n4630), .A(n6135), .ZN(n4631) );
  OAI21_X1 U5176 ( .B1(n6141), .B2(n6696), .A(n4635), .ZN(U2956) );
  INV_X1 U5177 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n6051) );
  NOR2_X2 U5178 ( .A1(n6053), .A2(n4636), .ZN(n6043) );
  NAND2_X1 U5179 ( .A1(n6106), .A2(n4637), .ZN(n4638) );
  NAND2_X1 U5180 ( .A1(n6043), .A2(n4638), .ZN(n6034) );
  INV_X1 U5181 ( .A(n4639), .ZN(n4641) );
  AOI22_X1 U5182 ( .A1(n6034), .A2(n4641), .B1(n5776), .B2(n4640), .ZN(n4644)
         );
  AOI21_X1 U5183 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6106), .A(n6029), 
        .ZN(n4642) );
  INV_X1 U5184 ( .A(n4642), .ZN(n4643) );
  XNOR2_X1 U5185 ( .A(n4644), .B(n4643), .ZN(n5806) );
  NAND2_X1 U5186 ( .A1(n7088), .A2(n5849), .ZN(n4814) );
  AOI21_X1 U5187 ( .B1(n4751), .B2(n6733), .A(n4814), .ZN(n4647) );
  NOR2_X1 U5188 ( .A1(n3600), .A2(n4939), .ZN(n4645) );
  NOR2_X1 U5189 ( .A1(n5854), .A2(n4645), .ZN(n4646) );
  MUX2_X1 U5190 ( .A(n4647), .B(n4646), .S(n4377), .Z(n4648) );
  INV_X1 U5191 ( .A(n4648), .ZN(n4660) );
  OR2_X1 U5192 ( .A1(n4841), .A2(n3604), .ZN(n4699) );
  INV_X1 U5193 ( .A(n4699), .ZN(n4658) );
  OR2_X1 U5194 ( .A1(n4649), .A2(n3443), .ZN(n4652) );
  NAND2_X1 U5195 ( .A1(n3444), .A2(n4733), .ZN(n4650) );
  NAND2_X1 U5196 ( .A1(n6741), .A2(n4650), .ZN(n4651) );
  NAND2_X1 U5197 ( .A1(n4652), .A2(n4651), .ZN(n4689) );
  NAND2_X1 U5198 ( .A1(n4662), .A2(n4689), .ZN(n4653) );
  NAND2_X1 U5199 ( .A1(n4653), .A2(n4258), .ZN(n4830) );
  OAI21_X1 U5200 ( .B1(n4751), .B2(n4727), .A(n4826), .ZN(n4655) );
  INV_X1 U5201 ( .A(n4655), .ZN(n4656) );
  NAND2_X1 U5202 ( .A1(n4654), .A2(n4656), .ZN(n4827) );
  NAND2_X1 U5203 ( .A1(n4830), .A2(n4827), .ZN(n4657) );
  AOI21_X1 U5204 ( .B1(n5854), .B2(n4658), .A(n4657), .ZN(n4659) );
  NAND2_X1 U5205 ( .A1(n4660), .A2(n4659), .ZN(n4661) );
  NAND2_X1 U5206 ( .A1(n4662), .A2(n5349), .ZN(n4815) );
  INV_X1 U5207 ( .A(n4815), .ZN(n5145) );
  NOR2_X1 U5208 ( .A1(n5145), .A2(n7034), .ZN(n5845) );
  INV_X1 U5209 ( .A(n4663), .ZN(n4664) );
  AOI22_X1 U5210 ( .A1(n4664), .A2(n3587), .B1(n4767), .B2(n4654), .ZN(n4665)
         );
  NAND3_X1 U5211 ( .A1(n5845), .A2(n4665), .A3(n5175), .ZN(n4666) );
  NAND2_X1 U5212 ( .A1(n4654), .A2(n5856), .ZN(n7052) );
  OAI21_X1 U5213 ( .B1(n4663), .B2(n3587), .A(n7052), .ZN(n4667) );
  MUX2_X1 U5214 ( .A(n4668), .B(n4268), .S(EBX_REG_25__SCAN_IN), .Z(n4670) );
  NOR2_X1 U5215 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4669)
         );
  NOR2_X1 U5216 ( .A1(n4670), .A2(n4669), .ZN(n5935) );
  INV_X1 U5217 ( .A(EBX_REG_26__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U5218 ( .A1(n4678), .A2(n4671), .ZN(n4674) );
  NAND2_X1 U5219 ( .A1(n4679), .A2(n6051), .ZN(n4672) );
  OAI211_X1 U5220 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5861), .A(n4672), .B(n5859), 
        .ZN(n4673) );
  AND2_X1 U5221 ( .A1(n4674), .A2(n4673), .ZN(n5920) );
  MUX2_X1 U5222 ( .A(n4675), .B(n5859), .S(EBX_REG_27__SCAN_IN), .Z(n4677) );
  NAND2_X1 U5223 ( .A1(n4823), .A2(n4637), .ZN(n4676) );
  NAND2_X1 U5224 ( .A1(n4677), .A2(n4676), .ZN(n5902) );
  OR2_X2 U5225 ( .A1(n5922), .A2(n5902), .ZN(n5904) );
  INV_X1 U5226 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U5227 ( .A1(n4678), .A2(n5968), .ZN(n4682) );
  INV_X1 U5228 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U5229 ( .A1(n4679), .A2(n5776), .ZN(n4680) );
  OAI211_X1 U5230 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5861), .A(n4680), .B(n5859), 
        .ZN(n4681) );
  AND2_X1 U5231 ( .A1(n4682), .A2(n4681), .ZN(n5784) );
  NOR2_X4 U5232 ( .A1(n5904), .A2(n5784), .ZN(n5819) );
  INV_X1 U5233 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5966) );
  AND2_X1 U5234 ( .A1(n3426), .A2(n5966), .ZN(n4684) );
  INV_X1 U5235 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4683) );
  AOI21_X1 U5236 ( .B1(n4823), .B2(n4683), .A(n4684), .ZN(n5820) );
  MUX2_X1 U5237 ( .A(n4684), .B(n5820), .S(n5859), .Z(n4685) );
  NAND2_X1 U5238 ( .A1(n5819), .A2(n4685), .ZN(n5858) );
  OR2_X1 U5239 ( .A1(n5819), .A2(n4685), .ZN(n4686) );
  NAND2_X1 U5240 ( .A1(n5858), .A2(n4686), .ZN(n5965) );
  INV_X1 U5241 ( .A(n5965), .ZN(n4704) );
  INV_X1 U5242 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6332) );
  NOR2_X1 U5243 ( .A1(n4480), .A2(n6332), .ZN(n5802) );
  NOR2_X1 U5244 ( .A1(n4258), .A2(n3604), .ZN(n5814) );
  INV_X1 U5245 ( .A(n6755), .ZN(n4697) );
  INV_X1 U5246 ( .A(n6858), .ZN(n5632) );
  NAND2_X1 U5247 ( .A1(n4939), .A2(n4751), .ZN(n5343) );
  OR2_X1 U5248 ( .A1(n5343), .A2(n4687), .ZN(n4829) );
  OAI21_X1 U5249 ( .B1(n3600), .B2(n4377), .A(n4829), .ZN(n4688) );
  INV_X1 U5250 ( .A(n4688), .ZN(n4690) );
  OAI211_X1 U5251 ( .C1(n4471), .C2(n4823), .A(n4690), .B(n4689), .ZN(n4691)
         );
  NOR2_X1 U5252 ( .A1(n4692), .A2(n4691), .ZN(n4840) );
  NAND2_X1 U5253 ( .A1(n4693), .A2(n3711), .ZN(n4695) );
  INV_X1 U5254 ( .A(n3630), .ZN(n4694) );
  OR2_X1 U5255 ( .A1(n4841), .A2(n4694), .ZN(n5154) );
  NAND3_X1 U5256 ( .A1(n4840), .A2(n4695), .A3(n5154), .ZN(n4696) );
  NAND2_X1 U5257 ( .A1(n4706), .A2(n4696), .ZN(n5622) );
  NAND2_X1 U5258 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6779) );
  NOR3_X1 U5259 ( .A1(n4427), .A2(n5598), .A3(n6779), .ZN(n5444) );
  NAND3_X1 U5260 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n5444), .ZN(n4700) );
  NAND2_X1 U5261 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6794) );
  NOR2_X1 U5262 ( .A1(n4700), .A2(n6794), .ZN(n5566) );
  NAND3_X1 U5263 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5566), .ZN(n5631) );
  NOR2_X1 U5264 ( .A1(n4698), .A2(n4699), .ZN(n5843) );
  AOI21_X1 U5265 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6795) );
  NOR2_X1 U5266 ( .A1(n6795), .A2(n4700), .ZN(n5563) );
  NAND3_X1 U5267 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n5563), .ZN(n5621) );
  NOR2_X1 U5268 ( .A1(n6798), .A2(n5621), .ZN(n5618) );
  NOR2_X1 U5269 ( .A1(n4457), .A2(n6830), .ZN(n5671) );
  NAND2_X1 U5270 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5671), .ZN(n5704) );
  NOR2_X1 U5271 ( .A1(n5703), .A2(n5704), .ZN(n5702) );
  NAND3_X1 U5272 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5702), .ZN(n6841) );
  NOR2_X1 U5273 ( .A1(n4462), .A2(n6841), .ZN(n6214) );
  NAND2_X1 U5274 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6214), .ZN(n4709) );
  INV_X1 U5275 ( .A(n4701), .ZN(n6151) );
  NOR2_X1 U5276 ( .A1(n6753), .A2(n6151), .ZN(n6155) );
  INV_X1 U5277 ( .A(n4702), .ZN(n4720) );
  NAND2_X1 U5278 ( .A1(n6155), .A2(n4720), .ZN(n6134) );
  INV_X1 U5279 ( .A(n4722), .ZN(n5788) );
  NOR3_X1 U5280 ( .A1(n6134), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5788), 
        .ZN(n4703) );
  AOI211_X1 U5281 ( .C1(n6860), .C2(n4704), .A(n5802), .B(n4703), .ZN(n4725)
         );
  INV_X1 U5282 ( .A(n4709), .ZN(n4705) );
  OR2_X1 U5283 ( .A1(n5567), .A2(n4705), .ZN(n4708) );
  INV_X1 U5284 ( .A(n5567), .ZN(n5441) );
  INV_X1 U5285 ( .A(n5622), .ZN(n4707) );
  INV_X1 U5286 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6855) );
  NOR2_X1 U5287 ( .A1(n6771), .A2(n4706), .ZN(n6857) );
  AOI21_X1 U5288 ( .B1(n4707), .B2(n6855), .A(n6857), .ZN(n5565) );
  INV_X1 U5289 ( .A(n5565), .ZN(n5440) );
  AOI21_X1 U5290 ( .B1(n5441), .B2(n5631), .A(n5440), .ZN(n5619) );
  AND2_X1 U5291 ( .A1(n4708), .A2(n5619), .ZN(n4713) );
  NOR2_X1 U5292 ( .A1(n5621), .A2(n4709), .ZN(n4710) );
  OR2_X1 U5293 ( .A1(n6798), .A2(n4710), .ZN(n4711) );
  NAND2_X1 U5294 ( .A1(n4713), .A2(n4711), .ZN(n6748) );
  INV_X1 U5295 ( .A(n6207), .ZN(n4712) );
  OR2_X1 U5296 ( .A1(n6748), .A2(n4712), .ZN(n4715) );
  NAND2_X1 U5297 ( .A1(n4713), .A2(n6754), .ZN(n4714) );
  NAND2_X1 U5298 ( .A1(n4715), .A2(n4714), .ZN(n6185) );
  OR2_X1 U5299 ( .A1(n6754), .A2(n6189), .ZN(n4716) );
  NAND2_X1 U5300 ( .A1(n6185), .A2(n4716), .ZN(n6179) );
  INV_X1 U5301 ( .A(n4717), .ZN(n4718) );
  AOI21_X1 U5302 ( .B1(n6790), .B2(n6798), .A(n4718), .ZN(n4719) );
  NAND2_X1 U5303 ( .A1(n6169), .A2(n6754), .ZN(n6122) );
  NAND2_X1 U5304 ( .A1(n6169), .A2(n4720), .ZN(n4721) );
  NOR2_X1 U5305 ( .A1(n6754), .A2(n4722), .ZN(n4723) );
  OAI21_X1 U5306 ( .B1(n6145), .B2(n4723), .A(INSTADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n4724) );
  OAI21_X1 U5307 ( .B1(n5806), .B2(n6800), .A(n4726), .ZN(U2989) );
  INV_X1 U5308 ( .A(n7052), .ZN(n4728) );
  OAI211_X1 U5309 ( .C1(n4728), .C2(n5814), .A(n4727), .B(n7047), .ZN(n4729)
         );
  AND2_X1 U5310 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4730), .ZN(n6570) );
  INV_X1 U5311 ( .A(n6570), .ZN(n6533) );
  AND2_X2 U5312 ( .A1(n6572), .A2(n6533), .ZN(n6569) );
  AND2_X1 U5313 ( .A1(n6569), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  INV_X1 U5314 ( .A(n4731), .ZN(n4732) );
  INV_X1 U5315 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n7098) );
  OAI211_X1 U5316 ( .C1(n4732), .C2(n7098), .A(n4750), .B(n6724), .ZN(U2788)
         );
  INV_X1 U5317 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4736) );
  INV_X1 U5318 ( .A(n6572), .ZN(n4734) );
  NAND2_X1 U5319 ( .A1(n4734), .A2(n4733), .ZN(n6537) );
  AOI22_X1 U5320 ( .A1(n6570), .A2(UWORD_REG_0__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4735) );
  OAI21_X1 U5321 ( .B1(n4736), .B2(n6537), .A(n4735), .ZN(U2907) );
  INV_X1 U5322 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4738) );
  AOI22_X1 U5323 ( .A1(n6570), .A2(UWORD_REG_4__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4737) );
  OAI21_X1 U5324 ( .B1(n4738), .B2(n6537), .A(n4737), .ZN(U2903) );
  INV_X1 U5325 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4740) );
  AOI22_X1 U5326 ( .A1(n6570), .A2(UWORD_REG_5__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4739) );
  OAI21_X1 U5327 ( .B1(n4740), .B2(n6537), .A(n4739), .ZN(U2902) );
  AOI22_X1 U5328 ( .A1(n6570), .A2(UWORD_REG_8__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4741) );
  OAI21_X1 U5329 ( .B1(n4180), .B2(n6537), .A(n4741), .ZN(U2899) );
  INV_X1 U5330 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4743) );
  AOI22_X1 U5331 ( .A1(n6570), .A2(UWORD_REG_11__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4742) );
  OAI21_X1 U5332 ( .B1(n4743), .B2(n6537), .A(n4742), .ZN(U2896) );
  INV_X1 U5333 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4745) );
  AOI22_X1 U5334 ( .A1(n6570), .A2(UWORD_REG_12__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4744) );
  OAI21_X1 U5335 ( .B1(n4745), .B2(n6537), .A(n4744), .ZN(U2895) );
  INV_X1 U5336 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4747) );
  AOI22_X1 U5337 ( .A1(n6570), .A2(UWORD_REG_2__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4746) );
  OAI21_X1 U5338 ( .B1(n4747), .B2(n6537), .A(n4746), .ZN(U2905) );
  AOI22_X1 U5339 ( .A1(n6570), .A2(UWORD_REG_3__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4748) );
  OAI21_X1 U5340 ( .B1(n4083), .B2(n6537), .A(n4748), .ZN(U2904) );
  AOI22_X1 U5341 ( .A1(n6570), .A2(UWORD_REG_14__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4749) );
  OAI21_X1 U5342 ( .B1(n4625), .B2(n6537), .A(n4749), .ZN(U2893) );
  NAND2_X1 U5343 ( .A1(n4754), .A2(n4751), .ZN(n4911) );
  NAND2_X1 U5344 ( .A1(n4876), .A2(DATAI_5_), .ZN(n4899) );
  OR2_X1 U5345 ( .A1(n7052), .A2(n7077), .ZN(n4752) );
  OR2_X1 U5346 ( .A1(n5854), .A2(n4752), .ZN(n4753) );
  INV_X2 U5347 ( .A(n4753), .ZN(n4909) );
  AOI22_X1 U5348 ( .A1(n4909), .A2(EAX_REG_5__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n4755) );
  NAND2_X1 U5349 ( .A1(n4899), .A2(n4755), .ZN(U2944) );
  NAND2_X1 U5350 ( .A1(n4876), .A2(DATAI_7_), .ZN(n4895) );
  AOI22_X1 U5351 ( .A1(n4909), .A2(EAX_REG_7__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U5352 ( .A1(n4895), .A2(n4756), .ZN(U2946) );
  INV_X1 U5353 ( .A(DATAI_12_), .ZN(n5610) );
  OR2_X1 U5354 ( .A1(n4911), .A2(n5610), .ZN(n4885) );
  AOI22_X1 U5355 ( .A1(n4909), .A2(EAX_REG_12__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n4757) );
  NAND2_X1 U5356 ( .A1(n4885), .A2(n4757), .ZN(U2951) );
  INV_X1 U5357 ( .A(DATAI_11_), .ZN(n5517) );
  OR2_X1 U5358 ( .A1(n4911), .A2(n5517), .ZN(n4887) );
  AOI22_X1 U5359 ( .A1(n4909), .A2(EAX_REG_11__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4758) );
  NAND2_X1 U5360 ( .A1(n4887), .A2(n4758), .ZN(U2950) );
  NAND2_X1 U5361 ( .A1(n4876), .A2(DATAI_10_), .ZN(n4889) );
  AOI22_X1 U5362 ( .A1(n4909), .A2(EAX_REG_10__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n4759) );
  NAND2_X1 U5363 ( .A1(n4889), .A2(n4759), .ZN(U2949) );
  NAND2_X1 U5364 ( .A1(n4876), .A2(DATAI_9_), .ZN(n4891) );
  AOI22_X1 U5365 ( .A1(n4909), .A2(EAX_REG_9__SCAN_IN), .B1(n4867), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4760) );
  NAND2_X1 U5366 ( .A1(n4891), .A2(n4760), .ZN(U2948) );
  NOR2_X1 U5367 ( .A1(n4763), .A2(n4762), .ZN(n4764) );
  NOR2_X1 U5368 ( .A1(n4761), .A2(n4764), .ZN(n6667) );
  INV_X1 U5369 ( .A(n6667), .ZN(n5028) );
  NAND2_X1 U5370 ( .A1(n5854), .A2(n5843), .ZN(n4834) );
  NOR2_X1 U5371 ( .A1(n3587), .A2(n7077), .ZN(n4766) );
  INV_X1 U5372 ( .A(n3700), .ZN(n6006) );
  AND3_X1 U5373 ( .A1(n4766), .A2(n6006), .A3(n4765), .ZN(n4816) );
  NAND3_X1 U5374 ( .A1(n4768), .A2(n4767), .A3(n4816), .ZN(n4769) );
  NAND2_X1 U5375 ( .A1(n6663), .A2(n3700), .ZN(n6001) );
  NOR2_X1 U5376 ( .A1(n4772), .A2(n4771), .ZN(n4773) );
  OR2_X1 U5377 ( .A1(n4800), .A2(n4773), .ZN(n6792) );
  INV_X1 U5378 ( .A(n6792), .ZN(n5348) );
  AOI22_X1 U5379 ( .A1(n6649), .A2(n5348), .B1(n5970), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4774) );
  OAI21_X1 U5380 ( .B1(n5028), .B2(n6001), .A(n4774), .ZN(U2857) );
  OAI21_X1 U5381 ( .B1(n4777), .B2(n4776), .A(n4775), .ZN(n5576) );
  XNOR2_X1 U5382 ( .A(n5362), .B(n5861), .ZN(n6758) );
  INV_X1 U5383 ( .A(n6758), .ZN(n4778) );
  AOI22_X1 U5384 ( .A1(n6649), .A2(n4778), .B1(n5970), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4779) );
  OAI21_X1 U5385 ( .B1(n6005), .B2(n5576), .A(n4779), .ZN(U2858) );
  INV_X1 U5386 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4781) );
  AOI22_X1 U5387 ( .A1(n6570), .A2(UWORD_REG_9__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4780) );
  OAI21_X1 U5388 ( .B1(n4781), .B2(n6537), .A(n4780), .ZN(U2898) );
  INV_X1 U5389 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4783) );
  AOI22_X1 U5390 ( .A1(n6570), .A2(UWORD_REG_10__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4782) );
  OAI21_X1 U5391 ( .B1(n4783), .B2(n6537), .A(n4782), .ZN(U2897) );
  INV_X1 U5392 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5393 ( .A1(n6570), .A2(UWORD_REG_1__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4784) );
  OAI21_X1 U5394 ( .B1(n4785), .B2(n6537), .A(n4784), .ZN(U2906) );
  INV_X1 U5395 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4787) );
  AOI22_X1 U5396 ( .A1(n6570), .A2(UWORD_REG_13__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4786) );
  OAI21_X1 U5397 ( .B1(n4787), .B2(n6537), .A(n4786), .ZN(U2894) );
  AOI22_X1 U5398 ( .A1(n6570), .A2(UWORD_REG_6__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4788) );
  OAI21_X1 U5399 ( .B1(n4163), .B2(n6537), .A(n4788), .ZN(U2901) );
  INV_X1 U5400 ( .A(n4789), .ZN(n4791) );
  NAND2_X1 U5401 ( .A1(n4761), .A2(n4798), .ZN(n4790) );
  NAND2_X1 U5402 ( .A1(n4791), .A2(n4790), .ZN(n4793) );
  AND2_X1 U5403 ( .A1(n4793), .A2(n4853), .ZN(n6875) );
  INV_X1 U5404 ( .A(n6875), .ZN(n4820) );
  NAND2_X1 U5405 ( .A1(n4802), .A2(n4794), .ZN(n4795) );
  NAND2_X1 U5406 ( .A1(n4855), .A2(n4795), .ZN(n6869) );
  INV_X1 U5407 ( .A(n6869), .ZN(n4796) );
  AOI22_X1 U5408 ( .A1(n6649), .A2(n4796), .B1(n5970), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4797) );
  OAI21_X1 U5409 ( .B1(n4820), .B2(n6005), .A(n4797), .ZN(U2855) );
  XNOR2_X1 U5410 ( .A(n4761), .B(n4798), .ZN(n6675) );
  OR2_X1 U5411 ( .A1(n4800), .A2(n4799), .ZN(n4801) );
  AND2_X1 U5412 ( .A1(n4802), .A2(n4801), .ZN(n6772) );
  AOI22_X1 U5413 ( .A1(n6649), .A2(n6772), .B1(n5970), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4803) );
  OAI21_X1 U5414 ( .B1(n6675), .B2(n6005), .A(n4803), .ZN(U2856) );
  INV_X1 U5415 ( .A(n4853), .ZN(n4805) );
  AOI21_X1 U5416 ( .B1(n4805), .B2(n4852), .A(n4804), .ZN(n4806) );
  OR2_X1 U5417 ( .A1(n5023), .A2(n4806), .ZN(n5477) );
  AND2_X1 U5418 ( .A1(n4857), .A2(n4807), .ZN(n4808) );
  OR2_X1 U5419 ( .A1(n4808), .A2(n5025), .ZN(n5600) );
  INV_X1 U5420 ( .A(n5600), .ZN(n4809) );
  AOI22_X1 U5421 ( .A1(n6649), .A2(n4809), .B1(n5970), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4810) );
  OAI21_X1 U5422 ( .B1(n5477), .B2(n6001), .A(n4810), .ZN(U2853) );
  OAI21_X1 U5423 ( .B1(n4813), .B2(n4812), .A(n4811), .ZN(n5399) );
  OAI22_X1 U5424 ( .A1(n5854), .A2(n4815), .B1(n4814), .B2(n5175), .ZN(n4836)
         );
  AOI22_X1 U5425 ( .A1(n4836), .A2(n7047), .B1(n4693), .B2(n4816), .ZN(n4817)
         );
  NAND2_X1 U5426 ( .A1(n3444), .A2(n3700), .ZN(n4818) );
  NAND2_X2 U5427 ( .A1(n6026), .A2(n4818), .ZN(n7100) );
  INV_X1 U5428 ( .A(n4818), .ZN(n4819) );
  INV_X1 U5429 ( .A(DATAI_0_), .ZN(n6489) );
  INV_X1 U5430 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6542) );
  OAI222_X1 U5431 ( .A1(n5399), .A2(n7100), .B1(n6027), .B2(n6489), .C1(n6026), 
        .C2(n6542), .ZN(U2891) );
  INV_X1 U5432 ( .A(DATAI_4_), .ZN(n6481) );
  INV_X1 U5433 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6550) );
  OAI222_X1 U5434 ( .A1(n4820), .A2(n7100), .B1(n6027), .B2(n6481), .C1(n6026), 
        .C2(n6550), .ZN(U2887) );
  INV_X1 U5435 ( .A(DATAI_3_), .ZN(n6484) );
  INV_X1 U5436 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6548) );
  OAI222_X1 U5437 ( .A1(n6675), .A2(n7100), .B1(n6027), .B2(n6484), .C1(n6026), 
        .C2(n6548), .ZN(U2888) );
  INV_X1 U5438 ( .A(n4821), .ZN(n4822) );
  AOI21_X1 U5439 ( .B1(n4823), .B2(n6855), .A(n4822), .ZN(n6859) );
  INV_X1 U5440 ( .A(n6859), .ZN(n4825) );
  INV_X1 U5441 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4824) );
  OAI222_X1 U5442 ( .A1(n4825), .A2(n6658), .B1(n6663), .B2(n4824), .C1(n5399), 
        .C2(n6005), .ZN(U2859) );
  INV_X1 U5443 ( .A(DATAI_6_), .ZN(n6431) );
  OAI222_X1 U5444 ( .A1(n5477), .A2(n7100), .B1(n6027), .B2(n6431), .C1(n6026), 
        .C2(n3862), .ZN(U2885) );
  INV_X1 U5445 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n7066) );
  NOR2_X1 U5446 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7066), .ZN(n7063) );
  NAND2_X1 U5447 ( .A1(n5814), .A2(n4826), .ZN(n4828) );
  AOI22_X1 U5448 ( .A1(n4828), .A2(n4827), .B1(n4254), .B2(n6733), .ZN(n4832)
         );
  NAND2_X1 U5449 ( .A1(n4830), .A2(n4829), .ZN(n4831) );
  NOR2_X1 U5450 ( .A1(n4832), .A2(n4831), .ZN(n4833) );
  NAND2_X1 U5451 ( .A1(n4834), .A2(n4833), .ZN(n4835) );
  INV_X1 U5452 ( .A(n5169), .ZN(n7026) );
  INV_X1 U5453 ( .A(FLUSH_REG_SCAN_IN), .ZN(n7037) );
  NOR2_X1 U5454 ( .A1(n6226), .A2(n7062), .ZN(n7058) );
  NAND2_X1 U5455 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n7058), .ZN(n7064) );
  OAI22_X1 U5456 ( .A1(n7026), .A2(n7077), .B1(n7037), .B2(n7064), .ZN(n7016)
         );
  NOR2_X1 U5457 ( .A1(n7063), .A2(n7016), .ZN(n5807) );
  NOR2_X1 U5458 ( .A1(n4654), .A2(n4693), .ZN(n4838) );
  AND2_X1 U5459 ( .A1(n4838), .A2(n5175), .ZN(n4839) );
  AND2_X1 U5460 ( .A1(n4840), .A2(n4839), .ZN(n5808) );
  INV_X1 U5461 ( .A(n4841), .ZN(n5809) );
  INV_X1 U5462 ( .A(n4842), .ZN(n4845) );
  INV_X1 U5463 ( .A(n4843), .ZN(n4844) );
  NAND2_X1 U5464 ( .A1(n4845), .A2(n4844), .ZN(n4848) );
  AOI22_X1 U5465 ( .A1(n5814), .A2(n3592), .B1(n5809), .B2(n4848), .ZN(n4846)
         );
  OAI21_X1 U5466 ( .B1(n5417), .B2(n5808), .A(n4846), .ZN(n7023) );
  INV_X1 U5467 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4847) );
  AOI22_X1 U5468 ( .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n6764), .B1(
        INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n4847), .ZN(n5766) );
  NOR2_X1 U5469 ( .A1(n7062), .A2(n6855), .ZN(n4849) );
  AOI222_X1 U5470 ( .A1(n7023), .A2(n7055), .B1(n5766), .B2(n4849), .C1(n4848), 
        .C2(n7069), .ZN(n4851) );
  NAND2_X1 U5471 ( .A1(n5807), .A2(n5137), .ZN(n4850) );
  OAI21_X1 U5472 ( .B1(n5807), .B2(n4851), .A(n4850), .ZN(U3460) );
  XNOR2_X1 U5473 ( .A(n4853), .B(n4852), .ZN(n6885) );
  INV_X1 U5474 ( .A(n6885), .ZN(n4859) );
  INV_X1 U5475 ( .A(DATAI_5_), .ZN(n6430) );
  INV_X1 U5476 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6552) );
  OAI222_X1 U5477 ( .A1(n7100), .A2(n4859), .B1(n6027), .B2(n6430), .C1(n6026), 
        .C2(n6552), .ZN(U2886) );
  NAND2_X1 U5478 ( .A1(n4855), .A2(n4854), .ZN(n4856) );
  AND2_X1 U5479 ( .A1(n4857), .A2(n4856), .ZN(n6879) );
  INV_X1 U5480 ( .A(n6879), .ZN(n6780) );
  INV_X1 U5481 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4858) );
  OAI222_X1 U5482 ( .A1(n6780), .A2(n6658), .B1(n6001), .B2(n4859), .C1(n4858), 
        .C2(n6663), .ZN(U2854) );
  OAI21_X1 U5483 ( .B1(n4861), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4860), 
        .ZN(n6852) );
  OAI21_X1 U5484 ( .B1(n6707), .B2(n4862), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4866) );
  INV_X1 U5485 ( .A(n5399), .ZN(n4864) );
  INV_X2 U5486 ( .A(n6121), .ZN(n6713) );
  NAND2_X1 U5487 ( .A1(n6771), .A2(REIP_REG_0__SCAN_IN), .ZN(n6863) );
  INV_X1 U5488 ( .A(n6863), .ZN(n4863) );
  AOI21_X1 U5489 ( .B1(n4864), .B2(n6713), .A(n4863), .ZN(n4865) );
  OAI211_X1 U5490 ( .C1(n6852), .C2(n6696), .A(n4866), .B(n4865), .ZN(U2986)
         );
  NAND2_X1 U5491 ( .A1(n4876), .A2(DATAI_14_), .ZN(n4879) );
  AOI22_X1 U5492 ( .A1(n4909), .A2(EAX_REG_14__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U5493 ( .A1(n4879), .A2(n4868), .ZN(U2953) );
  NAND2_X1 U5494 ( .A1(n4876), .A2(DATAI_8_), .ZN(n4893) );
  AOI22_X1 U5495 ( .A1(n4909), .A2(EAX_REG_8__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4869) );
  NAND2_X1 U5496 ( .A1(n4893), .A2(n4869), .ZN(U2947) );
  NAND2_X1 U5497 ( .A1(n4876), .A2(DATAI_6_), .ZN(n4897) );
  AOI22_X1 U5498 ( .A1(n4909), .A2(EAX_REG_6__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n4870) );
  NAND2_X1 U5499 ( .A1(n4897), .A2(n4870), .ZN(U2945) );
  NAND2_X1 U5500 ( .A1(n4876), .A2(DATAI_13_), .ZN(n4883) );
  AOI22_X1 U5501 ( .A1(n4909), .A2(EAX_REG_13__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n4871) );
  NAND2_X1 U5502 ( .A1(n4883), .A2(n4871), .ZN(U2952) );
  NAND2_X1 U5503 ( .A1(n4876), .A2(DATAI_4_), .ZN(n4881) );
  AOI22_X1 U5504 ( .A1(n4909), .A2(EAX_REG_4__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4872) );
  NAND2_X1 U5505 ( .A1(n4881), .A2(n4872), .ZN(U2943) );
  NAND2_X1 U5506 ( .A1(n4876), .A2(DATAI_3_), .ZN(n4903) );
  AOI22_X1 U5507 ( .A1(n4909), .A2(EAX_REG_3__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U5508 ( .A1(n4903), .A2(n4873), .ZN(U2942) );
  NAND2_X1 U5509 ( .A1(n4876), .A2(DATAI_2_), .ZN(n4905) );
  AOI22_X1 U5510 ( .A1(n4909), .A2(EAX_REG_2__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4874) );
  NAND2_X1 U5511 ( .A1(n4905), .A2(n4874), .ZN(U2941) );
  NAND2_X1 U5512 ( .A1(n4876), .A2(DATAI_1_), .ZN(n4907) );
  AOI22_X1 U5513 ( .A1(n4909), .A2(EAX_REG_1__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4875) );
  NAND2_X1 U5514 ( .A1(n4907), .A2(n4875), .ZN(U2940) );
  NAND2_X1 U5515 ( .A1(n4876), .A2(DATAI_0_), .ZN(n4901) );
  AOI22_X1 U5516 ( .A1(n4909), .A2(EAX_REG_0__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U5517 ( .A1(n4901), .A2(n4877), .ZN(U2939) );
  AOI22_X1 U5518 ( .A1(n4909), .A2(EAX_REG_30__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U5519 ( .A1(n4879), .A2(n4878), .ZN(U2938) );
  AOI22_X1 U5520 ( .A1(n4909), .A2(EAX_REG_20__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5521 ( .A1(n4881), .A2(n4880), .ZN(U2928) );
  AOI22_X1 U5522 ( .A1(n4909), .A2(EAX_REG_29__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n4882) );
  NAND2_X1 U5523 ( .A1(n4883), .A2(n4882), .ZN(U2937) );
  AOI22_X1 U5524 ( .A1(n4909), .A2(EAX_REG_28__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U5525 ( .A1(n4885), .A2(n4884), .ZN(U2936) );
  AOI22_X1 U5526 ( .A1(n4909), .A2(EAX_REG_27__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4886) );
  NAND2_X1 U5527 ( .A1(n4887), .A2(n4886), .ZN(U2935) );
  AOI22_X1 U5528 ( .A1(n4909), .A2(EAX_REG_26__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n4888) );
  NAND2_X1 U5529 ( .A1(n4889), .A2(n4888), .ZN(U2934) );
  AOI22_X1 U5530 ( .A1(n4909), .A2(EAX_REG_25__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4890) );
  NAND2_X1 U5531 ( .A1(n4891), .A2(n4890), .ZN(U2933) );
  AOI22_X1 U5532 ( .A1(n4909), .A2(EAX_REG_24__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4892) );
  NAND2_X1 U5533 ( .A1(n4893), .A2(n4892), .ZN(U2932) );
  AOI22_X1 U5534 ( .A1(n4909), .A2(EAX_REG_23__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4894) );
  NAND2_X1 U5535 ( .A1(n4895), .A2(n4894), .ZN(U2931) );
  AOI22_X1 U5536 ( .A1(n4909), .A2(EAX_REG_22__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4896) );
  NAND2_X1 U5537 ( .A1(n4897), .A2(n4896), .ZN(U2930) );
  AOI22_X1 U5538 ( .A1(n4909), .A2(EAX_REG_21__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4898) );
  NAND2_X1 U5539 ( .A1(n4899), .A2(n4898), .ZN(U2929) );
  AOI22_X1 U5540 ( .A1(n4909), .A2(EAX_REG_16__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4900) );
  NAND2_X1 U5541 ( .A1(n4901), .A2(n4900), .ZN(U2924) );
  AOI22_X1 U5542 ( .A1(n4909), .A2(EAX_REG_19__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4902) );
  NAND2_X1 U5543 ( .A1(n4903), .A2(n4902), .ZN(U2927) );
  AOI22_X1 U5544 ( .A1(n4909), .A2(EAX_REG_18__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4904) );
  NAND2_X1 U5545 ( .A1(n4905), .A2(n4904), .ZN(U2926) );
  AOI22_X1 U5546 ( .A1(n4909), .A2(EAX_REG_17__SCAN_IN), .B1(n4908), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4906) );
  NAND2_X1 U5547 ( .A1(n4907), .A2(n4906), .ZN(U2925) );
  INV_X1 U5548 ( .A(DATAI_15_), .ZN(n6460) );
  AOI22_X1 U5549 ( .A1(n4909), .A2(EAX_REG_15__SCAN_IN), .B1(n4908), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n4910) );
  OAI21_X1 U5550 ( .B1(n4911), .B2(n6460), .A(n4910), .ZN(U2954) );
  OR2_X1 U5551 ( .A1(n4924), .A2(n6226), .ZN(n5036) );
  NAND2_X1 U5552 ( .A1(n4974), .A2(n5036), .ZN(n6260) );
  NOR2_X1 U5553 ( .A1(n4913), .A2(n7132), .ZN(n6266) );
  INV_X1 U5554 ( .A(n6266), .ZN(n5064) );
  INV_X1 U5555 ( .A(n5344), .ZN(n4915) );
  NAND2_X1 U5556 ( .A1(n4915), .A2(n5417), .ZN(n5106) );
  NAND2_X1 U5557 ( .A1(n5106), .A2(n7146), .ZN(n5055) );
  NAND2_X1 U5558 ( .A1(n5185), .A2(n4386), .ZN(n4916) );
  NOR2_X2 U5559 ( .A1(n6230), .A2(n4916), .ZN(n6254) );
  INV_X1 U5560 ( .A(n6254), .ZN(n4919) );
  NOR2_X1 U5561 ( .A1(n5210), .A2(n4386), .ZN(n4918) );
  AND2_X1 U5562 ( .A1(n4918), .A2(n5415), .ZN(n5054) );
  NAND2_X1 U5563 ( .A1(n5054), .A2(n4403), .ZN(n7124) );
  AOI21_X1 U5564 ( .B1(n4919), .B2(n7124), .A(n7080), .ZN(n4920) );
  AOI21_X1 U5565 ( .B1(n5064), .B2(n5055), .A(n4920), .ZN(n4922) );
  NAND3_X1 U5566 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5523), .ZN(n6225) );
  NOR2_X1 U5567 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6225), .ZN(n5430)
         );
  INV_X1 U5568 ( .A(n5521), .ZN(n5060) );
  NAND2_X1 U5569 ( .A1(n5063), .A2(n5060), .ZN(n4981) );
  NAND2_X1 U5570 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4981), .ZN(n4975) );
  OAI21_X1 U5571 ( .B1(n5430), .B2(n7066), .A(n4975), .ZN(n4921) );
  AND2_X1 U5572 ( .A1(n6713), .A2(DATAI_25_), .ZN(n7156) );
  INV_X1 U5573 ( .A(n7156), .ZN(n5227) );
  NOR2_X2 U5574 ( .A1(n5252), .A2(n3604), .ZN(n7155) );
  NAND2_X1 U5575 ( .A1(n7155), .A2(n5430), .ZN(n4928) );
  NAND2_X1 U5576 ( .A1(n6713), .A2(DATAI_17_), .ZN(n6281) );
  INV_X1 U5577 ( .A(n6281), .ZN(n7154) );
  INV_X1 U5578 ( .A(DATAI_1_), .ZN(n5029) );
  NOR2_X1 U5579 ( .A1(n5029), .A2(n5253), .ZN(n6279) );
  INV_X1 U5580 ( .A(n5106), .ZN(n6221) );
  NAND2_X1 U5581 ( .A1(n5031), .A2(n6221), .ZN(n4926) );
  NAND2_X1 U5582 ( .A1(n4924), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6271) );
  OR2_X1 U5583 ( .A1(n4981), .A2(n6271), .ZN(n4925) );
  NAND2_X1 U5584 ( .A1(n4926), .A2(n4925), .ZN(n5431) );
  AOI22_X1 U5585 ( .A1(n6254), .A2(n7154), .B1(n6279), .B2(n5431), .ZN(n4927)
         );
  OAI211_X1 U5586 ( .C1(n7124), .C2(n5227), .A(n4928), .B(n4927), .ZN(n4929)
         );
  AOI21_X1 U5587 ( .B1(n5435), .B2(INSTQUEUE_REG_12__1__SCAN_IN), .A(n4929), 
        .ZN(n4930) );
  INV_X1 U5588 ( .A(n4930), .ZN(U3117) );
  AND2_X1 U5589 ( .A1(n6713), .A2(DATAI_31_), .ZN(n7208) );
  INV_X1 U5590 ( .A(n7208), .ZN(n5235) );
  NOR2_X2 U5591 ( .A1(n5252), .A2(n6006), .ZN(n7210) );
  NAND2_X1 U5592 ( .A1(n7210), .A2(n5430), .ZN(n4932) );
  NAND2_X1 U5593 ( .A1(n6713), .A2(DATAI_23_), .ZN(n6320) );
  INV_X1 U5594 ( .A(n6320), .ZN(n7212) );
  INV_X1 U5595 ( .A(DATAI_7_), .ZN(n6476) );
  NOR2_X1 U5596 ( .A1(n6476), .A2(n5253), .ZN(n6316) );
  AOI22_X1 U5597 ( .A1(n6254), .A2(n7212), .B1(n6316), .B2(n5431), .ZN(n4931)
         );
  OAI211_X1 U5598 ( .C1(n7124), .C2(n5235), .A(n4932), .B(n4931), .ZN(n4933)
         );
  AOI21_X1 U5599 ( .B1(n5435), .B2(INSTQUEUE_REG_12__7__SCAN_IN), .A(n4933), 
        .ZN(n4934) );
  INV_X1 U5600 ( .A(n4934), .ZN(U3123) );
  AND2_X1 U5601 ( .A1(n6713), .A2(DATAI_29_), .ZN(n7188) );
  INV_X1 U5602 ( .A(n7188), .ZN(n5239) );
  NOR2_X2 U5603 ( .A1(n5252), .A2(n5734), .ZN(n7187) );
  NAND2_X1 U5604 ( .A1(n7187), .A2(n5430), .ZN(n4936) );
  NAND2_X1 U5605 ( .A1(n6713), .A2(DATAI_21_), .ZN(n6305) );
  INV_X1 U5606 ( .A(n6305), .ZN(n7186) );
  NOR2_X1 U5607 ( .A1(n6430), .A2(n5253), .ZN(n6303) );
  AOI22_X1 U5608 ( .A1(n6254), .A2(n7186), .B1(n6303), .B2(n5431), .ZN(n4935)
         );
  OAI211_X1 U5609 ( .C1(n7124), .C2(n5239), .A(n4936), .B(n4935), .ZN(n4937)
         );
  AOI21_X1 U5610 ( .B1(n5435), .B2(INSTQUEUE_REG_12__5__SCAN_IN), .A(n4937), 
        .ZN(n4938) );
  INV_X1 U5611 ( .A(n4938), .ZN(U3121) );
  AND2_X1 U5612 ( .A1(n6713), .A2(DATAI_24_), .ZN(n7138) );
  INV_X1 U5613 ( .A(n7138), .ZN(n5243) );
  NOR2_X2 U5614 ( .A1(n5252), .A2(n4939), .ZN(n7139) );
  NAND2_X1 U5615 ( .A1(n7139), .A2(n5430), .ZN(n4941) );
  NAND2_X1 U5616 ( .A1(n6713), .A2(DATAI_16_), .ZN(n6275) );
  INV_X1 U5617 ( .A(n6275), .ZN(n7148) );
  NOR2_X1 U5618 ( .A1(n6489), .A2(n5253), .ZN(n6273) );
  AOI22_X1 U5619 ( .A1(n6254), .A2(n7148), .B1(n6273), .B2(n5431), .ZN(n4940)
         );
  OAI211_X1 U5620 ( .C1(n7124), .C2(n5243), .A(n4941), .B(n4940), .ZN(n4942)
         );
  AOI21_X1 U5621 ( .B1(n5435), .B2(INSTQUEUE_REG_12__0__SCAN_IN), .A(n4942), 
        .ZN(n4943) );
  INV_X1 U5622 ( .A(n4943), .ZN(U3116) );
  AND2_X1 U5623 ( .A1(n6713), .A2(DATAI_27_), .ZN(n7172) );
  INV_X1 U5624 ( .A(n7172), .ZN(n5231) );
  NOR2_X2 U5625 ( .A1(n5252), .A2(n4944), .ZN(n7171) );
  NAND2_X1 U5626 ( .A1(n7171), .A2(n5430), .ZN(n4946) );
  NAND2_X1 U5627 ( .A1(n6713), .A2(DATAI_19_), .ZN(n6293) );
  INV_X1 U5628 ( .A(n6293), .ZN(n7170) );
  NOR2_X1 U5629 ( .A1(n6484), .A2(n5253), .ZN(n6291) );
  AOI22_X1 U5630 ( .A1(n6254), .A2(n7170), .B1(n6291), .B2(n5431), .ZN(n4945)
         );
  OAI211_X1 U5631 ( .C1(n7124), .C2(n5231), .A(n4946), .B(n4945), .ZN(n4947)
         );
  AOI21_X1 U5632 ( .B1(n5435), .B2(INSTQUEUE_REG_12__3__SCAN_IN), .A(n4947), 
        .ZN(n4948) );
  INV_X1 U5633 ( .A(n4948), .ZN(U3119) );
  INV_X1 U5634 ( .A(n5800), .ZN(n5811) );
  NOR2_X1 U5635 ( .A1(n5344), .A2(n5417), .ZN(n6269) );
  NOR2_X1 U5636 ( .A1(n4949), .A2(n4200), .ZN(n5258) );
  AOI21_X1 U5637 ( .B1(n7122), .B2(n6269), .A(n5258), .ZN(n4953) );
  AND3_X1 U5638 ( .A1(n5210), .A2(n5185), .A3(n5415), .ZN(n4952) );
  NOR2_X1 U5639 ( .A1(n7132), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5212) );
  INV_X1 U5640 ( .A(n5212), .ZN(n5519) );
  OAI21_X1 U5641 ( .B1(n4952), .B2(n6121), .A(n5519), .ZN(n4950) );
  NAND3_X1 U5642 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6259) );
  AOI22_X1 U5643 ( .A1(n4953), .A2(n4950), .B1(n7132), .B2(n6259), .ZN(n4951)
         );
  INV_X1 U5644 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4957) );
  NAND2_X1 U5645 ( .A1(n4952), .A2(n4386), .ZN(n6319) );
  OAI22_X1 U5646 ( .A1(n4953), .A2(n7132), .B1(n6259), .B2(n6226), .ZN(n5254)
         );
  AOI22_X1 U5647 ( .A1(n5255), .A2(n7170), .B1(n6291), .B2(n5254), .ZN(n4954)
         );
  OAI21_X1 U5648 ( .B1(n5231), .B2(n6319), .A(n4954), .ZN(n4955) );
  AOI21_X1 U5649 ( .B1(n7171), .B2(n5258), .A(n4955), .ZN(n4956) );
  OAI21_X1 U5650 ( .B1(n5261), .B2(n4957), .A(n4956), .ZN(U3143) );
  INV_X1 U5651 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U5652 ( .A1(n5255), .A2(n7148), .B1(n6273), .B2(n5254), .ZN(n4958)
         );
  OAI21_X1 U5653 ( .B1(n5243), .B2(n6319), .A(n4958), .ZN(n4959) );
  AOI21_X1 U5654 ( .B1(n7139), .B2(n5258), .A(n4959), .ZN(n4960) );
  OAI21_X1 U5655 ( .B1(n5261), .B2(n4961), .A(n4960), .ZN(U3140) );
  INV_X1 U5656 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U5657 ( .A1(n5255), .A2(n7186), .B1(n6303), .B2(n5254), .ZN(n4962)
         );
  OAI21_X1 U5658 ( .B1(n5239), .B2(n6319), .A(n4962), .ZN(n4963) );
  AOI21_X1 U5659 ( .B1(n7187), .B2(n5258), .A(n4963), .ZN(n4964) );
  OAI21_X1 U5660 ( .B1(n5261), .B2(n4965), .A(n4964), .ZN(U3145) );
  INV_X1 U5661 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4969) );
  AOI22_X1 U5662 ( .A1(n5255), .A2(n7212), .B1(n6316), .B2(n5254), .ZN(n4966)
         );
  OAI21_X1 U5663 ( .B1(n5235), .B2(n6319), .A(n4966), .ZN(n4967) );
  AOI21_X1 U5664 ( .B1(n7210), .B2(n5258), .A(n4967), .ZN(n4968) );
  OAI21_X1 U5665 ( .B1(n5261), .B2(n4969), .A(n4968), .ZN(U3147) );
  INV_X1 U5666 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U5667 ( .A1(n5255), .A2(n7154), .B1(n6279), .B2(n5254), .ZN(n4970)
         );
  OAI21_X1 U5668 ( .B1(n5227), .B2(n6319), .A(n4970), .ZN(n4971) );
  AOI21_X1 U5669 ( .B1(n7155), .B2(n5258), .A(n4971), .ZN(n4972) );
  OAI21_X1 U5670 ( .B1(n5261), .B2(n4973), .A(n4972), .ZN(U3141) );
  NOR2_X1 U5671 ( .A1(n5210), .A2(n5415), .ZN(n5030) );
  NAND2_X1 U5672 ( .A1(n5030), .A2(n4403), .ZN(n5087) );
  NAND3_X1 U5673 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5181), .A3(n5523), .ZN(n5084) );
  NOR2_X1 U5674 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5084), .ZN(n5336)
         );
  NAND2_X1 U5675 ( .A1(n4974), .A2(n6271), .ZN(n5527) );
  OAI211_X1 U5676 ( .C1(n5336), .C2(n7066), .A(n5217), .B(n4975), .ZN(n4980)
         );
  NAND2_X1 U5677 ( .A1(n5344), .A2(n5417), .ZN(n5092) );
  NAND2_X1 U5678 ( .A1(n5092), .A2(n7146), .ZN(n5033) );
  NAND2_X1 U5679 ( .A1(n5210), .A2(n6229), .ZN(n5184) );
  INV_X1 U5680 ( .A(n5184), .ZN(n4977) );
  AND2_X1 U5681 ( .A1(n5415), .A2(n5209), .ZN(n4976) );
  NAND2_X1 U5682 ( .A1(n4977), .A2(n4976), .ZN(n7147) );
  AOI21_X1 U5683 ( .B1(n5339), .B2(n7147), .A(n7080), .ZN(n4978) );
  AOI21_X1 U5684 ( .B1(n5064), .B2(n5033), .A(n4978), .ZN(n4979) );
  NAND2_X1 U5685 ( .A1(n5333), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4987) );
  INV_X1 U5686 ( .A(n5092), .ZN(n5080) );
  NAND2_X1 U5687 ( .A1(n5031), .A2(n5080), .ZN(n4984) );
  INV_X1 U5688 ( .A(n5036), .ZN(n5522) );
  INV_X1 U5689 ( .A(n4981), .ZN(n4982) );
  NAND2_X1 U5690 ( .A1(n5522), .A2(n4982), .ZN(n4983) );
  OAI22_X1 U5691 ( .A1(n7147), .A2(n5239), .B1(n5334), .B2(n7191), .ZN(n4985)
         );
  AOI21_X1 U5692 ( .B1(n7187), .B2(n5336), .A(n4985), .ZN(n4986) );
  OAI211_X1 U5693 ( .C1(n5339), .C2(n6305), .A(n4987), .B(n4986), .ZN(U3089)
         );
  NAND2_X1 U5694 ( .A1(n5333), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4990) );
  OAI22_X1 U5695 ( .A1(n7147), .A2(n5231), .B1(n5334), .B2(n7175), .ZN(n4988)
         );
  AOI21_X1 U5696 ( .B1(n7171), .B2(n5336), .A(n4988), .ZN(n4989) );
  OAI211_X1 U5697 ( .C1(n5339), .C2(n6293), .A(n4990), .B(n4989), .ZN(U3087)
         );
  NAND2_X1 U5698 ( .A1(n5333), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4993) );
  OAI22_X1 U5699 ( .A1(n7147), .A2(n5235), .B1(n5334), .B2(n7216), .ZN(n4991)
         );
  AOI21_X1 U5700 ( .B1(n7210), .B2(n5336), .A(n4991), .ZN(n4992) );
  OAI211_X1 U5701 ( .C1(n5339), .C2(n6320), .A(n4993), .B(n4992), .ZN(U3091)
         );
  NAND2_X1 U5702 ( .A1(n5333), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4996) );
  OAI22_X1 U5703 ( .A1(n7147), .A2(n5227), .B1(n5334), .B2(n7159), .ZN(n4994)
         );
  AOI21_X1 U5704 ( .B1(n7155), .B2(n5336), .A(n4994), .ZN(n4995) );
  OAI211_X1 U5705 ( .C1(n5339), .C2(n6281), .A(n4996), .B(n4995), .ZN(U3085)
         );
  INV_X1 U5706 ( .A(n7139), .ZN(n6233) );
  NOR3_X1 U5707 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5181), .A3(n5523), 
        .ZN(n7145) );
  NAND2_X1 U5708 ( .A1(n7020), .A2(n7145), .ZN(n5414) );
  NAND2_X1 U5709 ( .A1(n5521), .A2(n4200), .ZN(n5222) );
  NAND2_X1 U5710 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n5222), .ZN(n5218) );
  INV_X1 U5711 ( .A(n5218), .ZN(n4997) );
  AOI211_X1 U5712 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5414), .A(n4997), .B(
        n6260), .ZN(n5001) );
  NOR2_X1 U5713 ( .A1(n6269), .A2(n7132), .ZN(n6265) );
  NAND2_X1 U5714 ( .A1(n5104), .A2(n6229), .ZN(n5053) );
  NOR2_X2 U5715 ( .A1(n5053), .A2(n4386), .ZN(n5411) );
  NAND2_X1 U5716 ( .A1(n5415), .A2(n4386), .ZN(n4998) );
  OAI21_X1 U5717 ( .B1(n5411), .B2(n7207), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4999) );
  OAI21_X1 U5718 ( .B1(n6265), .B2(n5031), .A(n4999), .ZN(n5000) );
  NAND2_X1 U5719 ( .A1(n5001), .A2(n5000), .ZN(n5407) );
  NAND2_X1 U5720 ( .A1(n5407), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n5005) );
  INV_X1 U5721 ( .A(n7207), .ZN(n5409) );
  NOR2_X1 U5722 ( .A1(n6271), .A2(n5222), .ZN(n5002) );
  AOI21_X1 U5723 ( .B1(n6266), .B2(n6269), .A(n5002), .ZN(n5408) );
  OAI22_X1 U5724 ( .A1(n5409), .A2(n6275), .B1(n5408), .B2(n7151), .ZN(n5003)
         );
  AOI21_X1 U5725 ( .B1(n5411), .B2(n7138), .A(n5003), .ZN(n5004) );
  OAI211_X1 U5726 ( .C1(n6233), .C2(n5414), .A(n5005), .B(n5004), .ZN(U3068)
         );
  INV_X1 U5727 ( .A(n7210), .ZN(n6258) );
  NAND2_X1 U5728 ( .A1(n5407), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5008) );
  OAI22_X1 U5729 ( .A1(n5409), .A2(n6320), .B1(n5408), .B2(n7216), .ZN(n5006)
         );
  AOI21_X1 U5730 ( .B1(n7208), .B2(n5411), .A(n5006), .ZN(n5007) );
  OAI211_X1 U5731 ( .C1(n5414), .C2(n6258), .A(n5008), .B(n5007), .ZN(U3075)
         );
  INV_X1 U5732 ( .A(n7187), .ZN(n6248) );
  NAND2_X1 U5733 ( .A1(n5407), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U5734 ( .A1(n5409), .A2(n6305), .B1(n5408), .B2(n7191), .ZN(n5009)
         );
  AOI21_X1 U5735 ( .B1(n7188), .B2(n5411), .A(n5009), .ZN(n5010) );
  OAI211_X1 U5736 ( .C1(n5414), .C2(n6248), .A(n5011), .B(n5010), .ZN(U3073)
         );
  INV_X1 U5737 ( .A(n7171), .ZN(n6242) );
  NAND2_X1 U5738 ( .A1(n5407), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5014) );
  OAI22_X1 U5739 ( .A1(n5409), .A2(n6293), .B1(n5408), .B2(n7175), .ZN(n5012)
         );
  AOI21_X1 U5740 ( .B1(n7172), .B2(n5411), .A(n5012), .ZN(n5013) );
  OAI211_X1 U5741 ( .C1(n5414), .C2(n6242), .A(n5014), .B(n5013), .ZN(U3071)
         );
  INV_X1 U5742 ( .A(n7155), .ZN(n6236) );
  NAND2_X1 U5743 ( .A1(n5407), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n5017) );
  OAI22_X1 U5744 ( .A1(n5409), .A2(n6281), .B1(n5408), .B2(n7159), .ZN(n5015)
         );
  AOI21_X1 U5745 ( .B1(n7156), .B2(n5411), .A(n5015), .ZN(n5016) );
  OAI211_X1 U5746 ( .C1(n5414), .C2(n6236), .A(n5017), .B(n5016), .ZN(U3069)
         );
  NAND2_X1 U5747 ( .A1(n5333), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n5020) );
  OAI22_X1 U5748 ( .A1(n7147), .A2(n5243), .B1(n5334), .B2(n7151), .ZN(n5018)
         );
  AOI21_X1 U5749 ( .B1(n7139), .B2(n5336), .A(n5018), .ZN(n5019) );
  OAI211_X1 U5750 ( .C1(n5339), .C2(n6275), .A(n5020), .B(n5019), .ZN(U3084)
         );
  OAI21_X1 U5751 ( .B1(n5023), .B2(n5022), .A(n5191), .ZN(n6890) );
  OR2_X1 U5752 ( .A1(n5025), .A2(n5024), .ZN(n5026) );
  AND2_X1 U5753 ( .A1(n5194), .A2(n5026), .ZN(n6892) );
  AOI22_X1 U5754 ( .A1(n6649), .A2(n6892), .B1(EBX_REG_7__SCAN_IN), .B2(n5970), 
        .ZN(n5027) );
  OAI21_X1 U5755 ( .B1(n6890), .B2(n6005), .A(n5027), .ZN(U2852) );
  INV_X1 U5756 ( .A(DATAI_2_), .ZN(n6483) );
  INV_X1 U5757 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6546) );
  OAI222_X1 U5758 ( .A1(n5028), .A2(n7100), .B1(n6027), .B2(n6483), .C1(n6026), 
        .C2(n6546), .ZN(U2889) );
  INV_X1 U5759 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6544) );
  OAI222_X1 U5760 ( .A1(n5576), .A2(n7100), .B1(n6027), .B2(n5029), .C1(n6026), 
        .C2(n6544), .ZN(U2890) );
  INV_X1 U5761 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6555) );
  OAI222_X1 U5762 ( .A1(n6890), .A2(n7100), .B1(n6027), .B2(n6476), .C1(n6026), 
        .C2(n6555), .ZN(U2884) );
  INV_X1 U5763 ( .A(n5031), .ZN(n6272) );
  AOI21_X1 U5764 ( .B1(n5326), .B2(n5321), .A(n7080), .ZN(n5032) );
  AOI21_X1 U5765 ( .B1(n6272), .B2(n5033), .A(n5032), .ZN(n5035) );
  NOR2_X1 U5766 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5216) );
  INV_X1 U5767 ( .A(n5216), .ZN(n5266) );
  OAI21_X1 U5768 ( .B1(n5521), .B2(n5063), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n5056) );
  OAI211_X1 U5769 ( .C1(n5323), .C2(n7066), .A(n5217), .B(n5056), .ZN(n5034)
         );
  NAND2_X1 U5770 ( .A1(n5319), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5040) );
  NOR3_X1 U5771 ( .A1(n5036), .A2(n5521), .A3(n5063), .ZN(n5037) );
  AOI21_X1 U5772 ( .B1(n6266), .B2(n5080), .A(n5037), .ZN(n5320) );
  OAI22_X1 U5773 ( .A1(n5321), .A2(n5235), .B1(n5320), .B2(n7216), .ZN(n5038)
         );
  AOI21_X1 U5774 ( .B1(n7210), .B2(n5323), .A(n5038), .ZN(n5039) );
  OAI211_X1 U5775 ( .C1(n6320), .C2(n5326), .A(n5040), .B(n5039), .ZN(U3027)
         );
  NAND2_X1 U5776 ( .A1(n5319), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5043) );
  OAI22_X1 U5777 ( .A1(n5321), .A2(n5227), .B1(n5320), .B2(n7159), .ZN(n5041)
         );
  AOI21_X1 U5778 ( .B1(n7155), .B2(n5323), .A(n5041), .ZN(n5042) );
  OAI211_X1 U5779 ( .C1(n6281), .C2(n5326), .A(n5043), .B(n5042), .ZN(U3021)
         );
  NAND2_X1 U5780 ( .A1(n5319), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5046) );
  OAI22_X1 U5781 ( .A1(n5321), .A2(n5243), .B1(n5320), .B2(n7151), .ZN(n5044)
         );
  AOI21_X1 U5782 ( .B1(n7139), .B2(n5323), .A(n5044), .ZN(n5045) );
  OAI211_X1 U5783 ( .C1(n5326), .C2(n6275), .A(n5046), .B(n5045), .ZN(U3020)
         );
  NAND2_X1 U5784 ( .A1(n5319), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U5785 ( .A1(n5321), .A2(n5231), .B1(n5320), .B2(n7175), .ZN(n5047)
         );
  AOI21_X1 U5786 ( .B1(n7171), .B2(n5323), .A(n5047), .ZN(n5048) );
  OAI211_X1 U5787 ( .C1(n6293), .C2(n5326), .A(n5049), .B(n5048), .ZN(U3023)
         );
  NAND2_X1 U5788 ( .A1(n5319), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5052) );
  OAI22_X1 U5789 ( .A1(n5321), .A2(n5239), .B1(n5320), .B2(n7191), .ZN(n5050)
         );
  AOI21_X1 U5790 ( .B1(n7187), .B2(n5323), .A(n5050), .ZN(n5051) );
  OAI211_X1 U5791 ( .C1(n6305), .C2(n5326), .A(n5052), .B(n5051), .ZN(U3025)
         );
  NOR2_X2 U5792 ( .A1(n5053), .A2(n5209), .ZN(n5390) );
  OAI21_X1 U5793 ( .B1(n5390), .B2(n5378), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5059) );
  NAND2_X1 U5794 ( .A1(n6272), .A2(n5055), .ZN(n5058) );
  NAND3_X1 U5795 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n4200), .A3(n5523), .ZN(n5110) );
  NOR2_X1 U5796 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5110), .ZN(n5379)
         );
  OAI21_X1 U5797 ( .B1(n5379), .B2(n7066), .A(n5056), .ZN(n5057) );
  AOI211_X2 U5798 ( .C1(n5059), .C2(n5058), .A(n5057), .B(n6260), .ZN(n5383)
         );
  INV_X1 U5799 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5067) );
  INV_X1 U5800 ( .A(n6271), .ZN(n5061) );
  NAND2_X1 U5801 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  OAI22_X1 U5802 ( .A1(n5064), .A2(n5106), .B1(n5063), .B2(n5062), .ZN(n5377)
         );
  AOI22_X1 U5803 ( .A1(n5390), .A2(n7154), .B1(n6279), .B2(n5377), .ZN(n5066)
         );
  AOI22_X1 U5804 ( .A1(n7155), .A2(n5379), .B1(n7156), .B2(n5378), .ZN(n5065)
         );
  OAI211_X1 U5805 ( .C1(n5383), .C2(n5067), .A(n5066), .B(n5065), .ZN(U3053)
         );
  INV_X1 U5806 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5070) );
  AOI22_X1 U5807 ( .A1(n5390), .A2(n7186), .B1(n6303), .B2(n5377), .ZN(n5069)
         );
  AOI22_X1 U5808 ( .A1(n7187), .A2(n5379), .B1(n7188), .B2(n5378), .ZN(n5068)
         );
  OAI211_X1 U5809 ( .C1(n5383), .C2(n5070), .A(n5069), .B(n5068), .ZN(U3057)
         );
  INV_X1 U5810 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5073) );
  AOI22_X1 U5811 ( .A1(n5390), .A2(n7148), .B1(n6273), .B2(n5377), .ZN(n5072)
         );
  AOI22_X1 U5812 ( .A1(n7139), .A2(n5379), .B1(n7138), .B2(n5378), .ZN(n5071)
         );
  OAI211_X1 U5813 ( .C1(n5383), .C2(n5073), .A(n5072), .B(n5071), .ZN(U3052)
         );
  INV_X1 U5814 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5076) );
  AOI22_X1 U5815 ( .A1(n5390), .A2(n7212), .B1(n6316), .B2(n5377), .ZN(n5075)
         );
  AOI22_X1 U5816 ( .A1(n7210), .A2(n5379), .B1(n7208), .B2(n5378), .ZN(n5074)
         );
  OAI211_X1 U5817 ( .C1(n5383), .C2(n5076), .A(n5075), .B(n5074), .ZN(U3059)
         );
  INV_X1 U5818 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5079) );
  AOI22_X1 U5819 ( .A1(n5390), .A2(n7170), .B1(n6291), .B2(n5377), .ZN(n5078)
         );
  AOI22_X1 U5820 ( .A1(n7171), .A2(n5379), .B1(n7172), .B2(n5378), .ZN(n5077)
         );
  OAI211_X1 U5821 ( .C1(n5383), .C2(n5079), .A(n5078), .B(n5077), .ZN(U3055)
         );
  INV_X1 U5822 ( .A(n5084), .ZN(n5083) );
  OAI21_X1 U5823 ( .B1(n5087), .B2(n7080), .A(n7146), .ZN(n5086) );
  INV_X1 U5824 ( .A(n5086), .ZN(n5081) );
  NOR2_X1 U5825 ( .A1(n7020), .A2(n5084), .ZN(n5310) );
  AOI21_X1 U5826 ( .B1(n7122), .B2(n5080), .A(n5310), .ZN(n5085) );
  NAND2_X1 U5827 ( .A1(n5081), .A2(n5085), .ZN(n5082) );
  OAI211_X1 U5828 ( .C1(n7146), .C2(n5083), .A(n7143), .B(n5082), .ZN(n5309)
         );
  OAI22_X1 U5829 ( .A1(n5086), .A2(n5085), .B1(n6226), .B2(n5084), .ZN(n5308)
         );
  AOI22_X1 U5830 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n5309), .B1(n6291), 
        .B2(n5308), .ZN(n5089) );
  AOI22_X1 U5831 ( .A1(n7171), .A2(n5310), .B1(n7170), .B2(n3425), .ZN(n5088)
         );
  OAI211_X1 U5832 ( .C1(n5231), .C2(n5339), .A(n5089), .B(n5088), .ZN(U3095)
         );
  INV_X1 U5833 ( .A(n5090), .ZN(n5091) );
  OAI21_X1 U5834 ( .B1(n5091), .B2(n7080), .A(n7146), .ZN(n5098) );
  NAND2_X1 U5835 ( .A1(n5214), .A2(n5811), .ZN(n7135) );
  OR2_X1 U5836 ( .A1(n7135), .A2(n5092), .ZN(n5094) );
  NAND2_X1 U5837 ( .A1(n5216), .A2(n5523), .ZN(n5097) );
  NOR2_X1 U5838 ( .A1(n7020), .A2(n5097), .ZN(n5305) );
  INV_X1 U5839 ( .A(n5305), .ZN(n5093) );
  AND2_X1 U5840 ( .A1(n5094), .A2(n5093), .ZN(n5099) );
  INV_X1 U5841 ( .A(n5099), .ZN(n5096) );
  NAND2_X1 U5842 ( .A1(n7132), .A2(n5097), .ZN(n5095) );
  OAI211_X1 U5843 ( .C1(n5098), .C2(n5096), .A(n7143), .B(n5095), .ZN(n5303)
         );
  OAI22_X1 U5844 ( .A1(n5099), .A2(n5098), .B1(n6226), .B2(n5097), .ZN(n5302)
         );
  AOI22_X1 U5845 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5303), .B1(n6273), 
        .B2(n5302), .ZN(n5101) );
  AOI22_X1 U5846 ( .A1(n7139), .A2(n5305), .B1(n7138), .B2(n5304), .ZN(n5100)
         );
  OAI211_X1 U5847 ( .C1(n5475), .C2(n6275), .A(n5101), .B(n5100), .ZN(U3028)
         );
  AOI22_X1 U5848 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5303), .B1(n6279), 
        .B2(n5302), .ZN(n5103) );
  AOI22_X1 U5849 ( .A1(n7155), .A2(n5305), .B1(n5304), .B2(n7156), .ZN(n5102)
         );
  OAI211_X1 U5850 ( .C1(n5475), .C2(n6281), .A(n5103), .B(n5102), .ZN(U3029)
         );
  OR2_X1 U5851 ( .A1(n7020), .A2(n5110), .ZN(n5393) );
  NAND3_X1 U5852 ( .A1(n5104), .A2(n6229), .A3(STATEBS16_REG_SCAN_IN), .ZN(
        n5105) );
  NAND2_X1 U5853 ( .A1(n5105), .A2(n7146), .ZN(n5111) );
  OR2_X1 U5854 ( .A1(n7135), .A2(n5106), .ZN(n5107) );
  AND2_X1 U5855 ( .A1(n5107), .A2(n5393), .ZN(n5112) );
  INV_X1 U5856 ( .A(n5112), .ZN(n5109) );
  NAND2_X1 U5857 ( .A1(n7132), .A2(n5110), .ZN(n5108) );
  OAI211_X1 U5858 ( .C1(n5111), .C2(n5109), .A(n7143), .B(n5108), .ZN(n5389)
         );
  OAI22_X1 U5859 ( .A1(n5112), .A2(n5111), .B1(n6226), .B2(n5110), .ZN(n5388)
         );
  AOI22_X1 U5860 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n5389), .B1(n6316), 
        .B2(n5388), .ZN(n5114) );
  AOI22_X1 U5861 ( .A1(n7212), .A2(n5411), .B1(n5390), .B2(n7208), .ZN(n5113)
         );
  OAI211_X1 U5862 ( .C1(n6258), .C2(n5393), .A(n5114), .B(n5113), .ZN(U3067)
         );
  AOI22_X1 U5863 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n5389), .B1(n6273), 
        .B2(n5388), .ZN(n5116) );
  AOI22_X1 U5864 ( .A1(n7148), .A2(n5411), .B1(n5390), .B2(n7138), .ZN(n5115)
         );
  OAI211_X1 U5865 ( .C1(n6233), .C2(n5393), .A(n5116), .B(n5115), .ZN(U3060)
         );
  AOI22_X1 U5866 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n5309), .B1(n6303), 
        .B2(n5308), .ZN(n5118) );
  AOI22_X1 U5867 ( .A1(n7187), .A2(n5310), .B1(n7186), .B2(n3425), .ZN(n5117)
         );
  OAI211_X1 U5868 ( .C1(n5239), .C2(n5339), .A(n5118), .B(n5117), .ZN(U3097)
         );
  AOI22_X1 U5869 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n5309), .B1(n6273), 
        .B2(n5308), .ZN(n5120) );
  AOI22_X1 U5870 ( .A1(n7139), .A2(n5310), .B1(n7148), .B2(n3425), .ZN(n5119)
         );
  OAI211_X1 U5871 ( .C1(n5243), .C2(n5339), .A(n5120), .B(n5119), .ZN(U3092)
         );
  AOI22_X1 U5872 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n5389), .B1(n6291), 
        .B2(n5388), .ZN(n5122) );
  AOI22_X1 U5873 ( .A1(n7170), .A2(n5411), .B1(n5390), .B2(n7172), .ZN(n5121)
         );
  OAI211_X1 U5874 ( .C1(n6242), .C2(n5393), .A(n5122), .B(n5121), .ZN(U3063)
         );
  AOI22_X1 U5875 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n5389), .B1(n6303), 
        .B2(n5388), .ZN(n5124) );
  AOI22_X1 U5876 ( .A1(n7186), .A2(n5411), .B1(n5390), .B2(n7188), .ZN(n5123)
         );
  OAI211_X1 U5877 ( .C1(n6248), .C2(n5393), .A(n5124), .B(n5123), .ZN(U3065)
         );
  AOI22_X1 U5878 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n5309), .B1(n6316), 
        .B2(n5308), .ZN(n5126) );
  AOI22_X1 U5879 ( .A1(n7210), .A2(n5310), .B1(n7212), .B2(n3425), .ZN(n5125)
         );
  OAI211_X1 U5880 ( .C1(n5235), .C2(n5339), .A(n5126), .B(n5125), .ZN(U3099)
         );
  AOI22_X1 U5881 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5303), .B1(n6291), 
        .B2(n5302), .ZN(n5128) );
  AOI22_X1 U5882 ( .A1(n7171), .A2(n5305), .B1(n5304), .B2(n7172), .ZN(n5127)
         );
  OAI211_X1 U5883 ( .C1(n5475), .C2(n6293), .A(n5128), .B(n5127), .ZN(U3031)
         );
  AOI22_X1 U5884 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5303), .B1(n6303), 
        .B2(n5302), .ZN(n5130) );
  AOI22_X1 U5885 ( .A1(n7187), .A2(n5305), .B1(n5304), .B2(n7188), .ZN(n5129)
         );
  OAI211_X1 U5886 ( .C1(n5475), .C2(n6305), .A(n5130), .B(n5129), .ZN(U3033)
         );
  AOI22_X1 U5887 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n5389), .B1(n6279), 
        .B2(n5388), .ZN(n5132) );
  AOI22_X1 U5888 ( .A1(n7154), .A2(n5411), .B1(n5390), .B2(n7156), .ZN(n5131)
         );
  OAI211_X1 U5889 ( .C1(n6236), .C2(n5393), .A(n5132), .B(n5131), .ZN(U3061)
         );
  AOI22_X1 U5890 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5303), .B1(n6316), 
        .B2(n5302), .ZN(n5134) );
  AOI22_X1 U5891 ( .A1(n7210), .A2(n5305), .B1(n5304), .B2(n7208), .ZN(n5133)
         );
  OAI211_X1 U5892 ( .C1(n5475), .C2(n6320), .A(n5134), .B(n5133), .ZN(U3035)
         );
  AOI22_X1 U5893 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n5309), .B1(n6279), 
        .B2(n5308), .ZN(n5136) );
  AOI22_X1 U5894 ( .A1(n7155), .A2(n5310), .B1(n7154), .B2(n3425), .ZN(n5135)
         );
  OAI211_X1 U5895 ( .C1(n5227), .C2(n5339), .A(n5136), .B(n5135), .ZN(U3093)
         );
  NAND2_X1 U5896 ( .A1(n5137), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5138) );
  XNOR2_X1 U5897 ( .A(n5138), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5144)
         );
  INV_X1 U5898 ( .A(n5154), .ZN(n5143) );
  CLKBUF_X1 U5899 ( .A(n5139), .Z(n5765) );
  INV_X1 U5900 ( .A(n5140), .ZN(n5141) );
  OAI211_X1 U5901 ( .C1(n5765), .C2(n5762), .A(n5142), .B(n5141), .ZN(n5760)
         );
  AOI22_X1 U5902 ( .A1(n5814), .A2(n5144), .B1(n5143), .B2(n5760), .ZN(n5151)
         );
  OR2_X1 U5903 ( .A1(n5843), .A2(n5145), .ZN(n5157) );
  INV_X1 U5904 ( .A(n5164), .ZN(n5149) );
  INV_X1 U5905 ( .A(n5146), .ZN(n5147) );
  MUX2_X1 U5906 ( .A(n5147), .B(n5762), .S(n5765), .Z(n5148) );
  NAND3_X1 U5907 ( .A1(n5157), .A2(n5149), .A3(n5148), .ZN(n5150) );
  OAI211_X1 U5908 ( .C1(n5214), .C2(n5808), .A(n5151), .B(n5150), .ZN(n5761)
         );
  MUX2_X1 U5909 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5761), .S(n5169), 
        .Z(n7031) );
  AND2_X1 U5910 ( .A1(n7062), .A2(n7031), .ZN(n5162) );
  OR2_X1 U5911 ( .A1(n5169), .A2(n3739), .ZN(n5160) );
  XNOR2_X1 U5912 ( .A(n5765), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5156)
         );
  XNOR2_X1 U5913 ( .A(n3592), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5152)
         );
  NAND2_X1 U5914 ( .A1(n5814), .A2(n5152), .ZN(n5153) );
  OAI21_X1 U5915 ( .B1(n5156), .B2(n5154), .A(n5153), .ZN(n5155) );
  AOI21_X1 U5916 ( .B1(n5157), .B2(n5156), .A(n5155), .ZN(n5158) );
  OAI21_X1 U5917 ( .B1(n5344), .B2(n5808), .A(n5158), .ZN(n5771) );
  NAND2_X1 U5918 ( .A1(n5169), .A2(n5771), .ZN(n5159) );
  INV_X1 U5919 ( .A(n7030), .ZN(n5161) );
  NAND2_X1 U5920 ( .A1(n5162), .A2(n5161), .ZN(n5166) );
  NOR2_X1 U5921 ( .A1(FLUSH_REG_SCAN_IN), .A2(n7062), .ZN(n5163) );
  NAND2_X1 U5922 ( .A1(n5164), .A2(n5163), .ZN(n5165) );
  NAND2_X1 U5923 ( .A1(n5166), .A2(n5165), .ZN(n7044) );
  INV_X1 U5924 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U5925 ( .A1(n7044), .A2(n5168), .ZN(n5179) );
  MUX2_X1 U5926 ( .A(n5169), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n5170) );
  INV_X1 U5927 ( .A(n5170), .ZN(n5178) );
  INV_X1 U5928 ( .A(n5172), .ZN(n5173) );
  NOR2_X1 U5929 ( .A1(n5171), .A2(n5173), .ZN(n5174) );
  XNOR2_X1 U5930 ( .A(n5174), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n7013)
         );
  INV_X1 U5931 ( .A(n5175), .ZN(n7015) );
  NAND2_X1 U5932 ( .A1(n7015), .A2(n7062), .ZN(n5176) );
  NOR2_X1 U5933 ( .A1(n7013), .A2(n5176), .ZN(n5177) );
  AOI21_X1 U5934 ( .B1(n5178), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(n5177), 
        .ZN(n7042) );
  NAND2_X1 U5935 ( .A1(n5179), .A2(n7042), .ZN(n5793) );
  INV_X1 U5936 ( .A(n7064), .ZN(n6738) );
  OAI21_X1 U5937 ( .B1(n5793), .B2(FLUSH_REG_SCAN_IN), .A(n6738), .ZN(n5180)
         );
  OAI21_X1 U5938 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n7062), .A(n5797), .ZN(
        n5799) );
  NAND2_X1 U5939 ( .A1(n5415), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5183) );
  NOR2_X1 U5940 ( .A1(n5210), .A2(n5183), .ZN(n7120) );
  AOI21_X1 U5941 ( .B1(n5210), .B2(n5183), .A(n7120), .ZN(n5182) );
  OAI222_X1 U5942 ( .A1(n5799), .A2(n5344), .B1(n5794), .B2(n5182), .C1(n5181), 
        .C2(n5797), .ZN(U3463) );
  NAND2_X1 U5943 ( .A1(n5210), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5187) );
  NOR2_X1 U5944 ( .A1(n5184), .A2(n5183), .ZN(n7133) );
  NAND2_X1 U5945 ( .A1(n5185), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5186) );
  NOR2_X1 U5946 ( .A1(n6230), .A2(n5186), .ZN(n6222) );
  AOI211_X1 U5947 ( .C1(n4403), .C2(n5187), .A(n7133), .B(n6222), .ZN(n5188)
         );
  OAI222_X1 U5948 ( .A1(n5799), .A2(n5214), .B1(n5797), .B2(n4200), .C1(n5794), 
        .C2(n5188), .ZN(U3462) );
  NAND2_X1 U5949 ( .A1(n5191), .A2(n5190), .ZN(n5192) );
  AND2_X1 U5950 ( .A1(n5189), .A2(n5192), .ZN(n5504) );
  NAND2_X1 U5951 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  NAND2_X1 U5952 ( .A1(n5419), .A2(n5195), .ZN(n5204) );
  INV_X1 U5953 ( .A(n5204), .ZN(n5448) );
  AOI22_X1 U5954 ( .A1(n6649), .A2(n5448), .B1(n5970), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n5196) );
  OAI21_X1 U5955 ( .B1(n5262), .B2(n6005), .A(n5196), .ZN(U2851) );
  NAND2_X1 U5956 ( .A1(n6998), .A2(n6904), .ZN(n5202) );
  NAND2_X1 U5957 ( .A1(n5826), .A2(n5202), .ZN(n6921) );
  AOI22_X1 U5958 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n6968), .B1(
        REIP_REG_8__SCAN_IN), .B2(n6921), .ZN(n5198) );
  INV_X1 U5959 ( .A(n6967), .ZN(n6944) );
  OAI211_X1 U5960 ( .C1(n6914), .C2(n5199), .A(n5198), .B(n6944), .ZN(n5200)
         );
  INV_X1 U5961 ( .A(n5200), .ZN(n5208) );
  INV_X1 U5962 ( .A(n5201), .ZN(n5203) );
  OAI22_X1 U5963 ( .A1(n7004), .A2(n5204), .B1(n5203), .B2(n5202), .ZN(n5205)
         );
  AOI21_X1 U5964 ( .B1(n5206), .B2(n6981), .A(n5205), .ZN(n5207) );
  OAI211_X1 U5965 ( .C1(n5262), .C2(n6978), .A(n5208), .B(n5207), .ZN(U2819)
         );
  INV_X1 U5966 ( .A(n5417), .ZN(n5364) );
  AND2_X1 U5967 ( .A1(n5344), .A2(n5364), .ZN(n7121) );
  NOR2_X1 U5968 ( .A1(n5210), .A2(n5209), .ZN(n5211) );
  AND2_X1 U5969 ( .A1(n5211), .A2(n5415), .ZN(n5518) );
  NAND2_X1 U5970 ( .A1(n5518), .A2(n5263), .ZN(n5220) );
  AOI21_X1 U5971 ( .B1(n5475), .B2(n5220), .A(n5212), .ZN(n5213) );
  AOI21_X1 U5972 ( .B1(n5214), .B2(n7121), .A(n5213), .ZN(n5215) );
  NOR2_X1 U5973 ( .A1(n5215), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U5974 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n5216), .ZN(n5271) );
  NOR2_X1 U5975 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5271), .ZN(n5221)
         );
  NAND2_X1 U5976 ( .A1(n5468), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5226) );
  INV_X1 U5977 ( .A(n5221), .ZN(n5470) );
  INV_X1 U5978 ( .A(n5222), .ZN(n5223) );
  AOI22_X1 U5979 ( .A1(n6266), .A2(n7121), .B1(n5223), .B2(n5522), .ZN(n5469)
         );
  OAI22_X1 U5980 ( .A1(n6236), .A2(n5470), .B1(n5469), .B2(n7159), .ZN(n5224)
         );
  AOI21_X1 U5981 ( .B1(n7154), .B2(n5472), .A(n5224), .ZN(n5225) );
  OAI211_X1 U5982 ( .C1(n5227), .C2(n5475), .A(n5226), .B(n5225), .ZN(U3037)
         );
  NAND2_X1 U5983 ( .A1(n5468), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5230) );
  OAI22_X1 U5984 ( .A1(n6242), .A2(n5470), .B1(n5469), .B2(n7175), .ZN(n5228)
         );
  AOI21_X1 U5985 ( .B1(n7170), .B2(n5472), .A(n5228), .ZN(n5229) );
  OAI211_X1 U5986 ( .C1(n5231), .C2(n5475), .A(n5230), .B(n5229), .ZN(U3039)
         );
  NAND2_X1 U5987 ( .A1(n5468), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5234) );
  OAI22_X1 U5988 ( .A1(n6258), .A2(n5470), .B1(n5469), .B2(n7216), .ZN(n5232)
         );
  AOI21_X1 U5989 ( .B1(n7212), .B2(n5472), .A(n5232), .ZN(n5233) );
  OAI211_X1 U5990 ( .C1(n5235), .C2(n5475), .A(n5234), .B(n5233), .ZN(U3043)
         );
  NAND2_X1 U5991 ( .A1(n5468), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5238) );
  OAI22_X1 U5992 ( .A1(n6248), .A2(n5470), .B1(n5469), .B2(n7191), .ZN(n5236)
         );
  AOI21_X1 U5993 ( .B1(n7186), .B2(n5472), .A(n5236), .ZN(n5237) );
  OAI211_X1 U5994 ( .C1(n5239), .C2(n5475), .A(n5238), .B(n5237), .ZN(U3041)
         );
  NAND2_X1 U5995 ( .A1(n5468), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U5996 ( .A1(n6233), .A2(n5470), .B1(n5469), .B2(n7151), .ZN(n5240)
         );
  AOI21_X1 U5997 ( .B1(n7148), .B2(n5472), .A(n5240), .ZN(n5241) );
  OAI211_X1 U5998 ( .C1(n5243), .C2(n5475), .A(n5242), .B(n5241), .ZN(U3036)
         );
  INV_X1 U5999 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5247) );
  NOR2_X2 U6000 ( .A1(n5252), .A2(n4377), .ZN(n7163) );
  AND2_X1 U6001 ( .A1(n6713), .A2(DATAI_26_), .ZN(n7162) );
  INV_X1 U6002 ( .A(n7162), .ZN(n5467) );
  NAND2_X1 U6003 ( .A1(n6713), .A2(DATAI_18_), .ZN(n6287) );
  INV_X1 U6004 ( .A(n6287), .ZN(n7164) );
  NOR2_X1 U6005 ( .A1(n6483), .A2(n5253), .ZN(n6285) );
  AOI22_X1 U6006 ( .A1(n5255), .A2(n7164), .B1(n6285), .B2(n5254), .ZN(n5244)
         );
  OAI21_X1 U6007 ( .B1(n5467), .B2(n6319), .A(n5244), .ZN(n5245) );
  AOI21_X1 U6008 ( .B1(n7163), .B2(n5258), .A(n5245), .ZN(n5246) );
  OAI21_X1 U6009 ( .B1(n5261), .B2(n5247), .A(n5246), .ZN(U3142) );
  INV_X1 U6010 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5251) );
  NOR2_X2 U6011 ( .A1(n5252), .A2(n3442), .ZN(n7195) );
  AND2_X1 U6012 ( .A1(n6713), .A2(DATAI_30_), .ZN(n7196) );
  INV_X1 U6013 ( .A(n7196), .ZN(n5463) );
  NAND2_X1 U6014 ( .A1(n6713), .A2(DATAI_22_), .ZN(n6311) );
  INV_X1 U6015 ( .A(n6311), .ZN(n7194) );
  NOR2_X1 U6016 ( .A1(n6431), .A2(n5253), .ZN(n6309) );
  AOI22_X1 U6017 ( .A1(n5255), .A2(n7194), .B1(n6309), .B2(n5254), .ZN(n5248)
         );
  OAI21_X1 U6018 ( .B1(n5463), .B2(n6319), .A(n5248), .ZN(n5249) );
  AOI21_X1 U6019 ( .B1(n7195), .B2(n5258), .A(n5249), .ZN(n5250) );
  OAI21_X1 U6020 ( .B1(n5261), .B2(n5251), .A(n5250), .ZN(U3146) );
  INV_X1 U6021 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5260) );
  NOR2_X2 U6022 ( .A1(n5252), .A2(n3594), .ZN(n7179) );
  AND2_X1 U6023 ( .A1(n6713), .A2(DATAI_28_), .ZN(n7178) );
  INV_X1 U6024 ( .A(n7178), .ZN(n5476) );
  NAND2_X1 U6025 ( .A1(n6713), .A2(DATAI_20_), .ZN(n6299) );
  INV_X1 U6026 ( .A(n6299), .ZN(n7180) );
  NOR2_X1 U6027 ( .A1(n6481), .A2(n5253), .ZN(n6297) );
  AOI22_X1 U6028 ( .A1(n5255), .A2(n7180), .B1(n6297), .B2(n5254), .ZN(n5256)
         );
  OAI21_X1 U6029 ( .B1(n5476), .B2(n6319), .A(n5256), .ZN(n5257) );
  AOI21_X1 U6030 ( .B1(n7179), .B2(n5258), .A(n5257), .ZN(n5259) );
  OAI21_X1 U6031 ( .B1(n5261), .B2(n5260), .A(n5259), .ZN(U3144) );
  INV_X1 U6032 ( .A(DATAI_8_), .ZN(n6474) );
  INV_X1 U6033 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6557) );
  OAI222_X1 U6034 ( .A1(n5262), .A2(n7100), .B1(n6027), .B2(n6474), .C1(n6026), 
        .C2(n6557), .ZN(U2883) );
  AOI21_X1 U6035 ( .B1(n7120), .B2(n5263), .A(n7132), .ZN(n5273) );
  INV_X1 U6036 ( .A(n7121), .ZN(n5268) );
  INV_X1 U6037 ( .A(n5264), .ZN(n5265) );
  NOR2_X1 U6038 ( .A1(n5266), .A2(n5265), .ZN(n5290) );
  INV_X1 U6039 ( .A(n5290), .ZN(n5267) );
  OAI21_X1 U6040 ( .B1(n7135), .B2(n5268), .A(n5267), .ZN(n5270) );
  INV_X1 U6041 ( .A(n5271), .ZN(n5269) );
  AOI22_X1 U6042 ( .A1(n5273), .A2(n5270), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5269), .ZN(n5293) );
  INV_X1 U6043 ( .A(n5270), .ZN(n5272) );
  AOI22_X1 U6044 ( .A1(n5273), .A2(n5272), .B1(n5271), .B2(n7132), .ZN(n5274)
         );
  NAND2_X1 U6045 ( .A1(n7143), .A2(n5274), .ZN(n5289) );
  AOI22_X1 U6046 ( .A1(n7139), .A2(n5290), .B1(INSTQUEUE_REG_3__0__SCAN_IN), 
        .B2(n5289), .ZN(n5276) );
  AOI22_X1 U6047 ( .A1(n5472), .A2(n7138), .B1(n5378), .B2(n7148), .ZN(n5275)
         );
  OAI211_X1 U6048 ( .C1(n5293), .C2(n7151), .A(n5276), .B(n5275), .ZN(U3044)
         );
  AOI22_X1 U6049 ( .A1(n7187), .A2(n5290), .B1(INSTQUEUE_REG_3__5__SCAN_IN), 
        .B2(n5289), .ZN(n5278) );
  AOI22_X1 U6050 ( .A1(n5472), .A2(n7188), .B1(n5378), .B2(n7186), .ZN(n5277)
         );
  OAI211_X1 U6051 ( .C1(n5293), .C2(n7191), .A(n5278), .B(n5277), .ZN(U3049)
         );
  AOI22_X1 U6052 ( .A1(n7210), .A2(n5290), .B1(INSTQUEUE_REG_3__7__SCAN_IN), 
        .B2(n5289), .ZN(n5280) );
  AOI22_X1 U6053 ( .A1(n5472), .A2(n7208), .B1(n5378), .B2(n7212), .ZN(n5279)
         );
  OAI211_X1 U6054 ( .C1(n5293), .C2(n7216), .A(n5280), .B(n5279), .ZN(U3051)
         );
  AOI22_X1 U6055 ( .A1(n7155), .A2(n5290), .B1(INSTQUEUE_REG_3__1__SCAN_IN), 
        .B2(n5289), .ZN(n5282) );
  AOI22_X1 U6056 ( .A1(n5472), .A2(n7156), .B1(n5378), .B2(n7154), .ZN(n5281)
         );
  OAI211_X1 U6057 ( .C1(n5293), .C2(n7159), .A(n5282), .B(n5281), .ZN(U3045)
         );
  AOI22_X1 U6058 ( .A1(n7171), .A2(n5290), .B1(INSTQUEUE_REG_3__3__SCAN_IN), 
        .B2(n5289), .ZN(n5284) );
  AOI22_X1 U6059 ( .A1(n5472), .A2(n7172), .B1(n5378), .B2(n7170), .ZN(n5283)
         );
  OAI211_X1 U6060 ( .C1(n5293), .C2(n7175), .A(n5284), .B(n5283), .ZN(U3047)
         );
  AOI22_X1 U6061 ( .A1(n7179), .A2(n5290), .B1(INSTQUEUE_REG_3__4__SCAN_IN), 
        .B2(n5289), .ZN(n5286) );
  AOI22_X1 U6062 ( .A1(n5472), .A2(n7178), .B1(n5378), .B2(n7180), .ZN(n5285)
         );
  OAI211_X1 U6063 ( .C1(n5293), .C2(n7183), .A(n5286), .B(n5285), .ZN(U3048)
         );
  AOI22_X1 U6064 ( .A1(n7195), .A2(n5290), .B1(INSTQUEUE_REG_3__6__SCAN_IN), 
        .B2(n5289), .ZN(n5288) );
  AOI22_X1 U6065 ( .A1(n5472), .A2(n7196), .B1(n5378), .B2(n7194), .ZN(n5287)
         );
  OAI211_X1 U6066 ( .C1(n5293), .C2(n7199), .A(n5288), .B(n5287), .ZN(U3050)
         );
  AOI22_X1 U6067 ( .A1(n7163), .A2(n5290), .B1(INSTQUEUE_REG_3__2__SCAN_IN), 
        .B2(n5289), .ZN(n5292) );
  AOI22_X1 U6068 ( .A1(n5472), .A2(n7162), .B1(n5378), .B2(n7164), .ZN(n5291)
         );
  OAI211_X1 U6069 ( .C1(n5293), .C2(n7167), .A(n5292), .B(n5291), .ZN(U3046)
         );
  AOI22_X1 U6070 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5303), .B1(n6309), 
        .B2(n5302), .ZN(n5295) );
  AOI22_X1 U6071 ( .A1(n7195), .A2(n5305), .B1(n5304), .B2(n7196), .ZN(n5294)
         );
  OAI211_X1 U6072 ( .C1(n5475), .C2(n6311), .A(n5295), .B(n5294), .ZN(U3034)
         );
  AOI22_X1 U6073 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5303), .B1(n6297), 
        .B2(n5302), .ZN(n5297) );
  AOI22_X1 U6074 ( .A1(n7179), .A2(n5305), .B1(n5304), .B2(n7178), .ZN(n5296)
         );
  OAI211_X1 U6075 ( .C1(n5475), .C2(n6299), .A(n5297), .B(n5296), .ZN(U3032)
         );
  AOI22_X1 U6076 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n5309), .B1(n6309), 
        .B2(n5308), .ZN(n5299) );
  AOI22_X1 U6077 ( .A1(n7195), .A2(n5310), .B1(n7194), .B2(n3425), .ZN(n5298)
         );
  OAI211_X1 U6078 ( .C1(n5463), .C2(n5339), .A(n5299), .B(n5298), .ZN(U3098)
         );
  AOI22_X1 U6079 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5309), .B1(n6297), 
        .B2(n5308), .ZN(n5301) );
  AOI22_X1 U6080 ( .A1(n7179), .A2(n5310), .B1(n7180), .B2(n3425), .ZN(n5300)
         );
  OAI211_X1 U6081 ( .C1(n5476), .C2(n5339), .A(n5301), .B(n5300), .ZN(U3096)
         );
  AOI22_X1 U6082 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5303), .B1(n6285), 
        .B2(n5302), .ZN(n5307) );
  AOI22_X1 U6083 ( .A1(n7163), .A2(n5305), .B1(n5304), .B2(n7162), .ZN(n5306)
         );
  OAI211_X1 U6084 ( .C1(n5475), .C2(n6287), .A(n5307), .B(n5306), .ZN(U3030)
         );
  AOI22_X1 U6085 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n5309), .B1(n6285), 
        .B2(n5308), .ZN(n5312) );
  AOI22_X1 U6086 ( .A1(n7163), .A2(n5310), .B1(n7164), .B2(n3425), .ZN(n5311)
         );
  OAI211_X1 U6087 ( .C1(n5467), .C2(n5339), .A(n5312), .B(n5311), .ZN(U3094)
         );
  NAND2_X1 U6088 ( .A1(n5319), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5315) );
  OAI22_X1 U6089 ( .A1(n5321), .A2(n5476), .B1(n5320), .B2(n7183), .ZN(n5313)
         );
  AOI21_X1 U6090 ( .B1(n7179), .B2(n5323), .A(n5313), .ZN(n5314) );
  OAI211_X1 U6091 ( .C1(n6299), .C2(n5326), .A(n5315), .B(n5314), .ZN(U3024)
         );
  NAND2_X1 U6092 ( .A1(n5319), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5318) );
  OAI22_X1 U6093 ( .A1(n5321), .A2(n5467), .B1(n5320), .B2(n7167), .ZN(n5316)
         );
  AOI21_X1 U6094 ( .B1(n7163), .B2(n5323), .A(n5316), .ZN(n5317) );
  OAI211_X1 U6095 ( .C1(n6287), .C2(n5326), .A(n5318), .B(n5317), .ZN(U3022)
         );
  NAND2_X1 U6096 ( .A1(n5319), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5325) );
  OAI22_X1 U6097 ( .A1(n5321), .A2(n5463), .B1(n5320), .B2(n7199), .ZN(n5322)
         );
  AOI21_X1 U6098 ( .B1(n7195), .B2(n5323), .A(n5322), .ZN(n5324) );
  OAI211_X1 U6099 ( .C1(n6311), .C2(n5326), .A(n5325), .B(n5324), .ZN(U3026)
         );
  NAND2_X1 U6100 ( .A1(n5333), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5329) );
  OAI22_X1 U6101 ( .A1(n7147), .A2(n5476), .B1(n5334), .B2(n7183), .ZN(n5327)
         );
  AOI21_X1 U6102 ( .B1(n7179), .B2(n5336), .A(n5327), .ZN(n5328) );
  OAI211_X1 U6103 ( .C1(n5339), .C2(n6299), .A(n5329), .B(n5328), .ZN(U3088)
         );
  NAND2_X1 U6104 ( .A1(n5333), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5332) );
  OAI22_X1 U6105 ( .A1(n7147), .A2(n5467), .B1(n5334), .B2(n7167), .ZN(n5330)
         );
  AOI21_X1 U6106 ( .B1(n7163), .B2(n5336), .A(n5330), .ZN(n5331) );
  OAI211_X1 U6107 ( .C1(n5339), .C2(n6287), .A(n5332), .B(n5331), .ZN(U3086)
         );
  NAND2_X1 U6108 ( .A1(n5333), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5338) );
  OAI22_X1 U6109 ( .A1(n7147), .A2(n5463), .B1(n5334), .B2(n7199), .ZN(n5335)
         );
  AOI21_X1 U6110 ( .B1(n7195), .B2(n5336), .A(n5335), .ZN(n5337) );
  OAI211_X1 U6111 ( .C1(n5339), .C2(n6311), .A(n5338), .B(n5337), .ZN(U3090)
         );
  INV_X1 U6112 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5342) );
  OAI211_X1 U6113 ( .C1(REIP_REG_1__SCAN_IN), .C2(REIP_REG_2__SCAN_IN), .A(
        n6998), .B(n5354), .ZN(n5341) );
  NAND2_X1 U6114 ( .A1(n6968), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5340)
         );
  OAI211_X1 U6115 ( .C1(n5342), .C2(n5826), .A(n5341), .B(n5340), .ZN(n5347)
         );
  INV_X1 U6116 ( .A(n5343), .ZN(n5855) );
  NAND2_X1 U6117 ( .A1(n5872), .A2(n5855), .ZN(n6865) );
  OAI22_X1 U6118 ( .A1(n6914), .A2(n5345), .B1(n5344), .B2(n6865), .ZN(n5346)
         );
  AOI211_X1 U6119 ( .C1(n6993), .C2(n5348), .A(n5347), .B(n5346), .ZN(n5352)
         );
  INV_X1 U6120 ( .A(n5349), .ZN(n5853) );
  OAI21_X1 U6121 ( .B1(n5853), .B2(n5350), .A(n6978), .ZN(n6886) );
  NAND2_X1 U6122 ( .A1(n6886), .A2(n6667), .ZN(n5351) );
  OAI211_X1 U6123 ( .C1(n7010), .C2(n6671), .A(n5352), .B(n5351), .ZN(U2825)
         );
  INV_X1 U6124 ( .A(n6886), .ZN(n5400) );
  INV_X1 U6125 ( .A(n6679), .ZN(n5360) );
  NAND2_X1 U6126 ( .A1(n5826), .A2(n6870), .ZN(n5353) );
  NAND2_X1 U6127 ( .A1(n5396), .A2(n5353), .ZN(n6866) );
  INV_X1 U6128 ( .A(n5354), .ZN(n5355) );
  AOI21_X1 U6129 ( .B1(n5826), .B2(n5355), .A(REIP_REG_3__SCAN_IN), .ZN(n5358)
         );
  AOI22_X1 U6130 ( .A1(n7003), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6968), .ZN(n5357) );
  INV_X1 U6131 ( .A(n6865), .ZN(n5365) );
  AOI22_X1 U6132 ( .A1(n5365), .A2(n4913), .B1(n6993), .B2(n6772), .ZN(n5356)
         );
  OAI211_X1 U6133 ( .C1(n6866), .C2(n5358), .A(n5357), .B(n5356), .ZN(n5359)
         );
  AOI21_X1 U6134 ( .B1(n5360), .B2(n6981), .A(n5359), .ZN(n5361) );
  OAI21_X1 U6135 ( .B1(n5400), .B2(n6675), .A(n5361), .ZN(U2824) );
  INV_X1 U6136 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5577) );
  NAND2_X1 U6137 ( .A1(n6981), .A2(n5577), .ZN(n5369) );
  AOI22_X1 U6138 ( .A1(n6993), .A2(n5362), .B1(n7003), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5368) );
  INV_X1 U6139 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6757) );
  OAI22_X1 U6140 ( .A1(n6999), .A2(n5577), .B1(n5826), .B2(n6757), .ZN(n5363)
         );
  AOI21_X1 U6141 ( .B1(n6998), .B2(n6757), .A(n5363), .ZN(n5367) );
  NAND2_X1 U6142 ( .A1(n5365), .A2(n5364), .ZN(n5366) );
  AND4_X1 U6143 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n5370)
         );
  OAI21_X1 U6144 ( .B1(n5400), .B2(n5576), .A(n5370), .ZN(U2826) );
  INV_X1 U6145 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5373) );
  AOI22_X1 U6146 ( .A1(n5390), .A2(n7164), .B1(n6285), .B2(n5377), .ZN(n5372)
         );
  AOI22_X1 U6147 ( .A1(n7163), .A2(n5379), .B1(n7162), .B2(n5378), .ZN(n5371)
         );
  OAI211_X1 U6148 ( .C1(n5383), .C2(n5373), .A(n5372), .B(n5371), .ZN(U3054)
         );
  INV_X1 U6149 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5376) );
  AOI22_X1 U6150 ( .A1(n5390), .A2(n7180), .B1(n6297), .B2(n5377), .ZN(n5375)
         );
  AOI22_X1 U6151 ( .A1(n7179), .A2(n5379), .B1(n7178), .B2(n5378), .ZN(n5374)
         );
  OAI211_X1 U6152 ( .C1(n5383), .C2(n5376), .A(n5375), .B(n5374), .ZN(U3056)
         );
  INV_X1 U6153 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5382) );
  AOI22_X1 U6154 ( .A1(n5390), .A2(n7194), .B1(n6309), .B2(n5377), .ZN(n5381)
         );
  AOI22_X1 U6155 ( .A1(n7195), .A2(n5379), .B1(n7196), .B2(n5378), .ZN(n5380)
         );
  OAI211_X1 U6156 ( .C1(n5383), .C2(n5382), .A(n5381), .B(n5380), .ZN(U3058)
         );
  INV_X1 U6157 ( .A(n7195), .ZN(n6251) );
  AOI22_X1 U6158 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n5389), .B1(n6309), 
        .B2(n5388), .ZN(n5385) );
  AOI22_X1 U6159 ( .A1(n7194), .A2(n5411), .B1(n5390), .B2(n7196), .ZN(n5384)
         );
  OAI211_X1 U6160 ( .C1(n6251), .C2(n5393), .A(n5385), .B(n5384), .ZN(U3066)
         );
  INV_X1 U6161 ( .A(n7163), .ZN(n6239) );
  AOI22_X1 U6162 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n5389), .B1(n6285), 
        .B2(n5388), .ZN(n5387) );
  AOI22_X1 U6163 ( .A1(n7164), .A2(n5411), .B1(n5390), .B2(n7162), .ZN(n5386)
         );
  OAI211_X1 U6164 ( .C1(n6239), .C2(n5393), .A(n5387), .B(n5386), .ZN(U3062)
         );
  INV_X1 U6165 ( .A(n7179), .ZN(n6245) );
  AOI22_X1 U6166 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n5389), .B1(n6297), 
        .B2(n5388), .ZN(n5392) );
  AOI22_X1 U6167 ( .A1(n7180), .A2(n5411), .B1(n5390), .B2(n7178), .ZN(n5391)
         );
  OAI211_X1 U6168 ( .C1(n6245), .C2(n5393), .A(n5392), .B(n5391), .ZN(U3064)
         );
  AOI22_X1 U6169 ( .A1(n6859), .A2(n6993), .B1(n7003), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5394) );
  OAI21_X1 U6170 ( .B1(n5800), .B2(n6865), .A(n5394), .ZN(n5395) );
  AOI21_X1 U6171 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5396), .A(n5395), .ZN(n5398)
         );
  OAI21_X1 U6172 ( .B1(n6981), .B2(n6968), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5397) );
  OAI211_X1 U6173 ( .C1(n5400), .C2(n5399), .A(n5398), .B(n5397), .ZN(U2827)
         );
  NAND2_X1 U6174 ( .A1(n5407), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5403) );
  OAI22_X1 U6175 ( .A1(n5409), .A2(n6311), .B1(n5408), .B2(n7199), .ZN(n5401)
         );
  AOI21_X1 U6176 ( .B1(n7196), .B2(n5411), .A(n5401), .ZN(n5402) );
  OAI211_X1 U6177 ( .C1(n5414), .C2(n6251), .A(n5403), .B(n5402), .ZN(U3074)
         );
  NAND2_X1 U6178 ( .A1(n5407), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5406) );
  OAI22_X1 U6179 ( .A1(n5409), .A2(n6287), .B1(n5408), .B2(n7167), .ZN(n5404)
         );
  AOI21_X1 U6180 ( .B1(n7162), .B2(n5411), .A(n5404), .ZN(n5405) );
  OAI211_X1 U6181 ( .C1(n5414), .C2(n6239), .A(n5406), .B(n5405), .ZN(U3070)
         );
  NAND2_X1 U6182 ( .A1(n5407), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5413) );
  OAI22_X1 U6183 ( .A1(n5409), .A2(n6299), .B1(n5408), .B2(n7183), .ZN(n5410)
         );
  AOI21_X1 U6184 ( .B1(n7178), .B2(n5411), .A(n5410), .ZN(n5412) );
  OAI211_X1 U6185 ( .C1(n5414), .C2(n6245), .A(n5413), .B(n5412), .ZN(U3072)
         );
  XNOR2_X1 U6186 ( .A(n5415), .B(STATEBS16_REG_SCAN_IN), .ZN(n5416) );
  OAI222_X1 U6187 ( .A1(n5799), .A2(n5417), .B1(n5794), .B2(n5416), .C1(n5523), 
        .C2(n5797), .ZN(U3464) );
  XNOR2_X1 U6188 ( .A(n5189), .B(n5418), .ZN(n6906) );
  AOI21_X1 U6189 ( .B1(n5420), .B2(n5419), .A(n5456), .ZN(n6903) );
  AOI22_X1 U6190 ( .A1(n6649), .A2(n6903), .B1(EBX_REG_9__SCAN_IN), .B2(n5970), 
        .ZN(n5421) );
  OAI21_X1 U6191 ( .B1(n6906), .B2(n6001), .A(n5421), .ZN(U2850) );
  NAND2_X1 U6192 ( .A1(n7179), .A2(n5430), .ZN(n5423) );
  AOI22_X1 U6193 ( .A1(n6254), .A2(n7180), .B1(n6297), .B2(n5431), .ZN(n5422)
         );
  OAI211_X1 U6194 ( .C1(n7124), .C2(n5476), .A(n5423), .B(n5422), .ZN(n5424)
         );
  AOI21_X1 U6195 ( .B1(n5435), .B2(INSTQUEUE_REG_12__4__SCAN_IN), .A(n5424), 
        .ZN(n5425) );
  INV_X1 U6196 ( .A(n5425), .ZN(U3120) );
  NAND2_X1 U6197 ( .A1(n7195), .A2(n5430), .ZN(n5427) );
  AOI22_X1 U6198 ( .A1(n6254), .A2(n7194), .B1(n6309), .B2(n5431), .ZN(n5426)
         );
  OAI211_X1 U6199 ( .C1(n7124), .C2(n5463), .A(n5427), .B(n5426), .ZN(n5428)
         );
  AOI21_X1 U6200 ( .B1(n5435), .B2(INSTQUEUE_REG_12__6__SCAN_IN), .A(n5428), 
        .ZN(n5429) );
  INV_X1 U6201 ( .A(n5429), .ZN(U3122) );
  NAND2_X1 U6202 ( .A1(n7163), .A2(n5430), .ZN(n5433) );
  AOI22_X1 U6203 ( .A1(n6254), .A2(n7164), .B1(n6285), .B2(n5431), .ZN(n5432)
         );
  OAI211_X1 U6204 ( .C1(n7124), .C2(n5467), .A(n5433), .B(n5432), .ZN(n5434)
         );
  AOI21_X1 U6205 ( .B1(n5435), .B2(INSTQUEUE_REG_12__2__SCAN_IN), .A(n5434), 
        .ZN(n5436) );
  INV_X1 U6206 ( .A(n5436), .ZN(U3118) );
  INV_X1 U6207 ( .A(DATAI_9_), .ZN(n6362) );
  INV_X1 U6208 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6559) );
  OAI222_X1 U6209 ( .A1(n7100), .A2(n6906), .B1(n6027), .B2(n6362), .C1(n6026), 
        .C2(n6559), .ZN(U2882) );
  XNOR2_X1 U6210 ( .A(n5439), .B(n5438), .ZN(n5506) );
  AOI21_X1 U6211 ( .B1(n5441), .B2(n6794), .A(n5440), .ZN(n6805) );
  INV_X1 U6212 ( .A(n6798), .ZN(n5669) );
  INV_X1 U6213 ( .A(n6805), .ZN(n5442) );
  AOI21_X1 U6214 ( .B1(n5669), .B2(n6795), .A(n5442), .ZN(n6778) );
  AOI22_X1 U6215 ( .A1(n6754), .A2(n6805), .B1(n5444), .B2(n6778), .ZN(n6808)
         );
  NAND2_X1 U6216 ( .A1(n6808), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n5450)
         );
  INV_X1 U6217 ( .A(n6795), .ZN(n5443) );
  OAI21_X1 U6218 ( .B1(n6790), .B2(n6794), .A(n6798), .ZN(n5560) );
  AND2_X1 U6219 ( .A1(n5443), .A2(n5560), .ZN(n6774) );
  NAND2_X1 U6220 ( .A1(n5444), .A2(n6774), .ZN(n6813) );
  AOI221_X1 U6221 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n5445), .C2(n6817), .A(n6813), 
        .ZN(n5447) );
  INV_X1 U6222 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U6223 ( .A1(n4480), .A2(n6584), .ZN(n5446) );
  AOI211_X1 U6224 ( .C1(n6860), .C2(n5448), .A(n5447), .B(n5446), .ZN(n5449)
         );
  OAI211_X1 U6225 ( .C1(n5506), .C2(n6800), .A(n5450), .B(n5449), .ZN(U3010)
         );
  NOR2_X1 U6226 ( .A1(n5452), .A2(n5453), .ZN(n5454) );
  OR2_X1 U6227 ( .A1(n5451), .A2(n5454), .ZN(n6919) );
  NOR2_X1 U6228 ( .A1(n5456), .A2(n5455), .ZN(n5457) );
  OR2_X1 U6229 ( .A1(n5491), .A2(n5457), .ZN(n6913) );
  INV_X1 U6230 ( .A(n6913), .ZN(n5458) );
  AOI22_X1 U6231 ( .A1(n6649), .A2(n5458), .B1(n5970), .B2(EBX_REG_10__SCAN_IN), .ZN(n5459) );
  OAI21_X1 U6232 ( .B1(n6919), .B2(n6005), .A(n5459), .ZN(U2849) );
  NAND2_X1 U6233 ( .A1(n5468), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5462) );
  OAI22_X1 U6234 ( .A1(n6251), .A2(n5470), .B1(n5469), .B2(n7199), .ZN(n5460)
         );
  AOI21_X1 U6235 ( .B1(n7194), .B2(n5472), .A(n5460), .ZN(n5461) );
  OAI211_X1 U6236 ( .C1(n5463), .C2(n5475), .A(n5462), .B(n5461), .ZN(U3042)
         );
  NAND2_X1 U6237 ( .A1(n5468), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5466) );
  OAI22_X1 U6238 ( .A1(n6239), .A2(n5470), .B1(n5469), .B2(n7167), .ZN(n5464)
         );
  AOI21_X1 U6239 ( .B1(n7164), .B2(n5472), .A(n5464), .ZN(n5465) );
  OAI211_X1 U6240 ( .C1(n5467), .C2(n5475), .A(n5466), .B(n5465), .ZN(U3038)
         );
  NAND2_X1 U6241 ( .A1(n5468), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5474) );
  OAI22_X1 U6242 ( .A1(n6245), .A2(n5470), .B1(n5469), .B2(n7183), .ZN(n5471)
         );
  AOI21_X1 U6243 ( .B1(n7180), .B2(n5472), .A(n5471), .ZN(n5473) );
  OAI211_X1 U6244 ( .C1(n5476), .C2(n5475), .A(n5474), .B(n5473), .ZN(U3040)
         );
  INV_X1 U6245 ( .A(n5477), .ZN(n5515) );
  OAI22_X1 U6246 ( .A1(n3860), .A2(n6999), .B1(n7004), .B2(n5600), .ZN(n5485)
         );
  INV_X1 U6247 ( .A(n5481), .ZN(n5478) );
  NOR3_X1 U6248 ( .A1(n6986), .A2(REIP_REG_6__SCAN_IN), .A3(n5478), .ZN(n6899)
         );
  NOR2_X1 U6249 ( .A1(n5479), .A2(n6914), .ZN(n5480) );
  NOR3_X1 U6250 ( .A1(n6899), .A2(n6967), .A3(n5480), .ZN(n5483) );
  OAI21_X1 U6251 ( .B1(n6986), .B2(n5481), .A(n5826), .ZN(n6898) );
  NAND2_X1 U6252 ( .A1(n6898), .A2(REIP_REG_6__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U6253 ( .C1(n7010), .C2(n5513), .A(n5483), .B(n5482), .ZN(n5484)
         );
  AOI211_X1 U6254 ( .C1(n5515), .C2(n7007), .A(n5485), .B(n5484), .ZN(n5486)
         );
  INV_X1 U6255 ( .A(n5486), .ZN(U2821) );
  INV_X1 U6256 ( .A(DATAI_10_), .ZN(n6464) );
  INV_X1 U6257 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6561) );
  OAI222_X1 U6258 ( .A1(n6919), .A2(n7100), .B1(n6027), .B2(n6464), .C1(n6026), 
        .C2(n6561), .ZN(U2881) );
  OAI21_X1 U6259 ( .B1(n5451), .B2(n5489), .A(n5488), .ZN(n5644) );
  OR2_X1 U6260 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  AND2_X1 U6261 ( .A1(n5628), .A2(n5492), .ZN(n6825) );
  AOI22_X1 U6262 ( .A1(n6649), .A2(n6825), .B1(EBX_REG_11__SCAN_IN), .B2(n5970), .ZN(n5493) );
  OAI21_X1 U6263 ( .B1(n5644), .B2(n6001), .A(n5493), .ZN(U2848) );
  INV_X1 U6264 ( .A(n5640), .ZN(n5496) );
  AOI22_X1 U6265 ( .A1(EBX_REG_11__SCAN_IN), .A2(n7003), .B1(n6993), .B2(n6825), .ZN(n5494) );
  OAI211_X1 U6266 ( .C1(n6999), .C2(n3939), .A(n5494), .B(n6944), .ZN(n5495)
         );
  AOI21_X1 U6267 ( .B1(n6981), .B2(n5496), .A(n5495), .ZN(n5500) );
  NOR2_X1 U6268 ( .A1(n6986), .A2(n5497), .ZN(n5685) );
  AND2_X1 U6269 ( .A1(n5498), .A2(n5826), .ZN(n6940) );
  NOR2_X1 U6270 ( .A1(n6941), .A2(n6940), .ZN(n6928) );
  OAI21_X1 U6271 ( .B1(REIP_REG_11__SCAN_IN), .B2(n5685), .A(n6928), .ZN(n5499) );
  OAI211_X1 U6272 ( .C1(n5644), .C2(n6978), .A(n5500), .B(n5499), .ZN(U2816)
         );
  AOI22_X1 U6273 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6771), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n5501) );
  OAI21_X1 U6274 ( .B1(n6717), .B2(n5502), .A(n5501), .ZN(n5503) );
  AOI21_X1 U6275 ( .B1(n5504), .B2(n6713), .A(n5503), .ZN(n5505) );
  OAI21_X1 U6276 ( .B1(n5506), .B2(n6696), .A(n5505), .ZN(U2978) );
  AND2_X1 U6277 ( .A1(n5508), .A2(n5507), .ZN(n5511) );
  XNOR2_X1 U6278 ( .A(n5509), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5510)
         );
  XNOR2_X1 U6279 ( .A(n5511), .B(n5510), .ZN(n5607) );
  NAND2_X1 U6280 ( .A1(n6771), .A2(REIP_REG_6__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U6281 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5512)
         );
  OAI211_X1 U6282 ( .C1(n6717), .C2(n5513), .A(n5599), .B(n5512), .ZN(n5514)
         );
  AOI21_X1 U6283 ( .B1(n5515), .B2(n6713), .A(n5514), .ZN(n5516) );
  OAI21_X1 U6284 ( .B1(n5607), .B2(n6696), .A(n5516), .ZN(U2980) );
  INV_X1 U6285 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6563) );
  OAI222_X1 U6286 ( .A1(n5644), .A2(n7100), .B1(n6027), .B2(n5517), .C1(n6026), 
        .C2(n6563), .ZN(U2880) );
  NAND2_X1 U6287 ( .A1(n5518), .A2(n4403), .ZN(n7129) );
  NAND2_X1 U6288 ( .A1(n7129), .A2(n7146), .ZN(n5520) );
  OAI21_X1 U6289 ( .B1(n3425), .B2(n5520), .A(n5519), .ZN(n5529) );
  AND2_X1 U6290 ( .A1(n7121), .A2(n4913), .ZN(n5525) );
  NAND2_X1 U6291 ( .A1(n5521), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6270) );
  INV_X1 U6292 ( .A(n6270), .ZN(n5526) );
  AOI22_X1 U6293 ( .A1(n5529), .A2(n5525), .B1(n5526), .B2(n5522), .ZN(n5558)
         );
  NOR3_X1 U6294 ( .A1(n4200), .A2(n5523), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n7128) );
  INV_X1 U6295 ( .A(n7128), .ZN(n5524) );
  NOR2_X1 U6296 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5524), .ZN(n5553)
         );
  INV_X1 U6297 ( .A(n5525), .ZN(n5528) );
  NOR2_X1 U6298 ( .A1(n5526), .A2(n6226), .ZN(n6261) );
  AOI211_X1 U6299 ( .C1(n5529), .C2(n5528), .A(n5527), .B(n6261), .ZN(n5530)
         );
  AOI22_X1 U6300 ( .A1(n7210), .A2(n5553), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5552), .ZN(n5531) );
  OAI21_X1 U6301 ( .B1(n6320), .B2(n7129), .A(n5531), .ZN(n5532) );
  AOI21_X1 U6302 ( .B1(n7208), .B2(n3425), .A(n5532), .ZN(n5533) );
  OAI21_X1 U6303 ( .B1(n5558), .B2(n7216), .A(n5533), .ZN(U3107) );
  AOI22_X1 U6304 ( .A1(n7195), .A2(n5553), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5552), .ZN(n5534) );
  OAI21_X1 U6305 ( .B1(n6311), .B2(n7129), .A(n5534), .ZN(n5535) );
  AOI21_X1 U6306 ( .B1(n7196), .B2(n3425), .A(n5535), .ZN(n5536) );
  OAI21_X1 U6307 ( .B1(n5558), .B2(n7199), .A(n5536), .ZN(U3106) );
  AOI22_X1 U6308 ( .A1(n7187), .A2(n5553), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5552), .ZN(n5537) );
  OAI21_X1 U6309 ( .B1(n6305), .B2(n7129), .A(n5537), .ZN(n5538) );
  AOI21_X1 U6310 ( .B1(n7188), .B2(n3425), .A(n5538), .ZN(n5539) );
  OAI21_X1 U6311 ( .B1(n5558), .B2(n7191), .A(n5539), .ZN(U3105) );
  AOI22_X1 U6312 ( .A1(n7171), .A2(n5553), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5552), .ZN(n5540) );
  OAI21_X1 U6313 ( .B1(n6293), .B2(n7129), .A(n5540), .ZN(n5541) );
  AOI21_X1 U6314 ( .B1(n7172), .B2(n3425), .A(n5541), .ZN(n5542) );
  OAI21_X1 U6315 ( .B1(n5558), .B2(n7175), .A(n5542), .ZN(U3103) );
  AOI22_X1 U6316 ( .A1(n7179), .A2(n5553), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5552), .ZN(n5543) );
  OAI21_X1 U6317 ( .B1(n6299), .B2(n7129), .A(n5543), .ZN(n5544) );
  AOI21_X1 U6318 ( .B1(n7178), .B2(n3425), .A(n5544), .ZN(n5545) );
  OAI21_X1 U6319 ( .B1(n5558), .B2(n7183), .A(n5545), .ZN(U3104) );
  AOI22_X1 U6320 ( .A1(n7139), .A2(n5553), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5552), .ZN(n5546) );
  OAI21_X1 U6321 ( .B1(n6275), .B2(n7129), .A(n5546), .ZN(n5547) );
  AOI21_X1 U6322 ( .B1(n7138), .B2(n3425), .A(n5547), .ZN(n5548) );
  OAI21_X1 U6323 ( .B1(n5558), .B2(n7151), .A(n5548), .ZN(U3100) );
  AOI22_X1 U6324 ( .A1(n7155), .A2(n5553), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5552), .ZN(n5549) );
  OAI21_X1 U6325 ( .B1(n6281), .B2(n7129), .A(n5549), .ZN(n5550) );
  AOI21_X1 U6326 ( .B1(n7156), .B2(n3425), .A(n5550), .ZN(n5551) );
  OAI21_X1 U6327 ( .B1(n5558), .B2(n7159), .A(n5551), .ZN(U3101) );
  AOI22_X1 U6328 ( .A1(n7163), .A2(n5553), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5552), .ZN(n5554) );
  OAI21_X1 U6329 ( .B1(n6287), .B2(n7129), .A(n5554), .ZN(n5555) );
  AOI21_X1 U6330 ( .B1(n7162), .B2(n3425), .A(n5555), .ZN(n5557) );
  OAI21_X1 U6331 ( .B1(n5558), .B2(n7167), .A(n5557), .ZN(U3102) );
  NAND2_X1 U6332 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5559) );
  OAI21_X1 U6333 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A(n5559), .ZN(n5573) );
  NAND2_X1 U6334 ( .A1(n5563), .A2(n5560), .ZN(n6823) );
  XNOR2_X1 U6335 ( .A(n6106), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5561)
         );
  XNOR2_X1 U6336 ( .A(n5562), .B(n5561), .ZN(n5593) );
  NAND2_X1 U6337 ( .A1(n5593), .A2(n6854), .ZN(n5572) );
  OR2_X1 U6338 ( .A1(n6798), .A2(n5563), .ZN(n5564) );
  OAI211_X1 U6339 ( .C1(n5567), .C2(n5566), .A(n5565), .B(n5564), .ZN(n6819)
         );
  INV_X1 U6340 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5568) );
  NOR2_X1 U6341 ( .A1(n4480), .A2(n5568), .ZN(n5595) );
  INV_X1 U6342 ( .A(n5595), .ZN(n5569) );
  OAI21_X1 U6343 ( .B1(n6793), .B2(n6913), .A(n5569), .ZN(n5570) );
  AOI21_X1 U6344 ( .B1(n6819), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5570), 
        .ZN(n5571) );
  OAI211_X1 U6345 ( .C1(n5573), .C2(n6823), .A(n5572), .B(n5571), .ZN(U3008)
         );
  XNOR2_X1 U6346 ( .A(n4860), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5574)
         );
  XNOR2_X1 U6347 ( .A(n5575), .B(n5574), .ZN(n6759) );
  NOR2_X1 U6348 ( .A1(n5576), .A2(n6121), .ZN(n5579) );
  OAI22_X1 U6349 ( .A1(n6101), .A2(n5577), .B1(n4480), .B2(n6757), .ZN(n5578)
         );
  AOI211_X1 U6350 ( .C1(n5577), .C2(n6693), .A(n5579), .B(n5578), .ZN(n5580)
         );
  OAI21_X1 U6351 ( .B1(n6759), .B2(n6696), .A(n5580), .ZN(U2985) );
  XOR2_X1 U6352 ( .A(n5582), .B(n5581), .Z(n6820) );
  NAND2_X1 U6353 ( .A1(n6820), .A2(n6714), .ZN(n5585) );
  NOR2_X1 U6354 ( .A1(n4480), .A2(n4356), .ZN(n6818) );
  NOR2_X1 U6355 ( .A1(n6717), .A2(n6907), .ZN(n5583) );
  AOI211_X1 U6356 ( .C1(n6707), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6818), 
        .B(n5583), .ZN(n5584) );
  OAI211_X1 U6357 ( .C1(n6906), .C2(n6121), .A(n5585), .B(n5584), .ZN(U2977)
         );
  CLKBUF_X1 U6358 ( .A(n5586), .Z(n5587) );
  INV_X1 U6359 ( .A(n5588), .ZN(n5589) );
  XNOR2_X1 U6360 ( .A(n5587), .B(n5589), .ZN(n6810) );
  NAND2_X1 U6361 ( .A1(n6810), .A2(n6714), .ZN(n5592) );
  NOR2_X1 U6362 ( .A1(n4480), .A2(n6582), .ZN(n6809) );
  NOR2_X1 U6363 ( .A1(n6717), .A2(n6902), .ZN(n5590) );
  AOI211_X1 U6364 ( .C1(n6707), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6809), 
        .B(n5590), .ZN(n5591) );
  OAI211_X1 U6365 ( .C1(n6121), .C2(n6890), .A(n5592), .B(n5591), .ZN(U2979)
         );
  NAND2_X1 U6366 ( .A1(n5593), .A2(n6714), .ZN(n5597) );
  AND2_X1 U6367 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5594)
         );
  AOI211_X1 U6368 ( .C1(n6693), .C2(n6917), .A(n5595), .B(n5594), .ZN(n5596)
         );
  OAI211_X1 U6369 ( .C1(n6121), .C2(n6919), .A(n5597), .B(n5596), .ZN(U2976)
         );
  NOR3_X1 U6370 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5598), .A3(n6779), 
        .ZN(n5605) );
  OAI21_X1 U6371 ( .B1(n6793), .B2(n5600), .A(n5599), .ZN(n5604) );
  INV_X1 U6372 ( .A(n6779), .ZN(n5601) );
  OAI21_X1 U6373 ( .B1(n6754), .B2(n5601), .A(n6778), .ZN(n6785) );
  NOR4_X1 U6374 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6790), .A3(n6779), 
        .A4(n6794), .ZN(n6786) );
  NOR2_X1 U6375 ( .A1(n6798), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6783)
         );
  NOR3_X1 U6376 ( .A1(n6785), .A2(n6786), .A3(n6783), .ZN(n5602) );
  NOR2_X1 U6377 ( .A1(n5602), .A2(n4427), .ZN(n5603) );
  AOI211_X1 U6378 ( .C1(n6774), .C2(n5605), .A(n5604), .B(n5603), .ZN(n5606)
         );
  OAI21_X1 U6379 ( .B1(n6800), .B2(n5607), .A(n5606), .ZN(U3012) );
  AOI21_X1 U6380 ( .B1(n5609), .B2(n5488), .A(n5608), .ZN(n6931) );
  INV_X1 U6381 ( .A(n6931), .ZN(n5613) );
  OAI222_X1 U6382 ( .A1(n5613), .A2(n7100), .B1(n6027), .B2(n5610), .C1(n6026), 
        .C2(n3945), .ZN(U2879) );
  XOR2_X1 U6383 ( .A(n5627), .B(n5628), .Z(n6929) );
  INV_X1 U6384 ( .A(n6929), .ZN(n5612) );
  OAI222_X1 U6385 ( .A1(n5613), .A2(n6005), .B1(n6658), .B2(n5612), .C1(n5611), 
        .C2(n6663), .ZN(U2847) );
  XOR2_X1 U6386 ( .A(n5615), .B(n5614), .Z(n5663) );
  NOR3_X1 U6387 ( .A1(n6855), .A2(n5622), .A3(n5631), .ZN(n5617) );
  OAI211_X1 U6388 ( .C1(n5618), .C2(n5617), .A(n5671), .B(n5616), .ZN(n5623)
         );
  INV_X1 U6389 ( .A(n5623), .ZN(n5625) );
  INV_X1 U6390 ( .A(n5619), .ZN(n5620) );
  AOI21_X1 U6391 ( .B1(n5669), .B2(n5621), .A(n5620), .ZN(n6831) );
  NAND2_X1 U6392 ( .A1(n5622), .A2(n6798), .ZN(n6856) );
  INV_X1 U6393 ( .A(n5671), .ZN(n5630) );
  AOI22_X1 U6394 ( .A1(n6858), .A2(n5704), .B1(n6856), .B2(n5630), .ZN(n5624)
         );
  NAND3_X1 U6395 ( .A1(n6831), .A2(n5624), .A3(n5623), .ZN(n5645) );
  OAI21_X1 U6396 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5625), .A(n5645), 
        .ZN(n5636) );
  OAI21_X1 U6397 ( .B1(n5628), .B2(n5627), .A(n5626), .ZN(n5629) );
  AND2_X1 U6398 ( .A1(n5629), .A2(n5650), .ZN(n6943) );
  NOR2_X1 U6399 ( .A1(n4480), .A2(n6949), .ZN(n5634) );
  NOR4_X1 U6400 ( .A1(n5632), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n5631), 
        .A4(n5630), .ZN(n5633) );
  AOI211_X1 U6401 ( .C1(n6860), .C2(n6943), .A(n5634), .B(n5633), .ZN(n5635)
         );
  OAI211_X1 U6402 ( .C1(n5663), .C2(n6800), .A(n5636), .B(n5635), .ZN(U3005)
         );
  OAI21_X1 U6403 ( .B1(n6830), .B2(n6106), .A(n5637), .ZN(n5639) );
  AOI21_X1 U6404 ( .B1(n4460), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5638), 
        .ZN(n5666) );
  XOR2_X1 U6405 ( .A(n5639), .B(n5666), .Z(n6827) );
  NAND2_X1 U6406 ( .A1(n6827), .A2(n6714), .ZN(n5643) );
  NOR2_X1 U6407 ( .A1(n4480), .A2(n6588), .ZN(n6824) );
  NOR2_X1 U6408 ( .A1(n6717), .A2(n5640), .ZN(n5641) );
  AOI211_X1 U6409 ( .C1(n6707), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6824), 
        .B(n5641), .ZN(n5642) );
  OAI211_X1 U6410 ( .C1(n6121), .C2(n5644), .A(n5643), .B(n5642), .ZN(U2975)
         );
  INV_X1 U6411 ( .A(n5645), .ZN(n5656) );
  OAI21_X1 U6412 ( .B1(n5648), .B2(n5647), .A(n5646), .ZN(n5676) );
  NAND2_X1 U6413 ( .A1(n5676), .A2(n6854), .ZN(n5655) );
  NOR2_X1 U6414 ( .A1(n6842), .A2(n5704), .ZN(n5653) );
  AND2_X1 U6415 ( .A1(n5650), .A2(n5649), .ZN(n5651) );
  OR2_X1 U6416 ( .A1(n5651), .A2(n5706), .ZN(n5693) );
  OAI22_X1 U6417 ( .A1(n6793), .A2(n5693), .B1(n6592), .B2(n4480), .ZN(n5652)
         );
  AOI21_X1 U6418 ( .B1(n5653), .B2(n5703), .A(n5652), .ZN(n5654) );
  OAI211_X1 U6419 ( .C1(n5703), .C2(n5656), .A(n5655), .B(n5654), .ZN(U3004)
         );
  XOR2_X1 U6420 ( .A(n5658), .B(n5657), .Z(n6938) );
  INV_X1 U6421 ( .A(n6938), .ZN(n5697) );
  AOI22_X1 U6422 ( .A1(n6649), .A2(n6943), .B1(EBX_REG_13__SCAN_IN), .B2(n5970), .ZN(n5659) );
  OAI21_X1 U6423 ( .B1(n5697), .B2(n6001), .A(n5659), .ZN(U2846) );
  AOI22_X1 U6424 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6771), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5660) );
  OAI21_X1 U6425 ( .B1(n6717), .B2(n6936), .A(n5660), .ZN(n5661) );
  AOI21_X1 U6426 ( .B1(n6938), .B2(n6713), .A(n5661), .ZN(n5662) );
  OAI21_X1 U6427 ( .B1(n5663), .B2(n6696), .A(n5662), .ZN(U2973) );
  NAND2_X1 U6428 ( .A1(n6106), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5665) );
  NAND3_X1 U6429 ( .A1(n5666), .A2(n4460), .A3(n6830), .ZN(n5664) );
  OAI21_X1 U6430 ( .B1(n5666), .B2(n5665), .A(n5664), .ZN(n5667) );
  XOR2_X1 U6431 ( .A(n4457), .B(n5667), .Z(n6697) );
  AOI22_X1 U6432 ( .A1(n6860), .A2(n6929), .B1(n6771), .B2(
        REIP_REG_12__SCAN_IN), .ZN(n5675) );
  NOR2_X1 U6433 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  OAI21_X1 U6434 ( .B1(n5671), .B2(n5670), .A(n6831), .ZN(n5673) );
  OAI21_X1 U6435 ( .B1(n6842), .B2(n6830), .A(n4457), .ZN(n5672) );
  NAND2_X1 U6436 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  OAI211_X1 U6437 ( .C1(n6697), .C2(n6800), .A(n5675), .B(n5674), .ZN(U3006)
         );
  INV_X1 U6438 ( .A(n5676), .ZN(n5682) );
  XOR2_X1 U6439 ( .A(n5678), .B(n5677), .Z(n5683) );
  AOI22_X1 U6440 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6771), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5679) );
  OAI21_X1 U6441 ( .B1(n6717), .B2(n5684), .A(n5679), .ZN(n5680) );
  AOI21_X1 U6442 ( .B1(n5683), .B2(n6713), .A(n5680), .ZN(n5681) );
  OAI21_X1 U6443 ( .B1(n5682), .B2(n6696), .A(n5681), .ZN(U2972) );
  INV_X1 U6444 ( .A(n5683), .ZN(n5696) );
  INV_X1 U6445 ( .A(n5684), .ZN(n5691) );
  NAND4_X1 U6446 ( .A1(REIP_REG_12__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n6953), .A4(n6592), .ZN(n5686) );
  OAI21_X1 U6447 ( .B1(n5693), .B2(n7004), .A(n5686), .ZN(n5690) );
  AOI21_X1 U6448 ( .B1(n5721), .B2(n6940), .A(n6941), .ZN(n5741) );
  AOI22_X1 U6449 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6968), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5741), .ZN(n5687) );
  OAI211_X1 U6450 ( .C1(n6914), .C2(n5688), .A(n5687), .B(n6944), .ZN(n5689)
         );
  AOI211_X1 U6451 ( .C1(n6981), .C2(n5691), .A(n5690), .B(n5689), .ZN(n5692)
         );
  OAI21_X1 U6452 ( .B1(n5696), .B2(n6978), .A(n5692), .ZN(U2813) );
  INV_X1 U6453 ( .A(n5693), .ZN(n5694) );
  AOI22_X1 U6454 ( .A1(n6649), .A2(n5694), .B1(n5970), .B2(EBX_REG_14__SCAN_IN), .ZN(n5695) );
  OAI21_X1 U6455 ( .B1(n5696), .B2(n6001), .A(n5695), .ZN(U2845) );
  INV_X1 U6456 ( .A(DATAI_14_), .ZN(n6364) );
  INV_X1 U6457 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6568) );
  OAI222_X1 U6458 ( .A1(n5696), .A2(n7100), .B1(n6027), .B2(n6364), .C1(n6026), 
        .C2(n6568), .ZN(U2877) );
  INV_X1 U6459 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6566) );
  INV_X1 U6460 ( .A(DATAI_13_), .ZN(n6465) );
  OAI222_X1 U6461 ( .A1(n6026), .A2(n6566), .B1(n6027), .B2(n6465), .C1(n7100), 
        .C2(n5697), .ZN(U2878) );
  OAI21_X1 U6462 ( .B1(n5698), .B2(n5700), .A(n5699), .ZN(n5701) );
  INV_X1 U6463 ( .A(n5701), .ZN(n5718) );
  OAI21_X1 U6464 ( .B1(n6754), .B2(n5702), .A(n6831), .ZN(n6834) );
  NOR3_X1 U6465 ( .A1(n6842), .A2(n5704), .A3(n5703), .ZN(n6836) );
  AOI22_X1 U6466 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6834), .B1(n6836), .B2(n6837), .ZN(n5709) );
  OAI21_X1 U6467 ( .B1(n5706), .B2(n5705), .A(n5956), .ZN(n6003) );
  INV_X1 U6468 ( .A(n6003), .ZN(n5720) );
  INV_X1 U6469 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5707) );
  NOR2_X1 U6470 ( .A1(n4480), .A2(n5707), .ZN(n5711) );
  AOI21_X1 U6471 ( .B1(n6860), .B2(n5720), .A(n5711), .ZN(n5708) );
  OAI211_X1 U6472 ( .C1(n5718), .C2(n6800), .A(n5709), .B(n5708), .ZN(U3003)
         );
  AND2_X1 U6473 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5710)
         );
  AOI211_X1 U6474 ( .C1(n6693), .C2(n5727), .A(n5711), .B(n5710), .ZN(n5717)
         );
  INV_X1 U6475 ( .A(n5712), .ZN(n5713) );
  AOI21_X1 U6476 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5719) );
  NAND2_X1 U6477 ( .A1(n5719), .A2(n6713), .ZN(n5716) );
  OAI211_X1 U6478 ( .C1(n5718), .C2(n6696), .A(n5717), .B(n5716), .ZN(U2971)
         );
  INV_X1 U6479 ( .A(n5719), .ZN(n6028) );
  AOI22_X1 U6480 ( .A1(n6993), .A2(n5720), .B1(REIP_REG_15__SCAN_IN), .B2(
        n5741), .ZN(n5724) );
  INV_X1 U6481 ( .A(n5721), .ZN(n5722) );
  INV_X1 U6482 ( .A(n6953), .ZN(n6942) );
  NOR3_X1 U6483 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5722), .A3(n6942), .ZN(n5742) );
  AOI211_X1 U6484 ( .C1(n7003), .C2(EBX_REG_15__SCAN_IN), .A(n6967), .B(n5742), 
        .ZN(n5723) );
  OAI211_X1 U6485 ( .C1(n5725), .C2(n6999), .A(n5724), .B(n5723), .ZN(n5726)
         );
  AOI21_X1 U6486 ( .B1(n5727), .B2(n6981), .A(n5726), .ZN(n5728) );
  OAI21_X1 U6487 ( .B1(n6028), .B2(n6978), .A(n5728), .ZN(U2812) );
  AND2_X1 U6488 ( .A1(n5712), .A2(n5729), .ZN(n5731) );
  OR2_X1 U6489 ( .A1(n5731), .A2(n5730), .ZN(n6120) );
  XNOR2_X1 U6490 ( .A(n5956), .B(n5952), .ZN(n6833) );
  AOI22_X1 U6491 ( .A1(n6833), .A2(n6649), .B1(n5970), .B2(EBX_REG_16__SCAN_IN), .ZN(n5732) );
  OAI21_X1 U6492 ( .B1(n6120), .B2(n6001), .A(n5732), .ZN(U2843) );
  NOR2_X2 U6493 ( .A1(n7116), .A2(n5733), .ZN(n7113) );
  AOI22_X1 U6494 ( .A1(n7113), .A2(DATAI_16_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n7116), .ZN(n5737) );
  AND2_X1 U6495 ( .A1(n5734), .A2(n3700), .ZN(n5735) );
  NAND2_X1 U6496 ( .A1(n7117), .A2(DATAI_0_), .ZN(n5736) );
  OAI211_X1 U6497 ( .C1(n6120), .C2(n7100), .A(n5737), .B(n5736), .ZN(U2875)
         );
  OR2_X1 U6498 ( .A1(n5738), .A2(n6942), .ZN(n5950) );
  AOI22_X1 U6499 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6968), .B1(
        EBX_REG_16__SCAN_IN), .B2(n7003), .ZN(n5739) );
  OAI211_X1 U6500 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5950), .A(n5739), .B(n6944), .ZN(n5740) );
  AOI221_X1 U6501 ( .B1(n5742), .B2(REIP_REG_16__SCAN_IN), .C1(n5741), .C2(
        REIP_REG_16__SCAN_IN), .A(n5740), .ZN(n5745) );
  INV_X1 U6502 ( .A(n6116), .ZN(n5743) );
  AOI22_X1 U6503 ( .A1(n6981), .A2(n5743), .B1(n6993), .B2(n6833), .ZN(n5744)
         );
  OAI211_X1 U6504 ( .C1(n6120), .C2(n6978), .A(n5745), .B(n5744), .ZN(U2811)
         );
  AOI22_X1 U6505 ( .A1(n7113), .A2(DATAI_22_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n7116), .ZN(n5747) );
  NAND2_X1 U6506 ( .A1(n7117), .A2(DATAI_6_), .ZN(n5746) );
  OAI211_X1 U6507 ( .C1(n5759), .C2(n7100), .A(n5747), .B(n5746), .ZN(U2869)
         );
  INV_X1 U6508 ( .A(n6198), .ZN(n5980) );
  XNOR2_X1 U6509 ( .A(n5980), .B(n5979), .ZN(n6187) );
  INV_X1 U6510 ( .A(n6187), .ZN(n5748) );
  AOI22_X1 U6511 ( .A1(n5748), .A2(n6649), .B1(n5970), .B2(EBX_REG_22__SCAN_IN), .ZN(n5749) );
  OAI21_X1 U6512 ( .B1(n5759), .B2(n6001), .A(n5749), .ZN(U2837) );
  NOR3_X1 U6513 ( .A1(n6986), .A2(REIP_REG_22__SCAN_IN), .A3(n5750), .ZN(n5751) );
  AOI21_X1 U6514 ( .B1(n6968), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n5751), 
        .ZN(n5752) );
  OAI21_X1 U6515 ( .B1(n6187), .B2(n7004), .A(n5752), .ZN(n5756) );
  INV_X1 U6516 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6601) );
  OAI21_X1 U6517 ( .B1(n6986), .B2(n6988), .A(n5826), .ZN(n6991) );
  AOI21_X1 U6518 ( .B1(n6998), .B2(n6601), .A(n6991), .ZN(n5754) );
  OAI22_X1 U6519 ( .A1(n5754), .A2(n6604), .B1(n5753), .B2(n6914), .ZN(n5755)
         );
  AOI211_X1 U6520 ( .C1(n6981), .C2(n5757), .A(n5756), .B(n5755), .ZN(n5758)
         );
  OAI21_X1 U6521 ( .B1(n5759), .B2(n6978), .A(n5758), .ZN(U2805) );
  AOI22_X1 U6522 ( .A1(n5761), .A2(n7055), .B1(n7069), .B2(n5760), .ZN(n5763)
         );
  MUX2_X1 U6523 ( .A(n5763), .B(n5762), .S(n5807), .Z(n5764) );
  INV_X1 U6524 ( .A(n5764), .ZN(U3456) );
  INV_X1 U6525 ( .A(n5765), .ZN(n5768) );
  AOI21_X1 U6526 ( .B1(n7069), .B2(n5768), .A(n5807), .ZN(n5773) );
  NOR3_X1 U6527 ( .A1(n7062), .A2(n6855), .A3(n5766), .ZN(n5770) );
  NOR3_X1 U6528 ( .A1(n5768), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5767), 
        .ZN(n5769) );
  AOI211_X1 U6529 ( .C1(n5771), .C2(n7055), .A(n5770), .B(n5769), .ZN(n5772)
         );
  OAI22_X1 U6530 ( .A1(n5773), .A2(n3739), .B1(n5807), .B2(n5772), .ZN(U3459)
         );
  NOR2_X1 U6531 ( .A1(n6106), .A2(n6051), .ZN(n6042) );
  NOR2_X1 U6532 ( .A1(n4640), .A2(n4637), .ZN(n5774) );
  NAND2_X1 U6533 ( .A1(n6034), .A2(n5775), .ZN(n5777) );
  XNOR2_X1 U6534 ( .A(n5777), .B(n3458), .ZN(n5791) );
  NAND2_X1 U6535 ( .A1(n6771), .A2(REIP_REG_28__SCAN_IN), .ZN(n5786) );
  OAI21_X1 U6536 ( .B1(n6101), .B2(n5891), .A(n5786), .ZN(n5782) );
  AND2_X2 U6537 ( .A1(n5917), .A2(n5778), .ZN(n5906) );
  OAI21_X4 U6538 ( .B1(n5906), .B2(n5780), .A(n5779), .ZN(n5889) );
  NOR2_X1 U6539 ( .A1(n5889), .A2(n6121), .ZN(n5781) );
  OAI21_X1 U6540 ( .B1(n5791), .B2(n6696), .A(n5783), .ZN(U2958) );
  AND2_X1 U6541 ( .A1(n5904), .A2(n5784), .ZN(n5785) );
  OR2_X1 U6542 ( .A1(n5785), .A2(n5819), .ZN(n5967) );
  OAI21_X1 U6543 ( .B1(n5967), .B2(n6793), .A(n5786), .ZN(n5787) );
  AOI21_X1 U6544 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n6145), .A(n5787), 
        .ZN(n5790) );
  INV_X1 U6545 ( .A(n6134), .ZN(n6146) );
  OAI211_X1 U6546 ( .C1(INSTADDRPOINTER_REG_28__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6146), .B(n5788), .ZN(n5789) );
  OAI211_X1 U6547 ( .C1(n5791), .C2(n6800), .A(n5790), .B(n5789), .ZN(U2990)
         );
  INV_X1 U6548 ( .A(n7058), .ZN(n5792) );
  NOR2_X1 U6549 ( .A1(n5793), .A2(n5792), .ZN(n7074) );
  NOR2_X1 U6550 ( .A1(n5797), .A2(n7020), .ZN(n5796) );
  NOR2_X1 U6551 ( .A1(n5794), .A2(n4386), .ZN(n5795) );
  AOI211_X1 U6552 ( .C1(n7074), .C2(n5797), .A(n5796), .B(n5795), .ZN(n5798)
         );
  OAI21_X1 U6553 ( .B1(n5800), .B2(n5799), .A(n5798), .ZN(U3465) );
  AOI21_X1 U6554 ( .B1(n5801), .B2(n5779), .A(n5868), .ZN(n5964) );
  AOI21_X1 U6555 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5802), 
        .ZN(n5803) );
  OAI21_X1 U6556 ( .B1(n5884), .B2(n6717), .A(n5803), .ZN(n5804) );
  AOI21_X1 U6557 ( .B1(n5964), .B2(n6713), .A(n5804), .ZN(n5805) );
  OAI21_X1 U6558 ( .B1(n5806), .B2(n6696), .A(n5805), .ZN(U2957) );
  INV_X1 U6559 ( .A(n5807), .ZN(n7018) );
  INV_X1 U6560 ( .A(n5808), .ZN(n5810) );
  AOI22_X1 U6561 ( .A1(n5811), .A2(n5810), .B1(n5809), .B2(n5818), .ZN(n7019)
         );
  INV_X1 U6562 ( .A(n7055), .ZN(n5813) );
  AOI22_X1 U6563 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6855), .B1(n5818), .B2(
        n7069), .ZN(n5812) );
  OAI21_X1 U6564 ( .B1(n7019), .B2(n5813), .A(n5812), .ZN(n5816) );
  INV_X1 U6565 ( .A(n5814), .ZN(n5815) );
  NOR2_X1 U6566 ( .A1(n5815), .A2(n5818), .ZN(n7021) );
  AOI22_X1 U6567 ( .A1(n7018), .A2(n5816), .B1(n7055), .B2(n7021), .ZN(n5817)
         );
  OAI21_X1 U6568 ( .B1(n5818), .B2(n7018), .A(n5817), .ZN(U3461) );
  AOI22_X1 U6569 ( .A1(n5858), .A2(n4268), .B1(n5820), .B2(n5819), .ZN(n5821)
         );
  OAI22_X1 U6570 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        EBX_REG_30__SCAN_IN), .B2(n5861), .ZN(n5860) );
  XNOR2_X1 U6571 ( .A(n5821), .B(n5860), .ZN(n6136) );
  INV_X1 U6572 ( .A(n6136), .ZN(n5837) );
  INV_X1 U6573 ( .A(n5822), .ZN(n5835) );
  NOR2_X1 U6574 ( .A1(n6608), .A2(n5823), .ZN(n5924) );
  NAND3_X1 U6575 ( .A1(REIP_REG_26__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        n5924), .ZN(n5909) );
  INV_X1 U6576 ( .A(n5909), .ZN(n5825) );
  NAND2_X1 U6577 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5825), .ZN(n5824) );
  NOR2_X1 U6578 ( .A1(n6986), .A2(n5824), .ZN(n5894) );
  NAND2_X1 U6579 ( .A1(n5894), .A2(REIP_REG_28__SCAN_IN), .ZN(n5883) );
  NOR2_X1 U6580 ( .A1(n5883), .A2(n6332), .ZN(n5832) );
  INV_X1 U6581 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6622) );
  NOR2_X1 U6582 ( .A1(n6622), .A2(n6332), .ZN(n5831) );
  AND2_X1 U6583 ( .A1(n5826), .A2(n5825), .ZN(n5827) );
  OR2_X1 U6584 ( .A1(n6941), .A2(n5827), .ZN(n5908) );
  INV_X1 U6585 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6615) );
  INV_X1 U6586 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U6587 ( .A1(n6615), .A2(n6613), .ZN(n5828) );
  OR2_X1 U6588 ( .A1(n6941), .A2(n5828), .ZN(n5829) );
  NAND2_X1 U6589 ( .A1(n5908), .A2(n5829), .ZN(n5893) );
  INV_X1 U6590 ( .A(n5893), .ZN(n5830) );
  OAI21_X1 U6591 ( .B1(n5831), .B2(n6986), .A(n5830), .ZN(n5877) );
  OAI21_X1 U6592 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5832), .A(n5877), .ZN(n5834) );
  AOI22_X1 U6593 ( .A1(n7003), .A2(EBX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6968), .ZN(n5833) );
  OAI211_X1 U6594 ( .C1(n7010), .C2(n5835), .A(n5834), .B(n5833), .ZN(n5836)
         );
  AOI21_X1 U6595 ( .B1(n5837), .B2(n6993), .A(n5836), .ZN(n5838) );
  OAI21_X1 U6596 ( .B1(n5841), .B2(n6978), .A(n5838), .ZN(U2797) );
  AOI22_X1 U6597 ( .A1(n7113), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n7116), .ZN(n5840) );
  NAND2_X1 U6598 ( .A1(n7117), .A2(DATAI_14_), .ZN(n5839) );
  OAI211_X1 U6599 ( .C1(n5841), .C2(n7100), .A(n5840), .B(n5839), .ZN(U2861)
         );
  INV_X1 U6600 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5842) );
  OAI222_X1 U6601 ( .A1(n5842), .A2(n6663), .B1(n6658), .B2(n6136), .C1(n6005), 
        .C2(n5841), .ZN(U2829) );
  INV_X1 U6602 ( .A(n5843), .ZN(n5844) );
  OR2_X1 U6603 ( .A1(n5854), .A2(n5844), .ZN(n5848) );
  NAND2_X1 U6604 ( .A1(n5845), .A2(n4254), .ZN(n5846) );
  NAND2_X1 U6605 ( .A1(n5854), .A2(n5846), .ZN(n5847) );
  OAI211_X1 U6606 ( .C1(n5849), .C2(n4258), .A(n5848), .B(n5847), .ZN(n7035)
         );
  INV_X1 U6607 ( .A(n5849), .ZN(n5850) );
  OAI21_X1 U6608 ( .B1(n5850), .B2(n4258), .A(n4254), .ZN(n5851) );
  INV_X1 U6609 ( .A(n5851), .ZN(n5852) );
  AOI21_X1 U6610 ( .B1(n5854), .B2(n5853), .A(n5852), .ZN(n6718) );
  OR2_X1 U6611 ( .A1(n5856), .A2(n5855), .ZN(n6727) );
  NAND2_X1 U6612 ( .A1(n6727), .A2(n6733), .ZN(n5857) );
  NAND2_X1 U6613 ( .A1(n5857), .A2(n7088), .ZN(n6743) );
  AND2_X1 U6614 ( .A1(n6718), .A2(n6743), .ZN(n7039) );
  NOR2_X1 U6615 ( .A1(n7039), .A2(n7077), .ZN(n7012) );
  MUX2_X1 U6616 ( .A(MORE_REG_SCAN_IN), .B(n7035), .S(n7012), .Z(U3471) );
  MUX2_X1 U6617 ( .A(n5860), .B(n5859), .S(n5858), .Z(n5864) );
  OAI22_X1 U6618 ( .A1(n5862), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5861), .ZN(n5863) );
  XNOR2_X2 U6619 ( .A(n5864), .B(n5863), .ZN(n6124) );
  AOI22_X1 U6620 ( .A1(n5866), .A2(EAX_REG_31__SCAN_IN), .B1(n5865), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5870) );
  NAND2_X1 U6621 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  XOR2_X1 U6622 ( .A(n5869), .B(n5870), .Z(n6040) );
  NAND2_X1 U6623 ( .A1(n6040), .A2(n7007), .ZN(n5879) );
  INV_X1 U6624 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6036) );
  NAND3_X1 U6625 ( .A1(REIP_REG_29__SCAN_IN), .A2(REIP_REG_30__SCAN_IN), .A3(
        n6036), .ZN(n5875) );
  NAND3_X1 U6626 ( .A1(n5872), .A2(EBX_REG_31__SCAN_IN), .A3(n5871), .ZN(n5874) );
  NAND2_X1 U6627 ( .A1(n6968), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5873)
         );
  OAI211_X1 U6628 ( .C1(n5883), .C2(n5875), .A(n5874), .B(n5873), .ZN(n5876)
         );
  AOI21_X1 U6629 ( .B1(n5877), .B2(REIP_REG_31__SCAN_IN), .A(n5876), .ZN(n5878) );
  OAI211_X1 U6630 ( .C1(n6124), .C2(n7004), .A(n5879), .B(n5878), .ZN(U2796)
         );
  NAND2_X1 U6631 ( .A1(n5964), .A2(n7007), .ZN(n5888) );
  NOR2_X1 U6632 ( .A1(n6999), .A2(n5880), .ZN(n5881) );
  AOI21_X1 U6633 ( .B1(n7003), .B2(EBX_REG_29__SCAN_IN), .A(n5881), .ZN(n5882)
         );
  OAI21_X1 U6634 ( .B1(n5883), .B2(REIP_REG_29__SCAN_IN), .A(n5882), .ZN(n5886) );
  NOR2_X1 U6635 ( .A1(n7010), .A2(n5884), .ZN(n5885) );
  AOI211_X1 U6636 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5893), .A(n5886), .B(n5885), .ZN(n5887) );
  OAI211_X1 U6637 ( .C1(n7004), .C2(n5965), .A(n5888), .B(n5887), .ZN(U2798)
         );
  INV_X1 U6638 ( .A(n5967), .ZN(n5900) );
  NAND2_X1 U6639 ( .A1(n6981), .A2(n5890), .ZN(n5898) );
  NOR2_X1 U6640 ( .A1(n6999), .A2(n5891), .ZN(n5892) );
  AOI21_X1 U6641 ( .B1(n7003), .B2(EBX_REG_28__SCAN_IN), .A(n5892), .ZN(n5897)
         );
  NAND2_X1 U6642 ( .A1(n5893), .A2(REIP_REG_28__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U6643 ( .A1(n5894), .A2(n6615), .ZN(n5895) );
  NAND4_X1 U6644 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n5899)
         );
  AOI21_X1 U6645 ( .B1(n5900), .B2(n6993), .A(n5899), .ZN(n5901) );
  OAI21_X1 U6646 ( .B1(n5889), .B2(n6978), .A(n5901), .ZN(U2799) );
  NAND2_X1 U6647 ( .A1(n5922), .A2(n5902), .ZN(n5903) );
  NAND2_X1 U6648 ( .A1(n5904), .A2(n5903), .ZN(n6142) );
  NAND2_X1 U6649 ( .A1(n5917), .A2(n5905), .ZN(n5918) );
  NAND2_X1 U6650 ( .A1(n6049), .A2(n7007), .ZN(n5915) );
  INV_X1 U6651 ( .A(n5908), .ZN(n5925) );
  INV_X1 U6652 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5969) );
  NOR3_X1 U6653 ( .A1(n6986), .A2(REIP_REG_27__SCAN_IN), .A3(n5909), .ZN(n5910) );
  AOI21_X1 U6654 ( .B1(n6968), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5910), 
        .ZN(n5911) );
  OAI21_X1 U6655 ( .B1(n6914), .B2(n5969), .A(n5911), .ZN(n5913) );
  NOR2_X1 U6656 ( .A1(n7010), .A2(n6047), .ZN(n5912) );
  AOI211_X1 U6657 ( .C1(n5925), .C2(REIP_REG_27__SCAN_IN), .A(n5913), .B(n5912), .ZN(n5914) );
  OAI211_X1 U6658 ( .C1(n7004), .C2(n6142), .A(n5915), .B(n5914), .ZN(U2800)
         );
  NAND2_X1 U6659 ( .A1(n5938), .A2(n5920), .ZN(n5921) );
  AND2_X1 U6660 ( .A1(n5922), .A2(n5921), .ZN(n6154) );
  INV_X1 U6661 ( .A(n5923), .ZN(n6056) );
  AOI22_X1 U6662 ( .A1(n7003), .A2(EBX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6968), .ZN(n5928) );
  NAND2_X1 U6663 ( .A1(n6998), .A2(n5924), .ZN(n5934) );
  INV_X1 U6664 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U6665 ( .A1(n5934), .A2(n6610), .ZN(n5926) );
  OAI21_X1 U6666 ( .B1(n5926), .B2(REIP_REG_26__SCAN_IN), .A(n5925), .ZN(n5927) );
  OAI211_X1 U6667 ( .C1(n7010), .C2(n6056), .A(n5928), .B(n5927), .ZN(n5929)
         );
  AOI21_X1 U6668 ( .B1(n6154), .B2(n6993), .A(n5929), .ZN(n5930) );
  OAI21_X1 U6669 ( .B1(n6054), .B2(n6978), .A(n5930), .ZN(U2801) );
  AOI21_X1 U6670 ( .B1(n5933), .B2(n5932), .A(n5931), .ZN(n6067) );
  INV_X1 U6671 ( .A(n6067), .ZN(n6021) );
  INV_X1 U6672 ( .A(n6065), .ZN(n5944) );
  OAI22_X1 U6673 ( .A1(REIP_REG_25__SCAN_IN), .A2(n5934), .B1(n4536), .B2(
        n6999), .ZN(n5943) );
  OR2_X1 U6674 ( .A1(n5936), .A2(n5935), .ZN(n5937) );
  NAND2_X1 U6675 ( .A1(n5938), .A2(n5937), .ZN(n6162) );
  AOI21_X1 U6676 ( .B1(n7000), .B2(n5939), .A(n6610), .ZN(n5940) );
  AOI21_X1 U6677 ( .B1(n7003), .B2(EBX_REG_25__SCAN_IN), .A(n5940), .ZN(n5941)
         );
  OAI21_X1 U6678 ( .B1(n6162), .B2(n7004), .A(n5941), .ZN(n5942) );
  AOI211_X1 U6679 ( .C1(n6981), .C2(n5944), .A(n5943), .B(n5942), .ZN(n5945)
         );
  OAI21_X1 U6680 ( .B1(n6021), .B2(n6978), .A(n5945), .ZN(U2802) );
  OR2_X1 U6681 ( .A1(n5730), .A2(n5948), .ZN(n5949) );
  AND2_X1 U6682 ( .A1(n5947), .A2(n5949), .ZN(n7101) );
  INV_X1 U6683 ( .A(n7101), .ZN(n6000) );
  OAI21_X1 U6684 ( .B1(n6594), .B2(n5950), .A(n6843), .ZN(n5961) );
  AOI21_X1 U6685 ( .B1(n6954), .B2(n6940), .A(n6941), .ZN(n6962) );
  INV_X1 U6686 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5951) );
  OAI22_X1 U6687 ( .A1(n5951), .A2(n6999), .B1(n6706), .B2(n7010), .ZN(n5960)
         );
  INV_X1 U6688 ( .A(n5952), .ZN(n5955) );
  INV_X1 U6689 ( .A(n5953), .ZN(n5954) );
  OAI21_X1 U6690 ( .B1(n5956), .B2(n5955), .A(n5954), .ZN(n5957) );
  NAND2_X1 U6691 ( .A1(n5957), .A2(n5995), .ZN(n6847) );
  AOI21_X1 U6692 ( .B1(n7003), .B2(EBX_REG_17__SCAN_IN), .A(n6967), .ZN(n5958)
         );
  OAI21_X1 U6693 ( .B1(n7004), .B2(n6847), .A(n5958), .ZN(n5959) );
  AOI211_X1 U6694 ( .C1(n5961), .C2(n6962), .A(n5960), .B(n5959), .ZN(n5962)
         );
  OAI21_X1 U6695 ( .B1(n6000), .B2(n6978), .A(n5962), .ZN(U2810) );
  OAI22_X1 U6696 ( .A1(n6124), .A2(n6658), .B1(n5963), .B2(n6663), .ZN(U2828)
         );
  INV_X1 U6697 ( .A(n5964), .ZN(n6011) );
  OAI222_X1 U6698 ( .A1(n5966), .A2(n6663), .B1(n6658), .B2(n5965), .C1(n6011), 
        .C2(n6005), .ZN(U2830) );
  OAI222_X1 U6699 ( .A1(n5968), .A2(n6663), .B1(n6658), .B2(n5967), .C1(n5889), 
        .C2(n6005), .ZN(U2831) );
  INV_X1 U6700 ( .A(n6049), .ZN(n6016) );
  OAI222_X1 U6701 ( .A1(n5969), .A2(n6663), .B1(n6658), .B2(n6142), .C1(n6016), 
        .C2(n6005), .ZN(U2832) );
  AOI22_X1 U6702 ( .A1(n6154), .A2(n6649), .B1(n5970), .B2(EBX_REG_26__SCAN_IN), .ZN(n5971) );
  OAI21_X1 U6703 ( .B1(n6054), .B2(n6001), .A(n5971), .ZN(U2833) );
  INV_X1 U6704 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5972) );
  OAI222_X1 U6705 ( .A1(n6162), .A2(n6658), .B1(n5972), .B2(n6663), .C1(n6021), 
        .C2(n6005), .ZN(U2834) );
  OAI222_X1 U6706 ( .A1(n6168), .A2(n6658), .B1(n6663), .B2(n4349), .C1(n6005), 
        .C2(n6073), .ZN(U2835) );
  INV_X1 U6707 ( .A(n7115), .ZN(n5984) );
  INV_X1 U6708 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5983) );
  AOI21_X1 U6709 ( .B1(n5980), .B2(n5979), .A(n5978), .ZN(n5982) );
  OR2_X1 U6710 ( .A1(n5982), .A2(n5981), .ZN(n7005) );
  OAI222_X1 U6711 ( .A1(n5984), .A2(n6005), .B1(n6663), .B2(n5983), .C1(n7005), 
        .C2(n6658), .ZN(U2836) );
  OR2_X1 U6712 ( .A1(n6657), .A2(n5985), .ZN(n5986) );
  NAND2_X1 U6713 ( .A1(n6196), .A2(n5986), .ZN(n6977) );
  AOI21_X1 U6715 ( .B1(n5990), .B2(n5987), .A(n5989), .ZN(n6103) );
  INV_X1 U6716 ( .A(n6103), .ZN(n6979) );
  OAI222_X1 U6717 ( .A1(n6658), .A2(n6977), .B1(n6663), .B2(n4333), .C1(n6979), 
        .C2(n6005), .ZN(U2839) );
  AOI21_X1 U6718 ( .B1(n5993), .B2(n5947), .A(n3441), .ZN(n7104) );
  AND2_X1 U6719 ( .A1(n5995), .A2(n5994), .ZN(n5996) );
  OR2_X1 U6720 ( .A1(n5996), .A2(n6655), .ZN(n6960) );
  OAI22_X1 U6721 ( .A1(n6960), .A2(n6658), .B1(n5997), .B2(n6663), .ZN(n5998)
         );
  AOI21_X1 U6722 ( .B1(n7104), .B2(n6660), .A(n5998), .ZN(n5999) );
  INV_X1 U6723 ( .A(n5999), .ZN(U2841) );
  INV_X1 U6724 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6002) );
  OAI222_X1 U6725 ( .A1(n6847), .A2(n6658), .B1(n6002), .B2(n6663), .C1(n6001), 
        .C2(n6000), .ZN(U2842) );
  INV_X1 U6726 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6004) );
  OAI222_X1 U6727 ( .A1(n6028), .A2(n6005), .B1(n6663), .B2(n6004), .C1(n6003), 
        .C2(n6658), .ZN(U2844) );
  NAND3_X1 U6728 ( .A1(n6040), .A2(n6006), .A3(n6026), .ZN(n6008) );
  AOI22_X1 U6729 ( .A1(n7113), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n7116), .ZN(n6007) );
  NAND2_X1 U6730 ( .A1(n6008), .A2(n6007), .ZN(U2860) );
  AOI22_X1 U6731 ( .A1(n7113), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n7116), .ZN(n6010) );
  NAND2_X1 U6732 ( .A1(n7117), .A2(DATAI_13_), .ZN(n6009) );
  OAI211_X1 U6733 ( .C1(n6011), .C2(n7100), .A(n6010), .B(n6009), .ZN(U2862)
         );
  AOI22_X1 U6734 ( .A1(n7113), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n7116), .ZN(n6013) );
  NAND2_X1 U6735 ( .A1(n7117), .A2(DATAI_12_), .ZN(n6012) );
  OAI211_X1 U6736 ( .C1(n5889), .C2(n7100), .A(n6013), .B(n6012), .ZN(U2863)
         );
  AOI22_X1 U6737 ( .A1(n7113), .A2(DATAI_27_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n7116), .ZN(n6015) );
  NAND2_X1 U6738 ( .A1(n7117), .A2(DATAI_11_), .ZN(n6014) );
  OAI211_X1 U6739 ( .C1(n6016), .C2(n7100), .A(n6015), .B(n6014), .ZN(U2864)
         );
  AOI22_X1 U6740 ( .A1(n7113), .A2(DATAI_26_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n7116), .ZN(n6018) );
  NAND2_X1 U6741 ( .A1(n7117), .A2(DATAI_10_), .ZN(n6017) );
  OAI211_X1 U6742 ( .C1(n6054), .C2(n7100), .A(n6018), .B(n6017), .ZN(U2865)
         );
  AOI22_X1 U6743 ( .A1(n7113), .A2(DATAI_25_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n7116), .ZN(n6020) );
  NAND2_X1 U6744 ( .A1(n7117), .A2(DATAI_9_), .ZN(n6019) );
  OAI211_X1 U6745 ( .C1(n6021), .C2(n7100), .A(n6020), .B(n6019), .ZN(U2866)
         );
  AOI22_X1 U6746 ( .A1(n7113), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n7116), .ZN(n6023) );
  NAND2_X1 U6747 ( .A1(n7117), .A2(DATAI_8_), .ZN(n6022) );
  OAI211_X1 U6748 ( .C1(n6073), .C2(n7100), .A(n6023), .B(n6022), .ZN(U2867)
         );
  AOI22_X1 U6749 ( .A1(n7113), .A2(DATAI_20_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n7116), .ZN(n6025) );
  NAND2_X1 U6750 ( .A1(n7117), .A2(DATAI_4_), .ZN(n6024) );
  OAI211_X1 U6751 ( .C1(n6979), .C2(n7100), .A(n6025), .B(n6024), .ZN(U2871)
         );
  INV_X1 U6752 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6573) );
  OAI222_X1 U6753 ( .A1(n6028), .A2(n7100), .B1(n6027), .B2(n6460), .C1(n6026), 
        .C2(n6573), .ZN(U2876) );
  NAND4_X1 U6754 ( .A1(n6106), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n6033) );
  INV_X1 U6755 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6132) );
  AND2_X1 U6756 ( .A1(n6029), .A2(n6132), .ZN(n6030) );
  NAND2_X1 U6757 ( .A1(n6031), .A2(n6030), .ZN(n6032) );
  OAI21_X1 U6758 ( .B1(n6034), .B2(n6033), .A(n6032), .ZN(n6035) );
  XNOR2_X1 U6759 ( .A(n6035), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n6130)
         );
  NOR2_X1 U6760 ( .A1(n4480), .A2(n6036), .ZN(n6126) );
  AOI21_X1 U6761 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n6126), 
        .ZN(n6037) );
  OAI21_X1 U6762 ( .B1(n6038), .B2(n6717), .A(n6037), .ZN(n6039) );
  OAI21_X1 U6763 ( .B1(n6130), .B2(n6696), .A(n6041), .ZN(U2955) );
  NOR2_X1 U6764 ( .A1(n6043), .A2(n6042), .ZN(n6045) );
  XNOR2_X1 U6765 ( .A(n6106), .B(n4637), .ZN(n6044) );
  XNOR2_X1 U6766 ( .A(n6045), .B(n6044), .ZN(n6149) );
  NOR2_X1 U6767 ( .A1(n4480), .A2(n6613), .ZN(n6144) );
  AOI21_X1 U6768 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n6144), 
        .ZN(n6046) );
  OAI21_X1 U6769 ( .B1(n6717), .B2(n6047), .A(n6046), .ZN(n6048) );
  AOI21_X1 U6770 ( .B1(n6049), .B2(n6713), .A(n6048), .ZN(n6050) );
  OAI21_X1 U6771 ( .B1(n6149), .B2(n6696), .A(n6050), .ZN(U2959) );
  XNOR2_X1 U6772 ( .A(n6106), .B(n6051), .ZN(n6052) );
  XNOR2_X1 U6773 ( .A(n6053), .B(n6052), .ZN(n6159) );
  INV_X1 U6774 ( .A(n6054), .ZN(n6058) );
  INV_X1 U6775 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6423) );
  NOR2_X1 U6776 ( .A1(n4480), .A2(n6423), .ZN(n6153) );
  AOI21_X1 U6777 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n6153), 
        .ZN(n6055) );
  OAI21_X1 U6778 ( .B1(n6717), .B2(n6056), .A(n6055), .ZN(n6057) );
  AOI21_X1 U6779 ( .B1(n6058), .B2(n6713), .A(n6057), .ZN(n6059) );
  OAI21_X1 U6780 ( .B1(n6159), .B2(n6696), .A(n6059), .ZN(U2960) );
  OAI21_X1 U6781 ( .B1(n6062), .B2(n6061), .A(n6060), .ZN(n6063) );
  INV_X1 U6782 ( .A(n6063), .ZN(n6167) );
  NOR2_X1 U6783 ( .A1(n4480), .A2(n6610), .ZN(n6160) );
  AOI21_X1 U6784 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6160), 
        .ZN(n6064) );
  OAI21_X1 U6785 ( .B1(n6717), .B2(n6065), .A(n6064), .ZN(n6066) );
  AOI21_X1 U6786 ( .B1(n6067), .B2(n6713), .A(n6066), .ZN(n6068) );
  OAI21_X1 U6787 ( .B1(n6167), .B2(n6696), .A(n6068), .ZN(U2961) );
  NAND4_X1 U6788 ( .A1(n6097), .A2(n6190), .A3(n4460), .A4(n6069), .ZN(n6083)
         );
  NAND4_X1 U6789 ( .A1(n6070), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .A4(n6106), .ZN(n6071) );
  OAI21_X1 U6790 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n6083), .A(n6071), 
        .ZN(n6072) );
  XNOR2_X1 U6791 ( .A(n6072), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n6176)
         );
  INV_X1 U6792 ( .A(n6074), .ZN(n6076) );
  NOR2_X1 U6793 ( .A1(n4480), .A2(n6608), .ZN(n6173) );
  AOI21_X1 U6794 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6173), 
        .ZN(n6075) );
  OAI21_X1 U6795 ( .B1(n6717), .B2(n6076), .A(n6075), .ZN(n6077) );
  AOI21_X1 U6796 ( .B1(n6078), .B2(n6713), .A(n6077), .ZN(n6079) );
  OAI21_X1 U6797 ( .B1(n6176), .B2(n6696), .A(n6079), .ZN(U2962) );
  NAND2_X1 U6798 ( .A1(n6106), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6702) );
  NOR2_X1 U6799 ( .A1(n6080), .A2(n6702), .ZN(n6107) );
  INV_X1 U6800 ( .A(n6081), .ZN(n6181) );
  NAND3_X1 U6801 ( .A1(n6107), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n6181), .ZN(n6082) );
  NAND2_X1 U6802 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  XNOR2_X1 U6803 ( .A(n6084), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6184)
         );
  INV_X1 U6804 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U6805 ( .A1(n4480), .A2(n6606), .ZN(n6178) );
  AOI21_X1 U6806 ( .B1(n6707), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6178), 
        .ZN(n6085) );
  OAI21_X1 U6807 ( .B1(n6717), .B2(n7011), .A(n6085), .ZN(n6086) );
  AOI21_X1 U6808 ( .B1(n7115), .B2(n6713), .A(n6086), .ZN(n6087) );
  OAI21_X1 U6809 ( .B1(n6184), .B2(n6696), .A(n6087), .ZN(U2963) );
  INV_X1 U6810 ( .A(n6097), .ZN(n6710) );
  OAI22_X1 U6811 ( .A1(n6710), .A2(n6088), .B1(n4460), .B2(n6207), .ZN(n6090)
         );
  XNOR2_X1 U6812 ( .A(n6090), .B(n6089), .ZN(n6205) );
  INV_X1 U6813 ( .A(n5989), .ZN(n6091) );
  AOI21_X1 U6814 ( .B1(n6092), .B2(n6091), .A(n5917), .ZN(n7110) );
  NAND2_X1 U6815 ( .A1(n6771), .A2(REIP_REG_21__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U6816 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n6093)
         );
  OAI211_X1 U6817 ( .C1(n6717), .C2(n6996), .A(n6199), .B(n6093), .ZN(n6094)
         );
  AOI21_X1 U6818 ( .B1(n7110), .B2(n6713), .A(n6094), .ZN(n6095) );
  OAI21_X1 U6819 ( .B1(n6205), .B2(n6696), .A(n6095), .ZN(U2965) );
  NOR2_X1 U6820 ( .A1(n4460), .A2(n6096), .ZN(n6098) );
  MUX2_X1 U6821 ( .A(n6098), .B(n4460), .S(n6097), .Z(n6099) );
  XNOR2_X1 U6822 ( .A(n6099), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6212)
         );
  NAND2_X1 U6823 ( .A1(n6693), .A2(n6982), .ZN(n6100) );
  OR2_X1 U6824 ( .A1(n4480), .A2(n6974), .ZN(n6206) );
  OAI211_X1 U6825 ( .C1(n6101), .C2(n6985), .A(n6100), .B(n6206), .ZN(n6102)
         );
  AOI21_X1 U6826 ( .B1(n6103), .B2(n6713), .A(n6102), .ZN(n6104) );
  OAI21_X1 U6827 ( .B1(n6212), .B2(n6696), .A(n6104), .ZN(U2966) );
  OAI21_X1 U6828 ( .B1(n6106), .B2(n6105), .A(n6080), .ZN(n6703) );
  NAND2_X1 U6829 ( .A1(n4460), .A2(n4462), .ZN(n6699) );
  NOR2_X1 U6830 ( .A1(n6703), .A2(n6699), .ZN(n6698) );
  NOR2_X1 U6831 ( .A1(n6698), .A2(n6107), .ZN(n6109) );
  XNOR2_X1 U6832 ( .A(n6109), .B(n6108), .ZN(n6219) );
  INV_X1 U6833 ( .A(n6957), .ZN(n6111) );
  NAND2_X1 U6834 ( .A1(n6707), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6110)
         );
  NAND2_X1 U6835 ( .A1(n6771), .A2(REIP_REG_18__SCAN_IN), .ZN(n6216) );
  OAI211_X1 U6836 ( .C1(n6717), .C2(n6111), .A(n6110), .B(n6216), .ZN(n6112)
         );
  AOI21_X1 U6837 ( .B1(n7104), .B2(n6713), .A(n6112), .ZN(n6113) );
  OAI21_X1 U6838 ( .B1(n6219), .B2(n6696), .A(n6113), .ZN(U2968) );
  XNOR2_X1 U6839 ( .A(n6106), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6114)
         );
  XNOR2_X1 U6840 ( .A(n6115), .B(n6114), .ZN(n6835) );
  NAND2_X1 U6841 ( .A1(n6835), .A2(n6714), .ZN(n6119) );
  NOR2_X1 U6842 ( .A1(n4480), .A2(n6594), .ZN(n6832) );
  NOR2_X1 U6843 ( .A1(n6717), .A2(n6116), .ZN(n6117) );
  AOI211_X1 U6844 ( .C1(n6707), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n6832), 
        .B(n6117), .ZN(n6118) );
  OAI211_X1 U6845 ( .C1(n6121), .C2(n6120), .A(n6119), .B(n6118), .ZN(U2970)
         );
  AOI211_X1 U6846 ( .C1(n6133), .C2(n6122), .A(n6132), .B(n6145), .ZN(n6131)
         );
  INV_X1 U6847 ( .A(n6122), .ZN(n6123) );
  NOR3_X1 U6848 ( .A1(n6131), .A2(n6123), .A3(n4847), .ZN(n6128) );
  NOR2_X1 U6849 ( .A1(n6124), .A2(n6793), .ZN(n6127) );
  NOR4_X1 U6850 ( .A1(n6134), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6132), 
        .A4(n6133), .ZN(n6125) );
  NOR4_X2 U6851 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n6129)
         );
  OAI21_X1 U6852 ( .B1(n6130), .B2(n6800), .A(n6129), .ZN(U2987) );
  INV_X1 U6853 ( .A(n6131), .ZN(n6139) );
  OAI21_X1 U6854 ( .B1(n6134), .B2(n6133), .A(n6132), .ZN(n6138) );
  OAI21_X1 U6855 ( .B1(n6136), .B2(n6793), .A(n6135), .ZN(n6137) );
  AOI21_X1 U6856 ( .B1(n6139), .B2(n6138), .A(n6137), .ZN(n6140) );
  OAI21_X1 U6857 ( .B1(n6141), .B2(n6800), .A(n6140), .ZN(U2988) );
  NOR2_X1 U6858 ( .A1(n6142), .A2(n6793), .ZN(n6143) );
  AOI211_X1 U6859 ( .C1(n6145), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n6144), .B(n6143), .ZN(n6148) );
  NAND2_X1 U6860 ( .A1(n6146), .A2(n4637), .ZN(n6147) );
  OAI211_X1 U6861 ( .C1(n6149), .C2(n6800), .A(n6148), .B(n6147), .ZN(U2991)
         );
  INV_X1 U6862 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6150) );
  NOR4_X1 U6863 ( .A1(n6753), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .A3(n6151), 
        .A4(n6150), .ZN(n6152) );
  AOI211_X1 U6864 ( .C1(n6860), .C2(n6154), .A(n6153), .B(n6152), .ZN(n6158)
         );
  INV_X1 U6865 ( .A(n6155), .ZN(n6156) );
  NOR2_X1 U6866 ( .A1(n6156), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6163)
         );
  INV_X1 U6867 ( .A(n6169), .ZN(n6165) );
  OAI21_X1 U6868 ( .B1(n6163), .B2(n6165), .A(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n6157) );
  OAI211_X1 U6869 ( .C1(n6159), .C2(n6800), .A(n6158), .B(n6157), .ZN(U2992)
         );
  INV_X1 U6870 ( .A(n6160), .ZN(n6161) );
  OAI21_X1 U6871 ( .B1(n6162), .B2(n6793), .A(n6161), .ZN(n6164) );
  AOI211_X1 U6872 ( .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n6165), .A(n6164), .B(n6163), .ZN(n6166) );
  OAI21_X1 U6873 ( .B1(n6167), .B2(n6800), .A(n6166), .ZN(U2993) );
  INV_X1 U6874 ( .A(n6168), .ZN(n6174) );
  INV_X1 U6875 ( .A(n6753), .ZN(n6188) );
  NAND3_X1 U6876 ( .A1(n6188), .A2(n6181), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n6170) );
  AOI21_X1 U6877 ( .B1(n6171), .B2(n6170), .A(n6169), .ZN(n6172) );
  AOI211_X1 U6878 ( .C1(n6860), .C2(n6174), .A(n6173), .B(n6172), .ZN(n6175)
         );
  OAI21_X1 U6879 ( .B1(n6176), .B2(n6800), .A(n6175), .ZN(U2994) );
  NOR2_X1 U6880 ( .A1(n7005), .A2(n6793), .ZN(n6177) );
  AOI211_X1 U6881 ( .C1(n6179), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n6178), .B(n6177), .ZN(n6183) );
  NAND3_X1 U6882 ( .A1(n6188), .A2(n6181), .A3(n6180), .ZN(n6182) );
  OAI211_X1 U6883 ( .C1(n6184), .C2(n6800), .A(n6183), .B(n6182), .ZN(U2995)
         );
  INV_X1 U6884 ( .A(n6185), .ZN(n6203) );
  OAI21_X1 U6885 ( .B1(n6187), .B2(n6793), .A(n6186), .ZN(n6192) );
  NAND2_X1 U6886 ( .A1(n6188), .A2(n6207), .ZN(n6200) );
  NOR3_X1 U6887 ( .A1(n6200), .A2(n6190), .A3(n6189), .ZN(n6191) );
  AOI211_X1 U6888 ( .C1(n6203), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n6192), .B(n6191), .ZN(n6193) );
  OAI21_X1 U6889 ( .B1(n6194), .B2(n6800), .A(n6193), .ZN(U2996) );
  NAND2_X1 U6890 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  NAND2_X1 U6891 ( .A1(n6198), .A2(n6197), .ZN(n6648) );
  OAI21_X1 U6892 ( .B1(n6648), .B2(n6793), .A(n6199), .ZN(n6202) );
  NOR2_X1 U6893 ( .A1(n6200), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6201)
         );
  AOI211_X1 U6894 ( .C1(n6203), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n6202), .B(n6201), .ZN(n6204) );
  OAI21_X1 U6895 ( .B1(n6205), .B2(n6800), .A(n6204), .ZN(U2997) );
  OAI21_X1 U6896 ( .B1(n6977), .B2(n6793), .A(n6206), .ZN(n6210) );
  NOR3_X1 U6897 ( .A1(n6753), .A2(n6208), .A3(n6207), .ZN(n6209) );
  AOI211_X1 U6898 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n6748), .A(n6210), .B(n6209), .ZN(n6211) );
  OAI21_X1 U6899 ( .B1(n6212), .B2(n6800), .A(n6211), .ZN(U2998) );
  OAI21_X1 U6900 ( .B1(n6754), .B2(n6214), .A(n6831), .ZN(n6849) );
  NOR2_X1 U6901 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6842), .ZN(n6213)
         );
  NAND2_X1 U6902 ( .A1(n6214), .A2(n6213), .ZN(n6215) );
  OAI211_X1 U6903 ( .C1(n6960), .C2(n6793), .A(n6216), .B(n6215), .ZN(n6217)
         );
  AOI21_X1 U6904 ( .B1(n6849), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6217), 
        .ZN(n6218) );
  OAI21_X1 U6905 ( .B1(n6219), .B2(n6800), .A(n6218), .ZN(U3000) );
  NOR2_X1 U6906 ( .A1(n7020), .A2(n6225), .ZN(n6220) );
  INV_X1 U6907 ( .A(n6220), .ZN(n6257) );
  AOI21_X1 U6908 ( .B1(n7122), .B2(n6221), .A(n6220), .ZN(n6228) );
  NOR2_X1 U6909 ( .A1(n6222), .A2(n7132), .ZN(n6224) );
  AOI22_X1 U6910 ( .A1(n6228), .A2(n6224), .B1(n7132), .B2(n6225), .ZN(n6223)
         );
  NAND2_X1 U6911 ( .A1(n7143), .A2(n6223), .ZN(n6253) );
  INV_X1 U6912 ( .A(n6224), .ZN(n6227) );
  OAI22_X1 U6913 ( .A1(n6228), .A2(n6227), .B1(n6226), .B2(n6225), .ZN(n6252)
         );
  AOI22_X1 U6914 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n6253), .B1(n6273), 
        .B2(n6252), .ZN(n6232) );
  NOR3_X4 U6915 ( .A1(n6230), .A2(n6229), .A3(n4386), .ZN(n6317) );
  AOI22_X1 U6916 ( .A1(n6317), .A2(n7148), .B1(n7138), .B2(n6254), .ZN(n6231)
         );
  OAI211_X1 U6917 ( .C1(n6233), .C2(n6257), .A(n6232), .B(n6231), .ZN(U3124)
         );
  AOI22_X1 U6918 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6253), .B1(n6279), 
        .B2(n6252), .ZN(n6235) );
  AOI22_X1 U6919 ( .A1(n6317), .A2(n7154), .B1(n7156), .B2(n6254), .ZN(n6234)
         );
  OAI211_X1 U6920 ( .C1(n6236), .C2(n6257), .A(n6235), .B(n6234), .ZN(U3125)
         );
  AOI22_X1 U6921 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n6253), .B1(n6285), 
        .B2(n6252), .ZN(n6238) );
  AOI22_X1 U6922 ( .A1(n6317), .A2(n7164), .B1(n7162), .B2(n6254), .ZN(n6237)
         );
  OAI211_X1 U6923 ( .C1(n6239), .C2(n6257), .A(n6238), .B(n6237), .ZN(U3126)
         );
  AOI22_X1 U6924 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6253), .B1(n6291), 
        .B2(n6252), .ZN(n6241) );
  AOI22_X1 U6925 ( .A1(n6317), .A2(n7170), .B1(n7172), .B2(n6254), .ZN(n6240)
         );
  OAI211_X1 U6926 ( .C1(n6242), .C2(n6257), .A(n6241), .B(n6240), .ZN(U3127)
         );
  AOI22_X1 U6927 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6253), .B1(n6297), 
        .B2(n6252), .ZN(n6244) );
  AOI22_X1 U6928 ( .A1(n6317), .A2(n7180), .B1(n7178), .B2(n6254), .ZN(n6243)
         );
  OAI211_X1 U6929 ( .C1(n6245), .C2(n6257), .A(n6244), .B(n6243), .ZN(U3128)
         );
  AOI22_X1 U6930 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6253), .B1(n6303), 
        .B2(n6252), .ZN(n6247) );
  AOI22_X1 U6931 ( .A1(n6317), .A2(n7186), .B1(n7188), .B2(n6254), .ZN(n6246)
         );
  OAI211_X1 U6932 ( .C1(n6248), .C2(n6257), .A(n6247), .B(n6246), .ZN(U3129)
         );
  AOI22_X1 U6933 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6253), .B1(n6309), 
        .B2(n6252), .ZN(n6250) );
  AOI22_X1 U6934 ( .A1(n6317), .A2(n7194), .B1(n7196), .B2(n6254), .ZN(n6249)
         );
  OAI211_X1 U6935 ( .C1(n6251), .C2(n6257), .A(n6250), .B(n6249), .ZN(U3130)
         );
  AOI22_X1 U6936 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6253), .B1(n6316), 
        .B2(n6252), .ZN(n6256) );
  AOI22_X1 U6937 ( .A1(n6317), .A2(n7212), .B1(n7208), .B2(n6254), .ZN(n6255)
         );
  OAI211_X1 U6938 ( .C1(n6258), .C2(n6257), .A(n6256), .B(n6255), .ZN(U3131)
         );
  NOR2_X1 U6939 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6259), .ZN(n6322)
         );
  INV_X1 U6940 ( .A(n6322), .ZN(n6262) );
  AOI211_X1 U6941 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6262), .A(n6261), .B(
        n6260), .ZN(n6268) );
  INV_X1 U6942 ( .A(n6319), .ZN(n6263) );
  OAI21_X1 U6943 ( .B1(n6317), .B2(n6263), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6264) );
  OAI21_X1 U6944 ( .B1(n6266), .B2(n6265), .A(n6264), .ZN(n6267) );
  INV_X1 U6945 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n6278) );
  INV_X1 U6946 ( .A(n6269), .ZN(n7134) );
  OAI22_X1 U6947 ( .A1(n6272), .A2(n7134), .B1(n6271), .B2(n6270), .ZN(n6315)
         );
  AOI22_X1 U6948 ( .A1(n6317), .A2(n7138), .B1(n6273), .B2(n6315), .ZN(n6274)
         );
  OAI21_X1 U6949 ( .B1(n6275), .B2(n6319), .A(n6274), .ZN(n6276) );
  AOI21_X1 U6950 ( .B1(n7139), .B2(n6322), .A(n6276), .ZN(n6277) );
  OAI21_X1 U6951 ( .B1(n6325), .B2(n6278), .A(n6277), .ZN(U3132) );
  INV_X1 U6952 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6284) );
  AOI22_X1 U6953 ( .A1(n6317), .A2(n7156), .B1(n6279), .B2(n6315), .ZN(n6280)
         );
  OAI21_X1 U6954 ( .B1(n6281), .B2(n6319), .A(n6280), .ZN(n6282) );
  AOI21_X1 U6955 ( .B1(n7155), .B2(n6322), .A(n6282), .ZN(n6283) );
  OAI21_X1 U6956 ( .B1(n6325), .B2(n6284), .A(n6283), .ZN(U3133) );
  INV_X1 U6957 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n6290) );
  AOI22_X1 U6958 ( .A1(n6317), .A2(n7162), .B1(n6285), .B2(n6315), .ZN(n6286)
         );
  OAI21_X1 U6959 ( .B1(n6287), .B2(n6319), .A(n6286), .ZN(n6288) );
  AOI21_X1 U6960 ( .B1(n7163), .B2(n6322), .A(n6288), .ZN(n6289) );
  OAI21_X1 U6961 ( .B1(n6325), .B2(n6290), .A(n6289), .ZN(U3134) );
  INV_X1 U6962 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n6296) );
  AOI22_X1 U6963 ( .A1(n6317), .A2(n7172), .B1(n6291), .B2(n6315), .ZN(n6292)
         );
  OAI21_X1 U6964 ( .B1(n6293), .B2(n6319), .A(n6292), .ZN(n6294) );
  AOI21_X1 U6965 ( .B1(n7171), .B2(n6322), .A(n6294), .ZN(n6295) );
  OAI21_X1 U6966 ( .B1(n6325), .B2(n6296), .A(n6295), .ZN(U3135) );
  INV_X1 U6967 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6302) );
  AOI22_X1 U6968 ( .A1(n6317), .A2(n7178), .B1(n6297), .B2(n6315), .ZN(n6298)
         );
  OAI21_X1 U6969 ( .B1(n6299), .B2(n6319), .A(n6298), .ZN(n6300) );
  AOI21_X1 U6970 ( .B1(n7179), .B2(n6322), .A(n6300), .ZN(n6301) );
  OAI21_X1 U6971 ( .B1(n6325), .B2(n6302), .A(n6301), .ZN(U3136) );
  INV_X1 U6972 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6308) );
  AOI22_X1 U6973 ( .A1(n6317), .A2(n7188), .B1(n6303), .B2(n6315), .ZN(n6304)
         );
  OAI21_X1 U6974 ( .B1(n6305), .B2(n6319), .A(n6304), .ZN(n6306) );
  AOI21_X1 U6975 ( .B1(n7187), .B2(n6322), .A(n6306), .ZN(n6307) );
  OAI21_X1 U6976 ( .B1(n6325), .B2(n6308), .A(n6307), .ZN(U3137) );
  INV_X1 U6977 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U6978 ( .A1(n6317), .A2(n7196), .B1(n6309), .B2(n6315), .ZN(n6310)
         );
  OAI21_X1 U6979 ( .B1(n6311), .B2(n6319), .A(n6310), .ZN(n6312) );
  AOI21_X1 U6980 ( .B1(n7195), .B2(n6322), .A(n6312), .ZN(n6313) );
  OAI21_X1 U6981 ( .B1(n6325), .B2(n6314), .A(n6313), .ZN(U3138) );
  INV_X1 U6982 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6324) );
  AOI22_X1 U6983 ( .A1(n6317), .A2(n7208), .B1(n6316), .B2(n6315), .ZN(n6318)
         );
  OAI21_X1 U6984 ( .B1(n6320), .B2(n6319), .A(n6318), .ZN(n6321) );
  AOI21_X1 U6985 ( .B1(n7210), .B2(n6322), .A(n6321), .ZN(n6323) );
  OAI21_X1 U6986 ( .B1(n6325), .B2(n6324), .A(n6323), .ZN(U3139) );
  INV_X1 U6987 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6639) );
  INV_X1 U6988 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6730) );
  AOI21_X1 U6989 ( .B1(n6730), .B2(STATE_REG_1__SCAN_IN), .A(n4357), .ZN(n6328) );
  NOR2_X1 U6990 ( .A1(n7099), .A2(n6328), .ZN(n7083) );
  INV_X1 U6991 ( .A(n7083), .ZN(n6326) );
  INV_X1 U6992 ( .A(BS16_N), .ZN(n6428) );
  NAND2_X1 U6993 ( .A1(n6730), .A2(n4357), .ZN(n6723) );
  AOI21_X1 U6994 ( .B1(n6428), .B2(n6723), .A(n6326), .ZN(n7079) );
  AOI21_X1 U6995 ( .B1(n6639), .B2(n6326), .A(n7079), .ZN(U3451) );
  AND2_X1 U6996 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6326), .ZN(U3180) );
  AND2_X1 U6997 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6326), .ZN(U3179) );
  AND2_X1 U6998 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6326), .ZN(U3178) );
  AND2_X1 U6999 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6326), .ZN(U3177) );
  AND2_X1 U7000 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6326), .ZN(U3176) );
  AND2_X1 U7001 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6326), .ZN(U3175) );
  AND2_X1 U7002 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6326), .ZN(U3174) );
  AND2_X1 U7003 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6326), .ZN(U3173) );
  AND2_X1 U7004 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6326), .ZN(U3172) );
  AND2_X1 U7005 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6326), .ZN(U3171) );
  AND2_X1 U7006 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6326), .ZN(U3170) );
  AND2_X1 U7007 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6326), .ZN(U3169) );
  AND2_X1 U7008 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6326), .ZN(U3168) );
  AND2_X1 U7009 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6326), .ZN(U3167) );
  AND2_X1 U7010 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6326), .ZN(U3166) );
  AND2_X1 U7011 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6326), .ZN(U3165) );
  AND2_X1 U7012 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6326), .ZN(U3164) );
  AND2_X1 U7013 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6326), .ZN(U3163) );
  AND2_X1 U7014 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6326), .ZN(U3162) );
  AND2_X1 U7015 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6326), .ZN(U3161) );
  AND2_X1 U7016 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6326), .ZN(U3160) );
  AND2_X1 U7017 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6326), .ZN(U3159) );
  AND2_X1 U7018 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6326), .ZN(U3158) );
  AND2_X1 U7019 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6326), .ZN(U3157) );
  AND2_X1 U7020 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6326), .ZN(U3156) );
  AND2_X1 U7021 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6326), .ZN(U3155) );
  AND2_X1 U7022 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6326), .ZN(U3154) );
  AND2_X1 U7023 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6326), .ZN(U3153) );
  AND2_X1 U7024 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6326), .ZN(U3152) );
  AND2_X1 U7025 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6326), .ZN(U3151) );
  AND2_X1 U7026 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n6327), .ZN(U3019)
         );
  INV_X1 U7027 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6499) );
  AOI21_X1 U7028 ( .B1(n6328), .B2(n6499), .A(n7099), .ZN(U2789) );
  AOI22_X1 U7029 ( .A1(REIP_REG_22__SCAN_IN), .A2(keyinput_60), .B1(n6606), 
        .B2(keyinput_59), .ZN(n6329) );
  OAI221_X1 U7030 ( .B1(REIP_REG_22__SCAN_IN), .B2(keyinput_60), .C1(n6606), 
        .C2(keyinput_59), .A(n6329), .ZN(n6417) );
  AOI22_X1 U7031 ( .A1(n6610), .A2(keyinput_57), .B1(n6423), .B2(keyinput_56), 
        .ZN(n6330) );
  OAI221_X1 U7032 ( .B1(n6610), .B2(keyinput_57), .C1(n6423), .C2(keyinput_56), 
        .A(n6330), .ZN(n6414) );
  OAI22_X1 U7033 ( .A1(n6332), .A2(keyinput_53), .B1(REIP_REG_28__SCAN_IN), 
        .B2(keyinput_54), .ZN(n6331) );
  AOI221_X1 U7034 ( .B1(n6332), .B2(keyinput_53), .C1(keyinput_54), .C2(
        REIP_REG_28__SCAN_IN), .A(n6331), .ZN(n6411) );
  INV_X1 U7035 ( .A(keyinput_49), .ZN(n6405) );
  INV_X1 U7036 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6515) );
  INV_X1 U7037 ( .A(keyinput_48), .ZN(n6403) );
  INV_X1 U7038 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6642) );
  INV_X1 U7039 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6504) );
  AOI22_X1 U7040 ( .A1(M_IO_N_REG_SCAN_IN), .A2(keyinput_40), .B1(
        CODEFETCH_REG_SCAN_IN), .B2(keyinput_39), .ZN(n6333) );
  OAI221_X1 U7041 ( .B1(M_IO_N_REG_SCAN_IN), .B2(keyinput_40), .C1(
        CODEFETCH_REG_SCAN_IN), .C2(keyinput_39), .A(n6333), .ZN(n6393) );
  OAI22_X1 U7042 ( .A1(HOLD), .A2(keyinput_36), .B1(keyinput_38), .B2(
        ADS_N_REG_SCAN_IN), .ZN(n6334) );
  AOI221_X1 U7043 ( .B1(HOLD), .B2(keyinput_36), .C1(ADS_N_REG_SCAN_IN), .C2(
        keyinput_38), .A(n6334), .ZN(n6390) );
  INV_X1 U7044 ( .A(NA_N), .ZN(n7090) );
  OAI22_X1 U7045 ( .A1(n7090), .A2(keyinput_33), .B1(BS16_N), .B2(keyinput_34), 
        .ZN(n6335) );
  AOI221_X1 U7046 ( .B1(n7090), .B2(keyinput_33), .C1(keyinput_34), .C2(BS16_N), .A(n6335), .ZN(n6387) );
  INV_X1 U7047 ( .A(keyinput_32), .ZN(n6385) );
  INV_X1 U7048 ( .A(keyinput_31), .ZN(n6383) );
  AOI22_X1 U7049 ( .A1(DATAI_5_), .A2(keyinput_26), .B1(n6431), .B2(
        keyinput_25), .ZN(n6336) );
  OAI221_X1 U7050 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(n6431), .C2(
        keyinput_25), .A(n6336), .ZN(n6376) );
  INV_X1 U7051 ( .A(keyinput_24), .ZN(n6374) );
  INV_X1 U7052 ( .A(DATAI_20_), .ZN(n6338) );
  OAI22_X1 U7053 ( .A1(n6338), .A2(keyinput_11), .B1(keyinput_10), .B2(
        DATAI_21_), .ZN(n6337) );
  AOI221_X1 U7054 ( .B1(n6338), .B2(keyinput_11), .C1(DATAI_21_), .C2(
        keyinput_10), .A(n6337), .ZN(n6359) );
  INV_X1 U7055 ( .A(keyinput_9), .ZN(n6353) );
  INV_X1 U7056 ( .A(DATAI_22_), .ZN(n6451) );
  INV_X1 U7057 ( .A(DATAI_28_), .ZN(n6436) );
  INV_X1 U7058 ( .A(DATAI_27_), .ZN(n6441) );
  INV_X1 U7059 ( .A(DATAI_25_), .ZN(n6340) );
  OAI22_X1 U7060 ( .A1(n6441), .A2(keyinput_4), .B1(n6340), .B2(keyinput_6), 
        .ZN(n6339) );
  AOI221_X1 U7061 ( .B1(n6441), .B2(keyinput_4), .C1(keyinput_6), .C2(n6340), 
        .A(n6339), .ZN(n6344) );
  INV_X1 U7062 ( .A(DATAI_26_), .ZN(n6435) );
  INV_X1 U7063 ( .A(DATAI_24_), .ZN(n6342) );
  OAI22_X1 U7064 ( .A1(n6435), .A2(keyinput_5), .B1(n6342), .B2(keyinput_7), 
        .ZN(n6341) );
  AOI221_X1 U7065 ( .B1(n6435), .B2(keyinput_5), .C1(keyinput_7), .C2(n6342), 
        .A(n6341), .ZN(n6343) );
  OAI211_X1 U7066 ( .C1(n6436), .C2(keyinput_3), .A(n6344), .B(n6343), .ZN(
        n6345) );
  AOI21_X1 U7067 ( .B1(n6436), .B2(keyinput_3), .A(n6345), .ZN(n6350) );
  INV_X1 U7068 ( .A(DATAI_29_), .ZN(n6444) );
  INV_X1 U7069 ( .A(keyinput_2), .ZN(n6348) );
  AOI22_X1 U7070 ( .A1(DATAI_30_), .A2(keyinput_1), .B1(DATAI_31_), .B2(
        keyinput_0), .ZN(n6346) );
  OAI221_X1 U7071 ( .B1(DATAI_30_), .B2(keyinput_1), .C1(DATAI_31_), .C2(
        keyinput_0), .A(n6346), .ZN(n6347) );
  OAI221_X1 U7072 ( .B1(DATAI_29_), .B2(keyinput_2), .C1(n6444), .C2(n6348), 
        .A(n6347), .ZN(n6349) );
  AOI22_X1 U7073 ( .A1(n6350), .A2(n6349), .B1(keyinput_8), .B2(DATAI_23_), 
        .ZN(n6351) );
  OAI21_X1 U7074 ( .B1(keyinput_8), .B2(DATAI_23_), .A(n6351), .ZN(n6352) );
  OAI221_X1 U7075 ( .B1(DATAI_22_), .B2(n6353), .C1(n6451), .C2(keyinput_9), 
        .A(n6352), .ZN(n6358) );
  XOR2_X1 U7076 ( .A(DATAI_18_), .B(keyinput_13), .Z(n6357) );
  INV_X1 U7077 ( .A(DATAI_17_), .ZN(n6355) );
  AOI22_X1 U7078 ( .A1(DATAI_19_), .A2(keyinput_12), .B1(n6355), .B2(
        keyinput_14), .ZN(n6354) );
  OAI221_X1 U7079 ( .B1(DATAI_19_), .B2(keyinput_12), .C1(n6355), .C2(
        keyinput_14), .A(n6354), .ZN(n6356) );
  AOI211_X1 U7080 ( .C1(n6359), .C2(n6358), .A(n6357), .B(n6356), .ZN(n6368)
         );
  INV_X1 U7081 ( .A(DATAI_16_), .ZN(n6461) );
  AOI22_X1 U7082 ( .A1(DATAI_15_), .A2(keyinput_16), .B1(n6461), .B2(
        keyinput_15), .ZN(n6360) );
  OAI221_X1 U7083 ( .B1(DATAI_15_), .B2(keyinput_16), .C1(n6461), .C2(
        keyinput_15), .A(n6360), .ZN(n6367) );
  OAI22_X1 U7084 ( .A1(n6464), .A2(keyinput_21), .B1(n6362), .B2(keyinput_22), 
        .ZN(n6361) );
  AOI221_X1 U7085 ( .B1(n6464), .B2(keyinput_21), .C1(keyinput_22), .C2(n6362), 
        .A(n6361), .ZN(n6366) );
  OAI22_X1 U7086 ( .A1(n6364), .A2(keyinput_17), .B1(n6465), .B2(keyinput_18), 
        .ZN(n6363) );
  AOI221_X1 U7087 ( .B1(n6364), .B2(keyinput_17), .C1(keyinput_18), .C2(n6465), 
        .A(n6363), .ZN(n6365) );
  OAI211_X1 U7088 ( .C1(n6368), .C2(n6367), .A(n6366), .B(n6365), .ZN(n6371)
         );
  AOI22_X1 U7089 ( .A1(DATAI_11_), .A2(keyinput_20), .B1(DATAI_12_), .B2(
        keyinput_19), .ZN(n6369) );
  OAI221_X1 U7090 ( .B1(DATAI_11_), .B2(keyinput_20), .C1(DATAI_12_), .C2(
        keyinput_19), .A(n6369), .ZN(n6370) );
  OAI22_X1 U7091 ( .A1(n6371), .A2(n6370), .B1(keyinput_23), .B2(DATAI_8_), 
        .ZN(n6372) );
  AOI21_X1 U7092 ( .B1(keyinput_23), .B2(DATAI_8_), .A(n6372), .ZN(n6373) );
  AOI221_X1 U7093 ( .B1(DATAI_7_), .B2(n6374), .C1(n6476), .C2(keyinput_24), 
        .A(n6373), .ZN(n6375) );
  OAI22_X1 U7094 ( .A1(n6376), .A2(n6375), .B1(keyinput_27), .B2(DATAI_4_), 
        .ZN(n6377) );
  AOI21_X1 U7095 ( .B1(keyinput_27), .B2(DATAI_4_), .A(n6377), .ZN(n6380) );
  AOI22_X1 U7096 ( .A1(DATAI_1_), .A2(keyinput_30), .B1(n6484), .B2(
        keyinput_28), .ZN(n6378) );
  OAI221_X1 U7097 ( .B1(DATAI_1_), .B2(keyinput_30), .C1(n6484), .C2(
        keyinput_28), .A(n6378), .ZN(n6379) );
  AOI211_X1 U7098 ( .C1(DATAI_2_), .C2(keyinput_29), .A(n6380), .B(n6379), 
        .ZN(n6381) );
  OAI21_X1 U7099 ( .B1(DATAI_2_), .B2(keyinput_29), .A(n6381), .ZN(n6382) );
  OAI221_X1 U7100 ( .B1(DATAI_0_), .B2(n6383), .C1(n6489), .C2(keyinput_31), 
        .A(n6382), .ZN(n6384) );
  OAI221_X1 U7101 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_32), .C1(n7098), 
        .C2(n6385), .A(n6384), .ZN(n6386) );
  AOI22_X1 U7102 ( .A1(keyinput_35), .A2(n7088), .B1(n6387), .B2(n6386), .ZN(
        n6388) );
  OAI21_X1 U7103 ( .B1(n7088), .B2(keyinput_35), .A(n6388), .ZN(n6389) );
  OAI211_X1 U7104 ( .C1(READREQUEST_REG_SCAN_IN), .C2(keyinput_37), .A(n6390), 
        .B(n6389), .ZN(n6391) );
  AOI21_X1 U7105 ( .B1(READREQUEST_REG_SCAN_IN), .B2(keyinput_37), .A(n6391), 
        .ZN(n6392) );
  OAI22_X1 U7106 ( .A1(n6393), .A2(n6392), .B1(n6504), .B2(keyinput_41), .ZN(
        n6394) );
  AOI21_X1 U7107 ( .B1(n6504), .B2(keyinput_41), .A(n6394), .ZN(n6401) );
  OAI22_X1 U7108 ( .A1(STATEBS16_REG_SCAN_IN), .A2(keyinput_43), .B1(
        REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_42), .ZN(n6395) );
  AOI221_X1 U7109 ( .B1(STATEBS16_REG_SCAN_IN), .B2(keyinput_43), .C1(
        keyinput_42), .C2(REQUESTPENDING_REG_SCAN_IN), .A(n6395), .ZN(n6400)
         );
  INV_X1 U7110 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U7111 ( .A1(n7037), .A2(keyinput_45), .B1(keyinput_47), .B2(n6647), 
        .ZN(n6396) );
  OAI221_X1 U7112 ( .B1(n7037), .B2(keyinput_45), .C1(n6647), .C2(keyinput_47), 
        .A(n6396), .ZN(n6399) );
  INV_X1 U7113 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6728) );
  INV_X1 U7114 ( .A(MORE_REG_SCAN_IN), .ZN(n7036) );
  AOI22_X1 U7115 ( .A1(n6728), .A2(keyinput_46), .B1(n7036), .B2(keyinput_44), 
        .ZN(n6397) );
  OAI221_X1 U7116 ( .B1(n6728), .B2(keyinput_46), .C1(n7036), .C2(keyinput_44), 
        .A(n6397), .ZN(n6398) );
  AOI211_X1 U7117 ( .C1(n6401), .C2(n6400), .A(n6399), .B(n6398), .ZN(n6402)
         );
  AOI221_X1 U7118 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6403), .C1(n6642), 
        .C2(keyinput_48), .A(n6402), .ZN(n6404) );
  AOI221_X1 U7119 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6405), .C1(n6515), 
        .C2(keyinput_49), .A(n6404), .ZN(n6408) );
  AOI22_X1 U7120 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_50), .B1(
        REIP_REG_30__SCAN_IN), .B2(keyinput_52), .ZN(n6406) );
  OAI221_X1 U7121 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_50), .C1(
        REIP_REG_30__SCAN_IN), .C2(keyinput_52), .A(n6406), .ZN(n6407) );
  AOI211_X1 U7122 ( .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_51), .A(n6408), 
        .B(n6407), .ZN(n6409) );
  OAI21_X1 U7123 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_51), .A(n6409), 
        .ZN(n6410) );
  OAI211_X1 U7124 ( .C1(n6613), .C2(keyinput_55), .A(n6411), .B(n6410), .ZN(
        n6412) );
  AOI21_X1 U7125 ( .B1(n6613), .B2(keyinput_55), .A(n6412), .ZN(n6413) );
  OAI22_X1 U7126 ( .A1(keyinput_58), .A2(n6608), .B1(n6414), .B2(n6413), .ZN(
        n6415) );
  AOI21_X1 U7127 ( .B1(keyinput_58), .B2(n6608), .A(n6415), .ZN(n6416) );
  OAI22_X1 U7128 ( .A1(n6417), .A2(n6416), .B1(REIP_REG_21__SCAN_IN), .B2(
        keyinput_61), .ZN(n6418) );
  AOI21_X1 U7129 ( .B1(REIP_REG_21__SCAN_IN), .B2(keyinput_61), .A(n6418), 
        .ZN(n6532) );
  INV_X1 U7130 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6598) );
  OAI22_X1 U7131 ( .A1(n6974), .A2(keyinput_62), .B1(n6598), .B2(keyinput_63), 
        .ZN(n6419) );
  AOI221_X1 U7132 ( .B1(n6974), .B2(keyinput_62), .C1(keyinput_63), .C2(n6598), 
        .A(n6419), .ZN(n6531) );
  AOI22_X1 U7133 ( .A1(n6974), .A2(keyinput_126), .B1(keyinput_127), .B2(n6598), .ZN(n6420) );
  OAI221_X1 U7134 ( .B1(n6974), .B2(keyinput_126), .C1(n6598), .C2(
        keyinput_127), .A(n6420), .ZN(n6530) );
  AOI22_X1 U7135 ( .A1(n6604), .A2(keyinput_124), .B1(n6606), .B2(keyinput_123), .ZN(n6421) );
  OAI221_X1 U7136 ( .B1(n6604), .B2(keyinput_124), .C1(n6606), .C2(
        keyinput_123), .A(n6421), .ZN(n6528) );
  AOI22_X1 U7137 ( .A1(REIP_REG_25__SCAN_IN), .A2(keyinput_121), .B1(n6423), 
        .B2(keyinput_120), .ZN(n6422) );
  OAI221_X1 U7138 ( .B1(REIP_REG_25__SCAN_IN), .B2(keyinput_121), .C1(n6423), 
        .C2(keyinput_120), .A(n6422), .ZN(n6524) );
  OAI22_X1 U7139 ( .A1(n6613), .A2(keyinput_119), .B1(keyinput_117), .B2(
        REIP_REG_29__SCAN_IN), .ZN(n6424) );
  AOI221_X1 U7140 ( .B1(n6613), .B2(keyinput_119), .C1(REIP_REG_29__SCAN_IN), 
        .C2(keyinput_117), .A(n6424), .ZN(n6521) );
  INV_X1 U7141 ( .A(keyinput_113), .ZN(n6514) );
  INV_X1 U7142 ( .A(keyinput_112), .ZN(n6512) );
  INV_X1 U7143 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n7097) );
  AOI22_X1 U7144 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput_103), .B1(n7097), 
        .B2(keyinput_104), .ZN(n6425) );
  OAI221_X1 U7145 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput_103), .C1(n7097), 
        .C2(keyinput_104), .A(n6425), .ZN(n6501) );
  INV_X1 U7146 ( .A(HOLD), .ZN(n6729) );
  OAI22_X1 U7147 ( .A1(n6729), .A2(keyinput_100), .B1(READREQUEST_REG_SCAN_IN), 
        .B2(keyinput_101), .ZN(n6426) );
  AOI221_X1 U7148 ( .B1(n6729), .B2(keyinput_100), .C1(keyinput_101), .C2(
        READREQUEST_REG_SCAN_IN), .A(n6426), .ZN(n6497) );
  OAI22_X1 U7149 ( .A1(n6428), .A2(keyinput_98), .B1(keyinput_97), .B2(NA_N), 
        .ZN(n6427) );
  AOI221_X1 U7150 ( .B1(n6428), .B2(keyinput_98), .C1(NA_N), .C2(keyinput_97), 
        .A(n6427), .ZN(n6494) );
  INV_X1 U7151 ( .A(keyinput_96), .ZN(n6492) );
  INV_X1 U7152 ( .A(keyinput_95), .ZN(n6490) );
  AOI22_X1 U7153 ( .A1(n6431), .A2(keyinput_89), .B1(keyinput_90), .B2(n6430), 
        .ZN(n6429) );
  OAI221_X1 U7154 ( .B1(n6431), .B2(keyinput_89), .C1(n6430), .C2(keyinput_90), 
        .A(n6429), .ZN(n6479) );
  INV_X1 U7155 ( .A(keyinput_88), .ZN(n6477) );
  INV_X1 U7156 ( .A(DATAI_21_), .ZN(n6433) );
  OAI22_X1 U7157 ( .A1(n6433), .A2(keyinput_74), .B1(DATAI_20_), .B2(
        keyinput_75), .ZN(n6432) );
  AOI221_X1 U7158 ( .B1(n6433), .B2(keyinput_74), .C1(keyinput_75), .C2(
        DATAI_20_), .A(n6432), .ZN(n6458) );
  INV_X1 U7159 ( .A(keyinput_73), .ZN(n6452) );
  INV_X1 U7160 ( .A(DATAI_23_), .ZN(n6449) );
  OAI22_X1 U7161 ( .A1(n6436), .A2(keyinput_67), .B1(n6435), .B2(keyinput_69), 
        .ZN(n6434) );
  AOI221_X1 U7162 ( .B1(n6436), .B2(keyinput_67), .C1(keyinput_69), .C2(n6435), 
        .A(n6434), .ZN(n6439) );
  OAI22_X1 U7163 ( .A1(DATAI_25_), .A2(keyinput_70), .B1(DATAI_24_), .B2(
        keyinput_71), .ZN(n6437) );
  AOI221_X1 U7164 ( .B1(DATAI_25_), .B2(keyinput_70), .C1(keyinput_71), .C2(
        DATAI_24_), .A(n6437), .ZN(n6438) );
  OAI211_X1 U7165 ( .C1(n6441), .C2(keyinput_68), .A(n6439), .B(n6438), .ZN(
        n6440) );
  AOI21_X1 U7166 ( .B1(n6441), .B2(keyinput_68), .A(n6440), .ZN(n6447) );
  INV_X1 U7167 ( .A(keyinput_66), .ZN(n6445) );
  AOI22_X1 U7168 ( .A1(DATAI_30_), .A2(keyinput_65), .B1(DATAI_31_), .B2(
        keyinput_64), .ZN(n6442) );
  OAI221_X1 U7169 ( .B1(DATAI_30_), .B2(keyinput_65), .C1(DATAI_31_), .C2(
        keyinput_64), .A(n6442), .ZN(n6443) );
  OAI221_X1 U7170 ( .B1(DATAI_29_), .B2(n6445), .C1(n6444), .C2(keyinput_66), 
        .A(n6443), .ZN(n6446) );
  AOI22_X1 U7171 ( .A1(keyinput_72), .A2(n6449), .B1(n6447), .B2(n6446), .ZN(
        n6448) );
  OAI21_X1 U7172 ( .B1(n6449), .B2(keyinput_72), .A(n6448), .ZN(n6450) );
  OAI221_X1 U7173 ( .B1(DATAI_22_), .B2(n6452), .C1(n6451), .C2(keyinput_73), 
        .A(n6450), .ZN(n6457) );
  XOR2_X1 U7174 ( .A(DATAI_17_), .B(keyinput_78), .Z(n6456) );
  INV_X1 U7175 ( .A(DATAI_18_), .ZN(n6454) );
  AOI22_X1 U7176 ( .A1(DATAI_19_), .A2(keyinput_76), .B1(n6454), .B2(
        keyinput_77), .ZN(n6453) );
  OAI221_X1 U7177 ( .B1(DATAI_19_), .B2(keyinput_76), .C1(n6454), .C2(
        keyinput_77), .A(n6453), .ZN(n6455) );
  AOI211_X1 U7178 ( .C1(n6458), .C2(n6457), .A(n6456), .B(n6455), .ZN(n6469)
         );
  AOI22_X1 U7179 ( .A1(n6461), .A2(keyinput_79), .B1(keyinput_80), .B2(n6460), 
        .ZN(n6459) );
  OAI221_X1 U7180 ( .B1(n6461), .B2(keyinput_79), .C1(n6460), .C2(keyinput_80), 
        .A(n6459), .ZN(n6468) );
  OAI22_X1 U7181 ( .A1(DATAI_14_), .A2(keyinput_81), .B1(DATAI_11_), .B2(
        keyinput_84), .ZN(n6462) );
  AOI221_X1 U7182 ( .B1(DATAI_14_), .B2(keyinput_81), .C1(keyinput_84), .C2(
        DATAI_11_), .A(n6462), .ZN(n6467) );
  OAI22_X1 U7183 ( .A1(n6465), .A2(keyinput_82), .B1(n6464), .B2(keyinput_85), 
        .ZN(n6463) );
  AOI221_X1 U7184 ( .B1(n6465), .B2(keyinput_82), .C1(keyinput_85), .C2(n6464), 
        .A(n6463), .ZN(n6466) );
  OAI211_X1 U7185 ( .C1(n6469), .C2(n6468), .A(n6467), .B(n6466), .ZN(n6472)
         );
  AOI22_X1 U7186 ( .A1(DATAI_9_), .A2(keyinput_86), .B1(DATAI_12_), .B2(
        keyinput_83), .ZN(n6470) );
  OAI221_X1 U7187 ( .B1(DATAI_9_), .B2(keyinput_86), .C1(DATAI_12_), .C2(
        keyinput_83), .A(n6470), .ZN(n6471) );
  OAI22_X1 U7188 ( .A1(keyinput_87), .A2(n6474), .B1(n6472), .B2(n6471), .ZN(
        n6473) );
  AOI21_X1 U7189 ( .B1(keyinput_87), .B2(n6474), .A(n6473), .ZN(n6475) );
  AOI221_X1 U7190 ( .B1(DATAI_7_), .B2(n6477), .C1(n6476), .C2(keyinput_88), 
        .A(n6475), .ZN(n6478) );
  OAI22_X1 U7191 ( .A1(keyinput_91), .A2(n6481), .B1(n6479), .B2(n6478), .ZN(
        n6480) );
  AOI21_X1 U7192 ( .B1(keyinput_91), .B2(n6481), .A(n6480), .ZN(n6486) );
  AOI22_X1 U7193 ( .A1(n6484), .A2(keyinput_92), .B1(keyinput_93), .B2(n6483), 
        .ZN(n6482) );
  OAI221_X1 U7194 ( .B1(n6484), .B2(keyinput_92), .C1(n6483), .C2(keyinput_93), 
        .A(n6482), .ZN(n6485) );
  AOI211_X1 U7195 ( .C1(DATAI_1_), .C2(keyinput_94), .A(n6486), .B(n6485), 
        .ZN(n6487) );
  OAI21_X1 U7196 ( .B1(DATAI_1_), .B2(keyinput_94), .A(n6487), .ZN(n6488) );
  OAI221_X1 U7197 ( .B1(DATAI_0_), .B2(n6490), .C1(n6489), .C2(keyinput_95), 
        .A(n6488), .ZN(n6491) );
  OAI221_X1 U7198 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_96), .C1(n7098), 
        .C2(n6492), .A(n6491), .ZN(n6493) );
  AOI22_X1 U7199 ( .A1(n6494), .A2(n6493), .B1(keyinput_99), .B2(READY_N), 
        .ZN(n6495) );
  OAI21_X1 U7200 ( .B1(keyinput_99), .B2(READY_N), .A(n6495), .ZN(n6496) );
  OAI211_X1 U7201 ( .C1(n6499), .C2(keyinput_102), .A(n6497), .B(n6496), .ZN(
        n6498) );
  AOI21_X1 U7202 ( .B1(n6499), .B2(keyinput_102), .A(n6498), .ZN(n6500) );
  OAI22_X1 U7203 ( .A1(n6501), .A2(n6500), .B1(n7080), .B2(keyinput_107), .ZN(
        n6502) );
  AOI21_X1 U7204 ( .B1(n7080), .B2(keyinput_107), .A(n6502), .ZN(n6510) );
  OAI22_X1 U7205 ( .A1(n6504), .A2(keyinput_105), .B1(keyinput_106), .B2(
        REQUESTPENDING_REG_SCAN_IN), .ZN(n6503) );
  AOI221_X1 U7206 ( .B1(n6504), .B2(keyinput_105), .C1(
        REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_106), .A(n6503), .ZN(n6509)
         );
  AOI22_X1 U7207 ( .A1(FLUSH_REG_SCAN_IN), .A2(keyinput_109), .B1(n6647), .B2(
        keyinput_111), .ZN(n6505) );
  OAI221_X1 U7208 ( .B1(FLUSH_REG_SCAN_IN), .B2(keyinput_109), .C1(n6647), 
        .C2(keyinput_111), .A(n6505), .ZN(n6508) );
  AOI22_X1 U7209 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput_110), .B1(
        MORE_REG_SCAN_IN), .B2(keyinput_108), .ZN(n6506) );
  OAI221_X1 U7210 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput_110), .C1(
        MORE_REG_SCAN_IN), .C2(keyinput_108), .A(n6506), .ZN(n6507) );
  AOI211_X1 U7211 ( .C1(n6510), .C2(n6509), .A(n6508), .B(n6507), .ZN(n6511)
         );
  AOI221_X1 U7212 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_112), .C1(
        n6642), .C2(n6512), .A(n6511), .ZN(n6513) );
  AOI221_X1 U7213 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_113), .C1(
        n6515), .C2(n6514), .A(n6513), .ZN(n6518) );
  AOI22_X1 U7214 ( .A1(BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_114), .B1(
        n6622), .B2(keyinput_116), .ZN(n6516) );
  OAI221_X1 U7215 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_114), .C1(
        n6622), .C2(keyinput_116), .A(n6516), .ZN(n6517) );
  AOI211_X1 U7216 ( .C1(REIP_REG_31__SCAN_IN), .C2(keyinput_115), .A(n6518), 
        .B(n6517), .ZN(n6519) );
  OAI21_X1 U7217 ( .B1(REIP_REG_31__SCAN_IN), .B2(keyinput_115), .A(n6519), 
        .ZN(n6520) );
  OAI211_X1 U7218 ( .C1(REIP_REG_28__SCAN_IN), .C2(keyinput_118), .A(n6521), 
        .B(n6520), .ZN(n6522) );
  AOI21_X1 U7219 ( .B1(REIP_REG_28__SCAN_IN), .B2(keyinput_118), .A(n6522), 
        .ZN(n6523) );
  OAI22_X1 U7220 ( .A1(keyinput_122), .A2(n6608), .B1(n6524), .B2(n6523), .ZN(
        n6525) );
  AOI21_X1 U7221 ( .B1(keyinput_122), .B2(n6608), .A(n6525), .ZN(n6527) );
  NAND2_X1 U7222 ( .A1(keyinput_125), .A2(REIP_REG_21__SCAN_IN), .ZN(n6526) );
  OAI221_X1 U7223 ( .B1(n6528), .B2(n6527), .C1(keyinput_125), .C2(
        REIP_REG_21__SCAN_IN), .A(n6526), .ZN(n6529) );
  AOI211_X1 U7224 ( .C1(n6532), .C2(n6531), .A(n6530), .B(n6529), .ZN(n6540)
         );
  INV_X1 U7225 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6536) );
  NAND2_X1 U7226 ( .A1(n6569), .A2(DATAO_REG_23__SCAN_IN), .ZN(n6535) );
  INV_X1 U7227 ( .A(n6533), .ZN(n7048) );
  NAND2_X1 U7228 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n7048), .ZN(n6534) );
  OAI211_X1 U7229 ( .C1(n6537), .C2(n6536), .A(n6535), .B(n6534), .ZN(n6538)
         );
  INV_X1 U7230 ( .A(n6538), .ZN(n6539) );
  XNOR2_X1 U7231 ( .A(n6540), .B(n6539), .ZN(U2900) );
  AOI22_X1 U7232 ( .A1(n7048), .A2(LWORD_REG_0__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6541) );
  OAI21_X1 U7233 ( .B1(n6542), .B2(n6572), .A(n6541), .ZN(U2923) );
  AOI22_X1 U7234 ( .A1(n7048), .A2(LWORD_REG_1__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6543) );
  OAI21_X1 U7235 ( .B1(n6544), .B2(n6572), .A(n6543), .ZN(U2922) );
  AOI22_X1 U7236 ( .A1(n7048), .A2(LWORD_REG_2__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6545) );
  OAI21_X1 U7237 ( .B1(n6546), .B2(n6572), .A(n6545), .ZN(U2921) );
  AOI22_X1 U7238 ( .A1(n7048), .A2(LWORD_REG_3__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U7239 ( .B1(n6548), .B2(n6572), .A(n6547), .ZN(U2920) );
  AOI22_X1 U7240 ( .A1(n7048), .A2(LWORD_REG_4__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6549) );
  OAI21_X1 U7241 ( .B1(n6550), .B2(n6572), .A(n6549), .ZN(U2919) );
  AOI22_X1 U7242 ( .A1(n7048), .A2(LWORD_REG_5__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6551) );
  OAI21_X1 U7243 ( .B1(n6552), .B2(n6572), .A(n6551), .ZN(U2918) );
  AOI22_X1 U7244 ( .A1(n7048), .A2(LWORD_REG_6__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6553) );
  OAI21_X1 U7245 ( .B1(n3862), .B2(n6572), .A(n6553), .ZN(U2917) );
  AOI22_X1 U7246 ( .A1(n7048), .A2(LWORD_REG_7__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6554) );
  OAI21_X1 U7247 ( .B1(n6555), .B2(n6572), .A(n6554), .ZN(U2916) );
  AOI22_X1 U7248 ( .A1(n7048), .A2(LWORD_REG_8__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U7249 ( .B1(n6557), .B2(n6572), .A(n6556), .ZN(U2915) );
  AOI22_X1 U7250 ( .A1(n7048), .A2(LWORD_REG_9__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6558) );
  OAI21_X1 U7251 ( .B1(n6559), .B2(n6572), .A(n6558), .ZN(U2914) );
  AOI22_X1 U7252 ( .A1(n7048), .A2(LWORD_REG_10__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6560) );
  OAI21_X1 U7253 ( .B1(n6561), .B2(n6572), .A(n6560), .ZN(U2913) );
  AOI22_X1 U7254 ( .A1(n7048), .A2(LWORD_REG_11__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6562) );
  OAI21_X1 U7255 ( .B1(n6563), .B2(n6572), .A(n6562), .ZN(U2912) );
  AOI22_X1 U7256 ( .A1(n6570), .A2(LWORD_REG_12__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6564) );
  OAI21_X1 U7257 ( .B1(n3945), .B2(n6572), .A(n6564), .ZN(U2911) );
  AOI22_X1 U7258 ( .A1(n6570), .A2(LWORD_REG_13__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6565) );
  OAI21_X1 U7259 ( .B1(n6566), .B2(n6572), .A(n6565), .ZN(U2910) );
  AOI22_X1 U7260 ( .A1(n6570), .A2(LWORD_REG_14__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6567) );
  OAI21_X1 U7261 ( .B1(n6568), .B2(n6572), .A(n6567), .ZN(U2909) );
  AOI22_X1 U7262 ( .A1(n6570), .A2(LWORD_REG_15__SCAN_IN), .B1(n6569), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6571) );
  OAI21_X1 U7263 ( .B1(n6573), .B2(n6572), .A(n6571), .ZN(U2908) );
  NAND2_X1 U7264 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7099), .ZN(n6621) );
  INV_X2 U7265 ( .A(n7099), .ZN(n7096) );
  NOR2_X2 U7266 ( .A1(STATE_REG_2__SCAN_IN), .A2(n7096), .ZN(n6619) );
  AOI22_X1 U7267 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n7096), .ZN(n6574) );
  OAI21_X1 U7268 ( .B1(n6757), .B2(n6621), .A(n6574), .ZN(U3184) );
  AOI22_X1 U7269 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n7096), .ZN(n6575) );
  OAI21_X1 U7270 ( .B1(n5342), .B2(n6621), .A(n6575), .ZN(U3185) );
  AOI22_X1 U7271 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n7096), .ZN(n6576) );
  OAI21_X1 U7272 ( .B1(n6577), .B2(n6621), .A(n6576), .ZN(U3186) );
  INV_X1 U7273 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6867) );
  AOI22_X1 U7274 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n7096), .ZN(n6578) );
  OAI21_X1 U7275 ( .B1(n6867), .B2(n6621), .A(n6578), .ZN(U3187) );
  AOI22_X1 U7276 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n7096), .ZN(n6579) );
  OAI21_X1 U7277 ( .B1(n6882), .B2(n6621), .A(n6579), .ZN(U3188) );
  INV_X1 U7278 ( .A(n6619), .ZN(n6618) );
  INV_X1 U7279 ( .A(n6621), .ZN(n6616) );
  AOI22_X1 U7280 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n7096), .ZN(n6580) );
  OAI21_X1 U7281 ( .B1(n6582), .B2(n6618), .A(n6580), .ZN(U3189) );
  AOI22_X1 U7282 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n7096), .ZN(n6581) );
  OAI21_X1 U7283 ( .B1(n6582), .B2(n6621), .A(n6581), .ZN(U3190) );
  AOI22_X1 U7284 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n7096), .ZN(n6583) );
  OAI21_X1 U7285 ( .B1(n6584), .B2(n6621), .A(n6583), .ZN(U3191) );
  AOI22_X1 U7286 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n7096), .ZN(n6585) );
  OAI21_X1 U7287 ( .B1(n5568), .B2(n6618), .A(n6585), .ZN(U3192) );
  AOI22_X1 U7288 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n7096), .ZN(n6586) );
  OAI21_X1 U7289 ( .B1(n6588), .B2(n6618), .A(n6586), .ZN(U3193) );
  AOI22_X1 U7290 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n7096), .ZN(n6587) );
  OAI21_X1 U7291 ( .B1(n6588), .B2(n6621), .A(n6587), .ZN(U3194) );
  AOI22_X1 U7292 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n7096), .ZN(n6589) );
  OAI21_X1 U7293 ( .B1(n6949), .B2(n6618), .A(n6589), .ZN(U3195) );
  AOI22_X1 U7294 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n7096), .ZN(n6590) );
  OAI21_X1 U7295 ( .B1(n6592), .B2(n6618), .A(n6590), .ZN(U3196) );
  AOI22_X1 U7296 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n7096), .ZN(n6591) );
  OAI21_X1 U7297 ( .B1(n6592), .B2(n6621), .A(n6591), .ZN(U3197) );
  AOI22_X1 U7298 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n7096), .ZN(n6593) );
  OAI21_X1 U7299 ( .B1(n6594), .B2(n6618), .A(n6593), .ZN(U3198) );
  AOI22_X1 U7300 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n7096), .ZN(n6595) );
  OAI21_X1 U7301 ( .B1(n6843), .B2(n6618), .A(n6595), .ZN(U3199) );
  AOI22_X1 U7302 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n7096), .ZN(n6596) );
  OAI21_X1 U7303 ( .B1(n6843), .B2(n6621), .A(n6596), .ZN(U3200) );
  AOI22_X1 U7304 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n7096), .ZN(n6597) );
  OAI21_X1 U7305 ( .B1(n6598), .B2(n6618), .A(n6597), .ZN(U3201) );
  AOI22_X1 U7306 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n7096), .ZN(n6599) );
  OAI21_X1 U7307 ( .B1(n6974), .B2(n6618), .A(n6599), .ZN(U3202) );
  AOI22_X1 U7308 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n7096), .ZN(n6600) );
  OAI21_X1 U7309 ( .B1(n6601), .B2(n6618), .A(n6600), .ZN(U3203) );
  AOI22_X1 U7310 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n7096), .ZN(n6602) );
  OAI21_X1 U7311 ( .B1(n6604), .B2(n6618), .A(n6602), .ZN(U3204) );
  AOI22_X1 U7312 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n7096), .ZN(n6603) );
  OAI21_X1 U7313 ( .B1(n6604), .B2(n6621), .A(n6603), .ZN(U3205) );
  AOI22_X1 U7314 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n7096), .ZN(n6605) );
  OAI21_X1 U7315 ( .B1(n6606), .B2(n6621), .A(n6605), .ZN(U3206) );
  AOI22_X1 U7316 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n7096), .ZN(n6607) );
  OAI21_X1 U7317 ( .B1(n6608), .B2(n6621), .A(n6607), .ZN(U3207) );
  AOI22_X1 U7318 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n7096), .ZN(n6609) );
  OAI21_X1 U7319 ( .B1(n6610), .B2(n6621), .A(n6609), .ZN(U3208) );
  AOI22_X1 U7320 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n7096), .ZN(n6611) );
  OAI21_X1 U7321 ( .B1(n6613), .B2(n6618), .A(n6611), .ZN(U3209) );
  AOI22_X1 U7322 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n7096), .ZN(n6612) );
  OAI21_X1 U7323 ( .B1(n6613), .B2(n6621), .A(n6612), .ZN(U3210) );
  AOI22_X1 U7324 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n7096), .ZN(n6614) );
  OAI21_X1 U7325 ( .B1(n6615), .B2(n6621), .A(n6614), .ZN(U3211) );
  AOI22_X1 U7326 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6616), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n7096), .ZN(n6617) );
  OAI21_X1 U7327 ( .B1(n6622), .B2(n6618), .A(n6617), .ZN(U3212) );
  AOI22_X1 U7328 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6619), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n7096), .ZN(n6620) );
  OAI21_X1 U7329 ( .B1(n6622), .B2(n6621), .A(n6620), .ZN(U3213) );
  MUX2_X1 U7330 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n7099), .Z(U3445) );
  NOR4_X1 U7331 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6632) );
  NOR4_X1 U7332 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n6631) );
  INV_X1 U7333 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n7082) );
  NOR4_X1 U7334 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_27__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6623) );
  OAI21_X1 U7335 ( .B1(n6639), .B2(n7082), .A(n6623), .ZN(n6629) );
  NOR4_X1 U7336 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_12__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(
        DATAWIDTH_REG_10__SCAN_IN), .ZN(n6627) );
  NOR4_X1 U7337 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_14__SCAN_IN), .ZN(n6626) );
  NOR4_X1 U7338 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(
        n6625) );
  NOR4_X1 U7339 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_6__SCAN_IN), .ZN(
        n6624) );
  NAND4_X1 U7340 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6628)
         );
  NOR4_X1 U7341 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(
        DATAWIDTH_REG_30__SCAN_IN), .A3(n6629), .A4(n6628), .ZN(n6630) );
  NAND3_X1 U7342 ( .A1(n6632), .A2(n6631), .A3(n6630), .ZN(n6646) );
  INV_X1 U7343 ( .A(n6646), .ZN(n6637) );
  INV_X1 U7344 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6633) );
  NOR2_X1 U7345 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6646), .ZN(n6643) );
  NAND2_X1 U7346 ( .A1(n6643), .A2(n7082), .ZN(n6640) );
  NOR2_X1 U7347 ( .A1(REIP_REG_0__SCAN_IN), .A2(n6646), .ZN(n6634) );
  NAND3_X1 U7348 ( .A1(n6634), .A2(n6639), .A3(n7082), .ZN(n6641) );
  OAI211_X1 U7349 ( .C1(n6637), .C2(n6633), .A(n6640), .B(n6641), .ZN(U2795)
         );
  MUX2_X1 U7350 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n7099), .Z(U3446) );
  NAND2_X1 U7351 ( .A1(n6634), .A2(n6757), .ZN(n6644) );
  AOI21_X1 U7352 ( .B1(REIP_REG_0__SCAN_IN), .B2(REIP_REG_1__SCAN_IN), .A(
        n6646), .ZN(n6635) );
  INV_X1 U7353 ( .A(n6635), .ZN(n6636) );
  OAI21_X1 U7354 ( .B1(BYTEENABLE_REG_2__SCAN_IN), .B2(n6637), .A(n6636), .ZN(
        n6638) );
  OAI221_X1 U7355 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6640), .C1(n6639), 
        .C2(n6644), .A(n6638), .ZN(U3468) );
  MUX2_X1 U7356 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n7099), .Z(U3447) );
  OAI221_X1 U7357 ( .B1(n6643), .B2(n6642), .C1(n6643), .C2(n6646), .A(n6641), 
        .ZN(U2794) );
  MUX2_X1 U7358 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n7099), .Z(U3448) );
  INV_X1 U7359 ( .A(n6644), .ZN(n6645) );
  AOI21_X1 U7360 ( .B1(n6647), .B2(n6646), .A(n6645), .ZN(U3469) );
  INV_X1 U7361 ( .A(n6648), .ZN(n6992) );
  AOI22_X1 U7362 ( .A1(n7110), .A2(n6660), .B1(n6649), .B2(n6992), .ZN(n6650)
         );
  OAI21_X1 U7363 ( .B1(n6663), .B2(n6651), .A(n6650), .ZN(U2838) );
  NAND2_X1 U7364 ( .A1(n5991), .A2(n6652), .ZN(n6653) );
  NOR2_X1 U7365 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  OR2_X1 U7366 ( .A1(n6657), .A2(n6656), .ZN(n6969) );
  NOR2_X1 U7367 ( .A1(n6969), .A2(n6658), .ZN(n6659) );
  AOI21_X1 U7368 ( .B1(n7107), .B2(n6660), .A(n6659), .ZN(n6661) );
  OAI21_X1 U7369 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(U2840) );
  AOI22_X1 U7370 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_2__SCAN_IN), .ZN(n6670) );
  XNOR2_X1 U7371 ( .A(n6664), .B(n6806), .ZN(n6665) );
  XNOR2_X1 U7372 ( .A(n6666), .B(n6665), .ZN(n6799) );
  INV_X1 U7373 ( .A(n6799), .ZN(n6668) );
  AOI22_X1 U7374 ( .A1(n6668), .A2(n6714), .B1(n6713), .B2(n6667), .ZN(n6669)
         );
  OAI211_X1 U7375 ( .C1(n6717), .C2(n6671), .A(n6670), .B(n6669), .ZN(U2984)
         );
  AOI22_X1 U7376 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_3__SCAN_IN), .ZN(n6678) );
  XNOR2_X1 U7377 ( .A(n6672), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6673)
         );
  XNOR2_X1 U7378 ( .A(n6674), .B(n6673), .ZN(n6773) );
  INV_X1 U7379 ( .A(n6675), .ZN(n6676) );
  AOI22_X1 U7380 ( .A1(n6714), .A2(n6773), .B1(n6676), .B2(n6713), .ZN(n6677)
         );
  OAI211_X1 U7381 ( .C1(n6717), .C2(n6679), .A(n6678), .B(n6677), .ZN(U2983)
         );
  AOI22_X1 U7382 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U7383 ( .A1(n6681), .A2(n6682), .ZN(n6683) );
  AND2_X1 U7384 ( .A1(n6680), .A2(n6683), .ZN(n6767) );
  AOI22_X1 U7385 ( .A1(n6767), .A2(n6714), .B1(n6713), .B2(n6875), .ZN(n6684)
         );
  OAI211_X1 U7386 ( .C1(n6717), .C2(n6878), .A(n6685), .B(n6684), .ZN(U2982)
         );
  AOI22_X1 U7387 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U7388 ( .A1(n6680), .A2(n6686), .ZN(n6689) );
  NAND2_X1 U7389 ( .A1(n6689), .A2(n6687), .ZN(n6688) );
  OAI21_X1 U7390 ( .B1(n6689), .B2(n6687), .A(n6688), .ZN(n6690) );
  INV_X1 U7391 ( .A(n6690), .ZN(n6784) );
  AOI22_X1 U7392 ( .A1(n6784), .A2(n6714), .B1(n6713), .B2(n6885), .ZN(n6691)
         );
  OAI211_X1 U7393 ( .C1(n6717), .C2(n6889), .A(n6692), .B(n6691), .ZN(U2981)
         );
  AOI22_X1 U7394 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n6695) );
  AOI22_X1 U7395 ( .A1(n6931), .A2(n6713), .B1(n6930), .B2(n6693), .ZN(n6694)
         );
  OAI211_X1 U7396 ( .C1(n6697), .C2(n6696), .A(n6695), .B(n6694), .ZN(U2974)
         );
  AOI22_X1 U7397 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_17__SCAN_IN), .ZN(n6705) );
  INV_X1 U7398 ( .A(n6698), .ZN(n6701) );
  NAND3_X1 U7399 ( .A1(n6703), .A2(n6702), .A3(n6699), .ZN(n6700) );
  OAI211_X1 U7400 ( .C1(n6703), .C2(n6702), .A(n6701), .B(n6700), .ZN(n6846)
         );
  AOI22_X1 U7401 ( .A1(n6846), .A2(n6714), .B1(n6713), .B2(n7101), .ZN(n6704)
         );
  OAI211_X1 U7402 ( .C1(n6717), .C2(n6706), .A(n6705), .B(n6704), .ZN(U2969)
         );
  AOI22_X1 U7403 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n6707), .B1(n6771), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6716) );
  INV_X1 U7404 ( .A(n6708), .ZN(n6712) );
  INV_X1 U7405 ( .A(n6709), .ZN(n6711) );
  OAI21_X1 U7406 ( .B1(n6712), .B2(n6711), .A(n6710), .ZN(n6750) );
  AOI22_X1 U7407 ( .A1(n6750), .A2(n6714), .B1(n6713), .B2(n7107), .ZN(n6715)
         );
  OAI211_X1 U7408 ( .C1(n6717), .C2(n6973), .A(n6716), .B(n6715), .ZN(U2967)
         );
  INV_X1 U7409 ( .A(n6718), .ZN(n6719) );
  OAI21_X1 U7410 ( .B1(n6719), .B2(n7077), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6720) );
  OAI21_X1 U7411 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6721), .A(n6720), .ZN(
        U2790) );
  NOR2_X1 U7412 ( .A1(n7099), .A2(D_C_N_REG_SCAN_IN), .ZN(n6722) );
  AOI22_X1 U7413 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(n7099), .B1(n6723), .B2(
        n6722), .ZN(U2791) );
  INV_X1 U7414 ( .A(n6724), .ZN(n6725) );
  NOR3_X1 U7415 ( .A1(n6739), .A2(n6725), .A3(READREQUEST_REG_SCAN_IN), .ZN(
        n6726) );
  AOI21_X1 U7416 ( .B1(n6739), .B2(n6727), .A(n6726), .ZN(U3474) );
  AOI22_X1 U7417 ( .A1(n7099), .A2(READREQUEST_REG_SCAN_IN), .B1(n6728), .B2(
        n7096), .ZN(U3470) );
  NOR2_X1 U7418 ( .A1(n6730), .A2(n6729), .ZN(n7085) );
  AOI22_X1 U7419 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        STATE_REG_0__SCAN_IN), .B2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6734) );
  NOR2_X1 U7420 ( .A1(n6731), .A2(n7088), .ZN(n7091) );
  INV_X1 U7421 ( .A(n7091), .ZN(n6732) );
  OAI211_X1 U7422 ( .C1(n7085), .C2(n6734), .A(n6733), .B(n6732), .ZN(U3182)
         );
  NOR2_X1 U7423 ( .A1(READY_N), .A2(n7072), .ZN(n6735) );
  AOI21_X1 U7424 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6735), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6737) );
  OAI21_X1 U7425 ( .B1(n6738), .B2(n6737), .A(n6736), .ZN(U3150) );
  INV_X1 U7426 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6747) );
  AOI211_X1 U7427 ( .C1(n7048), .C2(n7088), .A(n6740), .B(n6739), .ZN(n6746)
         );
  OAI21_X1 U7428 ( .B1(n6741), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n6742) );
  OAI21_X1 U7429 ( .B1(n6743), .B2(n6742), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n6745) );
  NOR2_X1 U7430 ( .A1(n6746), .A2(n7070), .ZN(n6744) );
  AOI22_X1 U7431 ( .A1(n6747), .A2(n6746), .B1(n6745), .B2(n6744), .ZN(U3472)
         );
  AOI22_X1 U7432 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n6748), .B1(n6771), .B2(REIP_REG_19__SCAN_IN), .ZN(n6752) );
  INV_X1 U7433 ( .A(n6969), .ZN(n6749) );
  AOI22_X1 U7434 ( .A1(n6750), .A2(n6854), .B1(n6860), .B2(n6749), .ZN(n6751)
         );
  OAI211_X1 U7435 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n6753), .A(n6752), .B(n6751), .ZN(U2999) );
  INV_X1 U7436 ( .A(n6754), .ZN(n6756) );
  NAND2_X1 U7437 ( .A1(n6756), .A2(n6755), .ZN(n6765) );
  AOI21_X1 U7438 ( .B1(n6855), .B2(n6856), .A(n6857), .ZN(n6763) );
  OAI22_X1 U7439 ( .A1(n6793), .A2(n6758), .B1(n6757), .B2(n4480), .ZN(n6761)
         );
  NOR2_X1 U7440 ( .A1(n6800), .A2(n6759), .ZN(n6760) );
  NOR2_X1 U7441 ( .A1(n6761), .A2(n6760), .ZN(n6762) );
  OAI221_X1 U7442 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6765), .C1(n6764), .C2(n6763), .A(n6762), .ZN(U3017) );
  OAI22_X1 U7443 ( .A1(n6793), .A2(n6869), .B1(n6867), .B2(n4480), .ZN(n6766)
         );
  AOI21_X1 U7444 ( .B1(n6767), .B2(n6854), .A(n6766), .ZN(n6769) );
  OAI211_X1 U7445 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6774), .B(n6779), .ZN(n6768) );
  OAI211_X1 U7446 ( .C1(n6778), .C2(n6770), .A(n6769), .B(n6768), .ZN(U3014)
         );
  AOI22_X1 U7447 ( .A1(n6860), .A2(n6772), .B1(n6771), .B2(REIP_REG_3__SCAN_IN), .ZN(n6776) );
  AOI22_X1 U7448 ( .A1(n6774), .A2(n6777), .B1(n6854), .B2(n6773), .ZN(n6775)
         );
  OAI211_X1 U7449 ( .C1(n6778), .C2(n6777), .A(n6776), .B(n6775), .ZN(U3015)
         );
  NOR2_X1 U7450 ( .A1(n6779), .A2(n6795), .ZN(n6782) );
  OAI22_X1 U7451 ( .A1(n6793), .A2(n6780), .B1(n6882), .B2(n4480), .ZN(n6781)
         );
  AOI21_X1 U7452 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(n6789) );
  AOI22_X1 U7453 ( .A1(n6785), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .B1(n6854), 
        .B2(n6784), .ZN(n6788) );
  INV_X1 U7454 ( .A(n6786), .ZN(n6787) );
  NAND3_X1 U7455 ( .A1(n6789), .A2(n6788), .A3(n6787), .ZN(U3013) );
  INV_X1 U7456 ( .A(n6790), .ZN(n6791) );
  NAND2_X1 U7457 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6791), .ZN(n6807)
         );
  OAI22_X1 U7458 ( .A1(n6793), .A2(n6792), .B1(n5342), .B2(n4480), .ZN(n6803)
         );
  INV_X1 U7459 ( .A(n6794), .ZN(n6796) );
  AOI21_X1 U7460 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6796), .A(n6795), 
        .ZN(n6797) );
  NOR2_X1 U7461 ( .A1(n6798), .A2(n6797), .ZN(n6802) );
  NOR2_X1 U7462 ( .A1(n6800), .A2(n6799), .ZN(n6801) );
  NOR3_X1 U7463 ( .A1(n6803), .A2(n6802), .A3(n6801), .ZN(n6804) );
  OAI221_X1 U7464 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n6807), .C1(n6806), .C2(n6805), .A(n6804), .ZN(U3016) );
  INV_X1 U7465 ( .A(n6808), .ZN(n6816) );
  AOI21_X1 U7466 ( .B1(n6860), .B2(n6892), .A(n6809), .ZN(n6812) );
  NAND2_X1 U7467 ( .A1(n6810), .A2(n6854), .ZN(n6811) );
  OAI211_X1 U7468 ( .C1(n6813), .C2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6812), 
        .B(n6811), .ZN(n6814) );
  INV_X1 U7469 ( .A(n6814), .ZN(n6815) );
  OAI21_X1 U7470 ( .B1(n6817), .B2(n6816), .A(n6815), .ZN(U3011) );
  AOI21_X1 U7471 ( .B1(n6860), .B2(n6903), .A(n6818), .ZN(n6822) );
  AOI22_X1 U7472 ( .A1(n6820), .A2(n6854), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6819), .ZN(n6821) );
  OAI211_X1 U7473 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6823), .A(n6822), 
        .B(n6821), .ZN(U3009) );
  AOI21_X1 U7474 ( .B1(n6860), .B2(n6825), .A(n6824), .ZN(n6829) );
  INV_X1 U7475 ( .A(n6842), .ZN(n6826) );
  AOI22_X1 U7476 ( .A1(n6827), .A2(n6854), .B1(n6830), .B2(n6826), .ZN(n6828)
         );
  OAI211_X1 U7477 ( .C1(n6831), .C2(n6830), .A(n6829), .B(n6828), .ZN(U3007)
         );
  AOI21_X1 U7478 ( .B1(n6860), .B2(n6833), .A(n6832), .ZN(n6840) );
  AOI22_X1 U7479 ( .A1(n6835), .A2(n6854), .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n6834), .ZN(n6839) );
  OAI221_X1 U7480 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .C1(n6105), .C2(n6837), .A(n6836), 
        .ZN(n6838) );
  NAND3_X1 U7481 ( .A1(n6840), .A2(n6839), .A3(n6838), .ZN(U3002) );
  NOR3_X1 U7482 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6842), .A3(n6841), 
        .ZN(n6845) );
  NOR2_X1 U7483 ( .A1(n4480), .A2(n6843), .ZN(n6844) );
  AOI211_X1 U7484 ( .C1(n6846), .C2(n6854), .A(n6845), .B(n6844), .ZN(n6851)
         );
  INV_X1 U7485 ( .A(n6847), .ZN(n6848) );
  AOI22_X1 U7486 ( .A1(n6849), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n6860), .B2(n6848), .ZN(n6850) );
  NAND2_X1 U7487 ( .A1(n6851), .A2(n6850), .ZN(U3001) );
  INV_X1 U7488 ( .A(n6852), .ZN(n6853) );
  AOI22_X1 U7489 ( .A1(n6856), .A2(n6855), .B1(n6854), .B2(n6853), .ZN(n6864)
         );
  OAI21_X1 U7490 ( .B1(n6858), .B2(n6857), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6862) );
  NAND2_X1 U7491 ( .A1(n6860), .A2(n6859), .ZN(n6861) );
  NAND4_X1 U7492 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(U3018)
         );
  OAI22_X1 U7493 ( .A1(n6867), .A2(n6866), .B1(n7013), .B2(n6865), .ZN(n6868)
         );
  AOI211_X1 U7494 ( .C1(n6968), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6967), 
        .B(n6868), .ZN(n6877) );
  NOR2_X1 U7495 ( .A1(n7004), .A2(n6869), .ZN(n6874) );
  NAND3_X1 U7496 ( .A1(n6998), .A2(n6870), .A3(n6867), .ZN(n6871) );
  OAI21_X1 U7497 ( .B1(n6914), .B2(n6872), .A(n6871), .ZN(n6873) );
  AOI211_X1 U7498 ( .C1(n6886), .C2(n6875), .A(n6874), .B(n6873), .ZN(n6876)
         );
  OAI211_X1 U7499 ( .C1(n6878), .C2(n7010), .A(n6877), .B(n6876), .ZN(U2823)
         );
  AOI22_X1 U7500 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6968), .B1(n6993), 
        .B2(n6879), .ZN(n6880) );
  INV_X1 U7501 ( .A(n6880), .ZN(n6881) );
  AOI211_X1 U7502 ( .C1(n7003), .C2(EBX_REG_5__SCAN_IN), .A(n6967), .B(n6881), 
        .ZN(n6888) );
  OAI21_X1 U7503 ( .B1(n6986), .B2(n6883), .A(n6882), .ZN(n6884) );
  AOI22_X1 U7504 ( .A1(n6886), .A2(n6885), .B1(n6898), .B2(n6884), .ZN(n6887)
         );
  OAI211_X1 U7505 ( .C1(n6889), .C2(n7010), .A(n6888), .B(n6887), .ZN(U2822)
         );
  INV_X1 U7506 ( .A(n6890), .ZN(n6897) );
  NOR3_X1 U7507 ( .A1(n6986), .A2(REIP_REG_7__SCAN_IN), .A3(n6891), .ZN(n6896)
         );
  INV_X1 U7508 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6894) );
  AOI22_X1 U7509 ( .A1(EBX_REG_7__SCAN_IN), .A2(n7003), .B1(n6993), .B2(n6892), 
        .ZN(n6893) );
  OAI211_X1 U7510 ( .C1(n6999), .C2(n6894), .A(n6893), .B(n6944), .ZN(n6895)
         );
  AOI211_X1 U7511 ( .C1(n7007), .C2(n6897), .A(n6896), .B(n6895), .ZN(n6901)
         );
  OAI21_X1 U7512 ( .B1(n6899), .B2(n6898), .A(REIP_REG_7__SCAN_IN), .ZN(n6900)
         );
  OAI211_X1 U7513 ( .C1(n7010), .C2(n6902), .A(n6901), .B(n6900), .ZN(U2820)
         );
  AOI22_X1 U7514 ( .A1(PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n6968), .B1(n6993), 
        .B2(n6903), .ZN(n6912) );
  NOR3_X1 U7515 ( .A1(n6986), .A2(REIP_REG_9__SCAN_IN), .A3(n6904), .ZN(n6922)
         );
  AND2_X1 U7516 ( .A1(n6921), .A2(REIP_REG_9__SCAN_IN), .ZN(n6905) );
  AOI211_X1 U7517 ( .C1(n7003), .C2(EBX_REG_9__SCAN_IN), .A(n6922), .B(n6905), 
        .ZN(n6911) );
  INV_X1 U7518 ( .A(n6906), .ZN(n6909) );
  INV_X1 U7519 ( .A(n6907), .ZN(n6908) );
  AOI22_X1 U7520 ( .A1(n6909), .A2(n7007), .B1(n6908), .B2(n6981), .ZN(n6910)
         );
  NAND4_X1 U7521 ( .A1(n6912), .A2(n6911), .A3(n6910), .A4(n6944), .ZN(U2818)
         );
  OAI22_X1 U7522 ( .A1(n6915), .A2(n6914), .B1(n7004), .B2(n6913), .ZN(n6916)
         );
  AOI211_X1 U7523 ( .C1(n6968), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6967), 
        .B(n6916), .ZN(n6927) );
  INV_X1 U7524 ( .A(n6917), .ZN(n6918) );
  OAI22_X1 U7525 ( .A1(n6919), .A2(n6978), .B1(n7010), .B2(n6918), .ZN(n6920)
         );
  INV_X1 U7526 ( .A(n6920), .ZN(n6926) );
  OAI21_X1 U7527 ( .B1(n6922), .B2(n6921), .A(REIP_REG_10__SCAN_IN), .ZN(n6925) );
  NAND3_X1 U7528 ( .A1(n6998), .A2(n6923), .A3(n5568), .ZN(n6924) );
  NAND4_X1 U7529 ( .A1(n6927), .A2(n6926), .A3(n6925), .A4(n6924), .ZN(U2817)
         );
  AOI22_X1 U7530 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6928), .B1(n6953), .B2(
        n6939), .ZN(n6935) );
  AOI22_X1 U7531 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6968), .B1(n6993), 
        .B2(n6929), .ZN(n6934) );
  AOI21_X1 U7532 ( .B1(n7003), .B2(EBX_REG_12__SCAN_IN), .A(n6967), .ZN(n6933)
         );
  AOI22_X1 U7533 ( .A1(n6931), .A2(n7007), .B1(n6930), .B2(n6981), .ZN(n6932)
         );
  NAND4_X1 U7534 ( .A1(n6935), .A2(n6934), .A3(n6933), .A4(n6932), .ZN(U2815)
         );
  INV_X1 U7535 ( .A(n6936), .ZN(n6937) );
  AOI22_X1 U7536 ( .A1(n6938), .A2(n7007), .B1(n6981), .B2(n6937), .ZN(n6952)
         );
  NOR2_X1 U7537 ( .A1(n6939), .A2(n6942), .ZN(n6950) );
  OAI22_X1 U7538 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6942), .B1(n6941), .B2(
        n6940), .ZN(n6948) );
  AOI22_X1 U7539 ( .A1(EBX_REG_13__SCAN_IN), .A2(n7003), .B1(n6993), .B2(n6943), .ZN(n6945) );
  OAI211_X1 U7540 ( .C1(n6999), .C2(n6946), .A(n6945), .B(n6944), .ZN(n6947)
         );
  AOI221_X1 U7541 ( .B1(n6950), .B2(n6949), .C1(n6948), .C2(
        REIP_REG_13__SCAN_IN), .A(n6947), .ZN(n6951) );
  NAND2_X1 U7542 ( .A1(n6952), .A2(n6951), .ZN(U2814) );
  NAND2_X1 U7543 ( .A1(n6954), .A2(n6953), .ZN(n6965) );
  AOI22_X1 U7544 ( .A1(EBX_REG_18__SCAN_IN), .A2(n7003), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6962), .ZN(n6955) );
  OAI21_X1 U7545 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6965), .A(n6955), .ZN(n6956) );
  AOI211_X1 U7546 ( .C1(n6968), .C2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6967), 
        .B(n6956), .ZN(n6959) );
  AOI22_X1 U7547 ( .A1(n7104), .A2(n7007), .B1(n6981), .B2(n6957), .ZN(n6958)
         );
  OAI211_X1 U7548 ( .C1(n7004), .C2(n6960), .A(n6959), .B(n6958), .ZN(U2809)
         );
  NAND2_X1 U7549 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n6961) );
  OAI21_X1 U7550 ( .B1(REIP_REG_18__SCAN_IN), .B2(REIP_REG_19__SCAN_IN), .A(
        n6961), .ZN(n6964) );
  AOI22_X1 U7551 ( .A1(EBX_REG_19__SCAN_IN), .A2(n7003), .B1(
        REIP_REG_19__SCAN_IN), .B2(n6962), .ZN(n6963) );
  OAI21_X1 U7552 ( .B1(n6965), .B2(n6964), .A(n6963), .ZN(n6966) );
  AOI211_X1 U7553 ( .C1(n6968), .C2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n6967), 
        .B(n6966), .ZN(n6972) );
  NOR2_X1 U7554 ( .A1(n6969), .A2(n7004), .ZN(n6970) );
  AOI21_X1 U7555 ( .B1(n7107), .B2(n7007), .A(n6970), .ZN(n6971) );
  OAI211_X1 U7556 ( .C1(n6973), .C2(n7010), .A(n6972), .B(n6971), .ZN(U2808)
         );
  OAI21_X1 U7557 ( .B1(n6986), .B2(n6975), .A(n6974), .ZN(n6976) );
  AOI22_X1 U7558 ( .A1(EBX_REG_20__SCAN_IN), .A2(n7003), .B1(n6991), .B2(n6976), .ZN(n6984) );
  OAI22_X1 U7559 ( .A1(n6979), .A2(n6978), .B1(n7004), .B2(n6977), .ZN(n6980)
         );
  AOI21_X1 U7560 ( .B1(n6982), .B2(n6981), .A(n6980), .ZN(n6983) );
  OAI211_X1 U7561 ( .C1(n6985), .C2(n6999), .A(n6984), .B(n6983), .ZN(U2807)
         );
  NOR2_X1 U7562 ( .A1(n6986), .A2(REIP_REG_21__SCAN_IN), .ZN(n6987) );
  AOI22_X1 U7563 ( .A1(EBX_REG_21__SCAN_IN), .A2(n7003), .B1(n6988), .B2(n6987), .ZN(n6989) );
  OAI21_X1 U7564 ( .B1(n4117), .B2(n6999), .A(n6989), .ZN(n6990) );
  AOI21_X1 U7565 ( .B1(REIP_REG_21__SCAN_IN), .B2(n6991), .A(n6990), .ZN(n6995) );
  AOI22_X1 U7566 ( .A1(n7110), .A2(n7007), .B1(n6993), .B2(n6992), .ZN(n6994)
         );
  OAI211_X1 U7567 ( .C1(n6996), .C2(n7010), .A(n6995), .B(n6994), .ZN(U2806)
         );
  AOI21_X1 U7568 ( .B1(n6998), .B2(n6997), .A(REIP_REG_23__SCAN_IN), .ZN(n7001) );
  OAI22_X1 U7569 ( .A1(n7001), .A2(n7000), .B1(n4145), .B2(n6999), .ZN(n7002)
         );
  AOI21_X1 U7570 ( .B1(EBX_REG_23__SCAN_IN), .B2(n7003), .A(n7002), .ZN(n7009)
         );
  NOR2_X1 U7571 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  AOI21_X1 U7572 ( .B1(n7115), .B2(n7007), .A(n7006), .ZN(n7008) );
  OAI211_X1 U7573 ( .C1(n7011), .C2(n7010), .A(n7009), .B(n7008), .ZN(U2804)
         );
  OAI21_X1 U7574 ( .B1(n7012), .B2(n7037), .A(n6696), .ZN(U2793) );
  INV_X1 U7575 ( .A(n7013), .ZN(n7014) );
  NAND4_X1 U7576 ( .A1(n7016), .A2(n7015), .A3(n7055), .A4(n7014), .ZN(n7017)
         );
  OAI21_X1 U7577 ( .B1(n7018), .B2(n4203), .A(n7017), .ZN(U3455) );
  INV_X1 U7578 ( .A(n7019), .ZN(n7022) );
  NOR3_X1 U7579 ( .A1(n7022), .A2(n7021), .A3(n7020), .ZN(n7024) );
  NAND2_X1 U7580 ( .A1(n7024), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n7028) );
  INV_X1 U7581 ( .A(n7023), .ZN(n7025) );
  OAI22_X1 U7582 ( .A1(n7026), .A2(n7025), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n7024), .ZN(n7027) );
  NAND2_X1 U7583 ( .A1(n7028), .A2(n7027), .ZN(n7029) );
  AOI222_X1 U7584 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n7030), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n7029), .C1(n7030), .C2(n7029), 
        .ZN(n7032) );
  AOI222_X1 U7585 ( .A1(n7032), .A2(n4200), .B1(n7032), .B2(n7031), .C1(n4200), 
        .C2(n7031), .ZN(n7033) );
  OR2_X1 U7586 ( .A1(n7033), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n7046)
         );
  NOR2_X1 U7587 ( .A1(n7035), .A2(n7034), .ZN(n7041) );
  NAND2_X1 U7588 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  NAND2_X1 U7589 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  NAND3_X1 U7590 ( .A1(n7042), .A2(n7041), .A3(n7040), .ZN(n7043) );
  NOR2_X1 U7591 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  NAND2_X1 U7592 ( .A1(n7078), .A2(n7047), .ZN(n7050) );
  NAND2_X1 U7593 ( .A1(READY_N), .A2(n7048), .ZN(n7049) );
  NAND2_X1 U7594 ( .A1(n7050), .A2(n7049), .ZN(n7054) );
  OR2_X1 U7595 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  AOI221_X1 U7596 ( .B1(n7067), .B2(n7088), .C1(n7067), .C2(
        STATE2_REG_2__SCAN_IN), .A(n7072), .ZN(n7071) );
  INV_X1 U7597 ( .A(n7071), .ZN(n7061) );
  NAND3_X1 U7598 ( .A1(n7055), .A2(STATE2_REG_0__SCAN_IN), .A3(n7088), .ZN(
        n7056) );
  NAND3_X1 U7599 ( .A1(n7056), .A2(n7077), .A3(n7067), .ZN(n7057) );
  OAI21_X1 U7600 ( .B1(n7058), .B2(n7067), .A(n7057), .ZN(n7060) );
  OAI211_X1 U7601 ( .C1(n7062), .C2(n7061), .A(n7060), .B(n7059), .ZN(U3149)
         );
  INV_X1 U7602 ( .A(n7063), .ZN(n7065) );
  OAI211_X1 U7603 ( .C1(n7067), .C2(n7066), .A(n7065), .B(n7064), .ZN(U3453)
         );
  AOI21_X1 U7604 ( .B1(n7070), .B2(n7069), .A(n7068), .ZN(n7073) );
  AOI221_X1 U7605 ( .B1(n7074), .B2(STATE2_REG_0__SCAN_IN), .C1(n7073), .C2(
        n7072), .A(n7071), .ZN(n7076) );
  OAI211_X1 U7606 ( .C1(n7078), .C2(n7077), .A(n7076), .B(n7075), .ZN(U3148)
         );
  INV_X1 U7607 ( .A(n7079), .ZN(n7081) );
  OAI21_X1 U7608 ( .B1(n7083), .B2(n7080), .A(n7081), .ZN(U2792) );
  OAI21_X1 U7609 ( .B1(n7083), .B2(n7082), .A(n7081), .ZN(U3452) );
  NAND2_X1 U7610 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n7087) );
  NAND2_X1 U7611 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_1__SCAN_IN), .ZN(
        n7084) );
  AOI221_X1 U7612 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n7090), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n7094) );
  AOI221_X1 U7613 ( .B1(n7085), .B2(n7084), .C1(n7091), .C2(n7084), .A(n7094), 
        .ZN(n7086) );
  OAI221_X1 U7614 ( .B1(n7099), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n7099), 
        .C2(n7087), .A(n7086), .ZN(U3181) );
  AOI221_X1 U7615 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n7088), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n7089) );
  AOI221_X1 U7616 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n7089), .C2(HOLD), .A(n4357), .ZN(n7095) );
  NAND4_X1 U7617 ( .A1(REQUESTPENDING_REG_SCAN_IN), .A2(STATE_REG_0__SCAN_IN), 
        .A3(n7091), .A4(n7090), .ZN(n7093) );
  NAND3_X1 U7618 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n7092) );
  OAI211_X1 U7619 ( .C1(n7095), .C2(n7094), .A(n7093), .B(n7092), .ZN(U3183)
         );
  AOI22_X1 U7620 ( .A1(n7099), .A2(n7098), .B1(n7097), .B2(n7096), .ZN(U3473)
         );
  INV_X1 U7621 ( .A(n7100), .ZN(n7114) );
  AOI22_X1 U7622 ( .A1(n7101), .A2(n7114), .B1(n7113), .B2(DATAI_17_), .ZN(
        n7103) );
  AOI22_X1 U7623 ( .A1(n7117), .A2(DATAI_1_), .B1(n7116), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n7102) );
  NAND2_X1 U7624 ( .A1(n7103), .A2(n7102), .ZN(U2874) );
  AOI22_X1 U7625 ( .A1(n7104), .A2(n7114), .B1(n7113), .B2(DATAI_18_), .ZN(
        n7106) );
  AOI22_X1 U7626 ( .A1(n7117), .A2(DATAI_2_), .B1(n7116), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n7105) );
  NAND2_X1 U7627 ( .A1(n7106), .A2(n7105), .ZN(U2873) );
  AOI22_X1 U7628 ( .A1(n7107), .A2(n7114), .B1(n7113), .B2(DATAI_19_), .ZN(
        n7109) );
  AOI22_X1 U7629 ( .A1(n7117), .A2(DATAI_3_), .B1(n7116), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n7108) );
  NAND2_X1 U7630 ( .A1(n7109), .A2(n7108), .ZN(U2872) );
  AOI22_X1 U7631 ( .A1(n7110), .A2(n7114), .B1(n7113), .B2(DATAI_21_), .ZN(
        n7112) );
  AOI22_X1 U7632 ( .A1(n7117), .A2(DATAI_5_), .B1(n7116), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n7111) );
  NAND2_X1 U7633 ( .A1(n7112), .A2(n7111), .ZN(U2870) );
  AOI22_X1 U7634 ( .A1(n7115), .A2(n7114), .B1(n7113), .B2(DATAI_23_), .ZN(
        n7119) );
  AOI22_X1 U7635 ( .A1(n7117), .A2(DATAI_7_), .B1(n7116), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n7118) );
  NAND2_X1 U7636 ( .A1(n7119), .A2(n7118), .ZN(U2868) );
  AOI21_X1 U7637 ( .B1(n7120), .B2(n4403), .A(n7132), .ZN(n7126) );
  AND2_X1 U7638 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n7128), .ZN(n7201)
         );
  AOI21_X1 U7639 ( .B1(n7122), .B2(n7121), .A(n7201), .ZN(n7125) );
  INV_X1 U7640 ( .A(n7125), .ZN(n7123) );
  AOI22_X1 U7641 ( .A1(n7126), .A2(n7123), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n7128), .ZN(n7206) );
  AOI22_X1 U7642 ( .A1(n7139), .A2(n7201), .B1(n7148), .B2(n7202), .ZN(n7131)
         );
  NAND2_X1 U7643 ( .A1(n7126), .A2(n7125), .ZN(n7127) );
  OAI211_X1 U7644 ( .C1(n7146), .C2(n7128), .A(n7127), .B(n7143), .ZN(n7203)
         );
  INV_X1 U7645 ( .A(n7129), .ZN(n7200) );
  AOI22_X1 U7646 ( .A1(n7203), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n7138), 
        .B2(n7200), .ZN(n7130) );
  OAI211_X1 U7647 ( .C1(n7206), .C2(n7151), .A(n7131), .B(n7130), .ZN(U3108)
         );
  NOR2_X1 U7648 ( .A1(n7133), .A2(n7132), .ZN(n7142) );
  OR2_X1 U7649 ( .A1(n7135), .A2(n7134), .ZN(n7136) );
  NAND2_X1 U7650 ( .A1(n7136), .A2(n7137), .ZN(n7140) );
  AOI22_X1 U7651 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n7145), .B1(n7142), .B2(
        n7140), .ZN(n7217) );
  INV_X1 U7652 ( .A(n7137), .ZN(n7209) );
  AOI22_X1 U7653 ( .A1(n7139), .A2(n7209), .B1(n7138), .B2(n7207), .ZN(n7150)
         );
  INV_X1 U7654 ( .A(n7140), .ZN(n7141) );
  NAND2_X1 U7655 ( .A1(n7142), .A2(n7141), .ZN(n7144) );
  OAI211_X1 U7656 ( .C1(n7146), .C2(n7145), .A(n7144), .B(n7143), .ZN(n7213)
         );
  AOI22_X1 U7657 ( .A1(n7213), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n7148), 
        .B2(n7211), .ZN(n7149) );
  OAI211_X1 U7658 ( .C1(n7217), .C2(n7151), .A(n7150), .B(n7149), .ZN(U3076)
         );
  AOI22_X1 U7659 ( .A1(n7155), .A2(n7201), .B1(n7156), .B2(n7200), .ZN(n7153)
         );
  AOI22_X1 U7660 ( .A1(n7203), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n7154), 
        .B2(n7202), .ZN(n7152) );
  OAI211_X1 U7661 ( .C1(n7206), .C2(n7159), .A(n7153), .B(n7152), .ZN(U3109)
         );
  AOI22_X1 U7662 ( .A1(n7155), .A2(n7209), .B1(n7154), .B2(n7211), .ZN(n7158)
         );
  AOI22_X1 U7663 ( .A1(n7213), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n7156), 
        .B2(n7207), .ZN(n7157) );
  OAI211_X1 U7664 ( .C1(n7217), .C2(n7159), .A(n7158), .B(n7157), .ZN(U3077)
         );
  AOI22_X1 U7665 ( .A1(n7163), .A2(n7201), .B1(n7162), .B2(n7200), .ZN(n7161)
         );
  AOI22_X1 U7666 ( .A1(n7203), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n7164), 
        .B2(n7202), .ZN(n7160) );
  OAI211_X1 U7667 ( .C1(n7206), .C2(n7167), .A(n7161), .B(n7160), .ZN(U3110)
         );
  AOI22_X1 U7668 ( .A1(n7163), .A2(n7209), .B1(n7162), .B2(n7207), .ZN(n7166)
         );
  AOI22_X1 U7669 ( .A1(n7213), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n7164), 
        .B2(n7211), .ZN(n7165) );
  OAI211_X1 U7670 ( .C1(n7217), .C2(n7167), .A(n7166), .B(n7165), .ZN(U3078)
         );
  AOI22_X1 U7671 ( .A1(n7171), .A2(n7201), .B1(n7172), .B2(n7200), .ZN(n7169)
         );
  AOI22_X1 U7672 ( .A1(n7203), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n7170), 
        .B2(n7202), .ZN(n7168) );
  OAI211_X1 U7673 ( .C1(n7206), .C2(n7175), .A(n7169), .B(n7168), .ZN(U3111)
         );
  AOI22_X1 U7674 ( .A1(n7171), .A2(n7209), .B1(n7170), .B2(n7211), .ZN(n7174)
         );
  AOI22_X1 U7675 ( .A1(n7213), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n7172), 
        .B2(n7207), .ZN(n7173) );
  OAI211_X1 U7676 ( .C1(n7217), .C2(n7175), .A(n7174), .B(n7173), .ZN(U3079)
         );
  AOI22_X1 U7677 ( .A1(n7179), .A2(n7201), .B1(n7180), .B2(n7202), .ZN(n7177)
         );
  AOI22_X1 U7678 ( .A1(n7203), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n7178), 
        .B2(n7200), .ZN(n7176) );
  OAI211_X1 U7679 ( .C1(n7206), .C2(n7183), .A(n7177), .B(n7176), .ZN(U3112)
         );
  AOI22_X1 U7680 ( .A1(n7179), .A2(n7209), .B1(n7178), .B2(n7207), .ZN(n7182)
         );
  AOI22_X1 U7681 ( .A1(n7213), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n7180), 
        .B2(n7211), .ZN(n7181) );
  OAI211_X1 U7682 ( .C1(n7217), .C2(n7183), .A(n7182), .B(n7181), .ZN(U3080)
         );
  AOI22_X1 U7683 ( .A1(n7187), .A2(n7201), .B1(n7188), .B2(n7200), .ZN(n7185)
         );
  AOI22_X1 U7684 ( .A1(n7203), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n7186), 
        .B2(n7202), .ZN(n7184) );
  OAI211_X1 U7685 ( .C1(n7206), .C2(n7191), .A(n7185), .B(n7184), .ZN(U3113)
         );
  AOI22_X1 U7686 ( .A1(n7187), .A2(n7209), .B1(n7186), .B2(n7211), .ZN(n7190)
         );
  AOI22_X1 U7687 ( .A1(n7213), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n7188), 
        .B2(n7207), .ZN(n7189) );
  OAI211_X1 U7688 ( .C1(n7217), .C2(n7191), .A(n7190), .B(n7189), .ZN(U3081)
         );
  AOI22_X1 U7689 ( .A1(n7195), .A2(n7201), .B1(n7194), .B2(n7202), .ZN(n7193)
         );
  AOI22_X1 U7690 ( .A1(n7203), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n7196), 
        .B2(n7200), .ZN(n7192) );
  OAI211_X1 U7691 ( .C1(n7206), .C2(n7199), .A(n7193), .B(n7192), .ZN(U3114)
         );
  AOI22_X1 U7692 ( .A1(n7195), .A2(n7209), .B1(n7194), .B2(n7211), .ZN(n7198)
         );
  AOI22_X1 U7693 ( .A1(n7213), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n7196), 
        .B2(n7207), .ZN(n7197) );
  OAI211_X1 U7694 ( .C1(n7217), .C2(n7199), .A(n7198), .B(n7197), .ZN(U3082)
         );
  AOI22_X1 U7695 ( .A1(n7210), .A2(n7201), .B1(n7208), .B2(n7200), .ZN(n7205)
         );
  AOI22_X1 U7696 ( .A1(n7203), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n7212), 
        .B2(n7202), .ZN(n7204) );
  OAI211_X1 U7697 ( .C1(n7206), .C2(n7216), .A(n7205), .B(n7204), .ZN(U3115)
         );
  AOI22_X1 U7698 ( .A1(n7210), .A2(n7209), .B1(n7208), .B2(n7207), .ZN(n7215)
         );
  AOI22_X1 U7699 ( .A1(n7213), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n7212), 
        .B2(n7211), .ZN(n7214) );
  OAI211_X1 U7700 ( .C1(n7217), .C2(n7216), .A(n7215), .B(n7214), .ZN(U3083)
         );
  BUF_X1 U3506 ( .A(n3799), .Z(n5185) );
  XNOR2_X1 U3495 ( .A(n4428), .B(n5598), .ZN(n6687) );
  CLKBUF_X1 U34700 ( .A(n3757), .Z(n4605) );
  NOR2_X1 U3479 ( .A1(n5189), .A2(n5418), .ZN(n3437) );
  CLKBUF_X1 U3485 ( .A(n4488), .Z(n6708) );
  CLKBUF_X1 U3487 ( .A(n5988), .Z(n5989) );
  CLKBUF_X1 U3499 ( .A(n4792), .Z(n4853) );
  CLKBUF_X1 U3749 ( .A(n4867), .Z(n4908) );
  CLKBUF_X1 U3793 ( .A(n3773), .Z(n5762) );
  AOI21_X1 U3798 ( .B1(n6040), .B2(n6713), .A(n6039), .ZN(n6041) );
  CLKBUF_X1 U4094 ( .A(n4837), .Z(n5417) );
  OR2_X1 U4108 ( .A1(n5087), .A2(n4386), .ZN(n7218) );
endmodule

