

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4403, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385;

  CLKBUF_X2 U4909 ( .A(n6613), .Z(n7735) );
  AND2_X1 U4910 ( .A1(n8091), .A2(n6598), .ZN(n8066) );
  NAND2_X1 U4911 ( .A1(n6946), .A2(n6944), .ZN(n6936) );
  CLKBUF_X2 U4912 ( .A(n8631), .Z(n6261) );
  BUF_X2 U4913 ( .A(n5835), .Z(n8757) );
  CLKBUF_X2 U4915 ( .A(n5836), .Z(n8756) );
  BUF_X2 U4916 ( .A(n5845), .Z(n8782) );
  CLKBUF_X2 U4917 ( .A(n5106), .Z(n7873) );
  NAND2_X1 U4918 ( .A1(n7922), .A2(n7923), .ZN(n5638) );
  XNOR2_X1 U4919 ( .A(n5734), .B(n10332), .ZN(n7602) );
  NAND2_X1 U4920 ( .A1(n5737), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5734) );
  OR2_X1 U4921 ( .A1(n5225), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5259) );
  AND2_X1 U4922 ( .A1(n7668), .A2(n7657), .ZN(n5277) );
  INV_X1 U4923 ( .A(n8066), .ZN(n8070) );
  INV_X1 U4924 ( .A(n7873), .ZN(n5398) );
  INV_X2 U4925 ( .A(n6234), .ZN(n8629) );
  BUF_X1 U4926 ( .A(n5048), .Z(n4497) );
  NAND2_X1 U4927 ( .A1(n5947), .A2(n5946), .ZN(n7306) );
  OR2_X1 U4928 ( .A1(n5716), .A2(n9562), .ZN(n5715) );
  NAND2_X1 U4929 ( .A1(n5718), .A2(n5719), .ZN(n9721) );
  NAND2_X1 U4931 ( .A1(n7698), .A2(n7697), .ZN(n7783) );
  INV_X1 U4932 ( .A(n8755), .ZN(n6212) );
  XNOR2_X2 U4933 ( .A(n7708), .B(n7706), .ZN(n7838) );
  NAND4_X2 U4934 ( .A1(n5099), .A2(n5098), .A3(n5097), .A4(n5096), .ZN(n8110)
         );
  INV_X2 U4935 ( .A(n9014), .ZN(n9131) );
  NAND2_X2 U4936 ( .A1(n5395), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5396) );
  INV_X2 U4937 ( .A(n6778), .ZN(n7926) );
  OAI211_X2 U4938 ( .C1(n5845), .C2(n6374), .A(n4968), .B(n4967), .ZN(n7047)
         );
  XNOR2_X1 U4939 ( .A(n5728), .B(n5727), .ZN(n9008) );
  AOI21_X1 U4942 ( .B1(n8661), .B2(n8732), .A(n8731), .ZN(n8733) );
  MUX2_X1 U4943 ( .A(n9515), .B(n9514), .S(n9927), .Z(n9516) );
  MUX2_X1 U4944 ( .A(n9436), .B(n9514), .S(n9932), .Z(n9437) );
  NAND2_X1 U4945 ( .A1(n7704), .A2(n7756), .ZN(n7758) );
  NAND2_X1 U4946 ( .A1(n7673), .A2(n7672), .ZN(n7857) );
  NAND2_X1 U4947 ( .A1(n4773), .A2(n4777), .ZN(n4772) );
  NAND2_X1 U4948 ( .A1(n6051), .A2(n6050), .ZN(n9555) );
  NAND2_X1 U4949 ( .A1(n8838), .A2(n8951), .ZN(n8797) );
  INV_X2 U4950 ( .A(n9648), .ZN(n9645) );
  NAND2_X1 U4951 ( .A1(n5917), .A2(n5916), .ZN(n7181) );
  INV_X2 U4952 ( .A(n9715), .ZN(n9887) );
  NAND2_X1 U4953 ( .A1(n8834), .A2(n8836), .ZN(n8796) );
  CLKBUF_X1 U4954 ( .A(n6603), .Z(n6779) );
  INV_X1 U4955 ( .A(n7705), .ZN(n6613) );
  BUF_X1 U4956 ( .A(n5052), .Z(n6693) );
  INV_X1 U4957 ( .A(n6878), .ZN(n9898) );
  NAND3_X1 U4958 ( .A1(n5042), .A2(n4809), .A3(n4807), .ZN(n5052) );
  CLKBUF_X2 U4959 ( .A(n5026), .Z(n5548) );
  NAND2_X1 U4960 ( .A1(n4810), .A2(n6377), .ZN(n4809) );
  INV_X8 U4961 ( .A(n6218), .ZN(n6194) );
  INV_X2 U4962 ( .A(n5490), .ZN(n7071) );
  INV_X2 U4963 ( .A(n5100), .ZN(n7872) );
  INV_X2 U4965 ( .A(n5826), .ZN(n8781) );
  AND2_X2 U4966 ( .A1(n6390), .A2(n6321), .ZN(P1_U3973) );
  NAND4_X1 U4967 ( .A1(n5799), .A2(n5798), .A3(n5797), .A4(n5796), .ZN(n5813)
         );
  NOR2_X1 U4968 ( .A1(n9008), .A2(n6708), .ZN(n5754) );
  NAND2_X1 U4969 ( .A1(n8577), .A2(n5023), .ZN(n7657) );
  NAND2_X1 U4970 ( .A1(n4495), .A2(n4494), .ZN(n5023) );
  NAND2_X1 U4971 ( .A1(n5024), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5025) );
  OR2_X1 U4972 ( .A1(n5591), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n5620) );
  NAND2_X2 U4973 ( .A1(n5731), .A2(n5758), .ZN(n9007) );
  INV_X2 U4974 ( .A(n8579), .ZN(n8588) );
  AND2_X1 U4975 ( .A1(n5610), .A2(n4464), .ZN(n5022) );
  INV_X2 U4976 ( .A(n8586), .ZN(n4406) );
  OR2_X1 U4977 ( .A1(n5729), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U4978 ( .A1(n4836), .A2(n4835), .ZN(n6510) );
  OR2_X1 U4979 ( .A1(n5148), .A2(n5013), .ZN(n5356) );
  INV_X2 U4980 ( .A(n5087), .ZN(n7868) );
  OR2_X1 U4981 ( .A1(n5735), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5737) );
  NOR2_X1 U4982 ( .A1(n5013), .A2(n5016), .ZN(n4826) );
  INV_X1 U4983 ( .A(n5148), .ZN(n4407) );
  NAND2_X1 U4984 ( .A1(n4696), .A2(n4695), .ZN(n5086) );
  NAND2_X1 U4985 ( .A1(n5334), .A2(n4432), .ZN(n5013) );
  NAND2_X1 U4986 ( .A1(n5066), .A2(n5067), .ZN(n5079) );
  INV_X1 U4987 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n10267) );
  NOR2_X1 U4988 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5823) );
  INV_X1 U4989 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5775) );
  NOR2_X1 U4990 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5702) );
  NOR2_X1 U4991 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5703) );
  NOR2_X1 U4992 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5704) );
  NOR2_X2 U4993 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5066) );
  NOR2_X1 U4994 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5010) );
  INV_X1 U4995 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5763) );
  NOR2_X1 U4996 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5009) );
  NOR2_X1 U4997 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5008) );
  INV_X4 U4998 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4999 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5768) );
  INV_X1 U5000 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6806) );
  INV_X2 U5001 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5002 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5007) );
  AOI21_X1 U5003 ( .B1(n4774), .B2(n4435), .A(n4772), .ZN(n7817) );
  INV_X1 U5004 ( .A(n7857), .ZN(n4774) );
  INV_X1 U5005 ( .A(n7657), .ZN(n5027) );
  NOR2_X1 U5006 ( .A1(n6983), .A2(n4848), .ZN(n4847) );
  NAND2_X1 U5007 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  NAND2_X1 U5008 ( .A1(n5028), .A2(n5027), .ZN(n5093) );
  AND2_X1 U5009 ( .A1(n7657), .A2(n5028), .ZN(n5074) );
  AND2_X1 U5010 ( .A1(n7669), .A2(n5745), .ZN(n5834) );
  AOI21_X1 U5011 ( .B1(n4538), .B2(n4537), .A(n4536), .ZN(n4535) );
  INV_X1 U5012 ( .A(n9274), .ZN(n4536) );
  NAND2_X1 U5013 ( .A1(n4448), .A2(n4668), .ZN(n4666) );
  NAND2_X1 U5014 ( .A1(n4668), .A2(n8045), .ZN(n4667) );
  INV_X1 U5015 ( .A(n5351), .ZN(n4721) );
  OR2_X1 U5016 ( .A1(n8501), .A2(n8272), .ZN(n8071) );
  CLKBUF_X1 U5017 ( .A(n5093), .Z(n5580) );
  NAND2_X1 U5018 ( .A1(n4506), .A2(n4508), .ZN(n4504) );
  INV_X1 U5019 ( .A(n6354), .ZN(n4508) );
  NAND2_X1 U5020 ( .A1(n4511), .A2(n4510), .ZN(n7153) );
  AOI21_X1 U5021 ( .B1(n4512), .B2(n4841), .A(n4441), .ZN(n4510) );
  NAND2_X1 U5022 ( .A1(n7524), .A2(n7496), .ZN(n4516) );
  NAND2_X1 U5023 ( .A1(n9975), .A2(n8104), .ZN(n7973) );
  NAND2_X1 U5024 ( .A1(n5048), .A2(n5087), .ZN(n5080) );
  NOR2_X1 U5025 ( .A1(n8299), .A2(n7843), .ZN(n8051) );
  NAND2_X1 U5026 ( .A1(n8299), .A2(n7843), .ZN(n8050) );
  OR2_X1 U5027 ( .A1(n8532), .A2(n8343), .ZN(n8037) );
  AND2_X1 U5028 ( .A1(n7812), .A2(n8367), .ZN(n8026) );
  OR2_X1 U5029 ( .A1(n8548), .A2(n7686), .ZN(n8021) );
  OR2_X1 U5030 ( .A1(n8553), .A2(n7749), .ZN(n4998) );
  OR2_X1 U5031 ( .A1(n8485), .A2(n8403), .ZN(n8016) );
  OR2_X1 U5032 ( .A1(n8445), .A2(n8432), .ZN(n7995) );
  NAND2_X1 U5033 ( .A1(n7622), .A2(n5305), .ZN(n4959) );
  INV_X1 U5034 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5067) );
  CLKBUF_X1 U5035 ( .A(n5066), .Z(n4496) );
  NAND2_X1 U5036 ( .A1(n4987), .A2(n4995), .ZN(n4986) );
  NAND2_X1 U5037 ( .A1(n4995), .A2(n4993), .ZN(n4988) );
  NAND2_X1 U5038 ( .A1(n6029), .A2(n6028), .ZN(n4995) );
  INV_X1 U5039 ( .A(n5754), .ZN(n5781) );
  OR2_X1 U5040 ( .A1(n9430), .A2(n8776), .ZN(n8920) );
  OR2_X1 U5041 ( .A1(n9226), .A2(n9202), .ZN(n9162) );
  OR2_X1 U5042 ( .A1(n9236), .A2(n8774), .ZN(n8915) );
  NAND2_X1 U5043 ( .A1(n9236), .A2(n8774), .ZN(n9160) );
  NOR2_X1 U5044 ( .A1(n9450), .A2(n9281), .ZN(n4682) );
  INV_X1 U5045 ( .A(n9195), .ZN(n4902) );
  NOR2_X1 U5046 ( .A1(n9534), .A2(n9188), .ZN(n9190) );
  NAND2_X1 U5047 ( .A1(n9009), .A2(n9014), .ZN(n6706) );
  NAND2_X1 U5048 ( .A1(n9325), .A2(n9534), .ZN(n9308) );
  NAND2_X1 U5049 ( .A1(n6926), .A2(n6884), .ZN(n6927) );
  OAI21_X1 U5050 ( .B1(n5577), .B2(n5576), .A(n5575), .ZN(n7659) );
  INV_X1 U5051 ( .A(n5570), .ZN(n5577) );
  OAI21_X1 U5052 ( .B1(n5372), .B2(n5371), .A(n5370), .ZN(n5389) );
  INV_X1 U5053 ( .A(n5311), .ZN(n4725) );
  NAND2_X1 U5054 ( .A1(n5292), .A2(n5291), .ZN(n5309) );
  INV_X1 U5055 ( .A(n5287), .ZN(n5288) );
  NAND2_X1 U5056 ( .A1(n5250), .A2(n5241), .ZN(n5251) );
  INV_X1 U5057 ( .A(n4676), .ZN(n4675) );
  INV_X1 U5058 ( .A(n5195), .ZN(n4677) );
  XNOR2_X1 U5059 ( .A(n5233), .B(SI_10_), .ZN(n5232) );
  OAI21_X1 U5060 ( .B1(n5185), .B2(n4677), .A(n4675), .ZN(n5219) );
  NAND2_X1 U5061 ( .A1(n4645), .A2(n4644), .ZN(n5182) );
  AOI21_X1 U5062 ( .B1(n4647), .B2(n4649), .A(n4449), .ZN(n4644) );
  INV_X1 U5063 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4964) );
  NAND2_X2 U5064 ( .A1(n8087), .A2(n8253), .ZN(n5048) );
  NAND2_X1 U5065 ( .A1(n5279), .A2(n5278), .ZN(n5299) );
  INV_X1 U5066 ( .A(n9965), .ZN(n7209) );
  CLKBUF_X1 U5067 ( .A(n5276), .Z(n7074) );
  INV_X1 U5068 ( .A(n7070), .ZN(n5603) );
  OR2_X1 U5069 ( .A1(n5093), .A2(n6608), .ZN(n5030) );
  NAND2_X1 U5070 ( .A1(n4522), .A2(n4521), .ZN(n4520) );
  INV_X1 U5071 ( .A(n7241), .ZN(n4521) );
  NOR2_X1 U5072 ( .A1(n7497), .A2(n9653), .ZN(n8133) );
  NAND2_X1 U5073 ( .A1(n4852), .A2(n4851), .ZN(n4850) );
  INV_X1 U5074 ( .A(n8137), .ZN(n4851) );
  NOR2_X1 U5075 ( .A1(n8160), .A2(n8159), .ZN(n8168) );
  NAND2_X1 U5076 ( .A1(n4563), .A2(n4562), .ZN(n4703) );
  INV_X1 U5077 ( .A(n8172), .ZN(n4562) );
  OR2_X1 U5078 ( .A1(n8490), .A2(n8419), .ZN(n8009) );
  AOI21_X1 U5079 ( .B1(n4947), .B2(n4949), .A(n4471), .ZN(n4946) );
  NOR2_X1 U5080 ( .A1(n4798), .A2(n5646), .ZN(n4797) );
  NAND2_X1 U5081 ( .A1(n5048), .A2(n7868), .ZN(n5106) );
  NAND2_X1 U5082 ( .A1(n6607), .A2(n6601), .ZN(n7917) );
  OR2_X1 U5083 ( .A1(n8467), .A2(n8329), .ZN(n5512) );
  OR2_X1 U5084 ( .A1(n8474), .A2(n8356), .ZN(n5476) );
  OR2_X1 U5085 ( .A1(n8474), .A2(n7808), .ZN(n8032) );
  OR2_X1 U5086 ( .A1(n6605), .A2(n8070), .ZN(n9640) );
  INV_X1 U5087 ( .A(n4497), .ZN(n5397) );
  AND2_X1 U5088 ( .A1(n5679), .A2(n5597), .ZN(n9637) );
  AND3_X1 U5089 ( .A1(n4407), .A2(n4825), .A3(n4824), .ZN(n5614) );
  NOR2_X1 U5090 ( .A1(n5016), .A2(n4827), .ZN(n4825) );
  INV_X1 U5091 ( .A(n5013), .ZN(n4824) );
  NAND2_X1 U5092 ( .A1(n8611), .A2(n8614), .ZN(n8612) );
  AOI21_X1 U5093 ( .B1(n9311), .B2(n6194), .A(n6181), .ZN(n8713) );
  NAND2_X1 U5094 ( .A1(n8601), .A2(n8602), .ZN(n4605) );
  AND2_X1 U5095 ( .A1(n7669), .A2(n9568), .ZN(n5835) );
  INV_X1 U5096 ( .A(n5971), .ZN(n5836) );
  INV_X1 U5097 ( .A(n9508), .ZN(n9137) );
  OR2_X1 U5098 ( .A1(n9236), .A2(n9201), .ZN(n4888) );
  NAND2_X1 U5099 ( .A1(n4890), .A2(n4889), .ZN(n9169) );
  OR2_X1 U5100 ( .A1(n4455), .A2(n7606), .ZN(n4889) );
  NOR2_X1 U5101 ( .A1(n8808), .A2(n4895), .ZN(n4894) );
  NOR2_X1 U5102 ( .A1(n9862), .A2(n4409), .ZN(n4895) );
  XNOR2_X1 U5103 ( .A(n9034), .B(n6874), .ZN(n8791) );
  NAND2_X1 U5104 ( .A1(n6155), .A2(n6154), .ZN(n9326) );
  NAND2_X1 U5105 ( .A1(n6070), .A2(n6069), .ZN(n9494) );
  XNOR2_X1 U5106 ( .A(n5744), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U5107 ( .A1(n5464), .A2(n5463), .ZN(n5479) );
  NAND2_X1 U5108 ( .A1(n5415), .A2(n5414), .ZN(n5430) );
  XNOR2_X1 U5109 ( .A(n4518), .B(n4517), .ZN(n7438) );
  INV_X1 U5110 ( .A(n7490), .ZN(n4517) );
  NAND2_X1 U5111 ( .A1(n4550), .A2(n4548), .ZN(n4547) );
  NAND2_X1 U5112 ( .A1(n8847), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U5113 ( .A1(n4546), .A2(n4545), .ZN(n4544) );
  NAND2_X1 U5114 ( .A1(n8846), .A2(n4549), .ZN(n4545) );
  AOI21_X1 U5115 ( .B1(n4544), .B2(n8857), .A(n4543), .ZN(n4542) );
  INV_X1 U5116 ( .A(n8858), .ZN(n4543) );
  AND2_X1 U5117 ( .A1(n4654), .A2(n7990), .ZN(n4653) );
  OR2_X1 U5118 ( .A1(n7986), .A2(n4655), .ZN(n4654) );
  INV_X1 U5119 ( .A(n9635), .ZN(n4655) );
  OAI21_X1 U5120 ( .B1(n8004), .B2(n8005), .A(n8416), .ZN(n4642) );
  NAND2_X1 U5121 ( .A1(n4558), .A2(n4556), .ZN(n8887) );
  OAI21_X1 U5122 ( .B1(n4422), .B2(n8977), .A(n4557), .ZN(n4556) );
  AOI21_X1 U5123 ( .B1(n4560), .B2(n4559), .A(n9385), .ZN(n4558) );
  NOR2_X1 U5124 ( .A1(n8972), .A2(n4549), .ZN(n4557) );
  NAND2_X1 U5125 ( .A1(n8901), .A2(n8902), .ZN(n4540) );
  OR2_X1 U5126 ( .A1(n8020), .A2(n8066), .ZN(n4635) );
  NAND2_X1 U5127 ( .A1(n8012), .A2(n4414), .ZN(n4631) );
  NOR2_X1 U5128 ( .A1(n4634), .A2(n4633), .ZN(n4632) );
  INV_X1 U5129 ( .A(n8023), .ZN(n4634) );
  INV_X1 U5130 ( .A(n8053), .ZN(n4668) );
  INV_X1 U5131 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4484) );
  INV_X1 U5132 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4485) );
  NAND2_X1 U5133 ( .A1(n4529), .A2(n4528), .ZN(n4527) );
  AOI21_X1 U5134 ( .B1(n8917), .B2(n4531), .A(n4530), .ZN(n4529) );
  OAI21_X1 U5135 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n4528) );
  AND2_X1 U5136 ( .A1(n8915), .A2(n4431), .ZN(n4531) );
  NOR2_X1 U5137 ( .A1(n9526), .A2(n9193), .ZN(n9195) );
  INV_X1 U5138 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4627) );
  INV_X1 U5139 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4626) );
  NAND2_X1 U5140 ( .A1(n7758), .A2(n4480), .ZN(n7708) );
  NAND2_X1 U5141 ( .A1(n7703), .A2(n7842), .ZN(n4480) );
  NAND2_X1 U5142 ( .A1(n4663), .A2(n4659), .ZN(n8078) );
  NAND2_X1 U5143 ( .A1(n4662), .A2(n4660), .ZN(n4659) );
  NAND2_X1 U5144 ( .A1(n4661), .A2(n8064), .ZN(n4660) );
  NAND2_X1 U5145 ( .A1(n6354), .A2(n4585), .ZN(n4505) );
  OR2_X1 U5146 ( .A1(n6664), .A2(n4508), .ZN(n4507) );
  NAND2_X1 U5147 ( .A1(n4577), .A2(n6771), .ZN(n4580) );
  NAND2_X1 U5148 ( .A1(n6660), .A2(n4583), .ZN(n4582) );
  INV_X1 U5149 ( .A(n6340), .ZN(n4584) );
  INV_X1 U5150 ( .A(n4948), .ZN(n4947) );
  OAI21_X1 U5151 ( .B1(n5368), .B2(n4949), .A(n5383), .ZN(n4948) );
  NOR2_X1 U5152 ( .A1(n4935), .A2(n4930), .ZN(n4929) );
  INV_X1 U5153 ( .A(n5216), .ZN(n4930) );
  INV_X1 U5154 ( .A(n4936), .ZN(n4935) );
  AOI21_X1 U5155 ( .B1(n4936), .B2(n4934), .A(n4933), .ZN(n4932) );
  INV_X1 U5156 ( .A(n4939), .ZN(n4934) );
  INV_X1 U5157 ( .A(n7973), .ZN(n7387) );
  NAND2_X1 U5158 ( .A1(n5208), .A2(n10288), .ZN(n5225) );
  INV_X1 U5159 ( .A(n5209), .ZN(n5208) );
  NAND2_X1 U5160 ( .A1(n8303), .A2(n5531), .ZN(n4956) );
  AND2_X1 U5161 ( .A1(n8548), .A2(n7686), .ZN(n5654) );
  OR2_X1 U5162 ( .A1(n8569), .A2(n8418), .ZN(n8003) );
  OR2_X1 U5163 ( .A1(n9631), .A2(n8101), .ZN(n7884) );
  OR2_X1 U5164 ( .A1(n7627), .A2(n9641), .ZN(n7997) );
  OR2_X1 U5165 ( .A1(n5220), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U5166 ( .A1(n4451), .A2(n4411), .ZN(n4976) );
  NAND2_X1 U5167 ( .A1(n6839), .A2(n4411), .ZN(n4977) );
  OR2_X1 U5168 ( .A1(n9445), .A2(n9200), .ZN(n8916) );
  NAND2_X1 U5169 ( .A1(n9445), .A2(n9200), .ZN(n9159) );
  OR2_X1 U5170 ( .A1(n9450), .A2(n9197), .ZN(n9158) );
  NOR2_X1 U5171 ( .A1(n4906), .A2(n9195), .ZN(n4900) );
  NOR2_X1 U5172 ( .A1(n9178), .A2(n4918), .ZN(n4917) );
  INV_X1 U5173 ( .A(n4920), .ZN(n4918) );
  INV_X1 U5174 ( .A(n4866), .ZN(n4864) );
  NOR2_X1 U5175 ( .A1(n7545), .A2(n4867), .ZN(n4866) );
  NOR2_X1 U5176 ( .A1(n9865), .A2(n9683), .ZN(n7553) );
  NOR2_X1 U5177 ( .A1(n7306), .A2(n9873), .ZN(n4691) );
  AND2_X1 U5178 ( .A1(n4881), .A2(n4463), .ZN(n4880) );
  NAND2_X1 U5179 ( .A1(n5516), .A2(n5515), .ZN(n5533) );
  INV_X1 U5180 ( .A(n4752), .ZN(n4751) );
  NAND2_X1 U5181 ( .A1(n5479), .A2(n5478), .ZN(n5497) );
  AND2_X1 U5182 ( .A1(n5498), .A2(n5483), .ZN(n5496) );
  AOI21_X1 U5183 ( .B1(n4742), .B2(n4744), .A(n4474), .ZN(n4741) );
  OAI21_X1 U5184 ( .B1(n5389), .B2(n5388), .A(n5387), .ZN(n5410) );
  NAND2_X1 U5185 ( .A1(n4720), .A2(n4718), .ZN(n5372) );
  AOI21_X1 U5186 ( .B1(n4719), .B2(n4722), .A(n4476), .ZN(n4718) );
  NAND2_X1 U5187 ( .A1(n5309), .A2(n4433), .ZN(n4720) );
  XNOR2_X1 U5188 ( .A(n5290), .B(SI_13_), .ZN(n5287) );
  AOI21_X1 U5189 ( .B1(n4729), .B2(n4418), .A(n4443), .ZN(n4728) );
  NAND2_X1 U5190 ( .A1(n5234), .A2(SI_10_), .ZN(n5235) );
  NOR2_X1 U5191 ( .A1(n5236), .A2(n4734), .ZN(n4733) );
  INV_X1 U5192 ( .A(n5232), .ZN(n5236) );
  NAND2_X1 U5193 ( .A1(n5195), .A2(n5189), .ZN(n5196) );
  INV_X1 U5194 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5720) );
  INV_X1 U5195 ( .A(SI_3_), .ZN(n10113) );
  NAND2_X1 U5196 ( .A1(n6722), .A2(n6721), .ZN(n6726) );
  OR2_X1 U5197 ( .A1(n7765), .A2(n7766), .ZN(n4775) );
  NAND2_X1 U5198 ( .A1(n7513), .A2(n8102), .ZN(n4765) );
  NOR2_X1 U5199 ( .A1(n7513), .A2(n8102), .ZN(n4766) );
  XNOR2_X1 U5200 ( .A(n6798), .B(n7705), .ZN(n6617) );
  OR2_X1 U5201 ( .A1(n7857), .A2(n7858), .ZN(n4783) );
  NAND2_X1 U5202 ( .A1(n7909), .A2(n5005), .ZN(n7910) );
  OAI211_X1 U5203 ( .C1(n4835), .C2(P2_REG1_REG_2__SCAN_IN), .A(n4834), .B(
        n4833), .ZN(n6502) );
  NAND2_X1 U5204 ( .A1(n4837), .A2(n4832), .ZN(n4833) );
  AND2_X1 U5205 ( .A1(n5067), .A2(n9995), .ZN(n4832) );
  NAND2_X1 U5206 ( .A1(n4568), .A2(n4567), .ZN(n4566) );
  INV_X1 U5207 ( .A(n6559), .ZN(n4567) );
  INV_X1 U5208 ( .A(n6338), .ZN(n4568) );
  NAND2_X1 U5209 ( .A1(n6338), .A2(n6559), .ZN(n6657) );
  NAND3_X1 U5210 ( .A1(n4580), .A2(n4578), .A3(n4582), .ZN(n6761) );
  NOR2_X1 U5211 ( .A1(n4579), .A2(n6764), .ZN(n4578) );
  INV_X1 U5212 ( .A(n4429), .ZN(n4579) );
  NAND2_X1 U5213 ( .A1(n6660), .A2(n6340), .ZN(n4581) );
  NOR2_X1 U5214 ( .A1(n6983), .A2(n4576), .ZN(n4574) );
  NAND2_X1 U5215 ( .A1(n6983), .A2(n4848), .ZN(n4842) );
  NAND3_X1 U5216 ( .A1(n4572), .A2(n4570), .A3(n4571), .ZN(n7036) );
  AND2_X1 U5217 ( .A1(n4575), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4570) );
  NAND2_X1 U5218 ( .A1(n4573), .A2(n6983), .ZN(n7034) );
  NAND2_X1 U5219 ( .A1(n6982), .A2(n6981), .ZN(n4573) );
  OR2_X1 U5220 ( .A1(n7153), .A2(n7249), .ZN(n4831) );
  NAND2_X1 U5221 ( .A1(n4829), .A2(n4830), .ZN(n4522) );
  OR2_X1 U5222 ( .A1(n7537), .A2(n7536), .ZN(n7539) );
  OR2_X1 U5223 ( .A1(n8133), .A2(n8134), .ZN(n4852) );
  INV_X1 U5224 ( .A(n4516), .ZN(n8131) );
  AND2_X1 U5225 ( .A1(n4850), .A2(n4849), .ZN(n8184) );
  NAND2_X1 U5226 ( .A1(n8158), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4849) );
  AND2_X1 U5227 ( .A1(n4703), .A2(n4702), .ZN(n8213) );
  NAND2_X1 U5228 ( .A1(n8204), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4702) );
  NAND2_X1 U5229 ( .A1(n5506), .A2(n5505), .ZN(n5524) );
  INV_X1 U5230 ( .A(n5507), .ZN(n5506) );
  OR2_X1 U5231 ( .A1(n5468), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5486) );
  OR2_X1 U5232 ( .A1(n5434), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5449) );
  AND2_X1 U5233 ( .A1(n4806), .A2(n8392), .ZN(n4805) );
  NAND2_X1 U5234 ( .A1(n8406), .A2(n8009), .ZN(n4806) );
  AND4_X1 U5235 ( .A1(n5406), .A2(n5405), .A3(n5404), .A4(n5403), .ZN(n8403)
         );
  OR2_X1 U5236 ( .A1(n5362), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5377) );
  OAI21_X1 U5237 ( .B1(n7357), .B2(n7387), .A(n7974), .ZN(n7401) );
  AND4_X1 U5238 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n7564)
         );
  NOR2_X1 U5239 ( .A1(n7891), .A2(n4795), .ZN(n4794) );
  INV_X1 U5240 ( .A(n7959), .ZN(n4795) );
  AND4_X1 U5241 ( .A1(n5165), .A2(n5164), .A3(n5163), .A4(n5162), .ZN(n7204)
         );
  NOR2_X1 U5242 ( .A1(n7945), .A2(n4787), .ZN(n4786) );
  INV_X1 U5243 ( .A(n7946), .ZN(n4787) );
  NAND2_X1 U5244 ( .A1(n6776), .A2(n5072), .ZN(n6802) );
  NAND2_X1 U5245 ( .A1(n7917), .A2(n7923), .ZN(n4801) );
  XNOR2_X1 U5246 ( .A(n5071), .B(n8112), .ZN(n6778) );
  NAND2_X1 U5247 ( .A1(n4803), .A2(n5639), .ZN(n6683) );
  INV_X1 U5248 ( .A(n7917), .ZN(n5639) );
  INV_X1 U5249 ( .A(n7913), .ZN(n4803) );
  OR2_X1 U5250 ( .A1(n8272), .A2(n8271), .ZN(n8502) );
  NAND2_X1 U5251 ( .A1(n5544), .A2(n5543), .ZN(n8299) );
  AOI21_X1 U5252 ( .B1(n4815), .B2(n4818), .A(n8047), .ZN(n4814) );
  OR2_X1 U5253 ( .A1(n8338), .A2(n4816), .ZN(n4812) );
  NOR2_X1 U5254 ( .A1(n4408), .A2(n8048), .ZN(n4815) );
  AOI21_X1 U5255 ( .B1(n4956), .B2(n4427), .A(n8291), .ZN(n8293) );
  AOI21_X1 U5256 ( .B1(n4408), .B2(n8033), .A(n4819), .ZN(n4818) );
  NAND2_X1 U5257 ( .A1(n8046), .A2(n4817), .ZN(n8302) );
  INV_X1 U5258 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5259 ( .B1(n8033), .B2(n8032), .A(n8037), .ZN(n4823) );
  NOR2_X1 U5260 ( .A1(n8029), .A2(n7882), .ZN(n8328) );
  AOI21_X1 U5261 ( .B1(n8350), .B2(n8024), .A(n8026), .ZN(n8338) );
  INV_X1 U5262 ( .A(n4943), .ZN(n4942) );
  OAI21_X1 U5263 ( .B1(n8376), .B2(n4944), .A(n8363), .ZN(n4943) );
  OAI21_X1 U5264 ( .B1(n8373), .B2(n4799), .A(n8018), .ZN(n8362) );
  INV_X1 U5265 ( .A(n4998), .ZN(n4799) );
  NAND2_X1 U5266 ( .A1(n8415), .A2(n5368), .ZN(n8421) );
  AND4_X1 U5267 ( .A1(n5382), .A2(n5381), .A3(n5380), .A4(n5379), .ZN(n8419)
         );
  AND2_X1 U5268 ( .A1(n7899), .A2(n5306), .ZN(n4958) );
  AND2_X1 U5269 ( .A1(n4643), .A2(n5224), .ZN(n9975) );
  NAND2_X1 U5270 ( .A1(n6464), .A2(n7872), .ZN(n4643) );
  AND3_X1 U5271 ( .A1(n5154), .A2(n5153), .A3(n5152), .ZN(n9955) );
  NAND2_X1 U5272 ( .A1(n5038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U5273 ( .A1(n5595), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5596) );
  OR2_X1 U5274 ( .A1(n5222), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5254) );
  NOR2_X1 U5275 ( .A1(n5901), .A2(n5900), .ZN(n5918) );
  NAND2_X1 U5276 ( .A1(n4974), .A2(n4976), .ZN(n7220) );
  OR2_X1 U5277 ( .A1(n6837), .A2(n4977), .ZN(n4974) );
  CLKBUF_X1 U5278 ( .A(n8612), .Z(n8613) );
  AND2_X1 U5279 ( .A1(n8702), .A2(n6136), .ZN(n4985) );
  INV_X1 U5280 ( .A(n8703), .ZN(n4983) );
  AND2_X1 U5281 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5877) );
  INV_X1 U5282 ( .A(n5890), .ZN(n5891) );
  AND2_X1 U5283 ( .A1(n8653), .A2(n4983), .ZN(n4982) );
  INV_X1 U5284 ( .A(n4985), .ZN(n4980) );
  NAND2_X1 U5285 ( .A1(n4607), .A2(n4606), .ZN(n4488) );
  NAND2_X1 U5286 ( .A1(n9687), .A2(n9686), .ZN(n4607) );
  XNOR2_X1 U5287 ( .A(n5812), .B(n6234), .ZN(n5815) );
  AOI21_X1 U5288 ( .B1(n5813), .B2(n8626), .A(n5814), .ZN(n5816) );
  OR2_X1 U5289 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  INV_X1 U5290 ( .A(n4973), .ZN(n4972) );
  OAI21_X1 U5291 ( .B1(n8693), .B2(n6221), .A(n8663), .ZN(n4973) );
  NAND2_X1 U5292 ( .A1(n4972), .A2(n6221), .ZN(n4970) );
  OAI21_X1 U5293 ( .B1(n8690), .B2(n6221), .A(n4972), .ZN(n8661) );
  AOI21_X1 U5294 ( .B1(n8927), .B2(n9137), .A(n8938), .ZN(n8928) );
  NAND2_X1 U5295 ( .A1(n9204), .A2(n9512), .ZN(n9145) );
  AND2_X1 U5296 ( .A1(n9295), .A2(n4426), .ZN(n9235) );
  AOI21_X1 U5297 ( .B1(n4906), .B2(n4904), .A(n4450), .ZN(n4903) );
  INV_X1 U5298 ( .A(n4911), .ZN(n4904) );
  NOR2_X1 U5299 ( .A1(n9190), .A2(n4914), .ZN(n4911) );
  OR2_X1 U5300 ( .A1(n4910), .A2(n9190), .ZN(n4909) );
  NAND2_X1 U5301 ( .A1(n4913), .A2(n9187), .ZN(n4910) );
  AND2_X1 U5302 ( .A1(n8825), .A2(n9155), .ZN(n9291) );
  NAND2_X1 U5303 ( .A1(n9356), .A2(n9541), .ZN(n9339) );
  NOR2_X1 U5304 ( .A1(n4922), .A2(n4921), .ZN(n4920) );
  NOR2_X1 U5305 ( .A1(n9552), .A2(n9174), .ZN(n4921) );
  NOR2_X1 U5306 ( .A1(n9175), .A2(n4926), .ZN(n4922) );
  NAND2_X1 U5307 ( .A1(n4925), .A2(n4924), .ZN(n4923) );
  INV_X1 U5308 ( .A(n9175), .ZN(n4925) );
  INV_X1 U5309 ( .A(n9406), .ZN(n4924) );
  AND2_X1 U5310 ( .A1(n8886), .A2(n8888), .ZN(n9372) );
  NAND2_X1 U5311 ( .A1(n9494), .A2(n9172), .ZN(n4926) );
  OAI21_X1 U5312 ( .B1(n9555), .B2(n9171), .A(n9170), .ZN(n9405) );
  OR2_X1 U5313 ( .A1(n9168), .A2(n9167), .ZN(n5000) );
  OR2_X1 U5314 ( .A1(n9405), .A2(n9406), .ZN(n4927) );
  AND2_X1 U5315 ( .A1(n8879), .A2(n8880), .ZN(n9406) );
  AOI21_X1 U5316 ( .B1(n4894), .B2(n4409), .A(n4446), .ZN(n4893) );
  NAND2_X1 U5317 ( .A1(n7553), .A2(n8600), .ZN(n7613) );
  AND2_X1 U5318 ( .A1(n8967), .A2(n8966), .ZN(n8808) );
  NAND2_X1 U5319 ( .A1(n7460), .A2(n8963), .ZN(n7461) );
  NAND2_X1 U5320 ( .A1(n7465), .A2(n7464), .ZN(n9863) );
  OR2_X1 U5321 ( .A1(n9693), .A2(n9026), .ZN(n7464) );
  OR2_X1 U5322 ( .A1(n4689), .A2(n9670), .ZN(n4999) );
  NAND2_X1 U5323 ( .A1(n6859), .A2(n6823), .ZN(n6846) );
  INV_X1 U5324 ( .A(n6827), .ZN(n4555) );
  NAND2_X1 U5325 ( .A1(n4555), .A2(n6860), .ZN(n6859) );
  XNOR2_X1 U5326 ( .A(n5813), .B(n6957), .ZN(n6827) );
  OR2_X1 U5327 ( .A1(n9000), .A2(n4403), .ZN(n6906) );
  NAND2_X1 U5328 ( .A1(n8763), .A2(n8762), .ZN(n9430) );
  INV_X1 U5329 ( .A(n9861), .ZN(n9915) );
  INV_X2 U5330 ( .A(n8782), .ZN(n6121) );
  AND2_X1 U5331 ( .A1(n5865), .A2(n4684), .ZN(n6884) );
  NOR2_X1 U5332 ( .A1(n4437), .A2(n4685), .ZN(n4684) );
  NOR2_X1 U5333 ( .A1(n6391), .A2(n9740), .ZN(n4685) );
  NAND2_X1 U5334 ( .A1(n7663), .A2(n7662), .ZN(n7867) );
  XNOR2_X1 U5335 ( .A(n7867), .B(n7866), .ZN(n8752) );
  AND2_X1 U5336 ( .A1(n5726), .A2(n5762), .ZN(n4868) );
  XNOR2_X1 U5337 ( .A(n5533), .B(n5532), .ZN(n7639) );
  XNOR2_X1 U5338 ( .A(n5497), .B(n5496), .ZN(n7590) );
  AOI21_X1 U5339 ( .B1(n5415), .B2(n4745), .A(n4744), .ZN(n5441) );
  OAI21_X1 U5340 ( .B1(n5309), .B2(n4723), .A(n4722), .ZN(n5352) );
  NAND2_X1 U5341 ( .A1(n4726), .A2(n5311), .ZN(n5331) );
  NAND2_X1 U5342 ( .A1(n5309), .A2(n5308), .ZN(n4726) );
  OR2_X1 U5343 ( .A1(n6031), .A2(n6030), .ZN(n6048) );
  OAI21_X1 U5344 ( .B1(n5219), .B2(n4410), .A(n4729), .ZN(n5270) );
  XNOR2_X1 U5345 ( .A(n5145), .B(SI_5_), .ZN(n5143) );
  NAND2_X1 U5346 ( .A1(n5126), .A2(n5125), .ZN(n5144) );
  NAND2_X1 U5347 ( .A1(n5124), .A2(SI_4_), .ZN(n5125) );
  NOR2_X1 U5348 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5708) );
  NOR2_X1 U5349 ( .A1(n9619), .A2(n10371), .ZN(n9620) );
  NAND2_X1 U5350 ( .A1(n7837), .A2(n4759), .ZN(n7734) );
  AND4_X1 U5351 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n7586)
         );
  AND2_X1 U5352 ( .A1(n5493), .A2(n5492), .ZN(n8343) );
  NAND2_X1 U5353 ( .A1(n7917), .A2(n6602), .ZN(n6615) );
  OR2_X1 U5354 ( .A1(n6613), .A2(n6601), .ZN(n6602) );
  AND4_X1 U5355 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n6607)
         );
  AND2_X1 U5356 ( .A1(n5530), .A2(n5529), .ZN(n8316) );
  AOI21_X1 U5357 ( .B1(n6997), .B2(n6996), .A(n6995), .ZN(n7825) );
  NAND2_X1 U5358 ( .A1(n7825), .A2(n7824), .ZN(n7823) );
  AND2_X1 U5359 ( .A1(n6538), .A2(n6537), .ZN(n7856) );
  INV_X1 U5360 ( .A(n5037), .ZN(n5039) );
  INV_X1 U5361 ( .A(n8343), .ZN(n8096) );
  OR2_X1 U5362 ( .A1(n6553), .A2(n10128), .ZN(n6667) );
  INV_X1 U5363 ( .A(n4518), .ZN(n7489) );
  AND2_X1 U5364 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  OR2_X1 U5365 ( .A1(n8168), .A2(n8169), .ZN(n4563) );
  INV_X1 U5366 ( .A(n4500), .ZN(n8189) );
  INV_X1 U5367 ( .A(n4703), .ZN(n8203) );
  AOI21_X1 U5368 ( .B1(n8211), .B2(n8226), .A(n4708), .ZN(n4707) );
  OR2_X1 U5369 ( .A1(n8210), .A2(n4709), .ZN(n4708) );
  OAI21_X1 U5370 ( .B1(n8259), .B2(n8208), .A(n8207), .ZN(n4709) );
  XNOR2_X1 U5371 ( .A(n8213), .B(n8231), .ZN(n8205) );
  NOR2_X1 U5372 ( .A1(n4857), .A2(n8234), .ZN(n4856) );
  INV_X1 U5373 ( .A(n8239), .ZN(n4857) );
  AND2_X1 U5374 ( .A1(n8236), .A2(n8235), .ZN(n4854) );
  NAND2_X1 U5375 ( .A1(n4589), .A2(n4587), .ZN(n4586) );
  INV_X1 U5376 ( .A(n8216), .ZN(n4587) );
  NOR2_X1 U5377 ( .A1(n4590), .A2(n4595), .ZN(n4589) );
  INV_X1 U5378 ( .A(n4592), .ZN(n4590) );
  AOI21_X1 U5379 ( .B1(n4595), .B2(n8242), .A(n8270), .ZN(n4592) );
  OAI21_X1 U5380 ( .B1(n5609), .B2(n9637), .A(n5608), .ZN(n5675) );
  INV_X1 U5381 ( .A(n5607), .ZN(n5608) );
  OAI22_X1 U5382 ( .A1(n8077), .A2(n9640), .B1(n8271), .B2(n7879), .ZN(n5607)
         );
  OR2_X1 U5383 ( .A1(n8514), .A2(n8448), .ZN(n4483) );
  NAND2_X1 U5384 ( .A1(n5467), .A2(n5466), .ZN(n8474) );
  NAND2_X1 U5385 ( .A1(n5244), .A2(n5243), .ZN(n7409) );
  INV_X1 U5386 ( .A(n8277), .ZN(n8444) );
  AOI21_X1 U5387 ( .B1(n8761), .B2(n7872), .A(n5579), .ZN(n5698) );
  NAND2_X1 U5388 ( .A1(n7875), .A2(n7874), .ZN(n8501) );
  NOR2_X1 U5389 ( .A1(n5675), .A2(n5674), .ZN(n5701) );
  AND2_X1 U5390 ( .A1(n5673), .A2(n9968), .ZN(n5674) );
  NAND2_X1 U5391 ( .A1(n8284), .A2(n8283), .ZN(n8285) );
  CLKBUF_X1 U5392 ( .A(n5024), .Z(n8577) );
  OR2_X1 U5393 ( .A1(n6837), .A2(n6838), .ZN(n6961) );
  OR2_X1 U5394 ( .A1(n8714), .A2(n8713), .ZN(n6182) );
  NAND2_X1 U5395 ( .A1(n5892), .A2(n5891), .ZN(n9709) );
  NAND2_X1 U5396 ( .A1(n6138), .A2(n6137), .ZN(n9342) );
  OR2_X1 U5397 ( .A1(n6391), .A2(n6640), .ZN(n4967) );
  OR2_X1 U5398 ( .A1(n5826), .A2(n6380), .ZN(n4968) );
  NAND4_X1 U5399 ( .A1(n5822), .A2(n5821), .A3(n5820), .A4(n5819), .ZN(n9034)
         );
  NAND2_X1 U5400 ( .A1(n5835), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5820) );
  NAND4_X1 U5401 ( .A1(n5788), .A2(n5787), .A3(n5786), .A4(n5785), .ZN(n6822)
         );
  AOI21_X1 U5402 ( .B1(n4884), .B2(n9233), .A(n4452), .ZN(n4883) );
  AOI21_X1 U5403 ( .B1(n9021), .B2(n9003), .A(n4877), .ZN(n4876) );
  NAND2_X1 U5404 ( .A1(n4879), .A2(n9402), .ZN(n4878) );
  NOR2_X1 U5405 ( .A1(n9166), .A2(n9165), .ZN(n4877) );
  AND2_X1 U5406 ( .A1(n9216), .A2(n9215), .ZN(n9433) );
  AND2_X1 U5407 ( .A1(n9220), .A2(n9219), .ZN(n9435) );
  NAND2_X1 U5408 ( .A1(n4886), .A2(n4884), .ZN(n9220) );
  NAND2_X1 U5409 ( .A1(n4886), .A2(n4888), .ZN(n9218) );
  AND2_X1 U5410 ( .A1(n8784), .A2(n8783), .ZN(n9508) );
  NAND2_X1 U5411 ( .A1(n4552), .A2(n4551), .ZN(n8864) );
  AND2_X1 U5412 ( .A1(n8860), .A2(n8958), .ZN(n4551) );
  AOI21_X1 U5413 ( .B1(n4653), .B2(n4655), .A(n4652), .ZN(n4651) );
  NAND2_X1 U5414 ( .A1(n8871), .A2(n8879), .ZN(n4560) );
  OAI21_X1 U5415 ( .B1(n4642), .B2(n8007), .A(n4641), .ZN(n4640) );
  AND2_X1 U5416 ( .A1(n8009), .A2(n5004), .ZN(n4641) );
  INV_X1 U5417 ( .A(n4642), .ZN(n4638) );
  INV_X1 U5418 ( .A(n8887), .ZN(n8885) );
  NAND2_X1 U5419 ( .A1(n4639), .A2(n4636), .ZN(n8015) );
  NAND2_X1 U5420 ( .A1(n4638), .A2(n4637), .ZN(n4636) );
  NAND2_X1 U5421 ( .A1(n4640), .A2(n8070), .ZN(n4639) );
  NOR2_X1 U5422 ( .A1(n8005), .A2(n8070), .ZN(n4637) );
  NOR2_X1 U5423 ( .A1(n8791), .A2(n4555), .ZN(n8795) );
  NAND2_X1 U5424 ( .A1(n4534), .A2(n4532), .ZN(n8914) );
  AOI21_X1 U5425 ( .B1(n4535), .B2(n4539), .A(n4533), .ZN(n4532) );
  INV_X1 U5426 ( .A(n8906), .ZN(n4533) );
  NAND2_X1 U5427 ( .A1(n4630), .A2(n8028), .ZN(n8036) );
  NAND2_X1 U5428 ( .A1(n8918), .A2(n9162), .ZN(n4530) );
  NAND2_X1 U5429 ( .A1(n4667), .A2(n4666), .ZN(n4661) );
  NOR2_X1 U5430 ( .A1(n8063), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5431 ( .A1(n4666), .A2(n8314), .ZN(n4665) );
  AND2_X1 U5432 ( .A1(n5017), .A2(n5018), .ZN(n4963) );
  INV_X1 U5433 ( .A(n4990), .ZN(n4987) );
  NAND2_X1 U5434 ( .A1(n9335), .A2(n4862), .ZN(n9154) );
  NOR2_X1 U5435 ( .A1(n4749), .A2(n4753), .ZN(n4748) );
  INV_X1 U5436 ( .A(n5478), .ZN(n4749) );
  OAI21_X1 U5437 ( .B1(n5496), .B2(n4753), .A(n5513), .ZN(n4752) );
  INV_X1 U5438 ( .A(n4743), .ZN(n4742) );
  OAI21_X1 U5439 ( .B1(n4745), .B2(n4744), .A(n4475), .ZN(n4743) );
  INV_X1 U5440 ( .A(n5349), .ZN(n5350) );
  NOR2_X1 U5441 ( .A1(n4724), .A2(n5351), .ZN(n4719) );
  INV_X1 U5442 ( .A(n4648), .ZN(n4647) );
  OAI21_X1 U5443 ( .B1(n5143), .B2(n4649), .A(n5167), .ZN(n4648) );
  INV_X1 U5444 ( .A(n5147), .ZN(n4649) );
  NAND2_X1 U5445 ( .A1(n7774), .A2(n4771), .ZN(n4780) );
  AND2_X1 U5446 ( .A1(n5698), .A2(n8282), .ZN(n7876) );
  INV_X1 U5447 ( .A(n4657), .ZN(n4656) );
  OAI21_X1 U5448 ( .B1(n4667), .B2(n8314), .A(n4666), .ZN(n4657) );
  NAND2_X1 U5449 ( .A1(n4566), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4565) );
  INV_X1 U5450 ( .A(n6981), .ZN(n4576) );
  AND2_X1 U5451 ( .A1(n7440), .A2(n7439), .ZN(n7473) );
  NOR2_X1 U5452 ( .A1(n8196), .A2(n4498), .ZN(n8230) );
  NOR2_X1 U5453 ( .A1(n8193), .A2(n8496), .ZN(n4498) );
  INV_X1 U5454 ( .A(n5531), .ZN(n4952) );
  INV_X1 U5455 ( .A(n5369), .ZN(n4949) );
  OR2_X1 U5456 ( .A1(n5259), .A2(n5258), .ZN(n5280) );
  NOR2_X1 U5457 ( .A1(n5249), .A2(n4940), .ZN(n4939) );
  INV_X1 U5458 ( .A(n5231), .ZN(n4940) );
  NOR2_X1 U5459 ( .A1(n4442), .A2(n4937), .ZN(n4936) );
  NOR2_X1 U5460 ( .A1(n5249), .A2(n4938), .ZN(n4937) );
  NAND2_X1 U5461 ( .A1(n7385), .A2(n5231), .ZN(n4938) );
  OR2_X1 U5462 ( .A1(n5174), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U5463 ( .A1(n5159), .A2(n5158), .ZN(n5174) );
  INV_X1 U5464 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5158) );
  INV_X1 U5465 ( .A(n5160), .ZN(n5159) );
  AND2_X1 U5466 ( .A1(n5617), .A2(n6410), .ZN(n5677) );
  AND2_X1 U5467 ( .A1(n8299), .A2(n8304), .ZN(n5556) );
  NAND2_X1 U5468 ( .A1(n4818), .A2(n4817), .ZN(n4816) );
  INV_X1 U5469 ( .A(n5654), .ZN(n8022) );
  INV_X1 U5470 ( .A(n4963), .ZN(n4827) );
  INV_X1 U5471 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4486) );
  NOR2_X1 U5472 ( .A1(n5190), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5335) );
  OR2_X1 U5473 ( .A1(n4496), .A2(n5021), .ZN(n4837) );
  NOR2_X1 U5474 ( .A1(n4615), .A2(n4613), .ZN(n4612) );
  INV_X1 U5475 ( .A(n9711), .ZN(n4613) );
  INV_X1 U5476 ( .A(n4976), .ZN(n4615) );
  NAND2_X1 U5477 ( .A1(n5892), .A2(n4614), .ZN(n4610) );
  AND2_X1 U5478 ( .A1(n4976), .A2(n5891), .ZN(n4614) );
  AOI21_X1 U5479 ( .B1(n4976), .B2(n4977), .A(n4434), .ZN(n4975) );
  AND2_X1 U5480 ( .A1(n6139), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n6156) );
  NOR2_X1 U5481 ( .A1(n6124), .A2(n10178), .ZN(n6139) );
  NOR2_X1 U5482 ( .A1(n6026), .A2(n4994), .ZN(n4993) );
  INV_X1 U5483 ( .A(n9673), .ZN(n4994) );
  INV_X1 U5484 ( .A(n9659), .ZN(n4608) );
  NAND2_X1 U5485 ( .A1(n5982), .A2(n5981), .ZN(n4609) );
  NAND2_X1 U5486 ( .A1(n4524), .A2(n8922), .ZN(n8926) );
  NAND2_X1 U5487 ( .A1(n4525), .A2(n9203), .ZN(n4524) );
  NAND2_X1 U5488 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  INV_X1 U5489 ( .A(n9022), .ZN(n9200) );
  AND2_X1 U5490 ( .A1(n9254), .A2(n4682), .ZN(n4681) );
  NOR2_X1 U5491 ( .A1(n6054), .A2(n6053), .ZN(n6071) );
  NAND2_X1 U5492 ( .A1(n8600), .A2(n7604), .ZN(n4896) );
  INV_X1 U5493 ( .A(n7606), .ZN(n4891) );
  INV_X1 U5494 ( .A(n6829), .ZN(n4871) );
  OAI21_X1 U5495 ( .B1(n7108), .B2(n9031), .A(n7102), .ZN(n7083) );
  AND2_X1 U5496 ( .A1(n5762), .A2(n5740), .ZN(n4561) );
  XNOR2_X1 U5497 ( .A(n7659), .B(n7660), .ZN(n7658) );
  NAND2_X1 U5498 ( .A1(n4713), .A2(n4711), .ZN(n5570) );
  AOI21_X1 U5499 ( .B1(n4715), .B2(n4717), .A(n4712), .ZN(n4711) );
  INV_X1 U5500 ( .A(n5557), .ZN(n4712) );
  NOR2_X1 U5501 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n4881) );
  INV_X1 U5502 ( .A(n4716), .ZN(n4715) );
  OAI21_X1 U5503 ( .B1(n5532), .B2(n4717), .A(n5539), .ZN(n4716) );
  INV_X1 U5504 ( .A(n5534), .ZN(n4717) );
  INV_X1 U5505 ( .A(n5498), .ZN(n4753) );
  AND2_X1 U5506 ( .A1(n4746), .A2(n5414), .ZN(n4745) );
  NAND2_X1 U5507 ( .A1(n5429), .A2(n10266), .ZN(n4746) );
  NOR2_X1 U5508 ( .A1(n5429), .A2(n10266), .ZN(n4744) );
  NAND2_X1 U5509 ( .A1(n5413), .A2(n5412), .ZN(n5415) );
  INV_X1 U5510 ( .A(n5411), .ZN(n5412) );
  INV_X1 U5511 ( .A(n5410), .ZN(n5413) );
  AOI21_X1 U5512 ( .B1(n5307), .B2(n4724), .A(n4473), .ZN(n4722) );
  INV_X1 U5513 ( .A(n5235), .ZN(n4731) );
  INV_X1 U5514 ( .A(n4730), .ZN(n4729) );
  OAI21_X1 U5515 ( .B1(n4733), .B2(n4410), .A(n5250), .ZN(n4730) );
  OR2_X1 U5516 ( .A1(n5944), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5968) );
  AND2_X1 U5517 ( .A1(n5218), .A2(n5201), .ZN(n5202) );
  NOR2_X1 U5518 ( .A1(n5196), .A2(n4679), .ZN(n4678) );
  INV_X1 U5519 ( .A(n5184), .ZN(n4679) );
  AND2_X1 U5520 ( .A1(n5721), .A2(n5720), .ZN(n4624) );
  XNOR2_X1 U5521 ( .A(n5183), .B(SI_7_), .ZN(n5180) );
  OAI211_X1 U5522 ( .C1(n4696), .C2(P2_DATAO_REG_1__SCAN_IN), .A(n4694), .B(
        n4692), .ZN(n5062) );
  INV_X1 U5523 ( .A(n7710), .ZN(n4761) );
  AND2_X1 U5524 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  NAND2_X1 U5525 ( .A1(n7795), .A2(n4479), .ZN(n7742) );
  AND2_X1 U5526 ( .A1(n7793), .A2(n7794), .ZN(n4479) );
  INV_X1 U5527 ( .A(n8104), .ZN(n7381) );
  INV_X1 U5528 ( .A(n7814), .ZN(n4777) );
  OR2_X1 U5529 ( .A1(n7775), .A2(n7858), .ZN(n4781) );
  INV_X1 U5530 ( .A(n7813), .ZN(n4778) );
  NAND2_X1 U5531 ( .A1(n4776), .A2(n4779), .ZN(n7815) );
  INV_X1 U5532 ( .A(n4780), .ZN(n4779) );
  OR2_X1 U5533 ( .A1(n7857), .A2(n4781), .ZN(n4776) );
  OR2_X1 U5534 ( .A1(n6522), .A2(n6322), .ZN(n6530) );
  AND3_X1 U5535 ( .A1(n5438), .A2(n5437), .A3(n5436), .ZN(n7686) );
  AND3_X1 U5536 ( .A1(n5427), .A2(n5426), .A3(n5425), .ZN(n7749) );
  NAND2_X1 U5537 ( .A1(n6506), .A2(n6505), .ZN(n6504) );
  NAND2_X1 U5538 ( .A1(n4564), .A2(n6657), .ZN(n6661) );
  INV_X1 U5539 ( .A(n4565), .ZN(n4564) );
  AND2_X1 U5540 ( .A1(n4504), .A2(n4503), .ZN(n4502) );
  OR2_X1 U5541 ( .A1(n4505), .A2(n6664), .ZN(n4503) );
  NAND2_X1 U5542 ( .A1(n4582), .A2(n4478), .ZN(n6763) );
  OR2_X1 U5543 ( .A1(n6760), .A2(n10279), .ZN(n6758) );
  OAI21_X1 U5544 ( .B1(n6353), .B2(n4508), .A(n4506), .ZN(n6357) );
  NAND2_X1 U5545 ( .A1(n6983), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5546 ( .A1(n6973), .A2(n4847), .ZN(n4846) );
  NAND2_X1 U5547 ( .A1(n6973), .A2(n6972), .ZN(n4839) );
  OR2_X1 U5548 ( .A1(n4845), .A2(n4844), .ZN(n7030) );
  NAND2_X1 U5549 ( .A1(n4846), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4845) );
  INV_X1 U5550 ( .A(n7029), .ZN(n4844) );
  AOI21_X1 U5551 ( .B1(n4840), .B2(n4419), .A(n4513), .ZN(n4512) );
  NOR2_X1 U5552 ( .A1(n6983), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U5553 ( .A1(n7036), .A2(n7034), .ZN(n7032) );
  NAND2_X1 U5554 ( .A1(n7141), .A2(n7249), .ZN(n4701) );
  OR2_X1 U5555 ( .A1(n7235), .A2(n4699), .ZN(n7236) );
  INV_X1 U5556 ( .A(n4701), .ZN(n4699) );
  NAND2_X1 U5557 ( .A1(n7236), .A2(n7237), .ZN(n7440) );
  NAND2_X1 U5558 ( .A1(n4520), .A2(n4519), .ZN(n4518) );
  NAND2_X1 U5559 ( .A1(n7443), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4519) );
  NOR2_X1 U5560 ( .A1(n4604), .A2(n4603), .ZN(n4596) );
  XNOR2_X1 U5561 ( .A(n4516), .B(n4515), .ZN(n7497) );
  OR2_X1 U5562 ( .A1(n8186), .A2(n8187), .ZN(n4500) );
  AND2_X1 U5563 ( .A1(n4500), .A2(n4499), .ZN(n8196) );
  INV_X1 U5564 ( .A(n8188), .ZN(n4499) );
  OAI21_X1 U5565 ( .B1(n8303), .B2(n4955), .A(n4950), .ZN(n5586) );
  AND2_X1 U5566 ( .A1(n4953), .A2(n4951), .ZN(n4950) );
  AOI21_X1 U5567 ( .B1(n4954), .B2(n5556), .A(n4417), .ZN(n4953) );
  NAND2_X1 U5568 ( .A1(n4954), .A2(n4952), .ZN(n4951) );
  NAND2_X1 U5569 ( .A1(n8057), .A2(n7878), .ZN(n5656) );
  NAND2_X1 U5570 ( .A1(n5523), .A2(n10055), .ZN(n5545) );
  NAND2_X1 U5571 ( .A1(n5448), .A2(n10179), .ZN(n5468) );
  NAND2_X1 U5572 ( .A1(n5422), .A2(n5421), .ZN(n5434) );
  INV_X1 U5573 ( .A(n5423), .ZN(n5422) );
  NAND2_X1 U5574 ( .A1(n5376), .A2(n5375), .ZN(n5401) );
  NAND2_X1 U5575 ( .A1(n5340), .A2(n5339), .ZN(n5362) );
  INV_X1 U5576 ( .A(n5341), .ZN(n5340) );
  NAND2_X1 U5577 ( .A1(n5298), .A2(n10192), .ZN(n5320) );
  AND2_X1 U5578 ( .A1(n7979), .A2(n4792), .ZN(n4791) );
  NAND2_X1 U5579 ( .A1(n4793), .A2(n7977), .ZN(n4792) );
  OAI21_X1 U5580 ( .B1(n7360), .B2(n7385), .A(n5231), .ZN(n7403) );
  CLKBUF_X1 U5581 ( .A(n7359), .Z(n7360) );
  AND2_X1 U5582 ( .A1(n7892), .A2(n5173), .ZN(n4961) );
  AND4_X1 U5583 ( .A1(n5214), .A2(n5213), .A3(n5212), .A4(n5211), .ZN(n7361)
         );
  NAND2_X1 U5584 ( .A1(n4962), .A2(n5173), .ZN(n7128) );
  OR2_X1 U5585 ( .A1(n5137), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5160) );
  NAND2_X1 U5586 ( .A1(n5114), .A2(n5113), .ZN(n5137) );
  INV_X1 U5587 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5113) );
  INV_X1 U5588 ( .A(n5115), .ZN(n5114) );
  NAND2_X1 U5589 ( .A1(n6806), .A2(n5094), .ZN(n5115) );
  INV_X1 U5590 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U5591 ( .A1(n6687), .A2(n6601), .ZN(n6686) );
  CLKBUF_X1 U5592 ( .A(n5638), .Z(n7913) );
  XNOR2_X1 U5593 ( .A(n8511), .B(n8295), .ZN(n8279) );
  INV_X1 U5594 ( .A(n8279), .ZN(n8280) );
  NAND2_X1 U5595 ( .A1(n5555), .A2(n8050), .ZN(n8291) );
  NAND2_X1 U5596 ( .A1(n5504), .A2(n5503), .ZN(n8467) );
  AND2_X1 U5597 ( .A1(n8032), .A2(n8323), .ZN(n8339) );
  NAND2_X1 U5598 ( .A1(n8021), .A2(n8022), .ZN(n8363) );
  INV_X1 U5599 ( .A(n5409), .ZN(n8377) );
  NAND2_X1 U5600 ( .A1(n8377), .A2(n8376), .ZN(n8375) );
  AND2_X1 U5601 ( .A1(n5004), .A2(n8008), .ZN(n8416) );
  AND4_X1 U5602 ( .A1(n5325), .A2(n5324), .A3(n5323), .A4(n5322), .ZN(n8432)
         );
  AND2_X1 U5603 ( .A1(n8003), .A2(n8006), .ZN(n8430) );
  NAND2_X1 U5604 ( .A1(n4959), .A2(n5306), .ZN(n7643) );
  INV_X1 U5605 ( .A(n9640), .ZN(n8388) );
  INV_X1 U5606 ( .A(n9642), .ZN(n8386) );
  INV_X1 U5607 ( .A(n9637), .ZN(n8391) );
  AND3_X1 U5608 ( .A1(n5133), .A2(n5132), .A3(n5131), .ZN(n9949) );
  INV_X1 U5609 ( .A(n6530), .ZN(n6407) );
  NAND2_X1 U5610 ( .A1(n5610), .A2(n5017), .ZN(n5611) );
  CLKBUF_X1 U5611 ( .A(n5148), .Z(n5149) );
  OR2_X1 U5612 ( .A1(n5149), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n5190) );
  INV_X1 U5613 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U5614 ( .A1(n5108), .A2(n5007), .ZN(n4698) );
  NAND2_X1 U5615 ( .A1(n4837), .A2(n5067), .ZN(n4836) );
  NAND2_X1 U5616 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4838) );
  NAND2_X1 U5617 ( .A1(n6822), .A2(n5755), .ZN(n4965) );
  NAND2_X1 U5618 ( .A1(n5877), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5901) );
  OR2_X1 U5619 ( .A1(n5951), .A2(n5747), .ZN(n5972) );
  NOR2_X1 U5620 ( .A1(n9678), .A2(n4991), .ZN(n4990) );
  AND2_X1 U5621 ( .A1(n6025), .A2(n9672), .ZN(n4991) );
  NAND2_X1 U5622 ( .A1(n9690), .A2(n4993), .ZN(n4992) );
  NOR2_X1 U5623 ( .A1(n5972), .A2(n9590), .ZN(n5990) );
  AND2_X1 U5624 ( .A1(n5990), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6008) );
  NAND2_X1 U5625 ( .A1(n4609), .A2(n5983), .ZN(n9658) );
  INV_X1 U5626 ( .A(n9027), .ZN(n7413) );
  XNOR2_X1 U5627 ( .A(n4620), .B(n6234), .ZN(n5829) );
  NAND2_X1 U5628 ( .A1(n5827), .A2(n4621), .ZN(n4620) );
  NAND2_X1 U5629 ( .A1(n8625), .A2(n9034), .ZN(n4621) );
  AND2_X1 U5630 ( .A1(n8785), .A2(n5801), .ZN(n9140) );
  AND2_X1 U5631 ( .A1(n9508), .A2(n9142), .ZN(n8995) );
  AND2_X1 U5632 ( .A1(n9137), .A2(n8822), .ZN(n8938) );
  OAI21_X1 U5633 ( .B1(n8931), .B2(n4403), .A(n4737), .ZN(n4736) );
  NAND2_X1 U5634 ( .A1(n8932), .A2(n9006), .ZN(n4737) );
  NAND2_X1 U5635 ( .A1(n5835), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5785) );
  XNOR2_X1 U5636 ( .A(n9164), .B(n9163), .ZN(n4879) );
  AOI21_X1 U5637 ( .B1(n9229), .B2(n9233), .A(n9161), .ZN(n9213) );
  INV_X1 U5638 ( .A(n6262), .ZN(n6299) );
  INV_X1 U5639 ( .A(n4888), .ZN(n4885) );
  OAI21_X1 U5640 ( .B1(n9246), .B2(n9243), .A(n9159), .ZN(n9229) );
  NAND2_X1 U5641 ( .A1(n9295), .A2(n4681), .ZN(n9249) );
  NAND2_X1 U5642 ( .A1(n9261), .A2(n9158), .ZN(n9246) );
  NAND2_X1 U5643 ( .A1(n8916), .A2(n9159), .ZN(n9243) );
  AND2_X1 U5644 ( .A1(n6225), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U5645 ( .A1(n9295), .A2(n9526), .ZN(n9278) );
  NAND2_X1 U5646 ( .A1(n4901), .A2(n4898), .ZN(n9257) );
  AOI21_X1 U5647 ( .B1(n4900), .B2(n4903), .A(n4899), .ZN(n4898) );
  NOR2_X1 U5648 ( .A1(n9281), .A2(n9194), .ZN(n4899) );
  AND2_X1 U5649 ( .A1(n9156), .A2(n9155), .ZN(n9273) );
  OR2_X1 U5650 ( .A1(n8773), .A2(n8895), .ZN(n4859) );
  AND2_X1 U5651 ( .A1(n4858), .A2(n9153), .ZN(n4860) );
  NAND2_X1 U5652 ( .A1(n4862), .A2(n4861), .ZN(n4858) );
  NAND2_X1 U5653 ( .A1(n8773), .A2(n8939), .ZN(n9335) );
  AOI21_X1 U5654 ( .B1(n4917), .B2(n4923), .A(n4423), .ZN(n4916) );
  AND2_X1 U5655 ( .A1(n8892), .A2(n8939), .ZN(n9355) );
  NOR2_X1 U5656 ( .A1(n9555), .A2(n7613), .ZN(n9407) );
  NAND2_X1 U5657 ( .A1(n9407), .A2(n9412), .ZN(n9408) );
  OAI211_X1 U5658 ( .C1(n9857), .C2(n4865), .A(n7608), .B(n4863), .ZN(n8769)
         );
  NAND2_X1 U5659 ( .A1(n6008), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U5660 ( .A1(n7333), .A2(n4689), .ZN(n4688) );
  INV_X1 U5661 ( .A(n4872), .ZN(n7298) );
  OAI21_X1 U5662 ( .B1(n7293), .B2(n8790), .A(n7297), .ZN(n4872) );
  NAND2_X1 U5663 ( .A1(n7298), .A2(n7299), .ZN(n7460) );
  NAND2_X1 U5664 ( .A1(n7271), .A2(n9704), .ZN(n7307) );
  OR2_X1 U5665 ( .A1(n7111), .A2(n8798), .ZN(n7293) );
  NAND2_X1 U5666 ( .A1(n4870), .A2(n4869), .ZN(n8835) );
  AND2_X1 U5667 ( .A1(n8830), .A2(n8946), .ZN(n4869) );
  NAND2_X1 U5668 ( .A1(n4870), .A2(n8946), .ZN(n8829) );
  NAND2_X1 U5669 ( .A1(n8754), .A2(n8753), .ZN(n9148) );
  NAND2_X1 U5670 ( .A1(n8584), .A2(n8781), .ZN(n6260) );
  NAND2_X1 U5671 ( .A1(n6224), .A2(n6223), .ZN(n9450) );
  NAND2_X1 U5672 ( .A1(n7596), .A2(n8781), .ZN(n6224) );
  NAND2_X1 U5673 ( .A1(n6123), .A2(n6122), .ZN(n9357) );
  NAND2_X1 U5674 ( .A1(n6090), .A2(n6089), .ZN(n9392) );
  INV_X1 U5675 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5740) );
  XNOR2_X1 U5676 ( .A(n5570), .B(n5571), .ZN(n8621) );
  NAND2_X1 U5677 ( .A1(n5558), .A2(n5541), .ZN(n8584) );
  OAI21_X1 U5678 ( .B1(n5533), .B2(n4717), .A(n4715), .ZN(n5558) );
  OR2_X1 U5679 ( .A1(n5540), .A2(n5539), .ZN(n5541) );
  NAND2_X1 U5680 ( .A1(n4714), .A2(n5534), .ZN(n5540) );
  XNOR2_X1 U5681 ( .A(n5514), .B(n5513), .ZN(n7596) );
  INV_X1 U5682 ( .A(n4750), .ZN(n5514) );
  AOI21_X1 U5683 ( .B1(n5497), .B2(n5496), .A(n4753), .ZN(n4750) );
  OAI21_X1 U5684 ( .B1(n5458), .B2(n5457), .A(n5456), .ZN(n5464) );
  AND2_X1 U5685 ( .A1(n5478), .A2(n5462), .ZN(n5463) );
  NAND2_X1 U5686 ( .A1(n4732), .A2(n5235), .ZN(n5252) );
  NAND2_X1 U5687 ( .A1(n5219), .A2(n4733), .ZN(n4732) );
  AOI21_X1 U5688 ( .B1(n4675), .B2(n4677), .A(n4734), .ZN(n4673) );
  OR2_X1 U5689 ( .A1(n5931), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5944) );
  AND2_X1 U5690 ( .A1(n5762), .A2(n5720), .ZN(n5893) );
  NAND2_X1 U5691 ( .A1(n5105), .A2(n5104), .ZN(n5122) );
  XNOR2_X1 U5692 ( .A(n5123), .B(SI_4_), .ZN(n5121) );
  NOR2_X1 U5693 ( .A1(n9621), .A2(n10374), .ZN(n9622) );
  NAND2_X1 U5694 ( .A1(n6726), .A2(n6725), .ZN(n6749) );
  NAND2_X1 U5695 ( .A1(n5400), .A2(n5399), .ZN(n8485) );
  AND2_X1 U5696 ( .A1(n5554), .A2(n5553), .ZN(n7843) );
  NAND2_X1 U5697 ( .A1(n4760), .A2(n4412), .ZN(n4755) );
  NAND2_X1 U5698 ( .A1(n7736), .A2(n4467), .ZN(n4756) );
  INV_X1 U5699 ( .A(n4775), .ZN(n4782) );
  NOR2_X1 U5700 ( .A1(n7516), .A2(n4763), .ZN(n4762) );
  INV_X1 U5701 ( .A(n4765), .ZN(n4763) );
  NAND2_X1 U5702 ( .A1(n4764), .A2(n4765), .ZN(n7515) );
  NAND2_X1 U5703 ( .A1(n5275), .A2(n5274), .ZN(n9631) );
  AND2_X1 U5704 ( .A1(n5447), .A2(n5446), .ZN(n7812) );
  NAND2_X1 U5705 ( .A1(n6620), .A2(n6619), .ZN(n6722) );
  OR2_X1 U5706 ( .A1(n6606), .A2(n6605), .ZN(n7841) );
  AND4_X1 U5707 ( .A1(n5346), .A2(n5345), .A3(n5344), .A4(n5343), .ZN(n8418)
         );
  OAI21_X1 U5708 ( .B1(n4671), .B2(n8083), .A(n4440), .ZN(n4670) );
  AOI21_X1 U5709 ( .B1(n7911), .B2(n6598), .A(n4421), .ZN(n4669) );
  NOR2_X1 U5710 ( .A1(n8062), .A2(n8061), .ZN(n4671) );
  AND2_X1 U5711 ( .A1(n7077), .A2(n7076), .ZN(n8272) );
  AND2_X1 U5712 ( .A1(n7077), .A2(n5606), .ZN(n7879) );
  INV_X1 U5713 ( .A(n8316), .ZN(n8095) );
  INV_X1 U5714 ( .A(n7686), .ZN(n8378) );
  INV_X1 U5715 ( .A(n7749), .ZN(n8387) );
  INV_X1 U5716 ( .A(n7564), .ZN(n8103) );
  INV_X1 U5717 ( .A(n7204), .ZN(n8107) );
  INV_X1 U5718 ( .A(n6603), .ZN(n8113) );
  INV_X1 U5719 ( .A(P2_U3893), .ZN(n8225) );
  INV_X1 U5720 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5051) );
  NAND2_X1 U5721 ( .A1(n6657), .A2(n4566), .ZN(n6551) );
  NAND2_X1 U5722 ( .A1(n6353), .A2(n6664), .ZN(n6669) );
  NAND2_X1 U5723 ( .A1(n6355), .A2(n6356), .ZN(n6973) );
  NAND2_X1 U5724 ( .A1(n4697), .A2(n6341), .ZN(n6982) );
  NAND2_X1 U5725 ( .A1(n7029), .A2(n4846), .ZN(n6975) );
  NAND2_X1 U5726 ( .A1(n4509), .A2(n4512), .ZN(n7152) );
  OR2_X1 U5727 ( .A1(n6355), .A2(n4841), .ZN(n4509) );
  NAND2_X1 U5728 ( .A1(n4829), .A2(n4831), .ZN(n7154) );
  NOR2_X1 U5729 ( .A1(n4830), .A2(n7239), .ZN(n7238) );
  NOR2_X1 U5730 ( .A1(n7142), .A2(n7323), .ZN(n7235) );
  NAND2_X1 U5731 ( .A1(n4700), .A2(n4701), .ZN(n7142) );
  OR2_X1 U5732 ( .A1(n7141), .A2(n7249), .ZN(n4700) );
  INV_X1 U5733 ( .A(n4522), .ZN(n7242) );
  INV_X1 U5734 ( .A(n4520), .ZN(n7437) );
  OR2_X1 U5735 ( .A1(n7527), .A2(n7526), .ZN(n7524) );
  NOR2_X1 U5736 ( .A1(n8115), .A2(n8116), .ZN(n8120) );
  AND2_X1 U5737 ( .A1(n7539), .A2(n7477), .ZN(n8114) );
  INV_X1 U5738 ( .A(n4852), .ZN(n8138) );
  INV_X1 U5739 ( .A(n4850), .ZN(n8145) );
  XNOR2_X1 U5740 ( .A(n8184), .B(n8185), .ZN(n8146) );
  NOR2_X1 U5741 ( .A1(n8146), .A2(n8147), .ZN(n8186) );
  OR2_X1 U5742 ( .A1(n4595), .A2(n8242), .ZN(n4593) );
  NAND2_X1 U5743 ( .A1(n9648), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n4491) );
  INV_X1 U5744 ( .A(n8518), .ZN(n4492) );
  NAND2_X1 U5745 ( .A1(n4960), .A2(n5495), .ZN(n8313) );
  NAND2_X1 U5746 ( .A1(n8404), .A2(n8009), .ZN(n8393) );
  NAND2_X1 U5747 ( .A1(n8421), .A2(n5369), .ZN(n8401) );
  NAND2_X1 U5748 ( .A1(n5374), .A2(n5373), .ZN(n8490) );
  NAND2_X1 U5749 ( .A1(n5319), .A2(n5318), .ZN(n8445) );
  NAND2_X1 U5750 ( .A1(n4790), .A2(n7977), .ZN(n7567) );
  OR2_X1 U5751 ( .A1(n7401), .A2(n4793), .ZN(n4790) );
  CLKBUF_X1 U5752 ( .A(n7357), .Z(n7358) );
  NAND2_X1 U5753 ( .A1(n4796), .A2(n7959), .ZN(n7315) );
  AND2_X1 U5754 ( .A1(n5193), .A2(n5192), .ZN(n9965) );
  CLKBUF_X1 U5755 ( .A(n7056), .Z(n7057) );
  INV_X1 U5756 ( .A(n9944), .ZN(n6954) );
  CLKBUF_X1 U5757 ( .A(n6942), .Z(n6943) );
  NAND2_X1 U5758 ( .A1(n5092), .A2(n5091), .ZN(n6948) );
  NAND2_X1 U5759 ( .A1(n6683), .A2(n7923), .ZN(n6773) );
  INV_X1 U5760 ( .A(n8501), .ZN(n8451) );
  AOI21_X1 U5761 ( .B1(n8752), .B2(n7872), .A(n7864), .ZN(n8454) );
  NAND2_X1 U5762 ( .A1(n5522), .A2(n5521), .ZN(n8523) );
  NAND2_X1 U5763 ( .A1(n7639), .A2(n7872), .ZN(n5522) );
  NAND2_X1 U5764 ( .A1(n4813), .A2(n4818), .ZN(n8301) );
  NAND2_X1 U5765 ( .A1(n8338), .A2(n4408), .ZN(n4813) );
  NAND2_X1 U5766 ( .A1(n4821), .A2(n4822), .ZN(n8310) );
  OR2_X1 U5767 ( .A1(n8338), .A2(n8033), .ZN(n4821) );
  NAND2_X1 U5768 ( .A1(n5485), .A2(n5484), .ZN(n8532) );
  AND2_X1 U5769 ( .A1(n8338), .A2(n8032), .ZN(n8325) );
  INV_X1 U5770 ( .A(n7812), .ZN(n8542) );
  NAND2_X1 U5771 ( .A1(n5433), .A2(n5432), .ZN(n8548) );
  NAND2_X1 U5772 ( .A1(n5418), .A2(n5417), .ZN(n8553) );
  NAND2_X1 U5773 ( .A1(n5361), .A2(n5360), .ZN(n8562) );
  NAND2_X1 U5774 ( .A1(n5338), .A2(n5337), .ZN(n8569) );
  NAND2_X1 U5775 ( .A1(n5297), .A2(n5296), .ZN(n7627) );
  NAND2_X1 U5776 ( .A1(n5020), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4494) );
  OAI21_X1 U5777 ( .B1(n5022), .B2(n5021), .A(P2_IR_REG_29__SCAN_IN), .ZN(
        n4495) );
  XNOR2_X1 U5778 ( .A(n4785), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7591) );
  INV_X1 U5779 ( .A(n5610), .ZN(n4828) );
  XNOR2_X1 U5780 ( .A(n5242), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7490) );
  INV_X1 U5781 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10294) );
  INV_X1 U5782 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6385) );
  INV_X1 U5783 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6373) );
  INV_X1 U5784 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6379) );
  XNOR2_X1 U5785 ( .A(n5109), .B(n5108), .ZN(n6674) );
  XNOR2_X1 U5786 ( .A(n4523), .B(n5007), .ZN(n6559) );
  NAND2_X1 U5787 ( .A1(n5079), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4523) );
  AND2_X1 U5788 ( .A1(n6276), .A2(n6298), .ZN(n4619) );
  NAND2_X1 U5789 ( .A1(n6186), .A2(n6185), .ZN(n9296) );
  OAI211_X1 U5790 ( .C1(n6391), .C2(n6438), .A(n5847), .B(n5846), .ZN(n6878)
         );
  OR2_X1 U5791 ( .A1(n5826), .A2(n6398), .ZN(n5847) );
  NAND2_X1 U5792 ( .A1(n8613), .A2(n4985), .ZN(n4984) );
  AOI21_X1 U5793 ( .B1(n9690), .B2(n9673), .A(n9672), .ZN(n9671) );
  INV_X1 U5794 ( .A(n9450), .ZN(n9259) );
  NAND2_X1 U5795 ( .A1(n8691), .A2(n6222), .ZN(n8662) );
  CLKBUF_X1 U5796 ( .A(n8681), .Z(n8682) );
  NAND2_X1 U5797 ( .A1(n4992), .A2(n4989), .ZN(n9679) );
  INV_X1 U5798 ( .A(n4991), .ZN(n4989) );
  AOI21_X1 U5799 ( .B1(n4982), .B2(n4980), .A(n4472), .ZN(n4979) );
  INV_X1 U5800 ( .A(n4982), .ZN(n4981) );
  NAND2_X1 U5801 ( .A1(n6169), .A2(n6168), .ZN(n9311) );
  NOR2_X1 U5802 ( .A1(n9658), .A2(n9659), .ZN(n9688) );
  INV_X1 U5803 ( .A(n4488), .ZN(n9690) );
  NAND2_X1 U5804 ( .A1(n9708), .A2(n9711), .ZN(n4616) );
  OR2_X1 U5805 ( .A1(n6313), .A2(n6308), .ZN(n9656) );
  AND2_X1 U5806 ( .A1(n4970), .A2(n6254), .ZN(n4969) );
  NAND2_X1 U5807 ( .A1(n8690), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U5808 ( .A1(n7639), .A2(n8781), .ZN(n6237) );
  AOI21_X1 U5809 ( .B1(n4738), .B2(n4735), .A(n9007), .ZN(n9018) );
  INV_X1 U5810 ( .A(n4739), .ZN(n4738) );
  NAND2_X1 U5811 ( .A1(n4736), .A2(n9131), .ZN(n4735) );
  OAI21_X1 U5812 ( .B1(n8933), .B2(n9131), .A(n8935), .ZN(n4739) );
  NAND4_X1 U5813 ( .A1(n5861), .A2(n5860), .A3(n5859), .A4(n5858), .ZN(n9033)
         );
  NAND2_X1 U5814 ( .A1(n5835), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U5815 ( .A1(n5834), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5798) );
  XNOR2_X1 U5816 ( .A(n9145), .B(n9137), .ZN(n4686) );
  NAND2_X1 U5817 ( .A1(n4897), .A2(n4903), .ZN(n9271) );
  OR2_X1 U5818 ( .A1(n9318), .A2(n4905), .ZN(n4897) );
  NAND2_X1 U5819 ( .A1(n4907), .A2(n4413), .ZN(n9289) );
  NAND2_X1 U5820 ( .A1(n9318), .A2(n4911), .ZN(n4907) );
  NAND2_X1 U5821 ( .A1(n4908), .A2(n4913), .ZN(n9304) );
  OR2_X1 U5822 ( .A1(n9318), .A2(n9187), .ZN(n4908) );
  NAND2_X1 U5823 ( .A1(n4919), .A2(n4920), .ZN(n9373) );
  OR2_X1 U5824 ( .A1(n9405), .A2(n4923), .ZN(n4919) );
  AND2_X1 U5825 ( .A1(n4927), .A2(n4926), .ZN(n9384) );
  NAND2_X1 U5826 ( .A1(n4892), .A2(n4893), .ZN(n7603) );
  NAND2_X1 U5827 ( .A1(n9863), .A2(n4894), .ZN(n4892) );
  NAND2_X1 U5828 ( .A1(n9857), .A2(n8862), .ZN(n7546) );
  NAND2_X1 U5829 ( .A1(n5725), .A2(n5724), .ZN(n9683) );
  AOI21_X1 U5830 ( .B1(n9863), .B2(n9862), .A(n4409), .ZN(n7552) );
  NAND2_X1 U5831 ( .A1(n6007), .A2(n6006), .ZN(n9861) );
  OR2_X1 U5832 ( .A1(n9904), .A2(n6908), .ZN(n9897) );
  NAND2_X1 U5833 ( .A1(n6866), .A2(n6829), .ZN(n6847) );
  NAND2_X1 U5834 ( .A1(n7046), .A2(n9874), .ZN(n9901) );
  NAND2_X1 U5835 ( .A1(n6864), .A2(n4555), .ZN(n6865) );
  NAND2_X1 U5836 ( .A1(n6859), .A2(n4553), .ZN(n6900) );
  NAND2_X1 U5837 ( .A1(n4554), .A2(n6827), .ZN(n4553) );
  INV_X1 U5838 ( .A(n6860), .ZN(n4554) );
  INV_X1 U5839 ( .A(n9897), .ZN(n9872) );
  INV_X1 U5840 ( .A(n9491), .ZN(n9503) );
  INV_X1 U5841 ( .A(n9148), .ZN(n9512) );
  NOR2_X1 U5842 ( .A1(n4874), .A2(n9429), .ZN(n4873) );
  NAND2_X1 U5843 ( .A1(n9430), .A2(n9495), .ZN(n4875) );
  AOI21_X1 U5844 ( .B1(n9435), .B2(n9924), .A(n9434), .ZN(n9514) );
  AOI211_X1 U5845 ( .C1(n9440), .C2(n9924), .A(n9439), .B(n9438), .ZN(n9518)
         );
  INV_X1 U5846 ( .A(n9296), .ZN(n9530) );
  INV_X1 U5847 ( .A(n9311), .ZN(n9534) );
  INV_X1 U5848 ( .A(n9326), .ZN(n9537) );
  INV_X1 U5849 ( .A(n9357), .ZN(n9545) );
  NAND2_X1 U5850 ( .A1(n6034), .A2(n6033), .ZN(n7605) );
  INV_X1 U5851 ( .A(n6884), .ZN(n7119) );
  NAND2_X1 U5852 ( .A1(n9927), .A2(n9495), .ZN(n9551) );
  XNOR2_X1 U5853 ( .A(n7871), .B(n7870), .ZN(n9559) );
  OAI21_X1 U5854 ( .B1(n7867), .B2(n7866), .A(n7865), .ZN(n7871) );
  INV_X1 U5855 ( .A(n5745), .ZN(n9568) );
  INV_X1 U5856 ( .A(n5716), .ZN(n5719) );
  OAI21_X1 U5857 ( .B1(n5732), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5717) );
  INV_X1 U5858 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10300) );
  INV_X1 U5859 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10281) );
  INV_X1 U5860 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U5861 ( .A1(n4646), .A2(n5147), .ZN(n5168) );
  NAND2_X1 U5862 ( .A1(n5144), .A2(n5143), .ZN(n4646) );
  INV_X1 U5863 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6375) );
  NAND2_X1 U5864 ( .A1(n5823), .A2(n5708), .ZN(n5862) );
  NOR2_X1 U5865 ( .A1(n10373), .A2(n10372), .ZN(n10371) );
  NOR2_X1 U5866 ( .A1(n10376), .A2(n10375), .ZN(n10374) );
  NOR2_X1 U5867 ( .A1(n10370), .A2(n10369), .ZN(n10368) );
  NOR2_X1 U5868 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  AOI21_X1 U5869 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10045), .ZN(n10044) );
  NOR2_X1 U5870 ( .A1(n10044), .A2(n10043), .ZN(n10042) );
  NAND2_X1 U5871 ( .A1(n7823), .A2(n7000), .ZN(n7003) );
  AND2_X1 U5872 ( .A1(n7717), .A2(n4469), .ZN(n4481) );
  INV_X1 U5873 ( .A(n4563), .ZN(n8173) );
  OAI21_X1 U5874 ( .B1(n8206), .B2(n8270), .A(n4705), .ZN(P2_U3199) );
  INV_X1 U5875 ( .A(n4706), .ZN(n4705) );
  OAI21_X1 U5876 ( .B1(n8212), .B2(n8237), .A(n4707), .ZN(n4706) );
  OAI211_X1 U5877 ( .C1(n8240), .C2(n8270), .A(n4855), .B(n4853), .ZN(P2_U3200) );
  OAI21_X1 U5878 ( .B1(n8246), .B2(n4854), .A(n8267), .ZN(n4853) );
  NOR2_X1 U5879 ( .A1(n8238), .A2(n4856), .ZN(n4855) );
  OAI211_X1 U5880 ( .C1(n8243), .C2(n4591), .A(n8269), .B(n4588), .ZN(P2_U3201) );
  NAND2_X1 U5881 ( .A1(n4592), .A2(n4593), .ZN(n4591) );
  OR2_X1 U5882 ( .A1(n8217), .A2(n4586), .ZN(n4588) );
  OAI21_X1 U5883 ( .B1(n5668), .B2(n8448), .A(n5667), .ZN(n5669) );
  NAND2_X1 U5884 ( .A1(n8289), .A2(n4438), .ZN(P2_U3205) );
  NAND2_X1 U5885 ( .A1(n4493), .A2(n4489), .ZN(P2_U3206) );
  AOI21_X1 U5886 ( .B1(n4492), .B2(n7137), .A(n4490), .ZN(n4489) );
  NAND2_X1 U5887 ( .A1(n8515), .A2(n9645), .ZN(n4493) );
  NAND2_X1 U5888 ( .A1(n8300), .A2(n4491), .ZN(n4490) );
  INV_X1 U5889 ( .A(n5699), .ZN(n5700) );
  OAI22_X1 U5890 ( .A1(n5698), .A2(n8460), .B1(n10012), .B2(n5697), .ZN(n5699)
         );
  AND2_X1 U5891 ( .A1(n5686), .A2(n5001), .ZN(n5687) );
  AND2_X1 U5892 ( .A1(n4822), .A2(n4820), .ZN(n4408) );
  AND2_X1 U5893 ( .A1(n9915), .A2(n7466), .ZN(n4409) );
  OR2_X1 U5894 ( .A1(n5251), .A2(n4731), .ZN(n4410) );
  INV_X1 U5895 ( .A(n8063), .ZN(n4662) );
  NAND2_X1 U5896 ( .A1(n6963), .A2(n5930), .ZN(n4411) );
  INV_X1 U5897 ( .A(n8295), .ZN(n8077) );
  NAND2_X1 U5898 ( .A1(n5569), .A2(n5568), .ZN(n8295) );
  INV_X1 U5899 ( .A(n4841), .ZN(n4840) );
  OAI21_X1 U5900 ( .B1(n4847), .B2(n10002), .A(n4842), .ZN(n4841) );
  NOR2_X1 U5901 ( .A1(n7736), .A2(n4467), .ZN(n4412) );
  AND2_X1 U5902 ( .A1(n4909), .A2(n4912), .ZN(n4413) );
  AND3_X1 U5903 ( .A1(n8021), .A2(n4998), .A3(n8066), .ZN(n4414) );
  NAND2_X1 U5904 ( .A1(n6104), .A2(n6103), .ZN(n9377) );
  INV_X1 U5905 ( .A(n9377), .ZN(n9548) );
  AND2_X1 U5906 ( .A1(n8291), .A2(n4427), .ZN(n4415) );
  NAND2_X1 U5907 ( .A1(n4868), .A2(n4436), .ZN(n5732) );
  AND2_X1 U5908 ( .A1(n6277), .A2(n6298), .ZN(n4416) );
  AND2_X1 U5909 ( .A1(n8511), .A2(n8295), .ZN(n4417) );
  AND2_X1 U5910 ( .A1(n4410), .A2(n5268), .ZN(n4418) );
  AND2_X1 U5911 ( .A1(n4984), .A2(n4983), .ZN(n8651) );
  OR2_X1 U5912 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(n5079), .ZN(n5107) );
  OR2_X1 U5913 ( .A1(n4843), .A2(n4514), .ZN(n4419) );
  NAND2_X1 U5914 ( .A1(n8108), .A2(n7831), .ZN(n4420) );
  INV_X1 U5915 ( .A(n5307), .ZN(n5308) );
  OR2_X1 U5916 ( .A1(n7910), .A2(n8084), .ZN(n4421) );
  AND2_X1 U5917 ( .A1(n8878), .A2(n8971), .ZN(n4422) );
  AND2_X1 U5918 ( .A1(n7997), .A2(n7994), .ZN(n7991) );
  INV_X1 U5919 ( .A(n7991), .ZN(n4652) );
  AND2_X1 U5920 ( .A1(n9548), .A2(n9176), .ZN(n4423) );
  NAND2_X1 U5921 ( .A1(n4597), .A2(n4704), .ZN(n4424) );
  AND2_X1 U5922 ( .A1(n7905), .A2(n5495), .ZN(n4425) );
  AND2_X1 U5923 ( .A1(n4681), .A2(n4680), .ZN(n4426) );
  INV_X1 U5924 ( .A(n7842), .ZN(n8329) );
  NAND2_X1 U5925 ( .A1(n8742), .A2(n8744), .ZN(n8743) );
  INV_X1 U5926 ( .A(n9021), .ZN(n9202) );
  INV_X1 U5927 ( .A(n5093), .ZN(n5073) );
  INV_X1 U5929 ( .A(n8376), .ZN(n8374) );
  OR2_X1 U5930 ( .A1(n8523), .A2(n8095), .ZN(n4427) );
  NAND2_X1 U5931 ( .A1(n6862), .A2(n8631), .ZN(n4428) );
  XNOR2_X1 U5932 ( .A(n5269), .B(n5253), .ZN(n5268) );
  OR2_X1 U5933 ( .A1(n6340), .A2(n4585), .ZN(n4429) );
  INV_X1 U5934 ( .A(n9226), .ZN(n9517) );
  NAND2_X1 U5935 ( .A1(n8624), .A2(n8623), .ZN(n9226) );
  INV_X1 U5936 ( .A(n6972), .ZN(n4848) );
  OAI21_X1 U5937 ( .B1(n8612), .B2(n4981), .A(n4979), .ZN(n8712) );
  AND2_X1 U5938 ( .A1(n8612), .A2(n6136), .ZN(n8701) );
  AND2_X1 U5939 ( .A1(n4963), .A2(n5019), .ZN(n4430) );
  NOR2_X1 U5940 ( .A1(n8467), .A2(n7842), .ZN(n8043) );
  INV_X1 U5941 ( .A(n8043), .ZN(n4820) );
  NAND2_X1 U5942 ( .A1(n5989), .A2(n5988), .ZN(n9693) );
  INV_X1 U5943 ( .A(n9693), .ZN(n4689) );
  AND2_X1 U5944 ( .A1(n8916), .A2(n8934), .ZN(n4431) );
  AND2_X1 U5945 ( .A1(n8915), .A2(n9160), .ZN(n9233) );
  NAND2_X1 U5946 ( .A1(n5070), .A2(n5069), .ZN(n6614) );
  AND4_X1 U5947 ( .A1(n5012), .A2(n4486), .A3(n4485), .A4(n4484), .ZN(n4432)
         );
  NAND2_X1 U5948 ( .A1(n5257), .A2(n5256), .ZN(n9991) );
  INV_X1 U5949 ( .A(n9991), .ZN(n4933) );
  INV_X1 U5950 ( .A(n8042), .ZN(n4819) );
  NAND2_X1 U5951 ( .A1(n8690), .A2(n8693), .ZN(n8691) );
  NAND2_X1 U5952 ( .A1(n4984), .A2(n4982), .ZN(n8652) );
  AND2_X1 U5953 ( .A1(n4722), .A2(n4721), .ZN(n4433) );
  AND2_X1 U5954 ( .A1(n7218), .A2(n9698), .ZN(n4434) );
  INV_X1 U5955 ( .A(n8901), .ZN(n4537) );
  INV_X1 U5956 ( .A(n7923), .ZN(n4802) );
  NOR2_X1 U5957 ( .A1(n4781), .A2(n4778), .ZN(n4435) );
  AND2_X1 U5958 ( .A1(n5713), .A2(n4881), .ZN(n4436) );
  NOR2_X1 U5959 ( .A1(n8782), .A2(n6375), .ZN(n4437) );
  OR2_X1 U5960 ( .A1(n9861), .A2(n7466), .ZN(n8862) );
  INV_X1 U5961 ( .A(n8862), .ZN(n4867) );
  INV_X1 U5962 ( .A(n7899), .ZN(n7992) );
  AND2_X1 U5963 ( .A1(n4483), .A2(n8288), .ZN(n4438) );
  INV_X1 U5964 ( .A(n9281), .ZN(n9526) );
  NAND2_X1 U5965 ( .A1(n6205), .A2(n6204), .ZN(n9281) );
  NAND2_X1 U5966 ( .A1(n9295), .A2(n4682), .ZN(n4683) );
  AND2_X1 U5967 ( .A1(n8523), .A2(n8316), .ZN(n8048) );
  INV_X1 U5968 ( .A(n8048), .ZN(n4817) );
  AND2_X1 U5969 ( .A1(n8920), .A2(n8921), .ZN(n9203) );
  INV_X1 U5970 ( .A(n4539), .ZN(n4538) );
  NAND2_X1 U5971 ( .A1(n8904), .A2(n4540), .ZN(n4539) );
  AND2_X1 U5972 ( .A1(n5453), .A2(n8024), .ZN(n8354) );
  INV_X1 U5973 ( .A(n8354), .ZN(n4633) );
  OR2_X1 U5974 ( .A1(n8511), .A2(n8295), .ZN(n4439) );
  OR2_X1 U5975 ( .A1(n8082), .A2(n8081), .ZN(n4440) );
  INV_X1 U5976 ( .A(n4914), .ZN(n4913) );
  NOR2_X1 U5977 ( .A1(n9537), .A2(n9186), .ZN(n4914) );
  NOR2_X1 U5978 ( .A1(n7151), .A2(n10004), .ZN(n4441) );
  NAND2_X1 U5979 ( .A1(n4960), .A2(n4425), .ZN(n8311) );
  INV_X1 U5980 ( .A(n4906), .ZN(n4905) );
  AND2_X1 U5981 ( .A1(n4413), .A2(n4454), .ZN(n4906) );
  NOR2_X1 U5982 ( .A1(n9981), .A2(n7564), .ZN(n4442) );
  INV_X1 U5983 ( .A(n4955), .ZN(n4954) );
  OAI21_X1 U5984 ( .B1(n4415), .B2(n5556), .A(n4439), .ZN(n4955) );
  NAND2_X1 U5985 ( .A1(n5199), .A2(n5198), .ZN(n5218) );
  INV_X1 U5986 ( .A(n5218), .ZN(n4734) );
  AND2_X1 U5987 ( .A1(n5269), .A2(SI_12_), .ZN(n4443) );
  AND2_X1 U5988 ( .A1(n4658), .A2(n4656), .ZN(n4444) );
  INV_X1 U5989 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10332) );
  AND2_X1 U5990 ( .A1(n4859), .A2(n4860), .ZN(n4445) );
  NOR2_X1 U5991 ( .A1(n9683), .A2(n9024), .ZN(n4446) );
  NAND2_X1 U5992 ( .A1(n7640), .A2(n4769), .ZN(n4447) );
  INV_X1 U5993 ( .A(n7905), .ZN(n8314) );
  INV_X1 U5994 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9562) );
  OR2_X1 U5995 ( .A1(n8049), .A2(n8291), .ZN(n4448) );
  AND2_X1 U5996 ( .A1(n5170), .A2(SI_6_), .ZN(n4449) );
  NOR2_X1 U5997 ( .A1(n9192), .A2(n9530), .ZN(n4450) );
  NAND2_X1 U5998 ( .A1(n6960), .A2(n5929), .ZN(n4451) );
  AND2_X1 U5999 ( .A1(n9226), .A2(n9021), .ZN(n4452) );
  INV_X1 U6000 ( .A(n4760), .ZN(n4759) );
  NAND2_X1 U6001 ( .A1(n7709), .A2(n4761), .ZN(n4760) );
  AND2_X1 U6002 ( .A1(n4903), .A2(n4902), .ZN(n4453) );
  OR2_X1 U6003 ( .A1(n8523), .A2(n8316), .ZN(n8046) );
  OR2_X1 U6004 ( .A1(n9296), .A2(n9191), .ZN(n4454) );
  AND2_X1 U6005 ( .A1(n4893), .A2(n4896), .ZN(n4455) );
  AND2_X1 U6006 ( .A1(n4894), .A2(n4891), .ZN(n4456) );
  AND2_X1 U6007 ( .A1(n9290), .A2(n8788), .ZN(n4457) );
  NOR2_X1 U6008 ( .A1(n9217), .A2(n4885), .ZN(n4884) );
  NOR2_X1 U6009 ( .A1(n6830), .A2(n4871), .ZN(n4458) );
  AND2_X1 U6010 ( .A1(n9686), .A2(n4608), .ZN(n4459) );
  AND2_X1 U6011 ( .A1(n8982), .A2(n9319), .ZN(n4862) );
  AND2_X1 U6012 ( .A1(n4878), .A2(n4876), .ZN(n4460) );
  AND2_X1 U6013 ( .A1(n7001), .A2(n7000), .ZN(n4461) );
  AND2_X1 U6014 ( .A1(n4729), .A2(n5268), .ZN(n4462) );
  AND2_X1 U6015 ( .A1(n5714), .A2(n4978), .ZN(n4463) );
  AND2_X1 U6016 ( .A1(n4430), .A2(n10341), .ZN(n4464) );
  AND2_X1 U6017 ( .A1(n4547), .A2(n8857), .ZN(n4465) );
  INV_X1 U6018 ( .A(n8364), .ZN(n4944) );
  INV_X1 U6019 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n5021) );
  INV_X1 U6020 ( .A(n9445), .ZN(n9254) );
  NAND2_X1 U6021 ( .A1(n6237), .A2(n6236), .ZN(n9445) );
  NAND2_X1 U6022 ( .A1(n6260), .A2(n6259), .ZN(n9236) );
  INV_X1 U6023 ( .A(n9236), .ZN(n4680) );
  AND2_X1 U6024 ( .A1(n7547), .A2(n8867), .ZN(n4466) );
  INV_X1 U6025 ( .A(n8102), .ZN(n9639) );
  XNOR2_X1 U6026 ( .A(n7658), .B(n5578), .ZN(n8761) );
  INV_X1 U6027 ( .A(n8939), .ZN(n4861) );
  AND2_X1 U6028 ( .A1(n7733), .A2(n8304), .ZN(n4467) );
  AND2_X1 U6029 ( .A1(n6065), .A2(n6066), .ZN(n8742) );
  AND2_X1 U6030 ( .A1(n4783), .A2(n4782), .ZN(n4468) );
  AND2_X1 U6031 ( .A1(n6153), .A2(n6152), .ZN(n8703) );
  OR2_X1 U6032 ( .A1(n8517), .A2(n7848), .ZN(n4469) );
  OR2_X1 U6033 ( .A1(n8405), .A2(n8406), .ZN(n8404) );
  NAND2_X1 U6034 ( .A1(n8743), .A2(n6066), .ZN(n8670) );
  INV_X1 U6035 ( .A(n4724), .ZN(n4723) );
  NOR2_X1 U6036 ( .A1(n5330), .A2(n4725), .ZN(n4724) );
  AND2_X1 U6037 ( .A1(n4992), .A2(n4990), .ZN(n4470) );
  AND2_X1 U6038 ( .A1(n8490), .A2(n8389), .ZN(n4471) );
  NOR2_X1 U6039 ( .A1(n6167), .A2(n6166), .ZN(n4472) );
  INV_X1 U6040 ( .A(n7536), .ZN(n4604) );
  AND2_X1 U6041 ( .A1(n5329), .A2(n5328), .ZN(n4473) );
  AND2_X1 U6042 ( .A1(n5440), .A2(SI_21_), .ZN(n4474) );
  OR2_X1 U6043 ( .A1(n5440), .A2(SI_21_), .ZN(n4475) );
  AND2_X1 U6044 ( .A1(n5350), .A2(SI_16_), .ZN(n4476) );
  NOR2_X1 U6045 ( .A1(n7477), .A2(n8132), .ZN(n4477) );
  INV_X1 U6046 ( .A(n4704), .ZN(n4603) );
  AND2_X1 U6047 ( .A1(n5560), .A2(n5559), .ZN(n8060) );
  INV_X1 U6048 ( .A(n8060), .ZN(n8511) );
  NAND2_X1 U6049 ( .A1(n4839), .A2(n6983), .ZN(n7029) );
  NAND2_X1 U6050 ( .A1(n4770), .A2(n7640), .ZN(n5618) );
  NAND2_X1 U6051 ( .A1(n4616), .A2(n9709), .ZN(n6837) );
  NAND2_X1 U6052 ( .A1(n4788), .A2(n7946), .ZN(n6935) );
  INV_X1 U6053 ( .A(n8270), .ZN(n4594) );
  NAND2_X1 U6054 ( .A1(n5970), .A2(n5969), .ZN(n9664) );
  INV_X1 U6055 ( .A(n4687), .ZN(n7418) );
  NOR2_X1 U6056 ( .A1(n4690), .A2(n9664), .ZN(n4687) );
  AND2_X1 U6057 ( .A1(n8785), .A2(n6636), .ZN(n9003) );
  AND2_X1 U6058 ( .A1(n4580), .A2(n4429), .ZN(n4478) );
  AND2_X1 U6059 ( .A1(n7153), .A2(n7249), .ZN(n7239) );
  INV_X1 U6060 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4978) );
  INV_X1 U6061 ( .A(n6376), .ZN(n4811) );
  INV_X1 U6062 ( .A(n8085), .ZN(n8084) );
  INV_X1 U6063 ( .A(n4403), .ZN(n8943) );
  INV_X1 U6064 ( .A(n6356), .ZN(n4514) );
  INV_X1 U6065 ( .A(n7028), .ZN(n4513) );
  INV_X1 U6066 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4769) );
  INV_X1 U6067 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4629) );
  INV_X1 U6068 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U6069 ( .A1(n4581), .A2(n6771), .ZN(n6342) );
  NOR2_X1 U6070 ( .A1(n4584), .A2(n6771), .ZN(n4583) );
  AND2_X1 U6071 ( .A1(n4507), .A2(n6771), .ZN(n4506) );
  INV_X1 U6072 ( .A(n6771), .ZN(n4585) );
  INV_X1 U6073 ( .A(n8132), .ZN(n4515) );
  NOR2_X1 U6074 ( .A1(n7536), .A2(n8132), .ZN(n4602) );
  AND2_X1 U6075 ( .A1(n7477), .A2(n8132), .ZN(n4704) );
  NAND2_X1 U6076 ( .A1(n8919), .A2(n8934), .ZN(n4526) );
  NOR2_X1 U6077 ( .A1(n8977), .A2(n8934), .ZN(n4559) );
  NAND2_X1 U6078 ( .A1(n8850), .A2(n8934), .ZN(n4550) );
  NAND2_X1 U6079 ( .A1(n8849), .A2(n8934), .ZN(n4546) );
  INV_X1 U6080 ( .A(n8934), .ZN(n4549) );
  NAND2_X1 U6081 ( .A1(n6942), .A2(n7939), .ZN(n4788) );
  NAND2_X1 U6082 ( .A1(n7055), .A2(n4797), .ZN(n4796) );
  OAI22_X1 U6083 ( .A1(n7880), .A2(n7881), .B1(n8451), .B2(n8068), .ZN(n7911)
         );
  AOI21_X2 U6084 ( .B1(n8290), .B2(n8050), .A(n8051), .ZN(n8278) );
  OAI21_X1 U6085 ( .B1(n8362), .B2(n5654), .A(n8021), .ZN(n8350) );
  OAI22_X1 U6086 ( .A1(n8278), .A2(n5655), .B1(n8077), .B2(n8511), .ZN(n7877)
         );
  AND2_X2 U6087 ( .A1(n4407), .A2(n4826), .ZN(n5610) );
  NAND3_X2 U6088 ( .A1(n5058), .A2(n5057), .A3(n5056), .ZN(n8112) );
  AND4_X2 U6089 ( .A1(n5011), .A2(n5008), .A3(n5009), .A4(n5010), .ZN(n5334)
         );
  NAND2_X1 U6090 ( .A1(n7060), .A2(n7957), .ZN(n4962) );
  NAND2_X1 U6091 ( .A1(n4931), .A2(n4936), .ZN(n7562) );
  NAND2_X1 U6092 ( .A1(n7645), .A2(n5326), .ZN(n8429) );
  NAND2_X1 U6093 ( .A1(n5454), .A2(n4633), .ZN(n8351) );
  NAND2_X1 U6094 ( .A1(n5638), .A2(n6686), .ZN(n6685) );
  NAND3_X1 U6095 ( .A1(n4784), .A2(n7783), .A3(n7808), .ZN(n7718) );
  NAND2_X1 U6096 ( .A1(n7742), .A2(n7685), .ZN(n7690) );
  NAND2_X1 U6097 ( .A1(n4482), .A2(n4481), .ZN(P2_U3154) );
  NAND2_X1 U6098 ( .A1(n7712), .A2(n7734), .ZN(n4482) );
  NAND2_X1 U6099 ( .A1(n5610), .A2(n4430), .ZN(n5038) );
  NAND2_X2 U6100 ( .A1(n8435), .A2(n5348), .ZN(n8415) );
  OR2_X1 U6101 ( .A1(n8462), .A2(n8461), .ZN(P2_U3486) );
  OR2_X1 U6102 ( .A1(n8520), .A2(n8519), .ZN(P2_U3454) );
  NAND2_X1 U6103 ( .A1(n4962), .A2(n4961), .ZN(n7130) );
  NAND2_X1 U6104 ( .A1(n8351), .A2(n5455), .ZN(n8340) );
  NAND2_X1 U6105 ( .A1(n4487), .A2(n5267), .ZN(n9636) );
  NAND2_X1 U6106 ( .A1(n7317), .A2(n5215), .ZN(n5217) );
  NAND2_X1 U6107 ( .A1(n7359), .A2(n4939), .ZN(n4931) );
  NAND2_X1 U6108 ( .A1(n5266), .A2(n4933), .ZN(n4487) );
  NAND2_X2 U6109 ( .A1(n8311), .A2(n5512), .ZN(n8303) );
  OR3_X1 U6110 ( .A1(n8293), .A2(n8292), .A3(n9637), .ZN(n8297) );
  NAND2_X1 U6111 ( .A1(n4941), .A2(n4942), .ZN(n8352) );
  NAND2_X1 U6112 ( .A1(n6184), .A2(n6183), .ZN(n8601) );
  NAND2_X1 U6113 ( .A1(n4622), .A2(n8672), .ZN(n8671) );
  OAI21_X2 U6114 ( .B1(n4488), .B2(n4988), .A(n4986), .ZN(n6044) );
  NAND2_X4 U6115 ( .A1(n9721), .A2(n5801), .ZN(n6391) );
  OAI22_X1 U6116 ( .A1(n9257), .A2(n9198), .B1(n9197), .B2(n9259), .ZN(n9244)
         );
  NAND2_X1 U6117 ( .A1(n9431), .A2(n4875), .ZN(n4874) );
  NAND2_X1 U6118 ( .A1(n4460), .A2(n4873), .ZN(n9513) );
  NAND2_X1 U6119 ( .A1(n5092), .A2(n4957), .ZN(n6946) );
  AND2_X4 U6120 ( .A1(n6600), .A2(n6599), .ZN(n7705) );
  AOI21_X2 U6121 ( .B1(n7349), .B2(n7348), .A(n7347), .ZN(n7380) );
  OR2_X2 U6122 ( .A1(n7514), .A2(n4766), .ZN(n4764) );
  NAND2_X2 U6123 ( .A1(n7838), .A2(n8316), .ZN(n7837) );
  XNOR2_X1 U6124 ( .A(n7705), .B(n5071), .ZN(n6723) );
  NAND2_X1 U6125 ( .A1(n7696), .A2(n7695), .ZN(n4784) );
  AOI21_X1 U6126 ( .B1(n7392), .B2(n4996), .A(n7391), .ZN(n7514) );
  NAND2_X1 U6127 ( .A1(n7726), .A2(n7725), .ZN(n7795) );
  NAND2_X1 U6128 ( .A1(n5652), .A2(n8008), .ZN(n8405) );
  INV_X1 U6129 ( .A(n5080), .ZN(n4808) );
  INV_X1 U6130 ( .A(n5106), .ZN(n4810) );
  AOI21_X1 U6131 ( .B1(n4670), .B2(n8084), .A(n4669), .ZN(n8086) );
  NAND2_X1 U6132 ( .A1(n6353), .A2(n4506), .ZN(n4501) );
  OAI211_X1 U6133 ( .C1(n6353), .C2(n4505), .A(n4502), .B(n4501), .ZN(n6760)
         );
  NAND2_X1 U6134 ( .A1(n6355), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U6135 ( .A1(n8903), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U6136 ( .A1(n8851), .A2(n4465), .ZN(n4541) );
  AOI21_X1 U6137 ( .B1(n8851), .B2(n4547), .A(n4544), .ZN(n8859) );
  NAND2_X1 U6138 ( .A1(n4541), .A2(n4542), .ZN(n4552) );
  AND4_X1 U6139 ( .A1(n4880), .A2(n5713), .A3(n5762), .A4(n5726), .ZN(n5716)
         );
  NAND4_X1 U6140 ( .A1(n4880), .A2(n4561), .A3(n5713), .A4(n5726), .ZN(n5743)
         );
  NOR2_X2 U6141 ( .A1(n5743), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U6142 ( .A1(n4565), .A2(n6657), .ZN(n6339) );
  INV_X1 U6143 ( .A(n6982), .ZN(n4569) );
  NAND2_X1 U6144 ( .A1(n6982), .A2(n4574), .ZN(n4571) );
  NAND2_X1 U6145 ( .A1(n4569), .A2(n6983), .ZN(n4572) );
  NAND3_X1 U6146 ( .A1(n4572), .A2(n4575), .A3(n4571), .ZN(n6984) );
  INV_X1 U6147 ( .A(n6660), .ZN(n4577) );
  NOR2_X1 U6148 ( .A1(n8217), .A2(n8216), .ZN(n8243) );
  INV_X1 U6149 ( .A(n8255), .ZN(n4595) );
  NOR2_X1 U6150 ( .A1(n7474), .A2(n7475), .ZN(n7537) );
  NAND2_X1 U6151 ( .A1(n4597), .A2(n4596), .ZN(n4600) );
  NAND2_X1 U6152 ( .A1(n7475), .A2(n4604), .ZN(n4597) );
  OAI211_X1 U6153 ( .C1(n7474), .C2(n4424), .A(n4601), .B(n4598), .ZN(n7478)
         );
  AOI21_X1 U6154 ( .B1(n7475), .B2(n4602), .A(n4477), .ZN(n4599) );
  NAND2_X1 U6155 ( .A1(n7474), .A2(n4602), .ZN(n4601) );
  NAND2_X2 U6156 ( .A1(n4605), .A2(n8603), .ZN(n8690) );
  NAND2_X1 U6157 ( .A1(n8722), .A2(n6119), .ZN(n8611) );
  NAND2_X1 U6158 ( .A1(n6118), .A2(n6117), .ZN(n8722) );
  NAND3_X1 U6159 ( .A1(n4609), .A2(n4459), .A3(n5983), .ZN(n4606) );
  NAND2_X1 U6160 ( .A1(n5979), .A2(n5980), .ZN(n5983) );
  NAND2_X1 U6161 ( .A1(n9708), .A2(n4612), .ZN(n4611) );
  NAND3_X1 U6162 ( .A1(n4611), .A2(n4610), .A3(n4975), .ZN(n5963) );
  NAND2_X1 U6163 ( .A1(n4618), .A2(n4617), .ZN(P1_U3214) );
  AOI21_X1 U6164 ( .B1(n8734), .B2(n4416), .A(n6319), .ZN(n4617) );
  NAND2_X1 U6165 ( .A1(n6273), .A2(n4619), .ZN(n4618) );
  NAND2_X1 U6166 ( .A1(n8734), .A2(n6277), .ZN(n8649) );
  INV_X2 U6167 ( .A(n6218), .ZN(n8625) );
  NAND2_X1 U6168 ( .A1(n8671), .A2(n6087), .ZN(n8680) );
  NAND2_X1 U6169 ( .A1(n4623), .A2(n6066), .ZN(n4622) );
  NAND2_X1 U6170 ( .A1(n6064), .A2(n6063), .ZN(n6066) );
  NAND2_X1 U6171 ( .A1(n6065), .A2(n8744), .ZN(n4623) );
  NAND2_X1 U6172 ( .A1(n5762), .A2(n4624), .ZN(n5931) );
  INV_X1 U6173 ( .A(n5931), .ZN(n4625) );
  NAND2_X1 U6174 ( .A1(n4625), .A2(n5726), .ZN(n5729) );
  NAND3_X1 U6175 ( .A1(n5726), .A2(n5762), .A3(n5713), .ZN(n5735) );
  NAND3_X1 U6176 ( .A1(n4626), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4695) );
  NAND3_X1 U6177 ( .A1(n4629), .A2(n4628), .A3(n4627), .ZN(n4696) );
  NAND3_X1 U6178 ( .A1(n4635), .A2(n4632), .A3(n4631), .ZN(n4630) );
  NAND2_X1 U6179 ( .A1(n5144), .A2(n4647), .ZN(n4645) );
  NAND2_X1 U6180 ( .A1(n7987), .A2(n4653), .ZN(n4650) );
  NAND2_X1 U6181 ( .A1(n4650), .A2(n4651), .ZN(n7993) );
  OR2_X1 U6182 ( .A1(n8041), .A2(n4667), .ZN(n4658) );
  NAND2_X1 U6183 ( .A1(n8041), .A2(n4664), .ZN(n4663) );
  NAND2_X1 U6184 ( .A1(n5185), .A2(n4675), .ZN(n4672) );
  NAND2_X1 U6185 ( .A1(n4672), .A2(n4673), .ZN(n5237) );
  NAND2_X1 U6186 ( .A1(n5185), .A2(n4678), .ZN(n4674) );
  NAND2_X1 U6187 ( .A1(n5185), .A2(n5184), .ZN(n5197) );
  NAND2_X1 U6188 ( .A1(n4674), .A2(n5195), .ZN(n5203) );
  OAI21_X1 U6189 ( .B1(n4678), .B2(n4677), .A(n5202), .ZN(n4676) );
  MUX2_X1 U6190 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n5087), .Z(n5103) );
  MUX2_X1 U6191 ( .A(n6375), .B(n6379), .S(n5087), .Z(n5123) );
  MUX2_X1 U6192 ( .A(n5127), .B(n6373), .S(n5087), .Z(n5145) );
  MUX2_X1 U6193 ( .A(n6383), .B(n6385), .S(n5087), .Z(n5169) );
  MUX2_X1 U6194 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n5087), .Z(n5183) );
  MUX2_X1 U6195 ( .A(n6406), .B(n10294), .S(n5087), .Z(n5187) );
  MUX2_X1 U6196 ( .A(n10281), .B(n6463), .S(n5087), .Z(n5199) );
  MUX2_X1 U6197 ( .A(n10259), .B(n5238), .S(n5087), .Z(n5239) );
  MUX2_X1 U6198 ( .A(n10300), .B(n6465), .S(n5087), .Z(n5233) );
  MUX2_X1 U6199 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n5087), .Z(n5269) );
  MUX2_X1 U6200 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n5087), .Z(n5290) );
  MUX2_X1 U6201 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n5087), .Z(n5310) );
  MUX2_X1 U6202 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n5087), .Z(n5327) );
  MUX2_X1 U6203 ( .A(n5332), .B(n10154), .S(n5087), .Z(n5349) );
  MUX2_X1 U6204 ( .A(n6897), .B(n6899), .S(n5087), .Z(n5353) );
  INV_X1 U6205 ( .A(n4683), .ZN(n9258) );
  NOR2_X2 U6206 ( .A1(n6927), .A2(n9715), .ZN(n7105) );
  NOR2_X2 U6207 ( .A1(n6850), .A2(n6878), .ZN(n6926) );
  NAND2_X1 U6208 ( .A1(n6874), .A2(n6861), .ZN(n6850) );
  NOR2_X2 U6209 ( .A1(n4686), .A2(n9410), .ZN(n9422) );
  NOR2_X2 U6210 ( .A1(n9223), .A2(n9430), .ZN(n9204) );
  NOR2_X2 U6211 ( .A1(n4690), .A2(n4688), .ZN(n9866) );
  NAND2_X1 U6212 ( .A1(n4691), .A2(n7271), .ZN(n4690) );
  NOR2_X2 U6213 ( .A1(n9339), .A2(n9326), .ZN(n9325) );
  NOR2_X2 U6214 ( .A1(n9374), .A2(n9357), .ZN(n9356) );
  INV_X1 U6215 ( .A(n4695), .ZN(n4693) );
  NAND2_X1 U6216 ( .A1(n4693), .A2(n6397), .ZN(n4692) );
  NAND3_X1 U6217 ( .A1(n4696), .A2(n4695), .A3(n6377), .ZN(n4694) );
  NAND2_X1 U6218 ( .A1(n6761), .A2(n6342), .ZN(n4697) );
  NOR2_X2 U6219 ( .A1(n5079), .A2(n4698), .ZN(n5128) );
  NOR2_X1 U6220 ( .A1(n7478), .A2(n9647), .ZN(n8115) );
  MUX2_X1 U6221 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6333), .S(n6510), .Z(n6506)
         );
  NAND2_X1 U6222 ( .A1(n4710), .A2(n5081), .ZN(n5085) );
  XNOR2_X1 U6223 ( .A(n4710), .B(n5081), .ZN(n6380) );
  NAND2_X1 U6224 ( .A1(n5065), .A2(n5064), .ZN(n4710) );
  NAND2_X1 U6225 ( .A1(n5533), .A2(n4715), .ZN(n4713) );
  NAND2_X1 U6226 ( .A1(n5533), .A2(n5532), .ZN(n4714) );
  NAND2_X1 U6227 ( .A1(n5219), .A2(n4462), .ZN(n4727) );
  NAND2_X1 U6228 ( .A1(n4727), .A2(n4728), .ZN(n5289) );
  NAND2_X1 U6229 ( .A1(n5415), .A2(n4742), .ZN(n4740) );
  NAND2_X1 U6230 ( .A1(n4740), .A2(n4741), .ZN(n5458) );
  NAND2_X1 U6231 ( .A1(n5479), .A2(n4748), .ZN(n4747) );
  NAND2_X1 U6232 ( .A1(n4747), .A2(n4751), .ZN(n5516) );
  NAND2_X1 U6233 ( .A1(n4754), .A2(n4412), .ZN(n4757) );
  INV_X1 U6234 ( .A(n7837), .ZN(n4754) );
  NAND2_X1 U6235 ( .A1(n7837), .A2(n7709), .ZN(n7711) );
  NAND4_X1 U6236 ( .A1(n4758), .A2(n4757), .A3(n4756), .A4(n4755), .ZN(n7741)
         );
  NAND3_X1 U6237 ( .A1(n7837), .A2(n7736), .A3(n4759), .ZN(n4758) );
  AND2_X2 U6238 ( .A1(n4764), .A2(n4762), .ZN(n7582) );
  OR2_X1 U6239 ( .A1(n5613), .A2(n7597), .ZN(n4770) );
  OAI21_X2 U6240 ( .B1(n4768), .B2(n5613), .A(n4767), .ZN(n6596) );
  NAND2_X1 U6241 ( .A1(n4447), .A2(n6408), .ZN(n4767) );
  NAND2_X1 U6242 ( .A1(n7599), .A2(n6408), .ZN(n4768) );
  NAND2_X1 U6243 ( .A1(n7823), .A2(n4461), .ZN(n7207) );
  NAND2_X1 U6244 ( .A1(n4775), .A2(n7677), .ZN(n4771) );
  NAND2_X1 U6245 ( .A1(n4780), .A2(n7813), .ZN(n4773) );
  INV_X1 U6246 ( .A(n4783), .ZN(n7855) );
  NAND2_X1 U6247 ( .A1(n6747), .A2(n6730), .ZN(n6734) );
  NAND3_X1 U6248 ( .A1(n6726), .A2(n6727), .A3(n6725), .ZN(n6747) );
  NAND2_X1 U6249 ( .A1(n4784), .A2(n7783), .ZN(n7719) );
  NAND2_X1 U6250 ( .A1(n4828), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4785) );
  AND2_X2 U6251 ( .A1(n8084), .A2(n8247), .ZN(n6597) );
  NAND2_X1 U6252 ( .A1(n4788), .A2(n4786), .ZN(n7013) );
  NAND2_X1 U6253 ( .A1(n4789), .A2(n4791), .ZN(n7568) );
  NAND2_X1 U6254 ( .A1(n7401), .A2(n7977), .ZN(n4789) );
  INV_X1 U6255 ( .A(n4997), .ZN(n4793) );
  NAND2_X1 U6256 ( .A1(n4796), .A2(n4794), .ZN(n7314) );
  NAND2_X1 U6257 ( .A1(n7059), .A2(n7962), .ZN(n7132) );
  INV_X1 U6258 ( .A(n7962), .ZN(n4798) );
  NAND2_X1 U6259 ( .A1(n5638), .A2(n7923), .ZN(n4800) );
  NAND3_X1 U6260 ( .A1(n4800), .A2(n4801), .A3(n7926), .ZN(n6772) );
  NAND2_X1 U6261 ( .A1(n8405), .A2(n8009), .ZN(n4804) );
  NAND2_X1 U6262 ( .A1(n4804), .A2(n4805), .ZN(n8395) );
  NAND2_X1 U6263 ( .A1(n4808), .A2(n4811), .ZN(n4807) );
  INV_X1 U6264 ( .A(n5052), .ZN(n6798) );
  NAND2_X1 U6265 ( .A1(n4812), .A2(n4814), .ZN(n8290) );
  NAND2_X1 U6266 ( .A1(n4831), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4830) );
  INV_X1 U6267 ( .A(n7239), .ZN(n4829) );
  NAND3_X1 U6268 ( .A1(n4836), .A2(n4835), .A3(P2_REG1_REG_2__SCAN_IN), .ZN(
        n4834) );
  OR2_X1 U6269 ( .A1(n4838), .A2(n4496), .ZN(n4835) );
  NAND2_X1 U6270 ( .A1(n6501), .A2(n6502), .ZN(n6500) );
  NAND3_X1 U6271 ( .A1(n4859), .A2(n4457), .A3(n4860), .ZN(n9305) );
  NAND2_X1 U6272 ( .A1(n4864), .A2(n8867), .ZN(n4863) );
  INV_X1 U6273 ( .A(n8867), .ZN(n4865) );
  NAND2_X1 U6274 ( .A1(n9857), .A2(n4866), .ZN(n7547) );
  NAND2_X1 U6275 ( .A1(n6866), .A2(n4458), .ZN(n4870) );
  NAND2_X1 U6276 ( .A1(n8835), .A2(n8833), .ZN(n6886) );
  NAND2_X1 U6277 ( .A1(n4882), .A2(n4883), .ZN(n4887) );
  NAND2_X1 U6278 ( .A1(n9234), .A2(n4884), .ZN(n4882) );
  OR2_X1 U6279 ( .A1(n9234), .A2(n9233), .ZN(n4886) );
  XNOR2_X1 U6280 ( .A(n4887), .B(n9203), .ZN(n9428) );
  NAND2_X1 U6281 ( .A1(n9863), .A2(n4456), .ZN(n4890) );
  NAND2_X1 U6282 ( .A1(n9318), .A2(n4453), .ZN(n4901) );
  OR2_X1 U6283 ( .A1(n9311), .A2(n9189), .ZN(n4912) );
  NAND2_X1 U6284 ( .A1(n9405), .A2(n4917), .ZN(n4915) );
  NAND2_X1 U6285 ( .A1(n4915), .A2(n4916), .ZN(n9354) );
  INV_X1 U6286 ( .A(n4927), .ZN(n9404) );
  NAND2_X2 U6287 ( .A1(n6798), .A2(n6603), .ZN(n7923) );
  NAND2_X2 U6288 ( .A1(n8113), .A2(n6693), .ZN(n7922) );
  AND4_X2 U6289 ( .A1(n5030), .A2(n5029), .A3(n5031), .A4(n5032), .ZN(n6603)
         );
  NAND2_X1 U6290 ( .A1(n5217), .A2(n4929), .ZN(n4928) );
  NAND2_X1 U6291 ( .A1(n5217), .A2(n5216), .ZN(n7359) );
  NAND2_X1 U6292 ( .A1(n4928), .A2(n4932), .ZN(n5265) );
  NAND2_X1 U6293 ( .A1(n5409), .A2(n8364), .ZN(n4941) );
  NAND2_X1 U6294 ( .A1(n8415), .A2(n4947), .ZN(n4945) );
  NAND2_X1 U6295 ( .A1(n4945), .A2(n4946), .ZN(n8385) );
  NOR2_X2 U6296 ( .A1(n8292), .A2(n5556), .ZN(n8281) );
  AND2_X2 U6297 ( .A1(n4956), .A2(n4415), .ZN(n8292) );
  AND2_X1 U6298 ( .A1(n5002), .A2(n5091), .ZN(n4957) );
  NAND2_X1 U6299 ( .A1(n4959), .A2(n4958), .ZN(n7645) );
  OR2_X2 U6300 ( .A1(n8327), .A2(n5494), .ZN(n4960) );
  AND3_X2 U6301 ( .A1(n5823), .A2(n5708), .A3(n4964), .ZN(n5762) );
  AND2_X1 U6302 ( .A1(n4428), .A2(n4965), .ZN(n4966) );
  NAND3_X1 U6303 ( .A1(n4428), .A2(n5793), .A3(n4965), .ZN(n6581) );
  NAND2_X1 U6304 ( .A1(n4966), .A2(n8629), .ZN(n5794) );
  NAND2_X1 U6305 ( .A1(n6391), .A2(n5087), .ZN(n5845) );
  NAND2_X2 U6306 ( .A1(n6391), .A2(n7868), .ZN(n5826) );
  NAND2_X2 U6307 ( .A1(n4971), .A2(n4969), .ZN(n8734) );
  NAND2_X1 U6308 ( .A1(n8297), .A2(n8296), .ZN(n8515) );
  INV_X1 U6309 ( .A(n6750), .ZN(n6727) );
  CLKBUF_X1 U6310 ( .A(n7055), .Z(n7059) );
  NAND2_X1 U6312 ( .A1(n8457), .A2(n8456), .ZN(n8459) );
  NAND2_X1 U6313 ( .A1(n6828), .A2(n8942), .ZN(n6823) );
  CLKBUF_X1 U6314 ( .A(n7649), .Z(n7650) );
  CLKBUF_X1 U6315 ( .A(n7620), .Z(n7621) );
  CLKBUF_X1 U6316 ( .A(n8690), .Z(n8692) );
  CLKBUF_X1 U6317 ( .A(n9628), .Z(n9629) );
  CLKBUF_X1 U6318 ( .A(n8413), .Z(n8414) );
  NAND2_X1 U6319 ( .A1(n5651), .A2(n5004), .ZN(n5652) );
  BUF_X4 U6320 ( .A(n5074), .Z(n7070) );
  CLKBUF_X1 U6321 ( .A(n5971), .Z(n6242) );
  NAND2_X4 U6322 ( .A1(n6706), .A2(n5781), .ZN(n6234) );
  NOR2_X1 U6323 ( .A1(n5048), .A2(n6510), .ZN(n5068) );
  NAND2_X1 U6324 ( .A1(n4497), .A2(n8589), .ZN(n5050) );
  NAND2_X1 U6325 ( .A1(n5746), .A2(n5745), .ZN(n5837) );
  NAND2_X1 U6326 ( .A1(n5746), .A2(n9568), .ZN(n5971) );
  INV_X1 U6327 ( .A(n5746), .ZN(n7669) );
  INV_X1 U6328 ( .A(n7668), .ZN(n5028) );
  OR2_X1 U6329 ( .A1(n5100), .A2(n6398), .ZN(n5089) );
  INV_X1 U6330 ( .A(n5277), .ZN(n5490) );
  OAI211_X2 U6331 ( .C1(n5809), .C2(n5801), .A(n5808), .B(n5807), .ZN(n6957)
         );
  INV_X1 U6332 ( .A(n10012), .ZN(n10010) );
  NOR2_X1 U6333 ( .A1(n7384), .A2(n7383), .ZN(n4996) );
  NAND2_X1 U6334 ( .A1(n7409), .A2(n7564), .ZN(n4997) );
  INV_X1 U6335 ( .A(n9641), .ZN(n8100) );
  AND4_X1 U6336 ( .A1(n5304), .A2(n5303), .A3(n5302), .A4(n5301), .ZN(n9641)
         );
  OR2_X1 U6337 ( .A1(n9993), .A2(n5685), .ZN(n5001) );
  OR2_X1 U6338 ( .A1(n8110), .A2(n6954), .ZN(n5002) );
  INV_X1 U6339 ( .A(n7808), .ZN(n8356) );
  AND2_X1 U6340 ( .A1(n5474), .A2(n5473), .ZN(n7808) );
  OAI21_X1 U6341 ( .B1(n8930), .B2(n8929), .A(n8928), .ZN(n8931) );
  OR2_X1 U6342 ( .A1(n9904), .A2(n9131), .ZN(n9345) );
  INV_X1 U6343 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U6344 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5003) );
  OR2_X1 U6345 ( .A1(n8562), .A2(n8433), .ZN(n5004) );
  INV_X1 U6346 ( .A(n8757), .ZN(n6052) );
  INV_X1 U6347 ( .A(n8406), .ZN(n5653) );
  NAND2_X1 U6348 ( .A1(n8501), .A2(n8272), .ZN(n5005) );
  AND2_X1 U6349 ( .A1(n5684), .A2(n5683), .ZN(n9994) );
  INV_X1 U6350 ( .A(n7916), .ZN(n6598) );
  NOR2_X1 U6351 ( .A1(n5080), .A2(n6380), .ZN(n5006) );
  INV_X1 U6352 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5012) );
  INV_X1 U6353 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5709) );
  INV_X1 U6354 ( .A(n8392), .ZN(n7902) );
  OR2_X1 U6355 ( .A1(n7218), .A2(n9698), .ZN(n5961) );
  INV_X1 U6356 ( .A(n8923), .ZN(n8924) );
  AND4_X1 U6357 ( .A1(n5712), .A2(n5711), .A3(n5710), .A4(n5709), .ZN(n5713)
         );
  INV_X1 U6358 ( .A(n7945), .ZN(n5642) );
  AND2_X1 U6359 ( .A1(n7221), .A2(n5961), .ZN(n5962) );
  INV_X1 U6360 ( .A(n8724), .ZN(n6117) );
  INV_X1 U6361 ( .A(n5280), .ZN(n5279) );
  OR2_X1 U6362 ( .A1(n7346), .A2(n7345), .ZN(n7347) );
  NOR2_X1 U6363 ( .A1(n5006), .A2(n5068), .ZN(n5070) );
  INV_X1 U6364 ( .A(n6818), .ZN(n5870) );
  NOR2_X1 U6365 ( .A1(n6187), .A2(n8606), .ZN(n6206) );
  AND2_X1 U6366 ( .A1(n6206), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n6225) );
  INV_X1 U6367 ( .A(n5327), .ZN(n5329) );
  INV_X1 U6368 ( .A(n5180), .ZN(n5181) );
  INV_X1 U6369 ( .A(n7004), .ZN(n7001) );
  INV_X1 U6370 ( .A(n5299), .ZN(n5298) );
  INV_X1 U6371 ( .A(n6735), .ZN(n6731) );
  INV_X1 U6372 ( .A(n5377), .ZN(n5376) );
  INV_X1 U6373 ( .A(n5524), .ZN(n5523) );
  INV_X1 U6374 ( .A(n5449), .ZN(n5448) );
  INV_X1 U6375 ( .A(n7957), .ZN(n5644) );
  OR2_X1 U6376 ( .A1(n5093), .A2(n5043), .ZN(n5046) );
  AND2_X1 U6377 ( .A1(n8070), .A2(n5634), .ZN(n5688) );
  NAND2_X1 U6378 ( .A1(n8304), .A2(n8388), .ZN(n8283) );
  INV_X1 U6379 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5589) );
  OR2_X1 U6380 ( .A1(n6171), .A2(n6170), .ZN(n6187) );
  NAND2_X1 U6381 ( .A1(n6156), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n6171) );
  INV_X1 U6382 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10288) );
  OR2_X1 U6383 ( .A1(n6108), .A2(n6107), .ZN(n6124) );
  OR2_X1 U6384 ( .A1(n6036), .A2(n6035), .ZN(n6054) );
  OR2_X1 U6385 ( .A1(n7181), .A2(n9030), .ZN(n7182) );
  AND2_X1 U6386 ( .A1(n7605), .A2(n9023), .ZN(n7606) );
  OR2_X1 U6387 ( .A1(n9664), .A2(n9027), .ZN(n7416) );
  INV_X1 U6388 ( .A(n6391), .ZN(n6120) );
  OR2_X1 U6389 ( .A1(n9033), .A2(n7119), .ZN(n6881) );
  OR2_X1 U6390 ( .A1(n7047), .A2(n9034), .ZN(n6824) );
  INV_X1 U6391 ( .A(SI_29_), .ZN(n5578) );
  NOR2_X1 U6392 ( .A1(n5329), .A2(n5328), .ZN(n5330) );
  NAND2_X1 U6393 ( .A1(n5239), .A2(n10151), .ZN(n5250) );
  OR2_X1 U6394 ( .A1(n5401), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5423) );
  AND2_X1 U6395 ( .A1(n7390), .A2(n7389), .ZN(n7391) );
  AND2_X1 U6396 ( .A1(n7675), .A2(n8099), .ZN(n7766) );
  AND2_X1 U6397 ( .A1(n7755), .A2(n7701), .ZN(n7784) );
  INV_X1 U6398 ( .A(n7074), .ZN(n5600) );
  OR2_X1 U6399 ( .A1(n5545), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5563) );
  OR2_X1 U6400 ( .A1(n5486), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5507) );
  AND2_X1 U6401 ( .A1(n8016), .A2(n8014), .ZN(n8392) );
  OR2_X1 U6402 ( .A1(n5320), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6403 ( .A1(n6071), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6108) );
  OR2_X1 U6404 ( .A1(n6429), .A2(n6430), .ZN(n9095) );
  AND2_X1 U6405 ( .A1(n9162), .A2(n8787), .ZN(n9217) );
  AND2_X1 U6406 ( .A1(n9157), .A2(n8905), .ZN(n9274) );
  INV_X1 U6407 ( .A(n9025), .ZN(n7466) );
  NAND2_X1 U6408 ( .A1(n5805), .A2(n5804), .ZN(n5808) );
  AND2_X1 U6409 ( .A1(n7434), .A2(n4403), .ZN(n6703) );
  AND2_X1 U6410 ( .A1(n6710), .A2(n6709), .ZN(n9854) );
  XNOR2_X1 U6411 ( .A(n5310), .B(SI_14_), .ZN(n5307) );
  NAND2_X1 U6412 ( .A1(n5146), .A2(SI_5_), .ZN(n5147) );
  AOI21_X1 U6413 ( .B1(n8419), .B2(n7681), .A(n7817), .ZN(n7726) );
  AND2_X1 U6414 ( .A1(n6604), .A2(n6605), .ZN(n7826) );
  INV_X1 U6415 ( .A(n7856), .ZN(n7839) );
  OR2_X1 U6416 ( .A1(n5663), .A2(n5580), .ZN(n7077) );
  AND4_X1 U6417 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n8433)
         );
  INV_X1 U6418 ( .A(n8264), .ZN(n8226) );
  AND3_X1 U6419 ( .A1(n5681), .A2(n5633), .A3(n5676), .ZN(n5696) );
  INV_X1 U6420 ( .A(n8516), .ZN(n8568) );
  AND2_X1 U6421 ( .A1(n5223), .A2(n5254), .ZN(n7248) );
  INV_X1 U6422 ( .A(n9660), .ZN(n6298) );
  NAND2_X1 U6423 ( .A1(n5918), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5951) );
  OR2_X1 U6424 ( .A1(n6011), .A2(n5748), .ZN(n6036) );
  INV_X1 U6425 ( .A(n9656), .ZN(n9713) );
  AND2_X1 U6426 ( .A1(n9158), .A2(n8907), .ZN(n9262) );
  OAI22_X1 U6427 ( .A1(n9354), .A2(n9181), .B1(n9180), .B2(n9545), .ZN(n9333)
         );
  INV_X1 U6428 ( .A(n9854), .ZN(n9402) );
  OR3_X1 U6429 ( .A1(n6904), .A2(n6901), .A3(n6701), .ZN(n6714) );
  AND2_X1 U6430 ( .A1(n6390), .A2(n6295), .ZN(n9004) );
  XNOR2_X1 U6431 ( .A(n5169), .B(SI_6_), .ZN(n5167) );
  XNOR2_X1 U6432 ( .A(n5103), .B(n10113), .ZN(n5101) );
  INV_X1 U6433 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10014) );
  NOR2_X1 U6434 ( .A1(n9617), .A2(n10361), .ZN(n9618) );
  AND2_X1 U6435 ( .A1(n5619), .A2(n7640), .ZN(n6522) );
  INV_X1 U6436 ( .A(n7861), .ZN(n7848) );
  INV_X1 U6437 ( .A(n7843), .ZN(n8304) );
  INV_X1 U6438 ( .A(n7586), .ZN(n8101) );
  INV_X1 U6439 ( .A(n8267), .ZN(n8237) );
  INV_X1 U6440 ( .A(n5669), .ZN(n5670) );
  OR2_X1 U6441 ( .A1(n9648), .A2(n9630), .ZN(n8448) );
  AND2_X1 U6442 ( .A1(n5662), .A2(n9632), .ZN(n9648) );
  XOR2_X1 U6443 ( .A(n8279), .B(n8278), .Z(n8514) );
  OR2_X1 U6444 ( .A1(n9994), .A2(n9986), .ZN(n8572) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6465) );
  INV_X1 U6446 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6463) );
  INV_X1 U6447 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6381) );
  OR2_X1 U6448 ( .A1(n6313), .A2(n6297), .ZN(n9660) );
  INV_X1 U6449 ( .A(n9728), .ZN(n9852) );
  AND2_X1 U6450 ( .A1(n6905), .A2(n9413), .ZN(n9421) );
  INV_X1 U6451 ( .A(n9416), .ZN(n9904) );
  NAND2_X1 U6452 ( .A1(n9932), .A2(n9495), .ZN(n9491) );
  OR2_X1 U6453 ( .A1(n6714), .A2(n6702), .ZN(n9929) );
  INV_X1 U6454 ( .A(n9342), .ZN(n9541) );
  OR2_X1 U6455 ( .A1(n6714), .A2(n6903), .ZN(n9557) );
  NAND2_X1 U6456 ( .A1(n9004), .A2(n6386), .ZN(n9906) );
  INV_X1 U6457 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10259) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6383) );
  INV_X1 U6459 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6374) );
  NOR2_X1 U6460 ( .A1(n10362), .A2(n6365), .ZN(n10361) );
  NOR2_X1 U6461 ( .A1(n9623), .A2(n10368), .ZN(n10047) );
  AND2_X1 U6462 ( .A1(n6412), .A2(n6522), .ZN(P2_U3893) );
  NAND2_X1 U6463 ( .A1(n5128), .A2(n5129), .ZN(n5148) );
  NOR2_X1 U6464 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5011) );
  NOR2_X1 U6465 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5015) );
  NOR2_X1 U6466 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5014) );
  NAND4_X1 U6467 ( .A1(n5015), .A2(n5014), .A3(n5589), .A4(n10267), .ZN(n5016)
         );
  INV_X1 U6468 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5017) );
  INV_X1 U6469 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5018) );
  NOR2_X1 U6470 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n5019) );
  INV_X1 U6471 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5020) );
  NAND2_X1 U6472 ( .A1(n5022), .A2(n5020), .ZN(n5024) );
  INV_X1 U6473 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8574) );
  XNOR2_X2 U6474 ( .A(n5025), .B(n8574), .ZN(n7668) );
  NAND2_X1 U6475 ( .A1(n5027), .A2(n7668), .ZN(n5276) );
  INV_X1 U6476 ( .A(n5276), .ZN(n5026) );
  NAND2_X1 U6477 ( .A1(n5026), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5032) );
  NAND2_X1 U6478 ( .A1(n5277), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5031) );
  INV_X1 U6479 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6608) );
  NAND2_X1 U6480 ( .A1(n5074), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5029) );
  INV_X1 U6481 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n10341) );
  XNOR2_X2 U6482 ( .A(n5033), .B(n10341), .ZN(n8087) );
  NAND2_X1 U6483 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n5034) );
  AOI22_X1 U6484 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n5021), .B1(n5034), .B2(
        P2_IR_REG_31__SCAN_IN), .ZN(n5035) );
  INV_X1 U6485 ( .A(n5035), .ZN(n5036) );
  OAI21_X1 U6486 ( .B1(n5614), .B2(n5003), .A(n5036), .ZN(n5037) );
  NAND2_X4 U6487 ( .A1(n5039), .A2(n5038), .ZN(n8253) );
  INV_X1 U6488 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6377) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6397) );
  XNOR2_X1 U6490 ( .A(n5062), .B(SI_1_), .ZN(n5061) );
  MUX2_X1 U6491 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(P2_DATAO_REG_0__SCAN_IN), 
        .S(n5086), .Z(n5040) );
  NAND2_X1 U6492 ( .A1(n5040), .A2(SI_0_), .ZN(n5059) );
  XNOR2_X1 U6493 ( .A(n5061), .B(n5059), .ZN(n6376) );
  NAND2_X1 U6494 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5041) );
  XNOR2_X1 U6495 ( .A(n5041), .B(P2_IR_REG_1__SCAN_IN), .ZN(n6347) );
  OR2_X1 U6496 ( .A1(n5048), .A2(n6347), .ZN(n5042) );
  NAND2_X1 U6497 ( .A1(n5074), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5047) );
  INV_X1 U6498 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5043) );
  NAND2_X1 U6499 ( .A1(n5026), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5045) );
  NAND2_X1 U6500 ( .A1(n5277), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5044) );
  INV_X1 U6501 ( .A(n6607), .ZN(n6687) );
  NAND2_X1 U6502 ( .A1(n5087), .A2(SI_0_), .ZN(n5049) );
  XNOR2_X1 U6503 ( .A(n5049), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8589) );
  OAI21_X2 U6504 ( .B1(n4497), .B2(n5051), .A(n5050), .ZN(n6601) );
  NAND2_X1 U6505 ( .A1(n6779), .A2(n6693), .ZN(n5053) );
  NAND2_X1 U6506 ( .A1(n6685), .A2(n5053), .ZN(n6777) );
  NAND2_X1 U6507 ( .A1(n5074), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5055) );
  NAND2_X1 U6508 ( .A1(n5277), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5054) );
  AND2_X1 U6509 ( .A1(n5055), .A2(n5054), .ZN(n5058) );
  NAND2_X1 U6510 ( .A1(n5026), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5057) );
  NAND2_X1 U6511 ( .A1(n5073), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5056) );
  INV_X1 U6512 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6513 ( .A1(n5061), .A2(n5060), .ZN(n5065) );
  INV_X1 U6514 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6515 ( .A1(n5063), .A2(SI_1_), .ZN(n5064) );
  MUX2_X1 U6516 ( .A(n6381), .B(n6374), .S(n5086), .Z(n5082) );
  XNOR2_X1 U6517 ( .A(n5082), .B(SI_2_), .ZN(n5081) );
  OR2_X1 U6518 ( .A1(n5106), .A2(n6381), .ZN(n5069) );
  INV_X2 U6519 ( .A(n6614), .ZN(n5071) );
  NAND2_X1 U6520 ( .A1(n6777), .A2(n6778), .ZN(n6776) );
  INV_X1 U6521 ( .A(n8112), .ZN(n6724) );
  NAND2_X1 U6522 ( .A1(n6724), .A2(n5071), .ZN(n5072) );
  NAND2_X1 U6523 ( .A1(n5277), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5078) );
  NAND2_X1 U6524 ( .A1(n5548), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U6525 ( .A1(n5073), .A2(n6806), .ZN(n5076) );
  NAND2_X1 U6526 ( .A1(n7070), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5075) );
  AND4_X2 U6527 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n6949)
         );
  INV_X1 U6528 ( .A(n6949), .ZN(n5640) );
  CLKBUF_X1 U6529 ( .A(n5640), .Z(n8111) );
  INV_X1 U6530 ( .A(n5082), .ZN(n5083) );
  NAND2_X1 U6531 ( .A1(n5083), .A2(SI_2_), .ZN(n5084) );
  NAND2_X1 U6532 ( .A1(n5085), .A2(n5084), .ZN(n5102) );
  INV_X4 U6533 ( .A(n5086), .ZN(n5087) );
  XNOR2_X1 U6534 ( .A(n5102), .B(n5101), .ZN(n6398) );
  INV_X1 U6535 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6370) );
  OR2_X1 U6536 ( .A1(n5106), .A2(n6370), .ZN(n5088) );
  OAI211_X1 U6537 ( .C1(n4497), .C2(n6559), .A(n5089), .B(n5088), .ZN(n9937)
         );
  NAND2_X1 U6538 ( .A1(n8111), .A2(n9937), .ZN(n5090) );
  NAND2_X1 U6539 ( .A1(n6802), .A2(n5090), .ZN(n5092) );
  INV_X1 U6540 ( .A(n9937), .ZN(n6746) );
  NAND2_X1 U6541 ( .A1(n6949), .A2(n6746), .ZN(n5091) );
  NAND2_X1 U6542 ( .A1(n5548), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6543 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5095) );
  NAND2_X1 U6544 ( .A1(n5115), .A2(n5095), .ZN(n6953) );
  NAND2_X1 U6545 ( .A1(n5547), .A2(n6953), .ZN(n5098) );
  NAND2_X1 U6546 ( .A1(n7070), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6547 ( .A1(n5277), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5096) );
  NAND2_X1 U6548 ( .A1(n5102), .A2(n5101), .ZN(n5105) );
  NAND2_X1 U6549 ( .A1(n5103), .A2(SI_3_), .ZN(n5104) );
  XNOR2_X1 U6550 ( .A(n5122), .B(n5121), .ZN(n6378) );
  OR2_X1 U6551 ( .A1(n5100), .A2(n6378), .ZN(n5112) );
  OR2_X1 U6552 ( .A1(n7873), .A2(n6379), .ZN(n5111) );
  NAND2_X1 U6553 ( .A1(n5107), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5109) );
  INV_X1 U6554 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5108) );
  OR2_X1 U6555 ( .A1(n4497), .A2(n6674), .ZN(n5110) );
  AND3_X2 U6556 ( .A1(n5112), .A2(n5111), .A3(n5110), .ZN(n9944) );
  NAND2_X1 U6557 ( .A1(n8110), .A2(n6954), .ZN(n6944) );
  NAND2_X1 U6558 ( .A1(n5548), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5120) );
  NAND2_X1 U6559 ( .A1(n5115), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6560 ( .A1(n5137), .A2(n5116), .ZN(n6938) );
  NAND2_X1 U6561 ( .A1(n5547), .A2(n6938), .ZN(n5119) );
  NAND2_X1 U6562 ( .A1(n7071), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U6563 ( .A1(n7070), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5117) );
  NAND4_X1 U6564 ( .A1(n5120), .A2(n5119), .A3(n5118), .A4(n5117), .ZN(n8109)
         );
  INV_X1 U6565 ( .A(n8109), .ZN(n7829) );
  NAND2_X1 U6566 ( .A1(n5122), .A2(n5121), .ZN(n5126) );
  INV_X1 U6567 ( .A(n5123), .ZN(n5124) );
  INV_X1 U6568 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5127) );
  XNOR2_X1 U6569 ( .A(n5144), .B(n5143), .ZN(n6372) );
  OR2_X1 U6570 ( .A1(n5100), .A2(n6372), .ZN(n5133) );
  OR2_X1 U6571 ( .A1(n7873), .A2(n6373), .ZN(n5132) );
  OR2_X1 U6572 ( .A1(n5128), .A2(n5021), .ZN(n5130) );
  XNOR2_X1 U6573 ( .A(n5130), .B(n5129), .ZN(n6771) );
  OR2_X1 U6574 ( .A1(n4497), .A2(n6771), .ZN(n5131) );
  NAND2_X1 U6575 ( .A1(n7829), .A2(n9949), .ZN(n5134) );
  NAND2_X1 U6576 ( .A1(n6936), .A2(n5134), .ZN(n5136) );
  INV_X1 U6577 ( .A(n9949), .ZN(n6939) );
  NAND2_X1 U6578 ( .A1(n8109), .A2(n6939), .ZN(n5135) );
  NAND2_X1 U6579 ( .A1(n5136), .A2(n5135), .ZN(n7016) );
  INV_X1 U6580 ( .A(n7016), .ZN(n5155) );
  NAND2_X1 U6581 ( .A1(n5548), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6582 ( .A1(n5137), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6583 ( .A1(n5160), .A2(n5138), .ZN(n7832) );
  NAND2_X1 U6584 ( .A1(n5547), .A2(n7832), .ZN(n5141) );
  NAND2_X1 U6585 ( .A1(n7071), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5140) );
  NAND2_X1 U6586 ( .A1(n7070), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5139) );
  NAND4_X1 U6587 ( .A1(n5142), .A2(n5141), .A3(n5140), .A4(n5139), .ZN(n8108)
         );
  INV_X1 U6588 ( .A(n5145), .ZN(n5146) );
  XNOR2_X1 U6589 ( .A(n5168), .B(n5167), .ZN(n6384) );
  OR2_X1 U6590 ( .A1(n5100), .A2(n6384), .ZN(n5154) );
  OR2_X1 U6591 ( .A1(n7873), .A2(n6385), .ZN(n5153) );
  NAND2_X1 U6592 ( .A1(n5149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5150) );
  MUX2_X1 U6593 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5150), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5151) );
  NAND2_X1 U6594 ( .A1(n5151), .A2(n5190), .ZN(n6980) );
  OR2_X1 U6595 ( .A1(n4497), .A2(n6980), .ZN(n5152) );
  INV_X1 U6596 ( .A(n9955), .ZN(n7831) );
  NAND2_X1 U6597 ( .A1(n5155), .A2(n4420), .ZN(n5157) );
  INV_X1 U6598 ( .A(n8108), .ZN(n7006) );
  NAND2_X1 U6599 ( .A1(n7006), .A2(n9955), .ZN(n5156) );
  NAND2_X1 U6600 ( .A1(n5157), .A2(n5156), .ZN(n7060) );
  NAND2_X1 U6601 ( .A1(n7071), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6602 ( .A1(n5548), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5164) );
  NAND2_X1 U6603 ( .A1(n5160), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6604 ( .A1(n5174), .A2(n5161), .ZN(n7005) );
  NAND2_X1 U6605 ( .A1(n5073), .A2(n7005), .ZN(n5163) );
  NAND2_X1 U6606 ( .A1(n7070), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6607 ( .A1(n5190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5166) );
  XNOR2_X1 U6608 ( .A(n5166), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7025) );
  AOI22_X1 U6609 ( .A1(n5398), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5397), .B2(
        n7025), .ZN(n5172) );
  INV_X1 U6610 ( .A(n5169), .ZN(n5170) );
  XNOR2_X1 U6611 ( .A(n5182), .B(n5180), .ZN(n6400) );
  NAND2_X1 U6612 ( .A1(n6400), .A2(n7872), .ZN(n5171) );
  NAND2_X1 U6613 ( .A1(n5172), .A2(n5171), .ZN(n7067) );
  NAND2_X1 U6614 ( .A1(n7204), .A2(n7067), .ZN(n7958) );
  INV_X1 U6615 ( .A(n7067), .ZN(n9959) );
  NAND2_X1 U6616 ( .A1(n8107), .A2(n9959), .ZN(n7962) );
  NAND2_X1 U6617 ( .A1(n7958), .A2(n7962), .ZN(n7957) );
  NAND2_X1 U6618 ( .A1(n7204), .A2(n9959), .ZN(n5173) );
  NAND2_X1 U6619 ( .A1(n5548), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U6620 ( .A1(n5174), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5175) );
  NAND2_X1 U6621 ( .A1(n5209), .A2(n5175), .ZN(n7210) );
  NAND2_X1 U6622 ( .A1(n5547), .A2(n7210), .ZN(n5178) );
  NAND2_X1 U6623 ( .A1(n7071), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6624 ( .A1(n7070), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5176) );
  NAND4_X1 U6625 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n8106)
         );
  INV_X1 U6626 ( .A(n8106), .ZN(n7340) );
  NAND2_X1 U6627 ( .A1(n5182), .A2(n5181), .ZN(n5185) );
  NAND2_X1 U6628 ( .A1(n5183), .A2(SI_7_), .ZN(n5184) );
  INV_X1 U6629 ( .A(SI_8_), .ZN(n5186) );
  NAND2_X1 U6630 ( .A1(n5187), .A2(n5186), .ZN(n5195) );
  INV_X1 U6631 ( .A(n5187), .ZN(n5188) );
  NAND2_X1 U6632 ( .A1(n5188), .A2(SI_8_), .ZN(n5189) );
  XNOR2_X1 U6633 ( .A(n5197), .B(n5196), .ZN(n6404) );
  NAND2_X1 U6634 ( .A1(n6404), .A2(n7872), .ZN(n5193) );
  OR2_X1 U6635 ( .A1(n5335), .A2(n5021), .ZN(n5191) );
  XNOR2_X1 U6636 ( .A(n5191), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7151) );
  AOI22_X1 U6637 ( .A1(n5398), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5397), .B2(
        n7151), .ZN(n5192) );
  NAND2_X1 U6638 ( .A1(n7340), .A2(n7209), .ZN(n7959) );
  AND2_X1 U6639 ( .A1(n9965), .A2(n8106), .ZN(n5646) );
  INV_X1 U6640 ( .A(n5646), .ZN(n7963) );
  NAND2_X1 U6641 ( .A1(n7959), .A2(n7963), .ZN(n7892) );
  INV_X1 U6642 ( .A(n7892), .ZN(n7127) );
  NAND2_X1 U6643 ( .A1(n7209), .A2(n8106), .ZN(n5194) );
  NAND2_X1 U6644 ( .A1(n7130), .A2(n5194), .ZN(n7317) );
  INV_X1 U6645 ( .A(SI_9_), .ZN(n5198) );
  INV_X1 U6646 ( .A(n5199), .ZN(n5200) );
  NAND2_X1 U6647 ( .A1(n5200), .A2(SI_9_), .ZN(n5201) );
  OR2_X1 U6648 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U6649 ( .A1(n5219), .A2(n5204), .ZN(n6460) );
  NAND2_X1 U6650 ( .A1(n6460), .A2(n7872), .ZN(n5207) );
  INV_X1 U6651 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U6652 ( .A1(n5335), .A2(n10342), .ZN(n5220) );
  NAND2_X1 U6653 ( .A1(n5220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6654 ( .A(n5205), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7158) );
  AOI22_X1 U6655 ( .A1(n5398), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5397), .B2(
        n7158), .ZN(n5206) );
  NAND2_X1 U6656 ( .A1(n5207), .A2(n5206), .ZN(n7325) );
  INV_X1 U6657 ( .A(n7325), .ZN(n9970) );
  NAND2_X1 U6658 ( .A1(n5548), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5214) );
  NAND2_X1 U6659 ( .A1(n7070), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6660 ( .A1(n5209), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6661 ( .A1(n5225), .A2(n5210), .ZN(n7321) );
  NAND2_X1 U6662 ( .A1(n5073), .A2(n7321), .ZN(n5212) );
  NAND2_X1 U6663 ( .A1(n7071), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5211) );
  NAND2_X1 U6664 ( .A1(n9970), .A2(n7361), .ZN(n5215) );
  INV_X1 U6665 ( .A(n7361), .ZN(n8105) );
  NAND2_X1 U6666 ( .A1(n8105), .A2(n7325), .ZN(n5216) );
  XNOR2_X1 U6667 ( .A(n5237), .B(n5232), .ZN(n6464) );
  NAND2_X1 U6668 ( .A1(n5222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5221) );
  MUX2_X1 U6669 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5221), .S(
        P2_IR_REG_10__SCAN_IN), .Z(n5223) );
  AOI22_X1 U6670 ( .A1(n5398), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5397), .B2(
        n7248), .ZN(n5224) );
  NAND2_X1 U6671 ( .A1(n5548), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6672 ( .A1(n5225), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6673 ( .A1(n5259), .A2(n5226), .ZN(n7350) );
  NAND2_X1 U6674 ( .A1(n5547), .A2(n7350), .ZN(n5229) );
  NAND2_X1 U6675 ( .A1(n7071), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5228) );
  NAND2_X1 U6676 ( .A1(n7070), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5227) );
  NAND4_X1 U6677 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n8104)
         );
  NOR2_X1 U6678 ( .A1(n9975), .A2(n7381), .ZN(n7385) );
  NAND2_X1 U6679 ( .A1(n9975), .A2(n7381), .ZN(n5231) );
  INV_X1 U6680 ( .A(n5233), .ZN(n5234) );
  INV_X1 U6681 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n5238) );
  INV_X1 U6682 ( .A(SI_11_), .ZN(n10151) );
  INV_X1 U6683 ( .A(n5239), .ZN(n5240) );
  NAND2_X1 U6684 ( .A1(n5240), .A2(SI_11_), .ZN(n5241) );
  XNOR2_X1 U6685 ( .A(n5252), .B(n5251), .ZN(n6488) );
  NAND2_X1 U6686 ( .A1(n6488), .A2(n7872), .ZN(n5244) );
  NAND2_X1 U6687 ( .A1(n5254), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5242) );
  AOI22_X1 U6688 ( .A1(n5398), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5397), .B2(
        n7490), .ZN(n5243) );
  NAND2_X1 U6689 ( .A1(n7071), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5248) );
  NAND2_X1 U6690 ( .A1(n5548), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5247) );
  INV_X2 U6691 ( .A(n5580), .ZN(n5547) );
  XNOR2_X1 U6692 ( .A(n5259), .B(P2_REG3_REG_11__SCAN_IN), .ZN(n7374) );
  NAND2_X1 U6693 ( .A1(n5547), .A2(n7374), .ZN(n5246) );
  NAND2_X1 U6694 ( .A1(n7070), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5245) );
  NOR2_X1 U6695 ( .A1(n7409), .A2(n8103), .ZN(n5249) );
  INV_X1 U6696 ( .A(n7409), .ZN(n9981) );
  INV_X1 U6697 ( .A(SI_12_), .ZN(n5253) );
  XNOR2_X1 U6698 ( .A(n5270), .B(n5268), .ZN(n6569) );
  NAND2_X1 U6699 ( .A1(n6569), .A2(n7872), .ZN(n5257) );
  NOR2_X1 U6700 ( .A1(n5254), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5272) );
  OR2_X1 U6701 ( .A1(n5272), .A2(n5021), .ZN(n5255) );
  XNOR2_X1 U6702 ( .A(n5255), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7542) );
  AOI22_X1 U6703 ( .A1(n5398), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5397), .B2(
        n7542), .ZN(n5256) );
  NAND2_X1 U6704 ( .A1(n5548), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5264) );
  OAI21_X1 U6705 ( .B1(n5259), .B2(P2_REG3_REG_11__SCAN_IN), .A(
        P2_REG3_REG_12__SCAN_IN), .ZN(n5260) );
  INV_X1 U6706 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10285) );
  INV_X1 U6707 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7395) );
  NAND2_X1 U6708 ( .A1(n10285), .A2(n7395), .ZN(n5258) );
  NAND2_X1 U6709 ( .A1(n5260), .A2(n5280), .ZN(n7394) );
  NAND2_X1 U6710 ( .A1(n5547), .A2(n7394), .ZN(n5263) );
  NAND2_X1 U6711 ( .A1(n7071), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6712 ( .A1(n7070), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5261) );
  NAND4_X1 U6713 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n8102)
         );
  NAND2_X1 U6714 ( .A1(n5265), .A2(n9639), .ZN(n5267) );
  INV_X1 U6715 ( .A(n7562), .ZN(n5266) );
  XNOR2_X1 U6716 ( .A(n5289), .B(n5287), .ZN(n6587) );
  NAND2_X1 U6717 ( .A1(n6587), .A2(n7872), .ZN(n5275) );
  INV_X1 U6718 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5271) );
  NAND2_X1 U6719 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  NAND2_X1 U6720 ( .A1(n5273), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5294) );
  XNOR2_X1 U6721 ( .A(n5294), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8132) );
  AOI22_X1 U6722 ( .A1(n5398), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5397), .B2(
        n8132), .ZN(n5274) );
  NAND2_X1 U6723 ( .A1(n5600), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5285) );
  NAND2_X1 U6724 ( .A1(n7071), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5284) );
  INV_X1 U6725 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6726 ( .A1(n5280), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6727 ( .A1(n5299), .A2(n5281), .ZN(n7517) );
  NAND2_X1 U6728 ( .A1(n5547), .A2(n7517), .ZN(n5283) );
  NAND2_X1 U6729 ( .A1(n7070), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6730 ( .A1(n9631), .A2(n8101), .ZN(n7883) );
  NAND2_X1 U6731 ( .A1(n9636), .A2(n7883), .ZN(n5286) );
  NAND2_X1 U6732 ( .A1(n5286), .A2(n7884), .ZN(n7622) );
  NAND2_X1 U6733 ( .A1(n5289), .A2(n5288), .ZN(n5292) );
  NAND2_X1 U6734 ( .A1(n5290), .A2(SI_13_), .ZN(n5291) );
  XNOR2_X1 U6735 ( .A(n5309), .B(n5307), .ZN(n6651) );
  NAND2_X1 U6736 ( .A1(n6651), .A2(n7872), .ZN(n5297) );
  INV_X1 U6737 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5293) );
  NAND2_X1 U6738 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  NAND2_X1 U6739 ( .A1(n5295), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5314) );
  XNOR2_X1 U6740 ( .A(n5314), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8136) );
  AOI22_X1 U6741 ( .A1(n8136), .A2(n5397), .B1(n5398), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6742 ( .A1(n7071), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5304) );
  NAND2_X1 U6743 ( .A1(n5548), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5303) );
  INV_X1 U6744 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10192) );
  NAND2_X1 U6745 ( .A1(n5299), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5300) );
  NAND2_X1 U6746 ( .A1(n5320), .A2(n5300), .ZN(n7631) );
  NAND2_X1 U6747 ( .A1(n5547), .A2(n7631), .ZN(n5302) );
  NAND2_X1 U6748 ( .A1(n7070), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5301) );
  NAND2_X1 U6749 ( .A1(n7627), .A2(n8100), .ZN(n5305) );
  OR2_X1 U6750 ( .A1(n7627), .A2(n8100), .ZN(n5306) );
  NAND2_X1 U6751 ( .A1(n5310), .A2(SI_14_), .ZN(n5311) );
  XNOR2_X1 U6752 ( .A(n5327), .B(SI_15_), .ZN(n5312) );
  XNOR2_X1 U6753 ( .A(n5331), .B(n5312), .ZN(n6718) );
  NAND2_X1 U6754 ( .A1(n6718), .A2(n7872), .ZN(n5319) );
  INV_X1 U6755 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5313) );
  NAND2_X1 U6756 ( .A1(n5314), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U6757 ( .A1(n5315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5316) );
  XNOR2_X1 U6758 ( .A(n5316), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8185) );
  INV_X1 U6759 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10242) );
  NOR2_X1 U6760 ( .A1(n7873), .A2(n10242), .ZN(n5317) );
  AOI21_X1 U6761 ( .B1(n8185), .B2(n5397), .A(n5317), .ZN(n5318) );
  NAND2_X1 U6762 ( .A1(n5600), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5325) );
  NAND2_X1 U6763 ( .A1(n7071), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6764 ( .A1(n5320), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6765 ( .A1(n5341), .A2(n5321), .ZN(n8442) );
  NAND2_X1 U6766 ( .A1(n5547), .A2(n8442), .ZN(n5323) );
  NAND2_X1 U6767 ( .A1(n7070), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5322) );
  NAND2_X1 U6768 ( .A1(n8445), .A2(n8432), .ZN(n7998) );
  NAND2_X1 U6769 ( .A1(n7995), .A2(n7998), .ZN(n7899) );
  INV_X1 U6770 ( .A(n8432), .ZN(n8099) );
  NAND2_X1 U6771 ( .A1(n8445), .A2(n8099), .ZN(n5326) );
  INV_X1 U6772 ( .A(SI_15_), .ZN(n5328) );
  INV_X1 U6773 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10154) );
  INV_X1 U6774 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5332) );
  XNOR2_X1 U6775 ( .A(n5349), .B(SI_16_), .ZN(n5333) );
  XNOR2_X1 U6776 ( .A(n5352), .B(n5333), .ZN(n6741) );
  NAND2_X1 U6777 ( .A1(n6741), .A2(n7872), .ZN(n5338) );
  NAND2_X1 U6778 ( .A1(n5335), .A2(n5334), .ZN(n5357) );
  NAND2_X1 U6779 ( .A1(n5357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5336) );
  XNOR2_X1 U6780 ( .A(n5336), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8193) );
  AOI22_X1 U6781 ( .A1(n5398), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5397), .B2(
        n8193), .ZN(n5337) );
  NAND2_X1 U6782 ( .A1(n7071), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5346) );
  NAND2_X1 U6783 ( .A1(n5600), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5345) );
  INV_X1 U6784 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6785 ( .A1(n5341), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5342) );
  NAND2_X1 U6786 ( .A1(n5362), .A2(n5342), .ZN(n8437) );
  NAND2_X1 U6787 ( .A1(n5547), .A2(n8437), .ZN(n5344) );
  NAND2_X1 U6788 ( .A1(n7070), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6789 ( .A1(n8569), .A2(n8418), .ZN(n8006) );
  INV_X1 U6790 ( .A(n8430), .ZN(n5347) );
  NAND2_X1 U6791 ( .A1(n8429), .A2(n5347), .ZN(n8435) );
  INV_X1 U6792 ( .A(n8418), .ZN(n8098) );
  NAND2_X1 U6793 ( .A1(n8569), .A2(n8098), .ZN(n5348) );
  NOR2_X1 U6794 ( .A1(n5350), .A2(SI_16_), .ZN(n5351) );
  INV_X1 U6795 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6899) );
  INV_X1 U6796 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6897) );
  INV_X1 U6797 ( .A(SI_17_), .ZN(n10106) );
  NAND2_X1 U6798 ( .A1(n5353), .A2(n10106), .ZN(n5370) );
  INV_X1 U6799 ( .A(n5353), .ZN(n5354) );
  NAND2_X1 U6800 ( .A1(n5354), .A2(SI_17_), .ZN(n5355) );
  NAND2_X1 U6801 ( .A1(n5370), .A2(n5355), .ZN(n5371) );
  XNOR2_X1 U6802 ( .A(n5372), .B(n5371), .ZN(n6896) );
  NAND2_X1 U6803 ( .A1(n6896), .A2(n7872), .ZN(n5361) );
  OAI21_X1 U6804 ( .B1(n5357), .B2(P2_IR_REG_16__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5358) );
  MUX2_X1 U6805 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5358), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5359) );
  AND2_X1 U6806 ( .A1(n5356), .A2(n5359), .ZN(n8231) );
  AOI22_X1 U6807 ( .A1(n5398), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5397), .B2(
        n8231), .ZN(n5360) );
  NAND2_X1 U6808 ( .A1(n5600), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5367) );
  NAND2_X1 U6809 ( .A1(n7070), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5366) );
  NAND2_X1 U6810 ( .A1(n5362), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6811 ( .A1(n5377), .A2(n5363), .ZN(n8424) );
  NAND2_X1 U6812 ( .A1(n5547), .A2(n8424), .ZN(n5365) );
  NAND2_X1 U6813 ( .A1(n7071), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6814 ( .A1(n8562), .A2(n8433), .ZN(n8008) );
  INV_X1 U6815 ( .A(n8416), .ZN(n5368) );
  INV_X1 U6816 ( .A(n8433), .ZN(n8097) );
  NAND2_X1 U6817 ( .A1(n8562), .A2(n8097), .ZN(n5369) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7021) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6992) );
  MUX2_X1 U6820 ( .A(n7021), .B(n6992), .S(n7868), .Z(n5385) );
  XNOR2_X1 U6821 ( .A(n5385), .B(SI_18_), .ZN(n5384) );
  XNOR2_X1 U6822 ( .A(n5389), .B(n5384), .ZN(n6991) );
  NAND2_X1 U6823 ( .A1(n6991), .A2(n7872), .ZN(n5374) );
  NAND2_X1 U6824 ( .A1(n5356), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6825 ( .A(n5394), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8251) );
  AOI22_X1 U6826 ( .A1(n5398), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5397), .B2(
        n8251), .ZN(n5373) );
  NAND2_X1 U6827 ( .A1(n7071), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U6828 ( .A1(n5600), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5381) );
  INV_X1 U6829 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5375) );
  NAND2_X1 U6830 ( .A1(n5377), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5378) );
  NAND2_X1 U6831 ( .A1(n5401), .A2(n5378), .ZN(n8408) );
  NAND2_X1 U6832 ( .A1(n5547), .A2(n8408), .ZN(n5380) );
  NAND2_X1 U6833 ( .A1(n7070), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5379) );
  INV_X1 U6834 ( .A(n8419), .ZN(n8389) );
  OR2_X1 U6835 ( .A1(n8490), .A2(n8389), .ZN(n5383) );
  INV_X1 U6836 ( .A(n5384), .ZN(n5388) );
  INV_X1 U6837 ( .A(n5385), .ZN(n5386) );
  NAND2_X1 U6838 ( .A1(n5386), .A2(SI_18_), .ZN(n5387) );
  INV_X1 U6839 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7173) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7175) );
  MUX2_X1 U6841 ( .A(n7173), .B(n7175), .S(n7868), .Z(n5391) );
  INV_X1 U6842 ( .A(SI_19_), .ZN(n5390) );
  NAND2_X1 U6843 ( .A1(n5391), .A2(n5390), .ZN(n5414) );
  INV_X1 U6844 ( .A(n5391), .ZN(n5392) );
  NAND2_X1 U6845 ( .A1(n5392), .A2(SI_19_), .ZN(n5393) );
  NAND2_X1 U6846 ( .A1(n5414), .A2(n5393), .ZN(n5411) );
  XNOR2_X1 U6847 ( .A(n5410), .B(n5411), .ZN(n7172) );
  NAND2_X1 U6848 ( .A1(n7172), .A2(n7872), .ZN(n5400) );
  NAND2_X1 U6849 ( .A1(n5394), .A2(n10267), .ZN(n5395) );
  XNOR2_X2 U6850 ( .A(n5396), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8262) );
  AOI22_X1 U6851 ( .A1(n5398), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8262), .B2(
        n5397), .ZN(n5399) );
  NAND2_X1 U6852 ( .A1(n7071), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6853 ( .A1(n5600), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6854 ( .A1(n5401), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5402) );
  NAND2_X1 U6855 ( .A1(n5423), .A2(n5402), .ZN(n8396) );
  NAND2_X1 U6856 ( .A1(n5073), .A2(n8396), .ZN(n5404) );
  NAND2_X1 U6857 ( .A1(n7070), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6858 ( .A1(n8485), .A2(n8403), .ZN(n8014) );
  NAND2_X1 U6859 ( .A1(n8385), .A2(n7902), .ZN(n5408) );
  INV_X1 U6860 ( .A(n8403), .ZN(n8379) );
  NAND2_X1 U6861 ( .A1(n8485), .A2(n8379), .ZN(n5407) );
  MUX2_X1 U6862 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7868), .Z(n5428) );
  INV_X1 U6863 ( .A(SI_20_), .ZN(n10266) );
  XNOR2_X1 U6864 ( .A(n5428), .B(n10266), .ZN(n5416) );
  XNOR2_X1 U6865 ( .A(n5430), .B(n5416), .ZN(n7258) );
  NAND2_X1 U6866 ( .A1(n7258), .A2(n7872), .ZN(n5418) );
  INV_X1 U6867 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7259) );
  OR2_X1 U6868 ( .A1(n7873), .A2(n7259), .ZN(n5417) );
  NAND2_X1 U6869 ( .A1(n5600), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5420) );
  NAND2_X1 U6870 ( .A1(n7071), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5419) );
  AND2_X1 U6871 ( .A1(n5420), .A2(n5419), .ZN(n5427) );
  INV_X1 U6872 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U6873 ( .A1(n5423), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5424) );
  NAND2_X1 U6874 ( .A1(n5434), .A2(n5424), .ZN(n8382) );
  NAND2_X1 U6875 ( .A1(n8382), .A2(n5547), .ZN(n5426) );
  NAND2_X1 U6876 ( .A1(n7070), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U6877 ( .A1(n8553), .A2(n7749), .ZN(n8018) );
  NAND2_X1 U6878 ( .A1(n4998), .A2(n8018), .ZN(n8376) );
  OR2_X1 U6879 ( .A1(n8553), .A2(n8387), .ZN(n8364) );
  INV_X1 U6880 ( .A(n5428), .ZN(n5429) );
  INV_X1 U6881 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10262) );
  INV_X1 U6882 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7338) );
  MUX2_X1 U6883 ( .A(n10262), .B(n7338), .S(n7868), .Z(n5439) );
  XNOR2_X1 U6884 ( .A(n5439), .B(SI_21_), .ZN(n5431) );
  XNOR2_X1 U6885 ( .A(n5441), .B(n5431), .ZN(n7337) );
  NAND2_X1 U6886 ( .A1(n7337), .A2(n7872), .ZN(n5433) );
  OR2_X1 U6887 ( .A1(n7873), .A2(n10262), .ZN(n5432) );
  NAND2_X1 U6888 ( .A1(n5434), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U6889 ( .A1(n5449), .A2(n5435), .ZN(n8370) );
  NAND2_X1 U6890 ( .A1(n8370), .A2(n5547), .ZN(n5438) );
  AOI22_X1 U6891 ( .A1(n7071), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n5548), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n5437) );
  NAND2_X1 U6892 ( .A1(n7070), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5436) );
  OR2_X1 U6893 ( .A1(n8548), .A2(n8378), .ZN(n8353) );
  NAND2_X1 U6894 ( .A1(n8352), .A2(n8353), .ZN(n5454) );
  INV_X1 U6895 ( .A(n5439), .ZN(n5440) );
  INV_X1 U6896 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7436) );
  INV_X1 U6897 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n10282) );
  MUX2_X1 U6898 ( .A(n7436), .B(n10282), .S(n7868), .Z(n5443) );
  INV_X1 U6899 ( .A(SI_22_), .ZN(n5442) );
  NAND2_X1 U6900 ( .A1(n5443), .A2(n5442), .ZN(n5456) );
  INV_X1 U6901 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U6902 ( .A1(n5444), .A2(SI_22_), .ZN(n5445) );
  NAND2_X1 U6903 ( .A1(n5456), .A2(n5445), .ZN(n5457) );
  XNOR2_X1 U6904 ( .A(n5458), .B(n5457), .ZN(n7433) );
  NAND2_X1 U6905 ( .A1(n7433), .A2(n7872), .ZN(n5447) );
  OR2_X1 U6906 ( .A1(n7873), .A2(n7436), .ZN(n5446) );
  INV_X1 U6907 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8358) );
  INV_X1 U6908 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U6909 ( .A1(n5449), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U6910 ( .A1(n5468), .A2(n5450), .ZN(n8359) );
  NAND2_X1 U6911 ( .A1(n8359), .A2(n5547), .ZN(n5452) );
  AOI22_X1 U6912 ( .A1(n7071), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n5600), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n5451) );
  OAI211_X1 U6913 ( .C1(n5603), .C2(n8358), .A(n5452), .B(n5451), .ZN(n8367)
         );
  INV_X1 U6914 ( .A(n8026), .ZN(n5453) );
  INV_X1 U6915 ( .A(n8367), .ZN(n8342) );
  NAND2_X1 U6916 ( .A1(n8542), .A2(n8342), .ZN(n8024) );
  NAND2_X1 U6917 ( .A1(n7812), .A2(n8342), .ZN(n5455) );
  INV_X1 U6918 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7511) );
  INV_X1 U6919 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7506) );
  MUX2_X1 U6920 ( .A(n7511), .B(n7506), .S(n7868), .Z(n5460) );
  INV_X1 U6921 ( .A(SI_23_), .ZN(n5459) );
  NAND2_X1 U6922 ( .A1(n5460), .A2(n5459), .ZN(n5478) );
  INV_X1 U6923 ( .A(n5460), .ZN(n5461) );
  NAND2_X1 U6924 ( .A1(n5461), .A2(SI_23_), .ZN(n5462) );
  OR2_X1 U6925 ( .A1(n5464), .A2(n5463), .ZN(n5465) );
  NAND2_X1 U6926 ( .A1(n5479), .A2(n5465), .ZN(n7507) );
  NAND2_X1 U6927 ( .A1(n7507), .A2(n7872), .ZN(n5467) );
  OR2_X1 U6928 ( .A1(n7873), .A2(n7511), .ZN(n5466) );
  NAND2_X1 U6929 ( .A1(n5468), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6930 ( .A1(n5486), .A2(n5469), .ZN(n8344) );
  NAND2_X1 U6931 ( .A1(n8344), .A2(n5547), .ZN(n5474) );
  INV_X1 U6932 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U6933 ( .A1(n7071), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6934 ( .A1(n7070), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U6935 ( .C1(n7074), .C2(n10283), .A(n5471), .B(n5470), .ZN(n5472)
         );
  INV_X1 U6936 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U6937 ( .A1(n8474), .A2(n8356), .ZN(n5475) );
  NAND2_X1 U6938 ( .A1(n8340), .A2(n5475), .ZN(n5477) );
  NAND2_X1 U6939 ( .A1(n5477), .A2(n5476), .ZN(n8327) );
  INV_X1 U6940 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n10061) );
  INV_X1 U6941 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7593) );
  MUX2_X1 U6942 ( .A(n10061), .B(n7593), .S(n7868), .Z(n5481) );
  INV_X1 U6943 ( .A(SI_24_), .ZN(n5480) );
  NAND2_X1 U6944 ( .A1(n5481), .A2(n5480), .ZN(n5498) );
  INV_X1 U6945 ( .A(n5481), .ZN(n5482) );
  NAND2_X1 U6946 ( .A1(n5482), .A2(SI_24_), .ZN(n5483) );
  NAND2_X1 U6947 ( .A1(n7590), .A2(n7872), .ZN(n5485) );
  OR2_X1 U6948 ( .A1(n7873), .A2(n10061), .ZN(n5484) );
  NAND2_X1 U6949 ( .A1(n5486), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6950 ( .A1(n5507), .A2(n5487), .ZN(n8334) );
  NAND2_X1 U6951 ( .A1(n8334), .A2(n5547), .ZN(n5493) );
  INV_X1 U6952 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n10190) );
  NAND2_X1 U6953 ( .A1(n5600), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U6954 ( .A1(n7070), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5488) );
  OAI211_X1 U6955 ( .C1(n10190), .C2(n5490), .A(n5489), .B(n5488), .ZN(n5491)
         );
  INV_X1 U6956 ( .A(n5491), .ZN(n5492) );
  NOR2_X1 U6957 ( .A1(n8532), .A2(n8096), .ZN(n5494) );
  NAND2_X1 U6958 ( .A1(n8532), .A2(n8096), .ZN(n5495) );
  INV_X1 U6959 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7598) );
  INV_X1 U6960 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7600) );
  MUX2_X1 U6961 ( .A(n7598), .B(n7600), .S(n7868), .Z(n5500) );
  INV_X1 U6962 ( .A(SI_25_), .ZN(n5499) );
  NAND2_X1 U6963 ( .A1(n5500), .A2(n5499), .ZN(n5515) );
  INV_X1 U6964 ( .A(n5500), .ZN(n5501) );
  NAND2_X1 U6965 ( .A1(n5501), .A2(SI_25_), .ZN(n5502) );
  AND2_X1 U6966 ( .A1(n5515), .A2(n5502), .ZN(n5513) );
  NAND2_X1 U6967 ( .A1(n7596), .A2(n7872), .ZN(n5504) );
  OR2_X1 U6968 ( .A1(n7873), .A2(n7598), .ZN(n5503) );
  INV_X1 U6969 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U6970 ( .A1(n5507), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U6971 ( .A1(n5524), .A2(n5508), .ZN(n8317) );
  INV_X1 U6972 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8468) );
  NAND2_X1 U6973 ( .A1(n7070), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U6974 ( .A1(n7071), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5509) );
  OAI211_X1 U6975 ( .C1(n7074), .C2(n8468), .A(n5510), .B(n5509), .ZN(n5511)
         );
  AOI21_X1 U6976 ( .B1(n8317), .B2(n5547), .A(n5511), .ZN(n7842) );
  NAND2_X1 U6977 ( .A1(n8467), .A2(n7842), .ZN(n8042) );
  NAND2_X1 U6978 ( .A1(n4820), .A2(n8042), .ZN(n7905) );
  INV_X1 U6979 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7641) );
  INV_X1 U6980 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9573) );
  MUX2_X1 U6981 ( .A(n7641), .B(n9573), .S(n7868), .Z(n5518) );
  INV_X1 U6982 ( .A(SI_26_), .ZN(n5517) );
  NAND2_X1 U6983 ( .A1(n5518), .A2(n5517), .ZN(n5534) );
  INV_X1 U6984 ( .A(n5518), .ZN(n5519) );
  NAND2_X1 U6985 ( .A1(n5519), .A2(SI_26_), .ZN(n5520) );
  AND2_X1 U6986 ( .A1(n5534), .A2(n5520), .ZN(n5532) );
  OR2_X1 U6987 ( .A1(n7873), .A2(n7641), .ZN(n5521) );
  INV_X1 U6988 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10055) );
  NAND2_X1 U6989 ( .A1(n5524), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5525) );
  NAND2_X1 U6990 ( .A1(n5545), .A2(n5525), .ZN(n8307) );
  NAND2_X1 U6991 ( .A1(n8307), .A2(n5547), .ZN(n5530) );
  INV_X1 U6992 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U6993 ( .A1(n7071), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5527) );
  NAND2_X1 U6994 ( .A1(n5600), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5526) );
  OAI211_X1 U6995 ( .C1(n8306), .C2(n5603), .A(n5527), .B(n5526), .ZN(n5528)
         );
  INV_X1 U6996 ( .A(n5528), .ZN(n5529) );
  NAND2_X1 U6997 ( .A1(n8523), .A2(n8095), .ZN(n5531) );
  INV_X1 U6998 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5542) );
  INV_X1 U6999 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10324) );
  MUX2_X1 U7000 ( .A(n5542), .B(n10324), .S(n7868), .Z(n5536) );
  INV_X1 U7001 ( .A(SI_27_), .ZN(n5535) );
  NAND2_X1 U7002 ( .A1(n5536), .A2(n5535), .ZN(n5557) );
  INV_X1 U7003 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7004 ( .A1(n5537), .A2(SI_27_), .ZN(n5538) );
  AND2_X1 U7005 ( .A1(n5557), .A2(n5538), .ZN(n5539) );
  NAND2_X1 U7006 ( .A1(n8584), .A2(n7872), .ZN(n5544) );
  OR2_X1 U7007 ( .A1(n7873), .A2(n5542), .ZN(n5543) );
  NAND2_X1 U7008 ( .A1(n5545), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n5546) );
  NAND2_X1 U7009 ( .A1(n5563), .A2(n5546), .ZN(n8298) );
  NAND2_X1 U7010 ( .A1(n8298), .A2(n5547), .ZN(n5554) );
  INV_X1 U7011 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7012 ( .A1(n5548), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7013 ( .A1(n7071), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5549) );
  OAI211_X1 U7014 ( .C1(n5603), .C2(n5551), .A(n5550), .B(n5549), .ZN(n5552)
         );
  INV_X1 U7015 ( .A(n5552), .ZN(n5553) );
  INV_X1 U7016 ( .A(n8051), .ZN(n5555) );
  MUX2_X1 U7017 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n7868), .Z(n5572) );
  INV_X1 U7018 ( .A(SI_28_), .ZN(n5573) );
  XNOR2_X1 U7019 ( .A(n5572), .B(n5573), .ZN(n5571) );
  NAND2_X1 U7020 ( .A1(n8621), .A2(n7872), .ZN(n5560) );
  INV_X1 U7021 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n10299) );
  OR2_X1 U7022 ( .A1(n7873), .A2(n10299), .ZN(n5559) );
  INV_X1 U7023 ( .A(n5563), .ZN(n5562) );
  INV_X1 U7024 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U7025 ( .A1(n5562), .A2(n5561), .ZN(n5663) );
  NAND2_X1 U7026 ( .A1(n5563), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5564) );
  NAND2_X1 U7027 ( .A1(n5663), .A2(n5564), .ZN(n8287) );
  NAND2_X1 U7028 ( .A1(n8287), .A2(n5073), .ZN(n5569) );
  INV_X1 U7029 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n10340) );
  NAND2_X1 U7030 ( .A1(n7071), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7031 ( .A1(n5600), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5565) );
  OAI211_X1 U7032 ( .C1(n10340), .C2(n5603), .A(n5566), .B(n5565), .ZN(n5567)
         );
  INV_X1 U7033 ( .A(n5567), .ZN(n5568) );
  INV_X1 U7034 ( .A(n5571), .ZN(n5576) );
  INV_X1 U7035 ( .A(n5572), .ZN(n5574) );
  NAND2_X1 U7036 ( .A1(n5574), .A2(n5573), .ZN(n5575) );
  MUX2_X1 U7037 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7868), .Z(n7660) );
  INV_X1 U7038 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7656) );
  NOR2_X1 U7039 ( .A1(n7873), .A2(n7656), .ZN(n5579) );
  INV_X1 U7040 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7041 ( .A1(n7071), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5582) );
  NAND2_X1 U7042 ( .A1(n5600), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5581) );
  OAI211_X1 U7043 ( .C1(n5665), .C2(n5603), .A(n5582), .B(n5581), .ZN(n5583)
         );
  INV_X1 U7044 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7045 ( .A1(n7077), .A2(n5584), .ZN(n8282) );
  INV_X1 U7046 ( .A(n7876), .ZN(n8057) );
  INV_X1 U7047 ( .A(n5698), .ZN(n8054) );
  INV_X1 U7048 ( .A(n8282), .ZN(n5585) );
  NAND2_X1 U7049 ( .A1(n8054), .A2(n5585), .ZN(n7878) );
  XNOR2_X1 U7050 ( .A(n5586), .B(n5656), .ZN(n5609) );
  INV_X1 U7051 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5587) );
  NAND2_X1 U7052 ( .A1(n10267), .A2(n5587), .ZN(n5588) );
  NOR2_X2 U7053 ( .A1(n5356), .A2(n5588), .ZN(n5594) );
  NAND2_X1 U7054 ( .A1(n5594), .A2(n5589), .ZN(n5591) );
  NAND2_X1 U7055 ( .A1(n5620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U7056 ( .A(n5590), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8091) );
  NAND2_X1 U7057 ( .A1(n8091), .A2(n8262), .ZN(n5679) );
  NAND2_X1 U7058 ( .A1(n5591), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5592) );
  MUX2_X1 U7059 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5592), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5593) );
  NAND2_X1 U7060 ( .A1(n5593), .A2(n5620), .ZN(n7916) );
  INV_X1 U7061 ( .A(n5594), .ZN(n5595) );
  XNOR2_X2 U7062 ( .A(n5596), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8085) );
  NAND2_X1 U7063 ( .A1(n6598), .A2(n8085), .ZN(n5597) );
  OR2_X1 U7064 ( .A1(n8087), .A2(n8253), .ZN(n5598) );
  NAND2_X1 U7065 ( .A1(n4497), .A2(n5598), .ZN(n6605) );
  NAND2_X1 U7066 ( .A1(n6605), .A2(n8066), .ZN(n9642) );
  AND2_X1 U7067 ( .A1(n4497), .A2(P2_B_REG_SCAN_IN), .ZN(n5599) );
  OR2_X1 U7068 ( .A1(n9642), .A2(n5599), .ZN(n8271) );
  INV_X1 U7069 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U7070 ( .A1(n7071), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U7071 ( .A1(n5600), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5601) );
  OAI211_X1 U7072 ( .C1(n5604), .C2(n5603), .A(n5602), .B(n5601), .ZN(n5605)
         );
  INV_X1 U7073 ( .A(n5605), .ZN(n5606) );
  XNOR2_X1 U7074 ( .A(n7591), .B(P2_B_REG_SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7075 ( .A1(n5611), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5612) );
  XNOR2_X1 U7076 ( .A(n5612), .B(P2_IR_REG_25__SCAN_IN), .ZN(n7597) );
  INV_X1 U7077 ( .A(n5614), .ZN(n5615) );
  NAND2_X1 U7078 ( .A1(n5615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5616) );
  XNOR2_X1 U7079 ( .A(n5616), .B(P2_IR_REG_26__SCAN_IN), .ZN(n7640) );
  OR2_X1 U7080 ( .A1(n5618), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5617) );
  OR2_X1 U7081 ( .A1(n7640), .A2(n7597), .ZN(n6410) );
  OR2_X1 U7082 ( .A1(n7640), .A2(n7591), .ZN(n6408) );
  NAND2_X1 U7083 ( .A1(n5677), .A2(n6596), .ZN(n5681) );
  AND2_X1 U7084 ( .A1(n7597), .A2(n7591), .ZN(n5619) );
  OAI21_X1 U7085 ( .B1(n5620), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5622) );
  INV_X1 U7086 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5621) );
  XNOR2_X1 U7087 ( .A(n5622), .B(n5621), .ZN(n7508) );
  NAND2_X1 U7088 ( .A1(n7508), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6322) );
  INV_X2 U7089 ( .A(n8262), .ZN(n8247) );
  INV_X1 U7090 ( .A(n6597), .ZN(n5658) );
  AND2_X1 U7091 ( .A1(n8066), .A2(n5658), .ZN(n6524) );
  NOR2_X1 U7092 ( .A1(n6530), .A2(n6524), .ZN(n5633) );
  NOR4_X1 U7093 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n10305) );
  NOR2_X1 U7094 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .ZN(
        n5625) );
  NOR4_X1 U7095 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5624) );
  NOR4_X1 U7096 ( .A1(P2_D_REG_30__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n5623) );
  NAND4_X1 U7097 ( .A1(n10305), .A2(n5625), .A3(n5624), .A4(n5623), .ZN(n5631)
         );
  NOR4_X1 U7098 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n5629) );
  NOR4_X1 U7099 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n5628) );
  NOR4_X1 U7100 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n5627) );
  NOR4_X1 U7101 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_11__SCAN_IN), .ZN(n5626) );
  NAND4_X1 U7102 ( .A1(n5629), .A2(n5628), .A3(n5627), .A4(n5626), .ZN(n5630)
         );
  NOR2_X1 U7103 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  OR2_X1 U7104 ( .A1(n5618), .A2(n5632), .ZN(n5676) );
  AND2_X1 U7105 ( .A1(n8091), .A2(n8247), .ZN(n5657) );
  NAND2_X1 U7106 ( .A1(n5657), .A2(n8085), .ZN(n5634) );
  INV_X1 U7107 ( .A(n5688), .ZN(n5692) );
  INV_X1 U7108 ( .A(n6596), .ZN(n5689) );
  NAND2_X1 U7109 ( .A1(n5692), .A2(n5689), .ZN(n5636) );
  INV_X1 U7110 ( .A(n5677), .ZN(n5691) );
  NAND2_X1 U7111 ( .A1(n5691), .A2(n5688), .ZN(n5635) );
  AND2_X1 U7112 ( .A1(n5636), .A2(n5635), .ZN(n5637) );
  NAND2_X1 U7113 ( .A1(n5696), .A2(n5637), .ZN(n5662) );
  OR2_X1 U7114 ( .A1(n8247), .A2(n8085), .ZN(n5661) );
  NOR2_X1 U7115 ( .A1(n8091), .A2(n5661), .ZN(n5672) );
  AND2_X1 U7116 ( .A1(n5672), .A2(n7916), .ZN(n5690) );
  NAND2_X1 U7117 ( .A1(n6407), .A2(n5690), .ZN(n9632) );
  NAND2_X1 U7118 ( .A1(n5675), .A2(n9645), .ZN(n5671) );
  NAND2_X1 U7119 ( .A1(n6724), .A2(n6614), .ZN(n7930) );
  NAND2_X1 U7120 ( .A1(n6772), .A2(n7930), .ZN(n6805) );
  NAND2_X1 U7121 ( .A1(n6949), .A2(n9937), .ZN(n7938) );
  NAND2_X1 U7122 ( .A1(n5640), .A2(n6746), .ZN(n7944) );
  AND2_X1 U7123 ( .A1(n7938), .A2(n7944), .ZN(n6804) );
  NAND2_X1 U7124 ( .A1(n6805), .A2(n6804), .ZN(n5641) );
  NAND2_X1 U7125 ( .A1(n5641), .A2(n7938), .ZN(n6942) );
  NAND2_X1 U7126 ( .A1(n8110), .A2(n9944), .ZN(n7939) );
  INV_X1 U7127 ( .A(n8110), .ZN(n6792) );
  NAND2_X1 U7128 ( .A1(n6792), .A2(n6954), .ZN(n7946) );
  NOR2_X1 U7129 ( .A1(n8109), .A2(n9949), .ZN(n7945) );
  NAND2_X1 U7130 ( .A1(n8108), .A2(n9955), .ZN(n7941) );
  NAND2_X1 U7131 ( .A1(n8109), .A2(n9949), .ZN(n7014) );
  AND2_X1 U7132 ( .A1(n7941), .A2(n7014), .ZN(n7951) );
  NAND2_X1 U7133 ( .A1(n7013), .A2(n7951), .ZN(n5643) );
  NAND2_X1 U7134 ( .A1(n7006), .A2(n7831), .ZN(n7949) );
  NAND2_X1 U7135 ( .A1(n5643), .A2(n7949), .ZN(n7056) );
  INV_X1 U7136 ( .A(n7056), .ZN(n5645) );
  NAND2_X1 U7137 ( .A1(n5645), .A2(n5644), .ZN(n7055) );
  OR2_X1 U7138 ( .A1(n7361), .A2(n7325), .ZN(n7964) );
  NAND2_X1 U7139 ( .A1(n7325), .A2(n7361), .ZN(n7960) );
  NAND2_X1 U7140 ( .A1(n7964), .A2(n7960), .ZN(n7891) );
  NAND2_X1 U7141 ( .A1(n7314), .A2(n7964), .ZN(n7357) );
  INV_X1 U7142 ( .A(n9975), .ZN(n7368) );
  NAND2_X1 U7143 ( .A1(n7368), .A2(n7381), .ZN(n7974) );
  OR2_X1 U7144 ( .A1(n7409), .A2(n7564), .ZN(n7977) );
  XNOR2_X1 U7145 ( .A(n9991), .B(n8102), .ZN(n7979) );
  OR2_X1 U7146 ( .A1(n9991), .A2(n9639), .ZN(n7982) );
  NAND2_X1 U7147 ( .A1(n7568), .A2(n7982), .ZN(n9628) );
  NAND2_X1 U7148 ( .A1(n9631), .A2(n7586), .ZN(n7989) );
  NAND2_X1 U7149 ( .A1(n9628), .A2(n7989), .ZN(n5647) );
  OR2_X1 U7150 ( .A1(n9631), .A2(n7586), .ZN(n7988) );
  NAND2_X1 U7151 ( .A1(n5647), .A2(n7988), .ZN(n7620) );
  NAND2_X1 U7152 ( .A1(n7627), .A2(n9641), .ZN(n7994) );
  NAND2_X1 U7153 ( .A1(n7620), .A2(n7991), .ZN(n5648) );
  NAND2_X1 U7154 ( .A1(n5648), .A2(n7997), .ZN(n7649) );
  NAND2_X1 U7155 ( .A1(n7649), .A2(n7998), .ZN(n5649) );
  NAND2_X1 U7156 ( .A1(n5649), .A2(n7995), .ZN(n8427) );
  NAND2_X1 U7157 ( .A1(n8427), .A2(n8006), .ZN(n5650) );
  NAND2_X1 U7158 ( .A1(n5650), .A2(n8003), .ZN(n8413) );
  INV_X1 U7159 ( .A(n8413), .ZN(n5651) );
  NAND2_X1 U7160 ( .A1(n8490), .A2(n8419), .ZN(n8013) );
  NAND2_X1 U7161 ( .A1(n8009), .A2(n8013), .ZN(n8406) );
  NAND2_X1 U7162 ( .A1(n8395), .A2(n8016), .ZN(n8373) );
  NAND2_X1 U7163 ( .A1(n8532), .A2(n8343), .ZN(n8030) );
  NAND2_X1 U7164 ( .A1(n8474), .A2(n7808), .ZN(n8323) );
  NAND2_X1 U7165 ( .A1(n8030), .A2(n8323), .ZN(n8033) );
  NOR2_X1 U7166 ( .A1(n8060), .A2(n8295), .ZN(n5655) );
  XNOR2_X1 U7167 ( .A(n7877), .B(n5656), .ZN(n5673) );
  INV_X1 U7168 ( .A(n5673), .ZN(n5668) );
  NAND2_X1 U7169 ( .A1(n8066), .A2(n6597), .ZN(n6541) );
  INV_X1 U7170 ( .A(n8091), .ZN(n7914) );
  NAND2_X1 U7171 ( .A1(n7914), .A2(n7916), .ZN(n9980) );
  AND2_X1 U7172 ( .A1(n6541), .A2(n9980), .ZN(n6561) );
  INV_X1 U7173 ( .A(n5657), .ZN(n5659) );
  NAND2_X1 U7174 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  NAND2_X1 U7175 ( .A1(n6561), .A2(n5660), .ZN(n7365) );
  INV_X1 U7176 ( .A(n5661), .ZN(n9634) );
  NAND2_X1 U7177 ( .A1(n9634), .A2(n6598), .ZN(n6775) );
  AND2_X1 U7178 ( .A1(n7365), .A2(n6775), .ZN(n9630) );
  OR2_X1 U7179 ( .A1(n9980), .A2(n9634), .ZN(n8331) );
  OR2_X1 U7180 ( .A1(n5662), .A2(n8331), .ZN(n8277) );
  INV_X1 U7181 ( .A(n5663), .ZN(n5664) );
  INV_X1 U7182 ( .A(n9632), .ZN(n8443) );
  NAND2_X1 U7183 ( .A1(n5664), .A2(n8443), .ZN(n8273) );
  OAI21_X1 U7184 ( .B1(n9645), .B2(n5665), .A(n8273), .ZN(n5666) );
  AOI21_X1 U7185 ( .B1(n8054), .B2(n8444), .A(n5666), .ZN(n5667) );
  NAND2_X1 U7186 ( .A1(n5671), .A2(n5670), .ZN(P2_U3204) );
  INV_X1 U7187 ( .A(n5672), .ZN(n9976) );
  NAND2_X1 U7188 ( .A1(n7365), .A2(n9976), .ZN(n9968) );
  INV_X1 U7189 ( .A(n5676), .ZN(n5680) );
  NOR2_X1 U7190 ( .A1(n5677), .A2(n5680), .ZN(n5678) );
  AND2_X1 U7191 ( .A1(n5678), .A2(n5689), .ZN(n6529) );
  AND2_X1 U7192 ( .A1(n6529), .A2(n6407), .ZN(n6543) );
  NAND2_X1 U7193 ( .A1(n7916), .A2(n8085), .ZN(n6594) );
  OR2_X1 U7194 ( .A1(n5679), .A2(n6594), .ZN(n6534) );
  NAND3_X1 U7195 ( .A1(n8070), .A2(n6534), .A3(n9980), .ZN(n6536) );
  NAND2_X1 U7196 ( .A1(n6536), .A2(n8331), .ZN(n6519) );
  NAND2_X1 U7197 ( .A1(n6543), .A2(n6519), .ZN(n5684) );
  NOR2_X1 U7198 ( .A1(n5681), .A2(n5680), .ZN(n6521) );
  NAND2_X1 U7199 ( .A1(n6521), .A2(n6407), .ZN(n6539) );
  AND2_X1 U7200 ( .A1(n6534), .A2(n6541), .ZN(n5682) );
  OR2_X1 U7201 ( .A1(n6539), .A2(n5682), .ZN(n5683) );
  INV_X2 U7202 ( .A(n9994), .ZN(n9993) );
  OR2_X1 U7203 ( .A1(n9994), .A2(n9980), .ZN(n8516) );
  NAND2_X1 U7204 ( .A1(n8054), .A2(n8568), .ZN(n5686) );
  INV_X1 U7205 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U7206 ( .B1(n5701), .B2(n9994), .A(n5687), .ZN(P2_U3456) );
  OAI21_X1 U7207 ( .B1(n5690), .B2(n5689), .A(n5688), .ZN(n5694) );
  NAND2_X1 U7208 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  AND2_X1 U7209 ( .A1(n5694), .A2(n5693), .ZN(n5695) );
  AND2_X2 U7210 ( .A1(n5696), .A2(n5695), .ZN(n10012) );
  INV_X1 U7211 ( .A(n9980), .ZN(n9992) );
  NAND2_X1 U7212 ( .A1(n10012), .A2(n9992), .ZN(n8460) );
  INV_X1 U7213 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5697) );
  OAI21_X1 U7214 ( .B1(n5701), .B2(n10010), .A(n5700), .ZN(P2_U3488) );
  NOR2_X1 U7215 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5705) );
  NAND4_X1 U7216 ( .A1(n5705), .A2(n5704), .A3(n5703), .A4(n5702), .ZN(n5707)
         );
  NAND4_X1 U7217 ( .A1(n5768), .A2(n5763), .A3(n5775), .A4(n5772), .ZN(n5706)
         );
  NOR2_X2 U7218 ( .A1(n5707), .A2(n5706), .ZN(n5726) );
  NOR2_X1 U7219 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5712) );
  NOR2_X1 U7220 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5711) );
  NOR2_X1 U7221 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5710) );
  INV_X1 U7222 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5714) );
  XNOR2_X2 U7223 ( .A(n5715), .B(n5740), .ZN(n5801) );
  MUX2_X1 U7224 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5717), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5718) );
  NAND2_X1 U7225 ( .A1(n6587), .A2(n8781), .ZN(n5725) );
  NOR2_X1 U7226 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5721) );
  INV_X1 U7227 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7228 ( .A1(n5768), .A2(n5984), .ZN(n5722) );
  OAI21_X1 U7229 ( .B1(n5968), .B2(n5722), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6005) );
  NAND2_X1 U7230 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), 
        .ZN(n10309) );
  NAND2_X1 U7231 ( .A1(n6005), .A2(n10309), .ZN(n6031) );
  INV_X1 U7232 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5723) );
  XNOR2_X1 U7233 ( .A(n6031), .B(n5723), .ZN(n9781) );
  AOI22_X1 U7234 ( .A1(n6121), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6120), .B2(
        n9781), .ZN(n5724) );
  NAND2_X1 U7235 ( .A1(n5758), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5728) );
  INV_X1 U7236 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7237 ( .A1(n5729), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5730) );
  MUX2_X1 U7238 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5730), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5731) );
  NAND2_X1 U7239 ( .A1(n5732), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5733) );
  XNOR2_X1 U7240 ( .A(n5733), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7241 ( .A1(n5735), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5736) );
  MUX2_X1 U7242 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5736), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5738) );
  NAND2_X1 U7243 ( .A1(n5738), .A2(n5737), .ZN(n7595) );
  NOR2_X1 U7244 ( .A1(n7602), .A2(n7595), .ZN(n5739) );
  NAND2_X1 U7245 ( .A1(n6289), .A2(n5739), .ZN(n6320) );
  AND2_X2 U7246 ( .A1(n5781), .A2(n6320), .ZN(n8631) );
  NAND2_X1 U7247 ( .A1(n9683), .A2(n6261), .ZN(n5757) );
  OR2_X2 U7248 ( .A1(n9560), .A2(n9562), .ZN(n5742) );
  INV_X1 U7249 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5741) );
  XNOR2_X2 U7250 ( .A(n5742), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U7251 ( .A1(n5743), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7252 ( .A1(n8755), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7253 ( .A1(n8756), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7254 ( .A1(n8757), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5751) );
  NAND2_X1 U7255 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n5747) );
  INV_X1 U7256 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9590) );
  INV_X1 U7257 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7258 ( .A1(n6011), .A2(n5748), .ZN(n5749) );
  NAND2_X1 U7259 ( .A1(n6036), .A2(n5749), .ZN(n9685) );
  OR2_X1 U7260 ( .A1(n8635), .A2(n9685), .ZN(n5750) );
  NAND4_X1 U7261 ( .A1(n5753), .A2(n5752), .A3(n5751), .A4(n5750), .ZN(n9024)
         );
  AND2_X1 U7262 ( .A1(n5754), .A2(n6320), .ZN(n5755) );
  INV_X2 U7263 ( .A(n5755), .ZN(n6218) );
  NAND2_X1 U7264 ( .A1(n9024), .A2(n6194), .ZN(n5756) );
  NAND2_X1 U7265 ( .A1(n5757), .A2(n5756), .ZN(n5782) );
  OAI21_X1 U7266 ( .B1(n5758), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5760) );
  INV_X1 U7267 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7268 ( .A1(n5760), .A2(n5759), .ZN(n6292) );
  OR2_X1 U7269 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  NAND2_X1 U7270 ( .A1(n6292), .A2(n5761), .ZN(n7434) );
  INV_X1 U7271 ( .A(n7434), .ZN(n9009) );
  NOR2_X1 U7272 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5766) );
  NOR2_X1 U7273 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5765) );
  NOR2_X1 U7274 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5764) );
  NAND4_X1 U7275 ( .A1(n5766), .A2(n5765), .A3(n5764), .A4(n5763), .ZN(n5770)
         );
  INV_X1 U7276 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10216) );
  INV_X1 U7277 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5767) );
  INV_X1 U7278 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6032) );
  NAND4_X1 U7279 ( .A1(n10216), .A2(n5768), .A3(n5767), .A4(n6032), .ZN(n5769)
         );
  NOR2_X1 U7280 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  NAND2_X1 U7281 ( .A1(n5762), .A2(n5771), .ZN(n6067) );
  INV_X1 U7282 ( .A(n6067), .ZN(n5773) );
  INV_X1 U7283 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U7284 ( .A1(n5773), .A2(n5772), .ZN(n5774) );
  NAND2_X1 U7285 ( .A1(n5774), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7286 ( .A1(n6088), .A2(n5775), .ZN(n5776) );
  NAND2_X1 U7287 ( .A1(n5776), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6102) );
  INV_X1 U7288 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U7289 ( .A1(n6102), .A2(n5777), .ZN(n5778) );
  NAND2_X1 U7290 ( .A1(n5778), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5780) );
  INV_X1 U7291 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5779) );
  XNOR2_X2 U7292 ( .A(n5780), .B(n5779), .ZN(n9014) );
  XNOR2_X1 U7293 ( .A(n5782), .B(n6234), .ZN(n6027) );
  INV_X1 U7294 ( .A(n6027), .ZN(n6029) );
  NAND2_X1 U7295 ( .A1(n9014), .A2(n9007), .ZN(n6705) );
  INV_X1 U7296 ( .A(n6705), .ZN(n9002) );
  NAND2_X1 U7297 ( .A1(n9002), .A2(n7434), .ZN(n5783) );
  NAND2_X1 U7298 ( .A1(n9131), .A2(n9007), .ZN(n9000) );
  AND3_X4 U7299 ( .A1(n6906), .A2(n5783), .A3(n6320), .ZN(n8626) );
  AOI22_X1 U7300 ( .A1(n9683), .A2(n6194), .B1(n8626), .B2(n9024), .ZN(n6028)
         );
  NAND2_X1 U7301 ( .A1(n5834), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5788) );
  INV_X1 U7302 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5784) );
  OR2_X1 U7303 ( .A1(n5837), .A2(n5784), .ZN(n5787) );
  INV_X1 U7304 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6920) );
  OR2_X1 U7305 ( .A1(n5971), .A2(n6920), .ZN(n5786) );
  NAND2_X1 U7306 ( .A1(n6822), .A2(n8626), .ZN(n5791) );
  NAND2_X1 U7307 ( .A1(n7868), .A2(SI_0_), .ZN(n5789) );
  XNOR2_X1 U7308 ( .A(n5789), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9577) );
  MUX2_X1 U7309 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9577), .S(n6391), .Z(n6862) );
  INV_X1 U7310 ( .A(n6320), .ZN(n5792) );
  AOI22_X1 U7311 ( .A1(n6862), .A2(n8625), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n5792), .ZN(n5790) );
  NAND2_X1 U7312 ( .A1(n5791), .A2(n5790), .ZN(n6580) );
  NAND2_X1 U7313 ( .A1(n5792), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7314 ( .A1(n6580), .A2(n6581), .ZN(n6583) );
  AND2_X1 U7315 ( .A1(n6583), .A2(n5794), .ZN(n6574) );
  NAND2_X1 U7316 ( .A1(n5836), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5797) );
  INV_X1 U7317 ( .A(n5837), .ZN(n5795) );
  NAND2_X1 U7318 ( .A1(n5795), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U7319 ( .A1(n5813), .A2(n5755), .ZN(n5811) );
  NOR2_X1 U7320 ( .A1(n7868), .A2(n6397), .ZN(n5800) );
  AOI21_X1 U7321 ( .B1(n6376), .B2(n7868), .A(n5800), .ZN(n5809) );
  INV_X1 U7322 ( .A(n6391), .ZN(n5805) );
  INV_X1 U7323 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7324 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5802) );
  XNOR2_X1 U7325 ( .A(n5803), .B(n5802), .ZN(n6433) );
  INV_X1 U7326 ( .A(n6433), .ZN(n5804) );
  INV_X1 U7327 ( .A(n9721), .ZN(n9138) );
  NAND2_X1 U7328 ( .A1(n5087), .A2(n6397), .ZN(n5806) );
  OAI211_X1 U7329 ( .C1(n6376), .C2(n5087), .A(n9138), .B(n5806), .ZN(n5807)
         );
  NAND2_X1 U7330 ( .A1(n6957), .A2(n8631), .ZN(n5810) );
  NAND2_X1 U7331 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  AND2_X1 U7332 ( .A1(n6957), .A2(n5755), .ZN(n5814) );
  XNOR2_X1 U7333 ( .A(n5815), .B(n5816), .ZN(n6572) );
  NAND2_X1 U7334 ( .A1(n6574), .A2(n6572), .ZN(n6573) );
  INV_X1 U7335 ( .A(n5815), .ZN(n5817) );
  NAND2_X1 U7336 ( .A1(n5817), .A2(n5816), .ZN(n5818) );
  NAND2_X1 U7337 ( .A1(n6573), .A2(n5818), .ZN(n6626) );
  NAND2_X1 U7338 ( .A1(n5834), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7339 ( .A1(n5836), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5821) );
  INV_X1 U7340 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6631) );
  OR2_X1 U7341 ( .A1(n5837), .A2(n6631), .ZN(n5819) );
  OR2_X1 U7342 ( .A1(n5823), .A2(n9562), .ZN(n5825) );
  INV_X1 U7343 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7344 ( .A1(n5825), .A2(n5824), .ZN(n5842) );
  OAI21_X1 U7345 ( .B1(n5825), .B2(n5824), .A(n5842), .ZN(n6640) );
  NAND2_X1 U7346 ( .A1(n7047), .A2(n8631), .ZN(n5827) );
  AND2_X1 U7347 ( .A1(n7047), .A2(n8625), .ZN(n5828) );
  AOI21_X1 U7348 ( .B1(n9034), .B2(n8626), .A(n5828), .ZN(n5830) );
  XNOR2_X1 U7349 ( .A(n5829), .B(n5830), .ZN(n6627) );
  NAND2_X1 U7350 ( .A1(n6626), .A2(n6627), .ZN(n5833) );
  INV_X1 U7351 ( .A(n5829), .ZN(n5831) );
  NAND2_X1 U7352 ( .A1(n5831), .A2(n5830), .ZN(n5832) );
  NAND2_X1 U7353 ( .A1(n5833), .A2(n5832), .ZN(n6675) );
  NAND2_X1 U7354 ( .A1(n5834), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7355 ( .A1(n5835), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5840) );
  NAND2_X1 U7356 ( .A1(n5836), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5839) );
  OR2_X1 U7357 ( .A1(n5837), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5838) );
  NAND4_X1 U7358 ( .A1(n5841), .A2(n5840), .A3(n5839), .A4(n5838), .ZN(n10048)
         );
  NAND2_X1 U7359 ( .A1(n10048), .A2(n6194), .ZN(n5849) );
  NAND2_X1 U7360 ( .A1(n5842), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5844) );
  INV_X1 U7361 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5843) );
  XNOR2_X1 U7362 ( .A(n5844), .B(n5843), .ZN(n6438) );
  INV_X1 U7363 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6399) );
  OR2_X1 U7364 ( .A1(n5845), .A2(n6399), .ZN(n5846) );
  NAND2_X1 U7365 ( .A1(n6878), .A2(n6261), .ZN(n5848) );
  NAND2_X1 U7366 ( .A1(n5849), .A2(n5848), .ZN(n5850) );
  XNOR2_X1 U7367 ( .A(n5850), .B(n6234), .ZN(n5852) );
  AND2_X1 U7368 ( .A1(n6878), .A2(n6194), .ZN(n5851) );
  AOI21_X1 U7369 ( .B1(n10048), .B2(n8626), .A(n5851), .ZN(n5853) );
  XNOR2_X1 U7370 ( .A(n5852), .B(n5853), .ZN(n6676) );
  NAND2_X1 U7371 ( .A1(n6675), .A2(n6676), .ZN(n5856) );
  INV_X1 U7372 ( .A(n5852), .ZN(n5854) );
  NAND2_X1 U7373 ( .A1(n5854), .A2(n5853), .ZN(n5855) );
  NAND2_X1 U7374 ( .A1(n5856), .A2(n5855), .ZN(n6817) );
  INV_X1 U7375 ( .A(n6817), .ZN(n5871) );
  NAND2_X1 U7376 ( .A1(n8757), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7377 ( .A1(n8755), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5860) );
  NOR2_X1 U7378 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5857) );
  NOR2_X1 U7379 ( .A1(n5877), .A2(n5857), .ZN(n7118) );
  NAND2_X1 U7380 ( .A1(n5795), .A2(n7118), .ZN(n5859) );
  NAND2_X1 U7381 ( .A1(n8756), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5858) );
  NAND2_X1 U7382 ( .A1(n9033), .A2(n6194), .ZN(n5867) );
  NAND2_X1 U7383 ( .A1(n5862), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5863) );
  MUX2_X1 U7384 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5863), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5864) );
  INV_X1 U7385 ( .A(n5762), .ZN(n5882) );
  NAND2_X1 U7386 ( .A1(n5864), .A2(n5882), .ZN(n9740) );
  OR2_X1 U7387 ( .A1(n6378), .A2(n5826), .ZN(n5865) );
  NAND2_X1 U7388 ( .A1(n7119), .A2(n6261), .ZN(n5866) );
  NAND2_X1 U7389 ( .A1(n5867), .A2(n5866), .ZN(n5868) );
  XNOR2_X1 U7390 ( .A(n5868), .B(n8629), .ZN(n5872) );
  AND2_X1 U7391 ( .A1(n7119), .A2(n6194), .ZN(n5869) );
  AOI21_X1 U7392 ( .B1(n9033), .B2(n8626), .A(n5869), .ZN(n5873) );
  XNOR2_X1 U7393 ( .A(n5872), .B(n5873), .ZN(n6818) );
  NAND2_X1 U7394 ( .A1(n5871), .A2(n5870), .ZN(n6815) );
  INV_X1 U7395 ( .A(n5872), .ZN(n5875) );
  INV_X1 U7396 ( .A(n5873), .ZN(n5874) );
  NAND2_X1 U7397 ( .A1(n5875), .A2(n5874), .ZN(n5876) );
  NAND2_X1 U7398 ( .A1(n6815), .A2(n5876), .ZN(n5889) );
  NAND2_X1 U7399 ( .A1(n8755), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U7400 ( .A1(n8756), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5880) );
  NAND2_X1 U7401 ( .A1(n8757), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5879) );
  OAI21_X1 U7402 ( .B1(n5877), .B2(P1_REG3_REG_5__SCAN_IN), .A(n5901), .ZN(
        n9883) );
  OR2_X1 U7403 ( .A1(n8635), .A2(n9883), .ZN(n5878) );
  NAND4_X1 U7404 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n9032)
         );
  NAND2_X1 U7405 ( .A1(n9032), .A2(n6194), .ZN(n5887) );
  OR2_X1 U7406 ( .A1(n6372), .A2(n5826), .ZN(n5885) );
  NAND2_X1 U7407 ( .A1(n5882), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  XNOR2_X1 U7408 ( .A(n5883), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9059) );
  AOI22_X1 U7409 ( .A1(n6121), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6120), .B2(
        n9059), .ZN(n5884) );
  NAND2_X1 U7410 ( .A1(n5885), .A2(n5884), .ZN(n9715) );
  NAND2_X1 U7411 ( .A1(n9715), .A2(n6261), .ZN(n5886) );
  NAND2_X1 U7412 ( .A1(n5887), .A2(n5886), .ZN(n5888) );
  XNOR2_X1 U7413 ( .A(n5888), .B(n6234), .ZN(n5890) );
  NAND2_X1 U7414 ( .A1(n5889), .A2(n5890), .ZN(n9708) );
  AOI22_X1 U7415 ( .A1(n9032), .A2(n8626), .B1(n6194), .B2(n9715), .ZN(n9711)
         );
  INV_X1 U7416 ( .A(n5889), .ZN(n5892) );
  OR2_X1 U7417 ( .A1(n6384), .A2(n5826), .ZN(n5899) );
  NOR2_X1 U7418 ( .A1(n5893), .A2(n9562), .ZN(n5894) );
  NAND2_X1 U7419 ( .A1(n5894), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5897) );
  INV_X1 U7420 ( .A(n5894), .ZN(n5896) );
  INV_X1 U7421 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7422 ( .A1(n5896), .A2(n5895), .ZN(n5914) );
  AND2_X1 U7423 ( .A1(n5897), .A2(n5914), .ZN(n9071) );
  AOI22_X1 U7424 ( .A1(n6121), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6120), .B2(
        n9071), .ZN(n5898) );
  NAND2_X1 U7425 ( .A1(n5899), .A2(n5898), .ZN(n7108) );
  NAND2_X1 U7426 ( .A1(n7108), .A2(n8631), .ZN(n5908) );
  NAND2_X1 U7427 ( .A1(n8757), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5906) );
  NAND2_X1 U7428 ( .A1(n8755), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U7429 ( .A1(n8756), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5904) );
  AND2_X1 U7430 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  OR2_X1 U7431 ( .A1(n5902), .A2(n5918), .ZN(n7106) );
  OR2_X1 U7432 ( .A1(n8635), .A2(n7106), .ZN(n5903) );
  NAND4_X1 U7433 ( .A1(n5906), .A2(n5905), .A3(n5904), .A4(n5903), .ZN(n9031)
         );
  NAND2_X1 U7434 ( .A1(n9031), .A2(n6194), .ZN(n5907) );
  NAND2_X1 U7435 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  XNOR2_X1 U7436 ( .A(n5909), .B(n8629), .ZN(n5910) );
  AOI22_X1 U7437 ( .A1(n7108), .A2(n6194), .B1(n9031), .B2(n8626), .ZN(n5911)
         );
  AND2_X1 U7438 ( .A1(n5910), .A2(n5911), .ZN(n6838) );
  INV_X1 U7439 ( .A(n5910), .ZN(n5913) );
  INV_X1 U7440 ( .A(n5911), .ZN(n5912) );
  NAND2_X1 U7441 ( .A1(n5913), .A2(n5912), .ZN(n6960) );
  NAND2_X1 U7442 ( .A1(n6400), .A2(n8781), .ZN(n5917) );
  NAND2_X1 U7443 ( .A1(n5914), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5915) );
  XNOR2_X1 U7444 ( .A(n5915), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9083) );
  AOI22_X1 U7445 ( .A1(n6121), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6120), .B2(
        n9083), .ZN(n5916) );
  NAND2_X1 U7446 ( .A1(n7181), .A2(n8631), .ZN(n5925) );
  NAND2_X1 U7447 ( .A1(n8755), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7448 ( .A1(n8757), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7449 ( .A1(n8756), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5921) );
  OR2_X1 U7450 ( .A1(n5918), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U7451 ( .A1(n5951), .A2(n5919), .ZN(n7094) );
  OR2_X1 U7452 ( .A1(n8635), .A2(n7094), .ZN(n5920) );
  NAND4_X1 U7453 ( .A1(n5923), .A2(n5922), .A3(n5921), .A4(n5920), .ZN(n9030)
         );
  NAND2_X1 U7454 ( .A1(n9030), .A2(n6194), .ZN(n5924) );
  NAND2_X1 U7455 ( .A1(n5925), .A2(n5924), .ZN(n5926) );
  XNOR2_X1 U7456 ( .A(n5926), .B(n8629), .ZN(n6963) );
  INV_X1 U7457 ( .A(n6963), .ZN(n5928) );
  AND2_X1 U7458 ( .A1(n9030), .A2(n8626), .ZN(n5927) );
  AOI21_X1 U7459 ( .B1(n7181), .B2(n6194), .A(n5927), .ZN(n5930) );
  INV_X1 U7460 ( .A(n5930), .ZN(n6962) );
  NAND2_X1 U7461 ( .A1(n5928), .A2(n6962), .ZN(n5929) );
  NAND2_X1 U7462 ( .A1(n6404), .A2(n8781), .ZN(n5935) );
  NAND2_X1 U7463 ( .A1(n5931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5932) );
  MUX2_X1 U7464 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5932), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5933) );
  AND2_X1 U7465 ( .A1(n5933), .A2(n5944), .ZN(n6449) );
  AOI22_X1 U7466 ( .A1(n6121), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6120), .B2(
        n6449), .ZN(n5934) );
  NAND2_X1 U7467 ( .A1(n5935), .A2(n5934), .ZN(n9873) );
  NAND2_X1 U7468 ( .A1(n9873), .A2(n8631), .ZN(n5941) );
  NAND2_X1 U7469 ( .A1(n8755), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5939) );
  NAND2_X1 U7470 ( .A1(n8757), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5938) );
  NAND2_X1 U7471 ( .A1(n8756), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5937) );
  INV_X1 U7472 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7473 ( .A(n5951), .B(n5950), .ZN(n9870) );
  OR2_X1 U7474 ( .A1(n8635), .A2(n9870), .ZN(n5936) );
  NAND4_X1 U7475 ( .A1(n5939), .A2(n5938), .A3(n5937), .A4(n5936), .ZN(n9029)
         );
  NAND2_X1 U7476 ( .A1(n9029), .A2(n8625), .ZN(n5940) );
  NAND2_X1 U7477 ( .A1(n5941), .A2(n5940), .ZN(n5942) );
  XNOR2_X1 U7478 ( .A(n5942), .B(n8629), .ZN(n7218) );
  AND2_X1 U7479 ( .A1(n9029), .A2(n8626), .ZN(n5943) );
  AOI21_X1 U7480 ( .B1(n9873), .B2(n6194), .A(n5943), .ZN(n9698) );
  NAND2_X1 U7481 ( .A1(n6460), .A2(n8781), .ZN(n5947) );
  NAND2_X1 U7482 ( .A1(n5944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5945) );
  XNOR2_X1 U7483 ( .A(n5945), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9107) );
  AOI22_X1 U7484 ( .A1(n6121), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6120), .B2(
        n9107), .ZN(n5946) );
  NAND2_X1 U7485 ( .A1(n7306), .A2(n6261), .ZN(n5958) );
  NAND2_X1 U7486 ( .A1(n8757), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5956) );
  INV_X1 U7487 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7488 ( .A1(n6212), .A2(n5948), .ZN(n5955) );
  NAND2_X1 U7489 ( .A1(n8756), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5954) );
  INV_X1 U7490 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5949) );
  OAI21_X1 U7491 ( .B1(n5951), .B2(n5950), .A(n5949), .ZN(n5952) );
  NAND2_X1 U7492 ( .A1(n5952), .A2(n5972), .ZN(n7230) );
  OR2_X1 U7493 ( .A1(n8635), .A2(n7230), .ZN(n5953) );
  NAND4_X1 U7494 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n9028)
         );
  NAND2_X1 U7495 ( .A1(n9028), .A2(n8625), .ZN(n5957) );
  NAND2_X1 U7496 ( .A1(n5958), .A2(n5957), .ZN(n5959) );
  XNOR2_X1 U7497 ( .A(n5959), .B(n6234), .ZN(n5966) );
  AND2_X1 U7498 ( .A1(n9028), .A2(n8626), .ZN(n5960) );
  AOI21_X1 U7499 ( .B1(n7306), .B2(n6194), .A(n5960), .ZN(n5964) );
  XNOR2_X1 U7500 ( .A(n5966), .B(n5964), .ZN(n7221) );
  NAND2_X1 U7501 ( .A1(n5963), .A2(n5962), .ZN(n7223) );
  INV_X1 U7502 ( .A(n5964), .ZN(n5965) );
  OR2_X1 U7503 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  NAND2_X1 U7504 ( .A1(n7223), .A2(n5967), .ZN(n5979) );
  NAND2_X1 U7505 ( .A1(n6464), .A2(n8781), .ZN(n5970) );
  NAND2_X1 U7506 ( .A1(n5968), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5985) );
  XNOR2_X1 U7507 ( .A(n5985), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9111) );
  AOI22_X1 U7508 ( .A1(n6121), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6120), .B2(
        n9111), .ZN(n5969) );
  NAND2_X1 U7509 ( .A1(n8755), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5977) );
  NAND2_X1 U7510 ( .A1(n8757), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5976) );
  INV_X1 U7511 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7308) );
  OR2_X1 U7512 ( .A1(n6242), .A2(n7308), .ZN(n5975) );
  AND2_X1 U7513 ( .A1(n5972), .A2(n9590), .ZN(n5973) );
  OR2_X1 U7514 ( .A1(n5973), .A2(n5990), .ZN(n9666) );
  OR2_X1 U7515 ( .A1(n8635), .A2(n9666), .ZN(n5974) );
  NAND4_X1 U7516 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n9027)
         );
  AOI22_X1 U7517 ( .A1(n9664), .A2(n8631), .B1(n6194), .B2(n9027), .ZN(n5978)
         );
  XNOR2_X1 U7518 ( .A(n5978), .B(n6234), .ZN(n5980) );
  INV_X1 U7519 ( .A(n5979), .ZN(n5982) );
  INV_X1 U7520 ( .A(n5980), .ZN(n5981) );
  INV_X1 U7521 ( .A(n9664), .ZN(n7333) );
  INV_X1 U7522 ( .A(n8626), .ZN(n6217) );
  OAI22_X1 U7523 ( .A1(n7333), .A2(n6218), .B1(n7413), .B2(n6217), .ZN(n9659)
         );
  INV_X1 U7524 ( .A(n5983), .ZN(n9687) );
  NAND2_X1 U7525 ( .A1(n6488), .A2(n8781), .ZN(n5989) );
  NAND2_X1 U7526 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U7527 ( .A1(n5986), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5987) );
  XNOR2_X1 U7528 ( .A(n5987), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9754) );
  AOI22_X1 U7529 ( .A1(n6121), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6120), .B2(
        n9754), .ZN(n5988) );
  NAND2_X1 U7530 ( .A1(n9693), .A2(n8631), .ZN(n5997) );
  NOR2_X1 U7531 ( .A1(n5990), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5991) );
  OR2_X1 U7532 ( .A1(n6008), .A2(n5991), .ZN(n9695) );
  OR2_X1 U7533 ( .A1(n8635), .A2(n9695), .ZN(n5995) );
  NAND2_X1 U7534 ( .A1(n8755), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5994) );
  NAND2_X1 U7535 ( .A1(n8757), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5993) );
  INV_X1 U7536 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7419) );
  OR2_X1 U7537 ( .A1(n6242), .A2(n7419), .ZN(n5992) );
  NAND4_X1 U7538 ( .A1(n5995), .A2(n5994), .A3(n5993), .A4(n5992), .ZN(n9026)
         );
  NAND2_X1 U7539 ( .A1(n9026), .A2(n6194), .ZN(n5996) );
  NAND2_X1 U7540 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7541 ( .A(n5998), .B(n8629), .ZN(n6000) );
  AND2_X1 U7542 ( .A1(n9026), .A2(n8626), .ZN(n5999) );
  AOI21_X1 U7543 ( .B1(n9693), .B2(n6194), .A(n5999), .ZN(n6001) );
  NAND2_X1 U7544 ( .A1(n6000), .A2(n6001), .ZN(n9673) );
  INV_X1 U7545 ( .A(n6000), .ZN(n6003) );
  INV_X1 U7546 ( .A(n6001), .ZN(n6002) );
  NAND2_X1 U7547 ( .A1(n6003), .A2(n6002), .ZN(n6004) );
  AND2_X1 U7548 ( .A1(n9673), .A2(n6004), .ZN(n9686) );
  NAND2_X1 U7549 ( .A1(n6569), .A2(n8781), .ZN(n6007) );
  XNOR2_X1 U7550 ( .A(P1_IR_REG_12__SCAN_IN), .B(n6005), .ZN(n9113) );
  AOI22_X1 U7551 ( .A1(n6121), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6120), .B2(
        n9113), .ZN(n6006) );
  NAND2_X1 U7552 ( .A1(n9861), .A2(n6261), .ZN(n6017) );
  NAND2_X1 U7553 ( .A1(n8755), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7554 ( .A1(n8756), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7555 ( .A1(n8757), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6013) );
  INV_X1 U7556 ( .A(n6008), .ZN(n6009) );
  INV_X1 U7557 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10087) );
  NAND2_X1 U7558 ( .A1(n6009), .A2(n10087), .ZN(n6010) );
  NAND2_X1 U7559 ( .A1(n6011), .A2(n6010), .ZN(n9859) );
  OR2_X1 U7560 ( .A1(n8635), .A2(n9859), .ZN(n6012) );
  NAND4_X1 U7561 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n9025)
         );
  NAND2_X1 U7562 ( .A1(n9025), .A2(n6194), .ZN(n6016) );
  NAND2_X1 U7563 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  XNOR2_X1 U7564 ( .A(n6018), .B(n8629), .ZN(n6020) );
  AND2_X1 U7565 ( .A1(n9025), .A2(n8626), .ZN(n6019) );
  AOI21_X1 U7566 ( .B1(n9861), .B2(n6194), .A(n6019), .ZN(n6021) );
  NAND2_X1 U7567 ( .A1(n6020), .A2(n6021), .ZN(n6025) );
  INV_X1 U7568 ( .A(n6020), .ZN(n6023) );
  INV_X1 U7569 ( .A(n6021), .ZN(n6022) );
  NAND2_X1 U7570 ( .A1(n6023), .A2(n6022), .ZN(n6024) );
  NAND2_X1 U7571 ( .A1(n6025), .A2(n6024), .ZN(n9672) );
  INV_X1 U7572 ( .A(n6025), .ZN(n6026) );
  XOR2_X1 U7573 ( .A(n6028), .B(n6027), .Z(n9678) );
  NAND2_X1 U7574 ( .A1(n6651), .A2(n8781), .ZN(n6034) );
  AND2_X1 U7575 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6030) );
  XNOR2_X1 U7576 ( .A(n6048), .B(n6032), .ZN(n9794) );
  AOI22_X1 U7577 ( .A1(n6121), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n9794), .B2(
        n6120), .ZN(n6033) );
  NAND2_X1 U7578 ( .A1(n8755), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7579 ( .A1(n8757), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6040) );
  INV_X1 U7580 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7581 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  NAND2_X1 U7582 ( .A1(n6054), .A2(n6037), .ZN(n8594) );
  OR2_X1 U7583 ( .A1(n8635), .A2(n8594), .ZN(n6039) );
  INV_X1 U7584 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7556) );
  OR2_X1 U7585 ( .A1(n6242), .A2(n7556), .ZN(n6038) );
  NAND4_X1 U7586 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9023)
         );
  AOI22_X1 U7587 ( .A1(n7605), .A2(n8631), .B1(n6194), .B2(n9023), .ZN(n6042)
         );
  XOR2_X1 U7588 ( .A(n6234), .B(n6042), .Z(n6043) );
  AND2_X1 U7589 ( .A1(n6044), .A2(n6043), .ZN(n6045) );
  NOR2_X2 U7590 ( .A1(n6044), .A2(n6043), .ZN(n6046) );
  NOR2_X2 U7591 ( .A1(n6045), .A2(n6046), .ZN(n8591) );
  AOI22_X1 U7592 ( .A1(n7605), .A2(n6194), .B1(n8626), .B2(n9023), .ZN(n8592)
         );
  NAND2_X1 U7593 ( .A1(n8591), .A2(n8592), .ZN(n8590) );
  INV_X1 U7594 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7595 ( .A1(n8590), .A2(n6047), .ZN(n6064) );
  INV_X1 U7596 ( .A(n6064), .ZN(n6062) );
  NAND2_X1 U7597 ( .A1(n6718), .A2(n8781), .ZN(n6051) );
  OAI21_X1 U7598 ( .B1(n6048), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6049) );
  XNOR2_X1 U7599 ( .A(n6049), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9806) );
  AOI22_X1 U7600 ( .A1(n9806), .A2(n6120), .B1(n6121), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n6050) );
  INV_X1 U7601 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n10168) );
  OR2_X1 U7602 ( .A1(n6052), .A2(n10168), .ZN(n6059) );
  INV_X1 U7603 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9799) );
  OR2_X1 U7604 ( .A1(n6212), .A2(n9799), .ZN(n6058) );
  NAND2_X1 U7605 ( .A1(n8756), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6057) );
  INV_X1 U7606 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6053) );
  INV_X1 U7607 ( .A(n6071), .ZN(n6073) );
  NAND2_X1 U7608 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  NAND2_X1 U7609 ( .A1(n6073), .A2(n6055), .ZN(n8746) );
  OR2_X1 U7610 ( .A1(n8635), .A2(n8746), .ZN(n6056) );
  NAND4_X1 U7611 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n9171)
         );
  AOI22_X1 U7612 ( .A1(n9555), .A2(n8631), .B1(n6194), .B2(n9171), .ZN(n6060)
         );
  XNOR2_X1 U7613 ( .A(n6060), .B(n6234), .ZN(n6063) );
  INV_X1 U7614 ( .A(n6063), .ZN(n6061) );
  NAND2_X1 U7615 ( .A1(n6062), .A2(n6061), .ZN(n6065) );
  AOI22_X1 U7616 ( .A1(n9555), .A2(n6194), .B1(n8626), .B2(n9171), .ZN(n8744)
         );
  NAND2_X1 U7617 ( .A1(n6741), .A2(n8781), .ZN(n6070) );
  NAND2_X1 U7618 ( .A1(n6067), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6068) );
  XNOR2_X1 U7619 ( .A(n6068), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9821) );
  AOI22_X1 U7620 ( .A1(n6121), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6120), .B2(
        n9821), .ZN(n6069) );
  NAND2_X1 U7621 ( .A1(n9494), .A2(n6261), .ZN(n6080) );
  NAND2_X1 U7622 ( .A1(n8755), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6078) );
  INV_X1 U7623 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10336) );
  OR2_X1 U7624 ( .A1(n6052), .A2(n10336), .ZN(n6077) );
  NAND2_X1 U7625 ( .A1(n8756), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6076) );
  INV_X1 U7626 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7627 ( .A1(n6073), .A2(n6072), .ZN(n6074) );
  NAND2_X1 U7628 ( .A1(n6108), .A2(n6074), .ZN(n9414) );
  OR2_X1 U7629 ( .A1(n8635), .A2(n9414), .ZN(n6075) );
  NAND4_X1 U7630 ( .A1(n6078), .A2(n6077), .A3(n6076), .A4(n6075), .ZN(n9172)
         );
  NAND2_X1 U7631 ( .A1(n9172), .A2(n6194), .ZN(n6079) );
  NAND2_X1 U7632 ( .A1(n6080), .A2(n6079), .ZN(n6081) );
  XNOR2_X1 U7633 ( .A(n6081), .B(n6234), .ZN(n6085) );
  NAND2_X1 U7634 ( .A1(n9494), .A2(n6194), .ZN(n6083) );
  NAND2_X1 U7635 ( .A1(n9172), .A2(n8626), .ZN(n6082) );
  NAND2_X1 U7636 ( .A1(n6083), .A2(n6082), .ZN(n6084) );
  NOR2_X1 U7637 ( .A1(n6085), .A2(n6084), .ZN(n6086) );
  AOI21_X1 U7638 ( .B1(n6085), .B2(n6084), .A(n6086), .ZN(n8672) );
  INV_X1 U7639 ( .A(n6086), .ZN(n6087) );
  NAND2_X1 U7640 ( .A1(n6896), .A2(n8781), .ZN(n6090) );
  XNOR2_X1 U7641 ( .A(n6088), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9831) );
  AOI22_X1 U7642 ( .A1(n6121), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6120), .B2(
        n9831), .ZN(n6089) );
  NAND2_X1 U7643 ( .A1(n9392), .A2(n6261), .ZN(n6096) );
  XNOR2_X1 U7644 ( .A(n6108), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9393) );
  NAND2_X1 U7645 ( .A1(n5795), .A2(n9393), .ZN(n6094) );
  NAND2_X1 U7646 ( .A1(n8755), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7647 ( .A1(n8756), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6092) );
  INV_X1 U7648 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n10051) );
  OR2_X1 U7649 ( .A1(n6052), .A2(n10051), .ZN(n6091) );
  NAND4_X1 U7650 ( .A1(n6094), .A2(n6093), .A3(n6092), .A4(n6091), .ZN(n9173)
         );
  NAND2_X1 U7651 ( .A1(n9173), .A2(n6194), .ZN(n6095) );
  NAND2_X1 U7652 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  XNOR2_X1 U7653 ( .A(n6097), .B(n6234), .ZN(n6100) );
  AOI22_X1 U7654 ( .A1(n9392), .A2(n6194), .B1(n8626), .B2(n9173), .ZN(n6098)
         );
  XNOR2_X1 U7655 ( .A(n6100), .B(n6098), .ZN(n8683) );
  NAND2_X1 U7656 ( .A1(n8680), .A2(n8683), .ZN(n8681) );
  INV_X1 U7657 ( .A(n6098), .ZN(n6099) );
  NAND2_X1 U7658 ( .A1(n8681), .A2(n6101), .ZN(n6116) );
  NAND2_X1 U7659 ( .A1(n6991), .A2(n8781), .ZN(n6104) );
  XNOR2_X1 U7660 ( .A(n6102), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9123) );
  AOI22_X1 U7661 ( .A1(n6121), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6120), .B2(
        n9123), .ZN(n6103) );
  INV_X1 U7662 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6106) );
  INV_X1 U7663 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6105) );
  OAI21_X1 U7664 ( .B1(n6108), .B2(n6106), .A(n6105), .ZN(n6109) );
  NAND2_X1 U7665 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n6107) );
  NAND2_X1 U7666 ( .A1(n6109), .A2(n6124), .ZN(n9365) );
  NAND2_X1 U7667 ( .A1(n8756), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7668 ( .B1(n9365), .B2(n8635), .A(n6110), .ZN(n6113) );
  INV_X1 U7669 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U7670 ( .A1(n8755), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7671 ( .B1(n6052), .B2(n10315), .A(n6111), .ZN(n6112) );
  OR2_X1 U7672 ( .A1(n6113), .A2(n6112), .ZN(n9177) );
  AOI22_X1 U7673 ( .A1(n9377), .A2(n8631), .B1(n6194), .B2(n9177), .ZN(n6114)
         );
  XNOR2_X1 U7674 ( .A(n6114), .B(n6234), .ZN(n6115) );
  NAND2_X1 U7675 ( .A1(n6116), .A2(n6115), .ZN(n6119) );
  OAI21_X1 U7676 ( .B1(n6116), .B2(n6115), .A(n6119), .ZN(n8721) );
  INV_X1 U7677 ( .A(n8721), .ZN(n6118) );
  INV_X1 U7678 ( .A(n9177), .ZN(n9176) );
  OAI22_X1 U7679 ( .A1(n9548), .A2(n6218), .B1(n9176), .B2(n6217), .ZN(n8724)
         );
  NAND2_X1 U7680 ( .A1(n7172), .A2(n8781), .ZN(n6123) );
  AOI22_X1 U7681 ( .A1(n6121), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n6120), .B2(
        n9131), .ZN(n6122) );
  NAND2_X1 U7682 ( .A1(n9357), .A2(n6261), .ZN(n6131) );
  INV_X1 U7683 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9359) );
  INV_X1 U7684 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10178) );
  INV_X1 U7685 ( .A(n6139), .ZN(n6141) );
  NAND2_X1 U7686 ( .A1(n6124), .A2(n10178), .ZN(n6125) );
  NAND2_X1 U7687 ( .A1(n6141), .A2(n6125), .ZN(n9358) );
  OR2_X1 U7688 ( .A1(n9358), .A2(n8635), .ZN(n6129) );
  NAND2_X1 U7689 ( .A1(n8757), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6127) );
  INV_X1 U7690 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10323) );
  OR2_X1 U7691 ( .A1(n6212), .A2(n10323), .ZN(n6126) );
  AND2_X1 U7692 ( .A1(n6127), .A2(n6126), .ZN(n6128) );
  OAI211_X1 U7693 ( .C1(n6242), .C2(n9359), .A(n6129), .B(n6128), .ZN(n9179)
         );
  NAND2_X1 U7694 ( .A1(n9179), .A2(n6194), .ZN(n6130) );
  NAND2_X1 U7695 ( .A1(n6131), .A2(n6130), .ZN(n6132) );
  XNOR2_X1 U7696 ( .A(n6132), .B(n6234), .ZN(n6133) );
  AOI22_X1 U7697 ( .A1(n9357), .A2(n6194), .B1(n8626), .B2(n9179), .ZN(n6134)
         );
  XNOR2_X1 U7698 ( .A(n6133), .B(n6134), .ZN(n8614) );
  INV_X1 U7699 ( .A(n6133), .ZN(n6135) );
  NAND2_X1 U7700 ( .A1(n6135), .A2(n6134), .ZN(n6136) );
  NAND2_X1 U7701 ( .A1(n7258), .A2(n8781), .ZN(n6138) );
  INV_X1 U7702 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7292) );
  OR2_X1 U7703 ( .A1(n8782), .A2(n7292), .ZN(n6137) );
  NAND2_X1 U7704 ( .A1(n9342), .A2(n8631), .ZN(n6146) );
  INV_X1 U7705 ( .A(n6156), .ZN(n6157) );
  INV_X1 U7706 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7707 ( .A1(n6141), .A2(n6140), .ZN(n6142) );
  NAND2_X1 U7708 ( .A1(n6157), .A2(n6142), .ZN(n9340) );
  AOI22_X1 U7709 ( .A1(n8755), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n8757), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7710 ( .A1(n8756), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6143) );
  OAI211_X1 U7711 ( .C1(n9340), .C2(n8635), .A(n6144), .B(n6143), .ZN(n9183)
         );
  NAND2_X1 U7712 ( .A1(n9183), .A2(n6194), .ZN(n6145) );
  NAND2_X1 U7713 ( .A1(n6146), .A2(n6145), .ZN(n6147) );
  XNOR2_X1 U7714 ( .A(n6147), .B(n6234), .ZN(n6153) );
  INV_X1 U7715 ( .A(n6153), .ZN(n6151) );
  NAND2_X1 U7716 ( .A1(n9342), .A2(n6194), .ZN(n6149) );
  NAND2_X1 U7717 ( .A1(n9183), .A2(n8626), .ZN(n6148) );
  NAND2_X1 U7718 ( .A1(n6149), .A2(n6148), .ZN(n6152) );
  INV_X1 U7719 ( .A(n6152), .ZN(n6150) );
  NAND2_X1 U7720 ( .A1(n6151), .A2(n6150), .ZN(n8702) );
  NAND2_X1 U7721 ( .A1(n7337), .A2(n8781), .ZN(n6155) );
  OR2_X1 U7722 ( .A1(n8782), .A2(n7338), .ZN(n6154) );
  NAND2_X1 U7723 ( .A1(n9326), .A2(n6261), .ZN(n6163) );
  INV_X1 U7724 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n6161) );
  INV_X1 U7725 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U7726 ( .A1(n6157), .A2(n8657), .ZN(n6158) );
  NAND2_X1 U7727 ( .A1(n6171), .A2(n6158), .ZN(n8655) );
  OR2_X1 U7728 ( .A1(n8655), .A2(n8635), .ZN(n6160) );
  AOI22_X1 U7729 ( .A1(n8755), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n8757), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7730 ( .C1(n6242), .C2(n6161), .A(n6160), .B(n6159), .ZN(n9185)
         );
  NAND2_X1 U7731 ( .A1(n9185), .A2(n6194), .ZN(n6162) );
  NAND2_X1 U7732 ( .A1(n6163), .A2(n6162), .ZN(n6164) );
  XNOR2_X1 U7733 ( .A(n6164), .B(n6234), .ZN(n6167) );
  AOI22_X1 U7734 ( .A1(n9326), .A2(n6194), .B1(n8626), .B2(n9185), .ZN(n6165)
         );
  XNOR2_X1 U7735 ( .A(n6167), .B(n6165), .ZN(n8653) );
  INV_X1 U7736 ( .A(n6165), .ZN(n6166) );
  NAND2_X1 U7737 ( .A1(n7433), .A2(n8781), .ZN(n6169) );
  OR2_X1 U7738 ( .A1(n8782), .A2(n10282), .ZN(n6168) );
  NAND2_X1 U7739 ( .A1(n9311), .A2(n6261), .ZN(n6179) );
  INV_X1 U7740 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n6170) );
  NAND2_X1 U7741 ( .A1(n6171), .A2(n6170), .ZN(n6172) );
  AND2_X1 U7742 ( .A1(n6187), .A2(n6172), .ZN(n9312) );
  NAND2_X1 U7743 ( .A1(n9312), .A2(n5795), .ZN(n6177) );
  INV_X1 U7744 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9466) );
  NAND2_X1 U7745 ( .A1(n8757), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6174) );
  NAND2_X1 U7746 ( .A1(n8756), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6173) );
  OAI211_X1 U7747 ( .C1(n6212), .C2(n9466), .A(n6174), .B(n6173), .ZN(n6175)
         );
  INV_X1 U7748 ( .A(n6175), .ZN(n6176) );
  NAND2_X1 U7749 ( .A1(n6177), .A2(n6176), .ZN(n9189) );
  NAND2_X1 U7750 ( .A1(n9189), .A2(n6194), .ZN(n6178) );
  NAND2_X1 U7751 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  XNOR2_X1 U7752 ( .A(n6180), .B(n8629), .ZN(n8714) );
  AND2_X1 U7753 ( .A1(n9189), .A2(n8626), .ZN(n6181) );
  NAND2_X1 U7754 ( .A1(n8712), .A2(n6182), .ZN(n6184) );
  NAND2_X1 U7755 ( .A1(n8714), .A2(n8713), .ZN(n6183) );
  NAND2_X1 U7756 ( .A1(n7507), .A2(n8781), .ZN(n6186) );
  OR2_X1 U7757 ( .A1(n8782), .A2(n7506), .ZN(n6185) );
  NAND2_X1 U7758 ( .A1(n9296), .A2(n6261), .ZN(n6196) );
  INV_X1 U7759 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8606) );
  INV_X1 U7760 ( .A(n6206), .ZN(n6207) );
  NAND2_X1 U7761 ( .A1(n6187), .A2(n8606), .ZN(n6188) );
  NAND2_X1 U7762 ( .A1(n6207), .A2(n6188), .ZN(n9297) );
  OR2_X1 U7763 ( .A1(n9297), .A2(n8635), .ZN(n6193) );
  INV_X1 U7764 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U7765 ( .A1(n8757), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7766 ( .A1(n8756), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n6189) );
  OAI211_X1 U7767 ( .C1(n6212), .C2(n9461), .A(n6190), .B(n6189), .ZN(n6191)
         );
  INV_X1 U7768 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7769 ( .A1(n6193), .A2(n6192), .ZN(n9191) );
  NAND2_X1 U7770 ( .A1(n9191), .A2(n6194), .ZN(n6195) );
  NAND2_X1 U7771 ( .A1(n6196), .A2(n6195), .ZN(n6197) );
  XNOR2_X1 U7772 ( .A(n6197), .B(n6234), .ZN(n6200) );
  NAND2_X1 U7773 ( .A1(n9296), .A2(n8625), .ZN(n6199) );
  NAND2_X1 U7774 ( .A1(n9191), .A2(n8626), .ZN(n6198) );
  NAND2_X1 U7775 ( .A1(n6199), .A2(n6198), .ZN(n6201) );
  NAND2_X1 U7776 ( .A1(n6200), .A2(n6201), .ZN(n8602) );
  INV_X1 U7777 ( .A(n6200), .ZN(n6203) );
  INV_X1 U7778 ( .A(n6201), .ZN(n6202) );
  NAND2_X1 U7779 ( .A1(n6203), .A2(n6202), .ZN(n8603) );
  NAND2_X1 U7780 ( .A1(n7590), .A2(n8781), .ZN(n6205) );
  OR2_X1 U7781 ( .A1(n8782), .A2(n7593), .ZN(n6204) );
  INV_X1 U7782 ( .A(n6225), .ZN(n6209) );
  INV_X1 U7783 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U7784 ( .A1(n6207), .A2(n8697), .ZN(n6208) );
  NAND2_X1 U7785 ( .A1(n6209), .A2(n6208), .ZN(n9282) );
  OR2_X1 U7786 ( .A1(n9282), .A2(n8635), .ZN(n6215) );
  INV_X1 U7787 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9456) );
  NAND2_X1 U7788 ( .A1(n8757), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7789 ( .A1(n8756), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n6210) );
  OAI211_X1 U7790 ( .C1(n6212), .C2(n9456), .A(n6211), .B(n6210), .ZN(n6213)
         );
  INV_X1 U7791 ( .A(n6213), .ZN(n6214) );
  NAND2_X1 U7792 ( .A1(n6215), .A2(n6214), .ZN(n9194) );
  AOI22_X1 U7793 ( .A1(n9281), .A2(n8631), .B1(n6194), .B2(n9194), .ZN(n6216)
         );
  XOR2_X1 U7794 ( .A(n6234), .B(n6216), .Z(n6220) );
  INV_X1 U7795 ( .A(n9194), .ZN(n9193) );
  OAI22_X1 U7796 ( .A1(n9526), .A2(n6218), .B1(n9193), .B2(n6217), .ZN(n6219)
         );
  NOR2_X1 U7797 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  AOI21_X1 U7798 ( .B1(n6220), .B2(n6219), .A(n6221), .ZN(n8693) );
  INV_X1 U7799 ( .A(n6221), .ZN(n6222) );
  OR2_X1 U7800 ( .A1(n8782), .A2(n7600), .ZN(n6223) );
  NAND2_X1 U7801 ( .A1(n9450), .A2(n6261), .ZN(n6233) );
  NOR2_X1 U7802 ( .A1(n6225), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7803 ( .A1(n6238), .A2(n6226), .ZN(n9267) );
  OR2_X1 U7804 ( .A1(n9267), .A2(n8635), .ZN(n6231) );
  INV_X1 U7805 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n10181) );
  NAND2_X1 U7806 ( .A1(n8755), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6228) );
  INV_X1 U7807 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10316) );
  OR2_X1 U7808 ( .A1(n6052), .A2(n10316), .ZN(n6227) );
  OAI211_X1 U7809 ( .C1(n10181), .C2(n6242), .A(n6228), .B(n6227), .ZN(n6229)
         );
  INV_X1 U7810 ( .A(n6229), .ZN(n6230) );
  NAND2_X1 U7811 ( .A1(n6231), .A2(n6230), .ZN(n9196) );
  NAND2_X1 U7812 ( .A1(n9196), .A2(n8625), .ZN(n6232) );
  NAND2_X1 U7813 ( .A1(n6233), .A2(n6232), .ZN(n6235) );
  XNOR2_X1 U7814 ( .A(n6235), .B(n6234), .ZN(n6253) );
  AOI22_X1 U7815 ( .A1(n9450), .A2(n6194), .B1(n8626), .B2(n9196), .ZN(n6251)
         );
  XNOR2_X1 U7816 ( .A(n6253), .B(n6251), .ZN(n8663) );
  OR2_X1 U7817 ( .A1(n8782), .A2(n9573), .ZN(n6236) );
  NAND2_X1 U7818 ( .A1(n9445), .A2(n6261), .ZN(n6248) );
  OR2_X1 U7819 ( .A1(n6238), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7820 ( .A1(n6238), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6262) );
  AND2_X1 U7821 ( .A1(n6239), .A2(n6262), .ZN(n9251) );
  NAND2_X1 U7822 ( .A1(n9251), .A2(n5795), .ZN(n6246) );
  INV_X1 U7823 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7824 ( .A1(n8755), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7825 ( .A1(n8757), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6240) );
  OAI211_X1 U7826 ( .C1(n6243), .C2(n6242), .A(n6241), .B(n6240), .ZN(n6244)
         );
  INV_X1 U7827 ( .A(n6244), .ZN(n6245) );
  NAND2_X1 U7828 ( .A1(n6246), .A2(n6245), .ZN(n9022) );
  NAND2_X1 U7829 ( .A1(n9022), .A2(n8625), .ZN(n6247) );
  NAND2_X1 U7830 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  XNOR2_X1 U7831 ( .A(n6249), .B(n8629), .ZN(n6255) );
  AND2_X1 U7832 ( .A1(n9022), .A2(n8626), .ZN(n6250) );
  AOI21_X1 U7833 ( .B1(n9445), .B2(n6194), .A(n6250), .ZN(n6256) );
  XNOR2_X1 U7834 ( .A(n6255), .B(n6256), .ZN(n8730) );
  INV_X1 U7835 ( .A(n6251), .ZN(n6252) );
  NOR2_X1 U7836 ( .A1(n6253), .A2(n6252), .ZN(n8729) );
  NOR2_X1 U7837 ( .A1(n8730), .A2(n8729), .ZN(n6254) );
  INV_X1 U7838 ( .A(n6255), .ZN(n6258) );
  INV_X1 U7839 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7840 ( .A1(n6258), .A2(n6257), .ZN(n6274) );
  NAND2_X1 U7841 ( .A1(n8734), .A2(n6274), .ZN(n6273) );
  OR2_X1 U7842 ( .A1(n8782), .A2(n10324), .ZN(n6259) );
  NAND2_X1 U7843 ( .A1(n9236), .A2(n6261), .ZN(n6268) );
  NAND2_X1 U7844 ( .A1(n8755), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6266) );
  NAND2_X1 U7845 ( .A1(n8757), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U7846 ( .A1(n8756), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7847 ( .A(P1_REG3_REG_27__SCAN_IN), .B(n6299), .ZN(n6316) );
  OR2_X1 U7848 ( .A1(n8635), .A2(n6316), .ZN(n6263) );
  NAND4_X1 U7849 ( .A1(n6266), .A2(n6265), .A3(n6264), .A4(n6263), .ZN(n9201)
         );
  NAND2_X1 U7850 ( .A1(n9201), .A2(n8625), .ZN(n6267) );
  NAND2_X1 U7851 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  XNOR2_X1 U7852 ( .A(n6269), .B(n8629), .ZN(n6272) );
  AND2_X1 U7853 ( .A1(n9201), .A2(n8626), .ZN(n6270) );
  AOI21_X1 U7854 ( .B1(n9236), .B2(n8625), .A(n6270), .ZN(n6271) );
  NAND2_X1 U7855 ( .A1(n6272), .A2(n6271), .ZN(n8643) );
  OAI21_X1 U7856 ( .B1(n6272), .B2(n6271), .A(n8643), .ZN(n6276) );
  INV_X1 U7857 ( .A(n6274), .ZN(n6275) );
  NOR2_X1 U7858 ( .A1(n6276), .A2(n6275), .ZN(n6277) );
  NOR4_X1 U7859 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U7860 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n6280) );
  NOR4_X1 U7861 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6279) );
  NOR4_X1 U7862 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6278) );
  NAND4_X1 U7863 ( .A1(n10306), .A2(n6280), .A3(n6279), .A4(n6278), .ZN(n6286)
         );
  NOR4_X1 U7864 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6284) );
  NOR4_X1 U7865 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6283) );
  NOR4_X1 U7866 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6282) );
  NOR4_X1 U7867 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6281) );
  NAND4_X1 U7868 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n6285)
         );
  NOR2_X1 U7869 ( .A1(n6286), .A2(n6285), .ZN(n6697) );
  NAND2_X1 U7870 ( .A1(n7602), .A2(P1_B_REG_SCAN_IN), .ZN(n6287) );
  MUX2_X1 U7871 ( .A(P1_B_REG_SCAN_IN), .B(n6287), .S(n7595), .Z(n6288) );
  NAND2_X1 U7872 ( .A1(n6288), .A2(n6289), .ZN(n6386) );
  INV_X1 U7873 ( .A(n6386), .ZN(n6291) );
  INV_X1 U7874 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6290) );
  INV_X1 U7875 ( .A(n6289), .ZN(n9576) );
  AND2_X1 U7876 ( .A1(n9576), .A2(n7595), .ZN(n6388) );
  AOI21_X1 U7877 ( .B1(n6291), .B2(n6290), .A(n6388), .ZN(n6903) );
  INV_X1 U7878 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6396) );
  AND2_X1 U7879 ( .A1(n9576), .A2(n7602), .ZN(n6394) );
  AOI21_X1 U7880 ( .B1(n6291), .B2(n6396), .A(n6394), .ZN(n6901) );
  OAI211_X1 U7881 ( .C1(n6697), .C2(n6386), .A(n6903), .B(n6901), .ZN(n6313)
         );
  NAND2_X1 U7882 ( .A1(n6292), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6294) );
  INV_X1 U7883 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6293) );
  XNOR2_X1 U7884 ( .A(n6294), .B(n6293), .ZN(n6390) );
  AND2_X1 U7885 ( .A1(n6320), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6295) );
  NOR2_X1 U7886 ( .A1(n7434), .A2(n4403), .ZN(n8785) );
  INV_X1 U7887 ( .A(n8785), .ZN(n6296) );
  AND2_X1 U7888 ( .A1(n6703), .A2(n6705), .ZN(n9495) );
  INV_X1 U7889 ( .A(n9495), .ZN(n9921) );
  NAND3_X1 U7890 ( .A1(n9004), .A2(n6296), .A3(n9921), .ZN(n6297) );
  INV_X1 U7891 ( .A(n5801), .ZN(n6636) );
  NAND2_X1 U7892 ( .A1(n8757), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6306) );
  NAND2_X1 U7893 ( .A1(n8755), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7894 ( .A1(n8756), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n6304) );
  NAND3_X1 U7895 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(P1_REG3_REG_27__SCAN_IN), 
        .A3(n6299), .ZN(n9205) );
  INV_X1 U7896 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7897 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(n6299), .ZN(n6300) );
  NAND2_X1 U7898 ( .A1(n6301), .A2(n6300), .ZN(n6302) );
  NAND2_X1 U7899 ( .A1(n9205), .A2(n6302), .ZN(n9221) );
  OR2_X1 U7900 ( .A1(n8635), .A2(n9221), .ZN(n6303) );
  NAND4_X1 U7901 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n9021)
         );
  AND2_X1 U7902 ( .A1(n9021), .A2(n9140), .ZN(n6307) );
  AOI21_X1 U7903 ( .B1(n9022), .B2(n9003), .A(n6307), .ZN(n9231) );
  INV_X1 U7904 ( .A(n9004), .ZN(n6389) );
  OR2_X1 U7905 ( .A1(n6389), .A2(n6705), .ZN(n6308) );
  INV_X1 U7906 ( .A(n9007), .ZN(n6708) );
  NAND2_X1 U7907 ( .A1(n6703), .A2(n6708), .ZN(n6908) );
  INV_X1 U7908 ( .A(n6908), .ZN(n6309) );
  NAND2_X1 U7909 ( .A1(n9004), .A2(n6309), .ZN(n6310) );
  OR2_X1 U7910 ( .A1(n6313), .A2(n6310), .ZN(n6311) );
  NAND2_X2 U7911 ( .A1(n6703), .A2(n9007), .ZN(n9410) );
  NOR2_X1 U7912 ( .A1(n9410), .A2(n9014), .ZN(n6701) );
  NAND2_X1 U7913 ( .A1(n6701), .A2(n9004), .ZN(n9413) );
  NAND2_X1 U7914 ( .A1(n6311), .A2(n9413), .ZN(n9716) );
  NAND2_X1 U7915 ( .A1(n9236), .A2(n9716), .ZN(n6318) );
  INV_X1 U7916 ( .A(n6701), .ZN(n6312) );
  NAND2_X1 U7917 ( .A1(n6313), .A2(n6312), .ZN(n6315) );
  NAND2_X1 U7918 ( .A1(n8785), .A2(n6705), .ZN(n6699) );
  AND3_X1 U7919 ( .A1(n6699), .A2(n6390), .A3(n6320), .ZN(n6314) );
  NAND2_X1 U7920 ( .A1(n6315), .A2(n6314), .ZN(n6571) );
  NAND2_X1 U7921 ( .A1(n6571), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9719) );
  INV_X1 U7922 ( .A(n9719), .ZN(n8737) );
  INV_X1 U7923 ( .A(n6316), .ZN(n9237) );
  AOI22_X1 U7924 ( .A1(n8737), .A2(n9237), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6317) );
  OAI211_X1 U7925 ( .C1(n9231), .C2(n9656), .A(n6318), .B(n6317), .ZN(n6319)
         );
  NOR2_X1 U7926 ( .A1(n6320), .A2(P1_U3086), .ZN(n6321) );
  INV_X1 U7927 ( .A(n6322), .ZN(n6412) );
  OAI21_X1 U7928 ( .B1(n6522), .B2(n8066), .A(n7508), .ZN(n6360) );
  NAND2_X1 U7929 ( .A1(n6360), .A2(n4497), .ZN(n6323) );
  NAND2_X1 U7930 ( .A1(n6323), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  MUX2_X1 U7931 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8253), .Z(n6329) );
  MUX2_X1 U7932 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8253), .Z(n6328) );
  MUX2_X1 U7933 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8253), .Z(n6327) );
  MUX2_X1 U7934 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8253), .Z(n6326) );
  MUX2_X1 U7935 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8253), .Z(n6325) );
  INV_X1 U7936 ( .A(n6347), .ZN(n6487) );
  XOR2_X1 U7937 ( .A(n6347), .B(n6325), .Z(n6472) );
  INV_X1 U7938 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6324) );
  INV_X1 U7939 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6566) );
  MUX2_X1 U7940 ( .A(n6324), .B(n6566), .S(n8253), .Z(n6490) );
  AND2_X1 U7941 ( .A1(n6490), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6492) );
  NOR2_X1 U7942 ( .A1(n6472), .A2(n6492), .ZN(n6471) );
  AOI21_X1 U7943 ( .B1(n6325), .B2(n6487), .A(n6471), .ZN(n6498) );
  XNOR2_X1 U7944 ( .A(n6326), .B(n6510), .ZN(n6499) );
  NOR2_X1 U7945 ( .A1(n6498), .A2(n6499), .ZN(n6497) );
  AOI21_X1 U7946 ( .B1(n6326), .B2(n6510), .A(n6497), .ZN(n6548) );
  XOR2_X1 U7947 ( .A(n6559), .B(n6327), .Z(n6547) );
  NAND2_X1 U7948 ( .A1(n6548), .A2(n6547), .ZN(n6546) );
  OAI21_X1 U7949 ( .B1(n6327), .B2(n6559), .A(n6546), .ZN(n6654) );
  XNOR2_X1 U7950 ( .A(n6328), .B(n6674), .ZN(n6655) );
  NOR2_X1 U7951 ( .A1(n6654), .A2(n6655), .ZN(n6653) );
  AOI21_X1 U7952 ( .B1(n6328), .B2(n6674), .A(n6653), .ZN(n6755) );
  XNOR2_X1 U7953 ( .A(n6329), .B(n6771), .ZN(n6756) );
  NOR2_X1 U7954 ( .A1(n6755), .A2(n6756), .ZN(n6754) );
  AOI21_X1 U7955 ( .B1(n6329), .B2(n6771), .A(n6754), .ZN(n6331) );
  MUX2_X1 U7956 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8253), .Z(n6977) );
  XOR2_X1 U7957 ( .A(n6980), .B(n6977), .Z(n6330) );
  NAND2_X1 U7958 ( .A1(n6331), .A2(n6330), .ZN(n6976) );
  OAI21_X1 U7959 ( .B1(n6331), .B2(n6330), .A(n6976), .ZN(n6332) );
  NAND2_X1 U7960 ( .A1(P2_U3893), .A2(n8087), .ZN(n8264) );
  AND2_X1 U7961 ( .A1(n6332), .A2(n8226), .ZN(n6369) );
  INV_X1 U7962 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6333) );
  NAND2_X1 U7963 ( .A1(n5051), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7964 ( .A1(n6347), .A2(n6334), .ZN(n6335) );
  NAND2_X1 U7965 ( .A1(n4496), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6336) );
  NAND2_X1 U7966 ( .A1(n6335), .A2(n6336), .ZN(n6475) );
  INV_X1 U7967 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6476) );
  OR2_X1 U7968 ( .A1(n6475), .A2(n6476), .ZN(n6473) );
  NAND2_X1 U7969 ( .A1(n6473), .A2(n6336), .ZN(n6505) );
  NAND2_X1 U7970 ( .A1(n6510), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6337) );
  NAND2_X1 U7971 ( .A1(n6504), .A2(n6337), .ZN(n6338) );
  INV_X1 U7972 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6808) );
  INV_X1 U7973 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6952) );
  XNOR2_X1 U7974 ( .A(n6674), .B(n6952), .ZN(n6658) );
  NAND2_X1 U7975 ( .A1(n6339), .A2(n6658), .ZN(n6660) );
  NAND2_X1 U7976 ( .A1(n6674), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6340) );
  INV_X1 U7977 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6764) );
  INV_X1 U7978 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10327) );
  MUX2_X1 U7979 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10327), .S(n6980), .Z(n6341)
         );
  INV_X1 U7980 ( .A(n6341), .ZN(n6343) );
  NAND3_X1 U7981 ( .A1(n6761), .A2(n6343), .A3(n6342), .ZN(n6345) );
  NOR2_X1 U7982 ( .A1(n8087), .A2(P2_U3151), .ZN(n8581) );
  AND2_X1 U7983 ( .A1(n6360), .A2(n8581), .ZN(n6493) );
  INV_X1 U7984 ( .A(n6493), .ZN(n6344) );
  OR2_X1 U7985 ( .A1(n6344), .A2(n8253), .ZN(n8270) );
  AOI21_X1 U7986 ( .B1(n6982), .B2(n6345), .A(n8270), .ZN(n6368) );
  INV_X1 U7987 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U7988 ( .A1(n5051), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6346) );
  NAND2_X1 U7989 ( .A1(n6347), .A2(n6346), .ZN(n6348) );
  NAND2_X1 U7990 ( .A1(n4496), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7991 ( .A1(n6348), .A2(n6349), .ZN(n6480) );
  INV_X1 U7992 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6692) );
  OR2_X1 U7993 ( .A1(n6480), .A2(n6692), .ZN(n6478) );
  NAND2_X1 U7994 ( .A1(n6478), .A2(n6349), .ZN(n6501) );
  NAND2_X1 U7995 ( .A1(n6510), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7996 ( .A1(n6500), .A2(n6350), .ZN(n6351) );
  NAND2_X1 U7997 ( .A1(n6351), .A2(n6559), .ZN(n6665) );
  OAI21_X1 U7998 ( .B1(n6351), .B2(n6559), .A(n6665), .ZN(n6553) );
  INV_X1 U7999 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10128) );
  NAND2_X1 U8000 ( .A1(n6667), .A2(n6665), .ZN(n6353) );
  INV_X1 U8001 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6352) );
  XNOR2_X1 U8002 ( .A(n6674), .B(n6352), .ZN(n6664) );
  NAND2_X1 U8003 ( .A1(n6674), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6354) );
  INV_X1 U8004 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10279) );
  NAND2_X1 U8005 ( .A1(n6758), .A2(n6357), .ZN(n6355) );
  INV_X1 U8006 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10000) );
  MUX2_X1 U8007 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10000), .S(n6980), .Z(n6356)
         );
  NAND3_X1 U8008 ( .A1(n6758), .A2(n4514), .A3(n6357), .ZN(n6358) );
  AND2_X1 U8009 ( .A1(n6493), .A2(n8253), .ZN(n8267) );
  AOI21_X1 U8010 ( .B1(n6973), .B2(n6358), .A(n8237), .ZN(n6367) );
  AND2_X1 U8011 ( .A1(n6522), .A2(n7508), .ZN(n6359) );
  OR2_X1 U8012 ( .A1(P2_U3150), .A2(n6359), .ZN(n8259) );
  INV_X1 U8013 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6365) );
  NOR2_X1 U8014 ( .A1(n8253), .A2(P2_U3151), .ZN(n8585) );
  AND2_X1 U8015 ( .A1(n6360), .A2(n8585), .ZN(n6361) );
  MUX2_X1 U8016 ( .A(P2_U3893), .B(n6361), .S(n8087), .Z(n8261) );
  INV_X1 U8017 ( .A(n6980), .ZN(n6362) );
  NAND2_X1 U8018 ( .A1(n8261), .A2(n6362), .ZN(n6364) );
  INV_X1 U8019 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6363) );
  OR2_X1 U8020 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6363), .ZN(n7827) );
  OAI211_X1 U8021 ( .C1(n8259), .C2(n6365), .A(n6364), .B(n7827), .ZN(n6366)
         );
  OR4_X1 U8022 ( .A1(n6369), .A2(n6368), .A3(n6367), .A4(n6366), .ZN(P2_U3188)
         );
  AND2_X1 U8023 ( .A1(n7868), .A2(P2_U3151), .ZN(n8586) );
  NOR2_X1 U8024 ( .A1(n7868), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8579) );
  OAI222_X1 U8025 ( .A1(n4406), .A2(n6370), .B1(n8588), .B2(n6398), .C1(
        P2_U3151), .C2(n6559), .ZN(P2_U3292) );
  NAND2_X1 U8026 ( .A1(n7868), .A2(P1_U3086), .ZN(n9575) );
  NOR2_X1 U8027 ( .A1(n7868), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9565) );
  AOI22_X1 U8028 ( .A1(n9059), .A2(P1_STATE_REG_SCAN_IN), .B1(n9565), .B2(
        P2_DATAO_REG_5__SCAN_IN), .ZN(n6371) );
  OAI21_X1 U8029 ( .B1(n6372), .B2(n9575), .A(n6371), .ZN(P1_U3350) );
  OAI222_X1 U8030 ( .A1(n4406), .A2(n6373), .B1(n8588), .B2(n6372), .C1(
        P2_U3151), .C2(n6771), .ZN(P2_U3290) );
  INV_X1 U8031 ( .A(n9565), .ZN(n9572) );
  OAI222_X1 U8032 ( .A1(n9572), .A2(n6374), .B1(n9575), .B2(n6380), .C1(
        P1_U3086), .C2(n6640), .ZN(P1_U3353) );
  OAI222_X1 U8033 ( .A1(n9572), .A2(n6375), .B1(n9575), .B2(n6378), .C1(
        P1_U3086), .C2(n9740), .ZN(P1_U3351) );
  OAI222_X1 U8034 ( .A1(n8588), .A2(n4811), .B1(n6487), .B2(P2_U3151), .C1(
        n6377), .C2(n4406), .ZN(P2_U3294) );
  OAI222_X1 U8035 ( .A1(n4406), .A2(n6379), .B1(n8588), .B2(n6378), .C1(
        P2_U3151), .C2(n6674), .ZN(P2_U3291) );
  OAI222_X1 U8036 ( .A1(n4406), .A2(n6381), .B1(n8588), .B2(n6380), .C1(
        P2_U3151), .C2(n6510), .ZN(P2_U3293) );
  INV_X1 U8037 ( .A(n9071), .ZN(n6382) );
  OAI222_X1 U8038 ( .A1(n9572), .A2(n6383), .B1(n9575), .B2(n6384), .C1(
        P1_U3086), .C2(n6382), .ZN(P1_U3349) );
  OAI222_X1 U8039 ( .A1(n4406), .A2(n6385), .B1(n8588), .B2(n6384), .C1(
        P2_U3151), .C2(n6980), .ZN(P2_U3289) );
  NAND2_X1 U8040 ( .A1(n9906), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6387) );
  OAI21_X1 U8041 ( .B1(n9906), .B2(n6388), .A(n6387), .ZN(P1_U3439) );
  OR2_X1 U8042 ( .A1(n6390), .A2(P1_U3086), .ZN(n9010) );
  NAND2_X1 U8043 ( .A1(n6389), .A2(n9010), .ZN(n6432) );
  NAND2_X1 U8044 ( .A1(n8785), .A2(n6390), .ZN(n6392) );
  AND2_X1 U8045 ( .A1(n6392), .A2(n6391), .ZN(n6431) );
  INV_X1 U8046 ( .A(n6431), .ZN(n6393) );
  AND2_X1 U8047 ( .A1(n6432), .A2(n6393), .ZN(n9728) );
  NOR2_X1 U8048 ( .A1(n9728), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8049 ( .A(n9906), .ZN(n9905) );
  OR2_X1 U8050 ( .A1(n9906), .A2(n6394), .ZN(n6395) );
  OAI21_X1 U8051 ( .B1(n9905), .B2(n6396), .A(n6395), .ZN(P1_U3440) );
  INV_X1 U8052 ( .A(n9575), .ZN(n7504) );
  INV_X1 U8053 ( .A(n7504), .ZN(n9571) );
  OAI222_X1 U8054 ( .A1(P1_U3086), .A2(n6433), .B1(n9571), .B2(n4811), .C1(
        n6397), .C2(n9572), .ZN(P1_U3354) );
  OAI222_X1 U8055 ( .A1(n9572), .A2(n6399), .B1(n9571), .B2(n6398), .C1(
        P1_U3086), .C2(n6438), .ZN(P1_U3352) );
  INV_X1 U8056 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10295) );
  INV_X1 U8057 ( .A(n6400), .ZN(n6402) );
  INV_X1 U8058 ( .A(n9083), .ZN(n6401) );
  OAI222_X1 U8059 ( .A1(n9572), .A2(n10295), .B1(n9575), .B2(n6402), .C1(
        P1_U3086), .C2(n6401), .ZN(P1_U3348) );
  INV_X1 U8060 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6403) );
  INV_X1 U8061 ( .A(n7025), .ZN(n6983) );
  OAI222_X1 U8062 ( .A1(n4406), .A2(n6403), .B1(n8588), .B2(n6402), .C1(
        P2_U3151), .C2(n6983), .ZN(P2_U3288) );
  INV_X1 U8063 ( .A(n6404), .ZN(n6405) );
  INV_X1 U8064 ( .A(n7151), .ZN(n7143) );
  OAI222_X1 U8065 ( .A1(n4406), .A2(n10294), .B1(n8588), .B2(n6405), .C1(
        P2_U3151), .C2(n7143), .ZN(P2_U3287) );
  INV_X1 U8066 ( .A(n6449), .ZN(n9601) );
  OAI222_X1 U8067 ( .A1(n9572), .A2(n6406), .B1(n9575), .B2(n6405), .C1(
        P1_U3086), .C2(n9601), .ZN(P1_U3347) );
  NAND2_X1 U8068 ( .A1(n6407), .A2(n5618), .ZN(n6458) );
  INV_X1 U8069 ( .A(n6408), .ZN(n6409) );
  AOI22_X1 U8070 ( .A1(n6458), .A2(n4769), .B1(n6412), .B2(n6409), .ZN(
        P2_U3376) );
  INV_X1 U8071 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6413) );
  INV_X1 U8072 ( .A(n6410), .ZN(n6411) );
  AOI22_X1 U8073 ( .A1(n6458), .A2(n6413), .B1(n6412), .B2(n6411), .ZN(
        P2_U3377) );
  AND2_X1 U8074 ( .A1(n6458), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8075 ( .A1(n6458), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8076 ( .A1(n6458), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8077 ( .A1(n6458), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8078 ( .A1(n6458), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8079 ( .A1(n6458), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8080 ( .A1(n6458), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8081 ( .A1(n6458), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8082 ( .A1(n6458), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8083 ( .A1(n6458), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8084 ( .A1(n6458), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8085 ( .A1(n6458), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8086 ( .A1(n6458), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8087 ( .A1(n6458), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8088 ( .A1(n6458), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8089 ( .A1(n6458), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8090 ( .A1(n6458), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8091 ( .A1(n6458), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8092 ( .A1(n6458), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8093 ( .A1(n6458), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8094 ( .A1(n6458), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8095 ( .A1(n6458), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8096 ( .A1(n6458), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8097 ( .A1(n6458), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8098 ( .A1(n6458), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  XNOR2_X1 U8099 ( .A(n9107), .B(P1_REG2_REG_9__SCAN_IN), .ZN(n6430) );
  INV_X1 U8100 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6414) );
  MUX2_X1 U8101 ( .A(n6414), .B(P1_REG2_REG_1__SCAN_IN), .S(n6433), .Z(n9040)
         );
  AND2_X1 U8102 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9039) );
  NAND2_X1 U8103 ( .A1(n9040), .A2(n9039), .ZN(n9038) );
  NAND2_X1 U8104 ( .A1(n5804), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8105 ( .A1(n9038), .A2(n6415), .ZN(n6645) );
  XNOR2_X1 U8106 ( .A(n6640), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8107 ( .A1(n6645), .A2(n6646), .ZN(n6644) );
  INV_X1 U8108 ( .A(n6640), .ZN(n6436) );
  NAND2_X1 U8109 ( .A1(n6436), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8110 ( .A1(n6644), .A2(n6416), .ZN(n9050) );
  XNOR2_X1 U8111 ( .A(n6438), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9051) );
  NAND2_X1 U8112 ( .A1(n9050), .A2(n9051), .ZN(n9049) );
  INV_X1 U8113 ( .A(n6438), .ZN(n9048) );
  NAND2_X1 U8114 ( .A1(n9048), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8115 ( .A1(n9049), .A2(n6417), .ZN(n9736) );
  INV_X1 U8116 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6418) );
  MUX2_X1 U8117 ( .A(n6418), .B(P1_REG2_REG_4__SCAN_IN), .S(n9740), .Z(n9737)
         );
  NAND2_X1 U8118 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  INV_X1 U8119 ( .A(n9740), .ZN(n6441) );
  NAND2_X1 U8120 ( .A1(n6441), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8121 ( .A1(n9735), .A2(n6419), .ZN(n9061) );
  INV_X1 U8122 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6420) );
  XNOR2_X1 U8123 ( .A(n9059), .B(n6420), .ZN(n9062) );
  NAND2_X1 U8124 ( .A1(n9061), .A2(n9062), .ZN(n9060) );
  NAND2_X1 U8125 ( .A1(n9059), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U8126 ( .A1(n9060), .A2(n6421), .ZN(n9076) );
  INV_X1 U8127 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6422) );
  MUX2_X1 U8128 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6422), .S(n9071), .Z(n9077)
         );
  NAND2_X1 U8129 ( .A1(n9076), .A2(n9077), .ZN(n9075) );
  NAND2_X1 U8130 ( .A1(n9071), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8131 ( .A1(n9075), .A2(n6423), .ZN(n9088) );
  INV_X1 U8132 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6424) );
  XNOR2_X1 U8133 ( .A(n9083), .B(n6424), .ZN(n9089) );
  NAND2_X1 U8134 ( .A1(n9088), .A2(n9089), .ZN(n9087) );
  NAND2_X1 U8135 ( .A1(n9083), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6425) );
  NAND2_X1 U8136 ( .A1(n9087), .A2(n6425), .ZN(n9597) );
  INV_X1 U8137 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6426) );
  XNOR2_X1 U8138 ( .A(n6449), .B(n6426), .ZN(n9598) );
  NAND2_X1 U8139 ( .A1(n9597), .A2(n9598), .ZN(n9596) );
  NAND2_X1 U8140 ( .A1(n6449), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6427) );
  NAND2_X1 U8141 ( .A1(n9596), .A2(n6427), .ZN(n6429) );
  INV_X1 U8142 ( .A(n9095), .ZN(n6428) );
  AOI21_X1 U8143 ( .B1(n6430), .B2(n6429), .A(n6428), .ZN(n6457) );
  NAND2_X1 U8144 ( .A1(n6432), .A2(n6431), .ZN(n9731) );
  OR3_X1 U8145 ( .A1(n9731), .A2(n5801), .A3(n9721), .ZN(n9816) );
  OR2_X1 U8146 ( .A1(n9731), .A2(n6636), .ZN(n9848) );
  INV_X1 U8147 ( .A(n9848), .ZN(n9830) );
  INV_X1 U8148 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10335) );
  NAND2_X1 U8149 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n7228) );
  OAI21_X1 U8150 ( .B1(n9852), .B2(n10335), .A(n7228), .ZN(n6455) );
  INV_X1 U8151 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6434) );
  MUX2_X1 U8152 ( .A(n6434), .B(P1_REG1_REG_1__SCAN_IN), .S(n6433), .Z(n9037)
         );
  AND2_X1 U8153 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9036) );
  NAND2_X1 U8154 ( .A1(n9037), .A2(n9036), .ZN(n9035) );
  NAND2_X1 U8155 ( .A1(n5804), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U8156 ( .A1(n9035), .A2(n6435), .ZN(n6642) );
  XNOR2_X1 U8157 ( .A(n6640), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8158 ( .A1(n6642), .A2(n6643), .ZN(n6641) );
  NAND2_X1 U8159 ( .A1(n6436), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8160 ( .A1(n6641), .A2(n6437), .ZN(n9053) );
  XNOR2_X1 U8161 ( .A(n6438), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9054) );
  NAND2_X1 U8162 ( .A1(n9053), .A2(n9054), .ZN(n9052) );
  NAND2_X1 U8163 ( .A1(n9048), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6439) );
  NAND2_X1 U8164 ( .A1(n9052), .A2(n6439), .ZN(n9733) );
  INV_X1 U8165 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6440) );
  MUX2_X1 U8166 ( .A(n6440), .B(P1_REG1_REG_4__SCAN_IN), .S(n9740), .Z(n9734)
         );
  NAND2_X1 U8167 ( .A1(n9733), .A2(n9734), .ZN(n9732) );
  NAND2_X1 U8168 ( .A1(n6441), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8169 ( .A1(n9732), .A2(n6442), .ZN(n9064) );
  INV_X1 U8170 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6443) );
  XNOR2_X1 U8171 ( .A(n9059), .B(n6443), .ZN(n9065) );
  NAND2_X1 U8172 ( .A1(n9064), .A2(n9065), .ZN(n9063) );
  NAND2_X1 U8173 ( .A1(n9059), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6444) );
  NAND2_X1 U8174 ( .A1(n9063), .A2(n6444), .ZN(n9073) );
  INV_X1 U8175 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10284) );
  MUX2_X1 U8176 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10284), .S(n9071), .Z(n9074)
         );
  NAND2_X1 U8177 ( .A1(n9073), .A2(n9074), .ZN(n9072) );
  NAND2_X1 U8178 ( .A1(n9071), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U8179 ( .A1(n9072), .A2(n6445), .ZN(n9085) );
  INV_X1 U8180 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6446) );
  XNOR2_X1 U8181 ( .A(n9083), .B(n6446), .ZN(n9086) );
  NAND2_X1 U8182 ( .A1(n9085), .A2(n9086), .ZN(n9084) );
  NAND2_X1 U8183 ( .A1(n9083), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8184 ( .A1(n9084), .A2(n6447), .ZN(n9594) );
  INV_X1 U8185 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6448) );
  XNOR2_X1 U8186 ( .A(n6449), .B(n6448), .ZN(n9595) );
  NAND2_X1 U8187 ( .A1(n9594), .A2(n9595), .ZN(n9593) );
  NAND2_X1 U8188 ( .A1(n6449), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U8189 ( .A1(n9593), .A2(n6450), .ZN(n6452) );
  MUX2_X1 U8190 ( .A(n5948), .B(P1_REG1_REG_9__SCAN_IN), .S(n9107), .Z(n6451)
         );
  OR2_X1 U8191 ( .A1(n6452), .A2(n6451), .ZN(n9109) );
  NAND2_X1 U8192 ( .A1(n6452), .A2(n6451), .ZN(n6453) );
  OR2_X1 U8193 ( .A1(n9731), .A2(n9138), .ZN(n9812) );
  AOI21_X1 U8194 ( .B1(n9109), .B2(n6453), .A(n9812), .ZN(n6454) );
  AOI211_X1 U8195 ( .C1(n9830), .C2(n9107), .A(n6455), .B(n6454), .ZN(n6456)
         );
  OAI21_X1 U8196 ( .B1(n6457), .B2(n9816), .A(n6456), .ZN(P1_U3252) );
  INV_X1 U8197 ( .A(n6458), .ZN(n6459) );
  INV_X1 U8198 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10138) );
  NOR2_X1 U8199 ( .A1(n6459), .A2(n10138), .ZN(P2_U3249) );
  INV_X1 U8200 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10175) );
  NOR2_X1 U8201 ( .A1(n6459), .A2(n10175), .ZN(P2_U3263) );
  INV_X1 U8202 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U8203 ( .A1(n6459), .A2(n10189), .ZN(P2_U3251) );
  INV_X1 U8204 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U8205 ( .A1(n6459), .A2(n10050), .ZN(P2_U3262) );
  INV_X1 U8206 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10118) );
  NOR2_X1 U8207 ( .A1(n6459), .A2(n10118), .ZN(P2_U3235) );
  INV_X1 U8208 ( .A(n6460), .ZN(n6462) );
  INV_X1 U8209 ( .A(n9107), .ZN(n6461) );
  OAI222_X1 U8210 ( .A1(n9572), .A2(n10281), .B1(n9571), .B2(n6462), .C1(
        P1_U3086), .C2(n6461), .ZN(P1_U3346) );
  INV_X1 U8211 ( .A(n7158), .ZN(n7249) );
  OAI222_X1 U8212 ( .A1(n4406), .A2(n6463), .B1(n8588), .B2(n6462), .C1(
        P2_U3151), .C2(n7249), .ZN(P2_U3286) );
  INV_X1 U8213 ( .A(n6464), .ZN(n6466) );
  INV_X1 U8214 ( .A(n7248), .ZN(n7443) );
  OAI222_X1 U8215 ( .A1(n8588), .A2(n6466), .B1(n7443), .B2(P2_U3151), .C1(
        n6465), .C2(n4406), .ZN(P2_U3285) );
  INV_X1 U8216 ( .A(n9111), .ZN(n9588) );
  OAI222_X1 U8217 ( .A1(n9572), .A2(n10300), .B1(n9571), .B2(n6466), .C1(n9588), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U8218 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U8219 ( .A1(n6687), .A2(P2_U3893), .ZN(n6467) );
  OAI21_X1 U8220 ( .B1(P2_U3893), .B2(n6468), .A(n6467), .ZN(P2_U3491) );
  INV_X1 U8221 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8222 ( .A1(n6822), .A2(P1_U3973), .ZN(n6469) );
  OAI21_X1 U8223 ( .B1(P1_U3973), .B2(n6470), .A(n6469), .ZN(P1_U3554) );
  INV_X1 U8224 ( .A(n8261), .ZN(n8224) );
  AOI211_X1 U8225 ( .C1(n6472), .C2(n6492), .A(n8264), .B(n6471), .ZN(n6485)
         );
  INV_X1 U8226 ( .A(n6473), .ZN(n6474) );
  AOI21_X1 U8227 ( .B1(n6476), .B2(n6475), .A(n6474), .ZN(n6477) );
  OAI22_X1 U8228 ( .A1(n8270), .A2(n6477), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6608), .ZN(n6484) );
  INV_X1 U8229 ( .A(n6478), .ZN(n6479) );
  AOI21_X1 U8230 ( .B1(n6692), .B2(n6480), .A(n6479), .ZN(n6482) );
  INV_X1 U8231 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6481) );
  OAI22_X1 U8232 ( .A1(n8237), .A2(n6482), .B1(n8259), .B2(n6481), .ZN(n6483)
         );
  NOR3_X1 U8233 ( .A1(n6485), .A2(n6484), .A3(n6483), .ZN(n6486) );
  OAI21_X1 U8234 ( .B1(n6487), .B2(n8224), .A(n6486), .ZN(P2_U3183) );
  INV_X1 U8235 ( .A(n6488), .ZN(n6518) );
  AOI22_X1 U8236 ( .A1(n7490), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n8586), .ZN(n6489) );
  OAI21_X1 U8237 ( .B1(n6518), .B2(n8588), .A(n6489), .ZN(P2_U3284) );
  INV_X1 U8238 ( .A(n8259), .ZN(n7038) );
  NOR2_X1 U8239 ( .A1(n6490), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6491) );
  OAI22_X1 U8240 ( .A1(n8226), .A2(n6493), .B1(n6492), .B2(n6491), .ZN(n6494)
         );
  OAI21_X1 U8241 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5043), .A(n6494), .ZN(n6495) );
  AOI21_X1 U8242 ( .B1(n7038), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6495), .ZN(
        n6496) );
  OAI21_X1 U8243 ( .B1(n5051), .B2(n8224), .A(n6496), .ZN(P2_U3182) );
  AOI211_X1 U8244 ( .C1(n6499), .C2(n6498), .A(n8264), .B(n6497), .ZN(n6512)
         );
  OAI21_X1 U8245 ( .B1(n6502), .B2(n6501), .A(n6500), .ZN(n6503) );
  AOI22_X1 U8246 ( .A1(n7038), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(n8267), .B2(
        n6503), .ZN(n6509) );
  OAI21_X1 U8247 ( .B1(n6506), .B2(n6505), .A(n6504), .ZN(n6507) );
  INV_X1 U8248 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6783) );
  AOI22_X1 U8249 ( .A1(n4594), .A2(n6507), .B1(P2_U3151), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6508) );
  OAI211_X1 U8250 ( .C1(n6510), .C2(n8224), .A(n6509), .B(n6508), .ZN(n6511)
         );
  OR2_X1 U8251 ( .A1(n6512), .A2(n6511), .ZN(P2_U3184) );
  NAND2_X1 U8252 ( .A1(n8755), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6515) );
  NAND2_X1 U8253 ( .A1(n8756), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6514) );
  NAND2_X1 U8254 ( .A1(n8757), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6513) );
  NAND3_X1 U8255 ( .A1(n6515), .A2(n6514), .A3(n6513), .ZN(n9142) );
  NAND2_X1 U8256 ( .A1(n9142), .A2(P1_U3973), .ZN(n6516) );
  OAI21_X1 U8257 ( .B1(P1_U3973), .B2(n8575), .A(n6516), .ZN(P1_U3585) );
  INV_X1 U8258 ( .A(n9754), .ZN(n6517) );
  OAI222_X1 U8259 ( .A1(n9572), .A2(n10259), .B1(n9571), .B2(n6518), .C1(
        P1_U3086), .C2(n6517), .ZN(P1_U3344) );
  INV_X1 U8260 ( .A(n6519), .ZN(n6520) );
  OR2_X1 U8261 ( .A1(n6521), .A2(n6520), .ZN(n6527) );
  INV_X1 U8262 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U8263 ( .A1(n6523), .A2(n7508), .ZN(n6525) );
  NOR2_X1 U8264 ( .A1(n6525), .A2(n6524), .ZN(n6526) );
  OAI211_X1 U8265 ( .C1(n6529), .C2(n6534), .A(n6527), .B(n6526), .ZN(n6528)
         );
  NAND2_X1 U8266 ( .A1(n6528), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6533) );
  INV_X1 U8267 ( .A(n6529), .ZN(n6531) );
  NOR2_X1 U8268 ( .A1(n6530), .A2(n6541), .ZN(n8089) );
  NAND2_X1 U8269 ( .A1(n6531), .A2(n8089), .ZN(n6532) );
  NAND2_X1 U8270 ( .A1(n6533), .A2(n6532), .ZN(n7851) );
  NOR2_X1 U8271 ( .A1(n7851), .A2(P2_U3151), .ZN(n6621) );
  INV_X1 U8272 ( .A(n6601), .ZN(n6593) );
  NAND2_X1 U8273 ( .A1(n6687), .A2(n6593), .ZN(n7915) );
  NAND2_X1 U8274 ( .A1(n7915), .A2(n7917), .ZN(n7885) );
  INV_X1 U8275 ( .A(n6534), .ZN(n6535) );
  NAND2_X1 U8276 ( .A1(n6543), .A2(n6535), .ZN(n6538) );
  OR2_X1 U8277 ( .A1(n6539), .A2(n6536), .ZN(n6537) );
  OR2_X1 U8278 ( .A1(n6539), .A2(n8331), .ZN(n6540) );
  NAND2_X1 U8279 ( .A1(n6540), .A2(n9632), .ZN(n7861) );
  AOI22_X1 U8280 ( .A1(n7885), .A2(n7839), .B1(n6601), .B2(n7861), .ZN(n6545)
         );
  INV_X1 U8281 ( .A(n6541), .ZN(n6542) );
  AND2_X1 U8282 ( .A1(n6543), .A2(n6542), .ZN(n6604) );
  NAND2_X1 U8283 ( .A1(n7826), .A2(n8113), .ZN(n6544) );
  OAI211_X1 U8284 ( .C1(n6621), .C2(n5043), .A(n6545), .B(n6544), .ZN(P2_U3172) );
  OAI21_X1 U8285 ( .B1(n6548), .B2(n6547), .A(n6546), .ZN(n6549) );
  NAND2_X1 U8286 ( .A1(n6549), .A2(n8226), .ZN(n6558) );
  INV_X1 U8287 ( .A(n6661), .ZN(n6550) );
  AOI21_X1 U8288 ( .B1(n6808), .B2(n6551), .A(n6550), .ZN(n6552) );
  NAND2_X1 U8289 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6744) );
  OAI21_X1 U8290 ( .B1(n8270), .B2(n6552), .A(n6744), .ZN(n6556) );
  NAND2_X1 U8291 ( .A1(n6553), .A2(n10128), .ZN(n6554) );
  AOI21_X1 U8292 ( .B1(n6667), .B2(n6554), .A(n8237), .ZN(n6555) );
  AOI211_X1 U8293 ( .C1(n7038), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6556), .B(
        n6555), .ZN(n6557) );
  OAI211_X1 U8294 ( .C1(n8224), .C2(n6559), .A(n6558), .B(n6557), .ZN(P2_U3185) );
  NOR2_X1 U8295 ( .A1(n9632), .A2(n5043), .ZN(n6560) );
  NOR2_X1 U8296 ( .A1(n6779), .A2(n9642), .ZN(n6564) );
  AOI211_X1 U8297 ( .C1(n6561), .C2(n7885), .A(n6560), .B(n6564), .ZN(n6563)
         );
  AOI22_X1 U8298 ( .A1(n8444), .A2(n6601), .B1(n9648), .B2(
        P2_REG2_REG_0__SCAN_IN), .ZN(n6562) );
  OAI21_X1 U8299 ( .B1(n6563), .B2(n9648), .A(n6562), .ZN(P2_U3233) );
  INV_X1 U8300 ( .A(n9968), .ZN(n9986) );
  NAND2_X1 U8301 ( .A1(n9986), .A2(n9637), .ZN(n6565) );
  AOI21_X1 U8302 ( .B1(n7885), .B2(n6565), .A(n6564), .ZN(n6591) );
  OAI22_X1 U8303 ( .A1(n8460), .A2(n6593), .B1(n10012), .B2(n6566), .ZN(n6567)
         );
  INV_X1 U8304 ( .A(n6567), .ZN(n6568) );
  OAI21_X1 U8305 ( .B1(n6591), .B2(n10010), .A(n6568), .ZN(P2_U3459) );
  INV_X1 U8306 ( .A(n6569), .ZN(n6579) );
  INV_X1 U8307 ( .A(n7542), .ZN(n7493) );
  INV_X1 U8308 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6570) );
  OAI222_X1 U8309 ( .A1(n8588), .A2(n6579), .B1(n7493), .B2(P2_U3151), .C1(
        n6570), .C2(n4406), .ZN(P2_U3283) );
  NOR2_X1 U8310 ( .A1(n6571), .A2(P1_U3086), .ZN(n6632) );
  INV_X1 U8311 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6909) );
  OAI21_X1 U8312 ( .B1(n6572), .B2(n6574), .A(n6573), .ZN(n6575) );
  NAND2_X1 U8313 ( .A1(n6575), .A2(n6298), .ZN(n6578) );
  INV_X1 U8314 ( .A(n9034), .ZN(n6677) );
  INV_X1 U8315 ( .A(n9140), .ZN(n9667) );
  INV_X1 U8316 ( .A(n6822), .ZN(n6576) );
  INV_X1 U8317 ( .A(n9003), .ZN(n9669) );
  OAI22_X1 U8318 ( .A1(n6677), .A2(n9667), .B1(n6576), .B2(n9669), .ZN(n6868)
         );
  AOI22_X1 U8319 ( .A1(n6868), .A2(n9713), .B1(n6957), .B2(n9716), .ZN(n6577)
         );
  OAI211_X1 U8320 ( .C1(n6632), .C2(n6909), .A(n6578), .B(n6577), .ZN(P1_U3222) );
  INV_X1 U8321 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10241) );
  INV_X1 U8322 ( .A(n9113), .ZN(n9767) );
  OAI222_X1 U8323 ( .A1(n9572), .A2(n10241), .B1(n9571), .B2(n6579), .C1(n9767), .C2(P1_U3086), .ZN(P1_U3343) );
  OR2_X1 U8324 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  NAND2_X1 U8325 ( .A1(n6583), .A2(n6582), .ZN(n6633) );
  INV_X1 U8326 ( .A(n6632), .ZN(n6585) );
  NAND2_X1 U8327 ( .A1(n5813), .A2(n9140), .ZN(n6915) );
  INV_X1 U8328 ( .A(n9716), .ZN(n9703) );
  INV_X1 U8329 ( .A(n6862), .ZN(n6922) );
  OAI22_X1 U8330 ( .A1(n6915), .A2(n9656), .B1(n9703), .B2(n6922), .ZN(n6584)
         );
  AOI21_X1 U8331 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n6585), .A(n6584), .ZN(
        n6586) );
  OAI21_X1 U8332 ( .B1(n6633), .B2(n9660), .A(n6586), .ZN(P1_U3232) );
  INV_X1 U8333 ( .A(n6587), .ZN(n6590) );
  AOI22_X1 U8334 ( .A1(n9781), .A2(P1_STATE_REG_SCAN_IN), .B1(n9565), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6588) );
  OAI21_X1 U8335 ( .B1(n6590), .B2(n9575), .A(n6588), .ZN(P1_U3342) );
  AOI22_X1 U8336 ( .A1(n8132), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n8586), .ZN(n6589) );
  OAI21_X1 U8337 ( .B1(n6590), .B2(n8588), .A(n6589), .ZN(P2_U3282) );
  INV_X1 U8338 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10308) );
  MUX2_X1 U8339 ( .A(n10308), .B(n6591), .S(n9993), .Z(n6592) );
  OAI21_X1 U8340 ( .B1(n6593), .B2(n8516), .A(n6592), .ZN(P2_U3390) );
  INV_X1 U8341 ( .A(n6594), .ZN(n6595) );
  NAND2_X1 U8342 ( .A1(n6596), .A2(n6595), .ZN(n6600) );
  AOI21_X2 U8343 ( .B1(n6598), .B2(n8084), .A(n6597), .ZN(n6599) );
  XNOR2_X1 U8344 ( .A(n6617), .B(n6779), .ZN(n6616) );
  XOR2_X1 U8345 ( .A(n6615), .B(n6616), .Z(n6612) );
  INV_X1 U8346 ( .A(n6604), .ZN(n6606) );
  OAI22_X1 U8347 ( .A1(n7848), .A2(n6693), .B1(n7841), .B2(n6607), .ZN(n6610)
         );
  NOR2_X1 U8348 ( .A1(n6621), .A2(n6608), .ZN(n6609) );
  AOI211_X1 U8349 ( .C1(n7826), .C2(n8112), .A(n6610), .B(n6609), .ZN(n6611)
         );
  OAI21_X1 U8350 ( .B1(n7856), .B2(n6612), .A(n6611), .ZN(P2_U3162) );
  XNOR2_X1 U8351 ( .A(n6723), .B(n8112), .ZN(n6721) );
  NAND2_X1 U8352 ( .A1(n6616), .A2(n6615), .ZN(n6620) );
  INV_X1 U8353 ( .A(n6617), .ZN(n6618) );
  NAND2_X1 U8354 ( .A1(n6779), .A2(n6618), .ZN(n6619) );
  XOR2_X1 U8355 ( .A(n6722), .B(n6721), .Z(n6625) );
  OAI22_X1 U8356 ( .A1(n7848), .A2(n5071), .B1(n7841), .B2(n6779), .ZN(n6623)
         );
  NOR2_X1 U8357 ( .A1(n6621), .A2(n6783), .ZN(n6622) );
  AOI211_X1 U8358 ( .C1(n7826), .C2(n8111), .A(n6623), .B(n6622), .ZN(n6624)
         );
  OAI21_X1 U8359 ( .B1(n7856), .B2(n6625), .A(n6624), .ZN(P2_U3177) );
  XNOR2_X1 U8360 ( .A(n6626), .B(n6627), .ZN(n6628) );
  NAND2_X1 U8361 ( .A1(n6628), .A2(n6298), .ZN(n6630) );
  INV_X1 U8362 ( .A(n5813), .ZN(n6828) );
  INV_X1 U8363 ( .A(n10048), .ZN(n6825) );
  OAI22_X1 U8364 ( .A1(n6828), .A2(n9669), .B1(n6825), .B2(n9667), .ZN(n6848)
         );
  AOI22_X1 U8365 ( .A1(n6848), .A2(n9713), .B1(n7047), .B2(n9716), .ZN(n6629)
         );
  OAI211_X1 U8366 ( .C1(n6632), .C2(n6631), .A(n6630), .B(n6629), .ZN(P1_U3237) );
  MUX2_X1 U8367 ( .A(n6633), .B(n9039), .S(n9138), .Z(n6637) );
  NOR2_X1 U8368 ( .A1(n9721), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6634) );
  OR2_X1 U8369 ( .A1(n6634), .A2(n5801), .ZN(n9720) );
  INV_X1 U8370 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U8371 ( .A1(n9720), .A2(n9723), .ZN(n9726) );
  NAND2_X1 U8372 ( .A1(P1_U3973), .A2(n9726), .ZN(n6635) );
  AOI21_X1 U8373 ( .B1(n6637), .B2(n6636), .A(n6635), .ZN(n9742) );
  NAND2_X1 U8374 ( .A1(n9728), .A2(P1_ADDR_REG_2__SCAN_IN), .ZN(n6639) );
  NAND2_X1 U8375 ( .A1(P1_U3086), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6638) );
  OAI211_X1 U8376 ( .C1(n9848), .C2(n6640), .A(n6639), .B(n6638), .ZN(n6650)
         );
  OAI21_X1 U8377 ( .B1(n6643), .B2(n6642), .A(n6641), .ZN(n6648) );
  OAI21_X1 U8378 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6647) );
  OAI22_X1 U8379 ( .A1(n9812), .A2(n6648), .B1(n9816), .B2(n6647), .ZN(n6649)
         );
  OR3_X1 U8380 ( .A1(n9742), .A2(n6650), .A3(n6649), .ZN(P1_U3245) );
  INV_X1 U8381 ( .A(n6651), .ZN(n6681) );
  AOI22_X1 U8382 ( .A1(n9794), .A2(P1_STATE_REG_SCAN_IN), .B1(n9565), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n6652) );
  OAI21_X1 U8383 ( .B1(n6681), .B2(n9575), .A(n6652), .ZN(P1_U3341) );
  AOI211_X1 U8384 ( .C1(n6655), .C2(n6654), .A(n8264), .B(n6653), .ZN(n6656)
         );
  INV_X1 U8385 ( .A(n6656), .ZN(n6673) );
  INV_X1 U8386 ( .A(n6657), .ZN(n6659) );
  NOR2_X1 U8387 ( .A1(n6659), .A2(n6658), .ZN(n6662) );
  AOI21_X1 U8388 ( .B1(n6662), .B2(n6661), .A(n4577), .ZN(n6663) );
  NAND2_X1 U8389 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6736) );
  OAI21_X1 U8390 ( .B1(n8270), .B2(n6663), .A(n6736), .ZN(n6671) );
  INV_X1 U8391 ( .A(n6664), .ZN(n6666) );
  NAND3_X1 U8392 ( .A1(n6667), .A2(n6666), .A3(n6665), .ZN(n6668) );
  AOI21_X1 U8393 ( .B1(n6669), .B2(n6668), .A(n8237), .ZN(n6670) );
  AOI211_X1 U8394 ( .C1(n7038), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6671), .B(
        n6670), .ZN(n6672) );
  OAI211_X1 U8395 ( .C1(n8224), .C2(n6674), .A(n6673), .B(n6672), .ZN(P2_U3186) );
  XOR2_X1 U8396 ( .A(n6675), .B(n6676), .Z(n6680) );
  INV_X1 U8397 ( .A(n9033), .ZN(n6887) );
  OAI22_X1 U8398 ( .A1(n6887), .A2(n9667), .B1(n6677), .B2(n9669), .ZN(n6831)
         );
  AOI22_X1 U8399 ( .A1(n6831), .A2(n9713), .B1(n6878), .B2(n9716), .ZN(n6679)
         );
  MUX2_X1 U8400 ( .A(n9719), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n6678) );
  OAI211_X1 U8401 ( .C1(n6680), .C2(n9660), .A(n6679), .B(n6678), .ZN(P1_U3218) );
  INV_X1 U8402 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6682) );
  INV_X1 U8403 ( .A(n8136), .ZN(n8158) );
  OAI222_X1 U8404 ( .A1(n4406), .A2(n6682), .B1(n8588), .B2(n6681), .C1(
        P2_U3151), .C2(n8158), .ZN(P2_U3281) );
  INV_X1 U8405 ( .A(n6683), .ZN(n6684) );
  AOI21_X1 U8406 ( .B1(n7913), .B2(n7917), .A(n6684), .ZN(n6801) );
  OAI21_X1 U8407 ( .B1(n6686), .B2(n7913), .A(n6685), .ZN(n6688) );
  AOI222_X1 U8408 ( .A1(n8391), .A2(n6688), .B1(n8112), .B2(n8386), .C1(n6687), 
        .C2(n8388), .ZN(n6797) );
  OAI21_X1 U8409 ( .B1(n9986), .B2(n6801), .A(n6797), .ZN(n6695) );
  INV_X1 U8410 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6689) );
  OAI22_X1 U8411 ( .A1(n6693), .A2(n8516), .B1(n9993), .B2(n6689), .ZN(n6690)
         );
  AOI21_X1 U8412 ( .B1(n6695), .B2(n9993), .A(n6690), .ZN(n6691) );
  INV_X1 U8413 ( .A(n6691), .ZN(P2_U3393) );
  OAI22_X1 U8414 ( .A1(n8460), .A2(n6693), .B1(n10012), .B2(n6692), .ZN(n6694)
         );
  AOI21_X1 U8415 ( .B1(n6695), .B2(n10012), .A(n6694), .ZN(n6696) );
  INV_X1 U8416 ( .A(n6696), .ZN(P2_U3460) );
  NAND2_X1 U8417 ( .A1(n9004), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8418 ( .A1(n9906), .A2(n6698), .ZN(n6700) );
  NAND2_X1 U8419 ( .A1(n6700), .A2(n6699), .ZN(n6904) );
  INV_X1 U8420 ( .A(n6903), .ZN(n6702) );
  INV_X2 U8421 ( .A(n9929), .ZN(n9932) );
  INV_X1 U8422 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10073) );
  INV_X1 U8423 ( .A(n6703), .ZN(n6712) );
  NAND2_X1 U8424 ( .A1(n8785), .A2(n9002), .ZN(n6704) );
  AND2_X1 U8425 ( .A1(n6704), .A2(n6712), .ZN(n6917) );
  NAND2_X1 U8426 ( .A1(n6706), .A2(n6705), .ZN(n6707) );
  NAND2_X1 U8427 ( .A1(n6917), .A2(n6707), .ZN(n7093) );
  AND2_X1 U8428 ( .A1(n9131), .A2(n7434), .ZN(n8934) );
  NAND2_X1 U8429 ( .A1(n8934), .A2(n9007), .ZN(n7272) );
  NAND2_X1 U8430 ( .A1(n7093), .A2(n7272), .ZN(n9924) );
  NAND2_X1 U8431 ( .A1(n9009), .A2(n9131), .ZN(n6710) );
  NAND2_X1 U8432 ( .A1(n8943), .A2(n6708), .ZN(n6709) );
  NOR2_X1 U8433 ( .A1(n6822), .A2(n6922), .ZN(n6863) );
  AND2_X1 U8434 ( .A1(n6822), .A2(n6922), .ZN(n8941) );
  NOR2_X1 U8435 ( .A1(n6863), .A2(n8941), .ZN(n8793) );
  INV_X1 U8436 ( .A(n8793), .ZN(n6918) );
  OAI21_X1 U8437 ( .B1(n9924), .B2(n9402), .A(n6918), .ZN(n6711) );
  OAI211_X1 U8438 ( .C1(n6712), .C2(n6922), .A(n6711), .B(n6915), .ZN(n6715)
         );
  NAND2_X1 U8439 ( .A1(n6715), .A2(n9932), .ZN(n6713) );
  OAI21_X1 U8440 ( .B1(n9932), .B2(n10073), .A(n6713), .ZN(P1_U3522) );
  INV_X2 U8441 ( .A(n9557), .ZN(n9927) );
  INV_X1 U8442 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6717) );
  NAND2_X1 U8443 ( .A1(n6715), .A2(n9927), .ZN(n6716) );
  OAI21_X1 U8444 ( .B1(n9927), .B2(n6717), .A(n6716), .ZN(P1_U3453) );
  INV_X1 U8445 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6719) );
  INV_X1 U8446 ( .A(n6718), .ZN(n6720) );
  INV_X1 U8447 ( .A(n9806), .ZN(n9119) );
  OAI222_X1 U8448 ( .A1(n9572), .A2(n6719), .B1(n9571), .B2(n6720), .C1(
        P1_U3086), .C2(n9119), .ZN(P1_U3340) );
  INV_X1 U8449 ( .A(n8185), .ZN(n8174) );
  OAI222_X1 U8450 ( .A1(n4406), .A2(n10242), .B1(n8588), .B2(n6720), .C1(
        P2_U3151), .C2(n8174), .ZN(P2_U3280) );
  XNOR2_X1 U8451 ( .A(n9944), .B(n6613), .ZN(n6787) );
  XNOR2_X1 U8452 ( .A(n6787), .B(n8110), .ZN(n6735) );
  NAND2_X1 U8453 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  XNOR2_X1 U8454 ( .A(n9937), .B(n6613), .ZN(n6728) );
  XNOR2_X1 U8455 ( .A(n6949), .B(n6728), .ZN(n6750) );
  INV_X1 U8456 ( .A(n6728), .ZN(n6729) );
  NAND2_X1 U8457 ( .A1(n8111), .A2(n6729), .ZN(n6730) );
  INV_X1 U8458 ( .A(n6734), .ZN(n6732) );
  NAND2_X1 U8459 ( .A1(n6732), .A2(n6731), .ZN(n6790) );
  INV_X1 U8460 ( .A(n6790), .ZN(n6733) );
  AOI21_X1 U8461 ( .B1(n6735), .B2(n6734), .A(n6733), .ZN(n6740) );
  INV_X1 U8462 ( .A(n7841), .ZN(n7850) );
  AOI22_X1 U8463 ( .A1(n7850), .A2(n8111), .B1(n7826), .B2(n8109), .ZN(n6737)
         );
  OAI211_X1 U8464 ( .C1(n9944), .C2(n7848), .A(n6737), .B(n6736), .ZN(n6738)
         );
  AOI21_X1 U8465 ( .B1(n6953), .B2(n7851), .A(n6738), .ZN(n6739) );
  OAI21_X1 U8466 ( .B1(n6740), .B2(n7856), .A(n6739), .ZN(P2_U3170) );
  INV_X1 U8467 ( .A(n6741), .ZN(n6743) );
  AOI22_X1 U8468 ( .A1(n9821), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9565), .ZN(n6742) );
  OAI21_X1 U8469 ( .B1(n6743), .B2(n9575), .A(n6742), .ZN(P1_U3339) );
  INV_X1 U8470 ( .A(n8193), .ZN(n8204) );
  OAI222_X1 U8471 ( .A1(n8588), .A2(n6743), .B1(n8204), .B2(P2_U3151), .C1(
        n10154), .C2(n4406), .ZN(P2_U3279) );
  AOI22_X1 U8472 ( .A1(n7850), .A2(n8112), .B1(n7826), .B2(n8110), .ZN(n6745)
         );
  OAI211_X1 U8473 ( .C1(n6746), .C2(n7848), .A(n6745), .B(n6744), .ZN(n6752)
         );
  INV_X1 U8474 ( .A(n6747), .ZN(n6748) );
  AOI211_X1 U8475 ( .C1(n6750), .C2(n6749), .A(n7856), .B(n6748), .ZN(n6751)
         );
  AOI211_X1 U8476 ( .C1(n6806), .C2(n7851), .A(n6752), .B(n6751), .ZN(n6753)
         );
  INV_X1 U8477 ( .A(n6753), .ZN(P2_U3158) );
  AOI211_X1 U8478 ( .C1(n6756), .C2(n6755), .A(n8264), .B(n6754), .ZN(n6757)
         );
  INV_X1 U8479 ( .A(n6757), .ZN(n6770) );
  NAND2_X1 U8480 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n6791) );
  INV_X1 U8481 ( .A(n6791), .ZN(n6768) );
  INV_X1 U8482 ( .A(n6758), .ZN(n6759) );
  AOI21_X1 U8483 ( .B1(n10279), .B2(n6760), .A(n6759), .ZN(n6766) );
  INV_X1 U8484 ( .A(n6761), .ZN(n6762) );
  AOI21_X1 U8485 ( .B1(n6764), .B2(n6763), .A(n6762), .ZN(n6765) );
  OAI22_X1 U8486 ( .A1(n8237), .A2(n6766), .B1(n6765), .B2(n8270), .ZN(n6767)
         );
  AOI211_X1 U8487 ( .C1(n7038), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6768), .B(
        n6767), .ZN(n6769) );
  OAI211_X1 U8488 ( .C1(n8224), .C2(n6771), .A(n6770), .B(n6769), .ZN(P2_U3187) );
  OAI21_X1 U8489 ( .B1(n6773), .B2(n7926), .A(n6772), .ZN(n6774) );
  INV_X1 U8490 ( .A(n6774), .ZN(n9933) );
  OR2_X1 U8491 ( .A1(n9648), .A2(n6775), .ZN(n7371) );
  OAI21_X1 U8492 ( .B1(n6778), .B2(n6777), .A(n6776), .ZN(n6781) );
  OAI22_X1 U8493 ( .A1(n6779), .A2(n9640), .B1(n6949), .B2(n9642), .ZN(n6780)
         );
  AOI21_X1 U8494 ( .B1(n6781), .B2(n8391), .A(n6780), .ZN(n6782) );
  OAI21_X1 U8495 ( .B1(n9933), .B2(n7365), .A(n6782), .ZN(n9935) );
  OAI22_X1 U8496 ( .A1(n5071), .A2(n8331), .B1(n6783), .B2(n9632), .ZN(n6784)
         );
  NOR2_X1 U8497 ( .A1(n9935), .A2(n6784), .ZN(n6785) );
  MUX2_X1 U8498 ( .A(n6333), .B(n6785), .S(n9645), .Z(n6786) );
  OAI21_X1 U8499 ( .B1(n9933), .B2(n7371), .A(n6786), .ZN(P2_U3231) );
  XNOR2_X1 U8500 ( .A(n9949), .B(n7705), .ZN(n6993) );
  XNOR2_X1 U8501 ( .A(n6993), .B(n8109), .ZN(n6996) );
  INV_X1 U8502 ( .A(n6787), .ZN(n6788) );
  NAND2_X1 U8503 ( .A1(n6792), .A2(n6788), .ZN(n6789) );
  NAND2_X1 U8504 ( .A1(n6790), .A2(n6789), .ZN(n6997) );
  XOR2_X1 U8505 ( .A(n6997), .B(n6996), .Z(n6796) );
  OAI21_X1 U8506 ( .B1(n7841), .B2(n6792), .A(n6791), .ZN(n6794) );
  INV_X1 U8507 ( .A(n7826), .ZN(n7854) );
  OAI22_X1 U8508 ( .A1(n7854), .A2(n7006), .B1(n9949), .B2(n7848), .ZN(n6793)
         );
  AOI211_X1 U8509 ( .C1(n6938), .C2(n7851), .A(n6794), .B(n6793), .ZN(n6795)
         );
  OAI21_X1 U8510 ( .B1(n6796), .B2(n7856), .A(n6795), .ZN(P2_U3167) );
  MUX2_X1 U8511 ( .A(n6476), .B(n6797), .S(n9645), .Z(n6800) );
  AOI22_X1 U8512 ( .A1(n8444), .A2(n6798), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8443), .ZN(n6799) );
  OAI211_X1 U8513 ( .C1(n8448), .C2(n6801), .A(n6800), .B(n6799), .ZN(P2_U3232) );
  INV_X1 U8514 ( .A(n6804), .ZN(n7886) );
  XNOR2_X1 U8515 ( .A(n6802), .B(n7886), .ZN(n6803) );
  AOI222_X1 U8516 ( .A1(n8391), .A2(n6803), .B1(n8112), .B2(n8388), .C1(n8110), 
        .C2(n8386), .ZN(n9940) );
  XNOR2_X1 U8517 ( .A(n6805), .B(n6804), .ZN(n9938) );
  INV_X1 U8518 ( .A(n8448), .ZN(n7137) );
  AOI22_X1 U8519 ( .A1(n8444), .A2(n9937), .B1(n8443), .B2(n6806), .ZN(n6807)
         );
  OAI21_X1 U8520 ( .B1(n6808), .B2(n9645), .A(n6807), .ZN(n6809) );
  AOI21_X1 U8521 ( .B1(n9938), .B2(n7137), .A(n6809), .ZN(n6810) );
  OAI21_X1 U8522 ( .B1(n9940), .B2(n9648), .A(n6810), .ZN(P2_U3230) );
  INV_X1 U8523 ( .A(n7118), .ZN(n6814) );
  NAND2_X1 U8524 ( .A1(n10048), .A2(n9003), .ZN(n6812) );
  NAND2_X1 U8525 ( .A1(n9032), .A2(n9140), .ZN(n6811) );
  NAND2_X1 U8526 ( .A1(n6812), .A2(n6811), .ZN(n6932) );
  NAND2_X1 U8527 ( .A1(n6932), .A2(n9713), .ZN(n6813) );
  NAND2_X1 U8528 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9743) );
  OAI211_X1 U8529 ( .C1(n9719), .C2(n6814), .A(n6813), .B(n9743), .ZN(n6820)
         );
  INV_X1 U8530 ( .A(n6815), .ZN(n6816) );
  AOI211_X1 U8531 ( .C1(n6818), .C2(n6817), .A(n9660), .B(n6816), .ZN(n6819)
         );
  AOI211_X1 U8532 ( .C1(n7119), .C2(n9716), .A(n6820), .B(n6819), .ZN(n6821)
         );
  INV_X1 U8533 ( .A(n6821), .ZN(P1_U3230) );
  INV_X1 U8534 ( .A(n6957), .ZN(n8942) );
  NAND2_X1 U8535 ( .A1(n6822), .A2(n6862), .ZN(n6860) );
  INV_X2 U8536 ( .A(n7047), .ZN(n6874) );
  NAND2_X1 U8537 ( .A1(n6846), .A2(n8791), .ZN(n6845) );
  NAND2_X1 U8538 ( .A1(n6845), .A2(n6824), .ZN(n6826) );
  NAND2_X1 U8539 ( .A1(n6825), .A2(n6878), .ZN(n8833) );
  NAND2_X1 U8540 ( .A1(n10048), .A2(n9898), .ZN(n8830) );
  NAND2_X1 U8541 ( .A1(n8833), .A2(n8830), .ZN(n8792) );
  NAND2_X1 U8542 ( .A1(n6826), .A2(n8792), .ZN(n6880) );
  OAI21_X1 U8543 ( .B1(n6826), .B2(n8792), .A(n6880), .ZN(n9900) );
  NOR2_X1 U8544 ( .A1(n6862), .A2(n6957), .ZN(n6861) );
  AOI211_X1 U8545 ( .C1(n6878), .C2(n6850), .A(n9410), .B(n6926), .ZN(n9892)
         );
  NAND2_X1 U8546 ( .A1(n6827), .A2(n6863), .ZN(n6866) );
  NAND2_X1 U8547 ( .A1(n6828), .A2(n6957), .ZN(n6829) );
  NOR2_X1 U8548 ( .A1(n9034), .A2(n6874), .ZN(n6830) );
  NAND2_X1 U8549 ( .A1(n9034), .A2(n6874), .ZN(n8946) );
  XNOR2_X1 U8550 ( .A(n8829), .B(n8792), .ZN(n6832) );
  AOI21_X1 U8551 ( .B1(n6832), .B2(n9402), .A(n6831), .ZN(n9903) );
  INV_X1 U8552 ( .A(n9903), .ZN(n6833) );
  AOI211_X1 U8553 ( .C1(n9924), .C2(n9900), .A(n9892), .B(n6833), .ZN(n6858)
         );
  INV_X1 U8554 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6834) );
  OAI22_X1 U8555 ( .A1(n9491), .A2(n9898), .B1(n9932), .B2(n6834), .ZN(n6835)
         );
  INV_X1 U8556 ( .A(n6835), .ZN(n6836) );
  OAI21_X1 U8557 ( .B1(n6858), .B2(n9929), .A(n6836), .ZN(P1_U3525) );
  INV_X1 U8558 ( .A(n6838), .ZN(n6839) );
  NAND2_X1 U8559 ( .A1(n6839), .A2(n6960), .ZN(n6840) );
  XNOR2_X1 U8560 ( .A(n6837), .B(n6840), .ZN(n6844) );
  NOR2_X1 U8561 ( .A1(n9719), .A2(n7106), .ZN(n6842) );
  AOI22_X1 U8562 ( .A1(n9003), .A2(n9032), .B1(n9030), .B2(n9140), .ZN(n7112)
         );
  OAI22_X1 U8563 ( .A1(n7112), .A2(n9656), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5900), .ZN(n6841) );
  AOI211_X1 U8564 ( .C1(n7108), .C2(n9716), .A(n6842), .B(n6841), .ZN(n6843)
         );
  OAI21_X1 U8565 ( .B1(n6844), .B2(n9660), .A(n6843), .ZN(P1_U3239) );
  INV_X1 U8566 ( .A(n9924), .ZN(n9498) );
  OAI21_X1 U8567 ( .B1(n6846), .B2(n8791), .A(n6845), .ZN(n7052) );
  INV_X1 U8568 ( .A(n7052), .ZN(n6851) );
  XOR2_X1 U8569 ( .A(n8791), .B(n6847), .Z(n6849) );
  AOI21_X1 U8570 ( .B1(n6849), .B2(n9402), .A(n6848), .ZN(n7054) );
  INV_X1 U8571 ( .A(n9410), .ZN(n9864) );
  OAI211_X1 U8572 ( .C1(n6861), .C2(n6874), .A(n6850), .B(n9864), .ZN(n7050)
         );
  OAI211_X1 U8573 ( .C1(n9498), .C2(n6851), .A(n7054), .B(n7050), .ZN(n6876)
         );
  INV_X1 U8574 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6852) );
  OAI22_X1 U8575 ( .A1(n9491), .A2(n6874), .B1(n9932), .B2(n6852), .ZN(n6853)
         );
  AOI21_X1 U8576 ( .B1(n6876), .B2(n9932), .A(n6853), .ZN(n6854) );
  INV_X1 U8577 ( .A(n6854), .ZN(P1_U3524) );
  INV_X1 U8578 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6855) );
  OAI22_X1 U8579 ( .A1(n9551), .A2(n9898), .B1(n9927), .B2(n6855), .ZN(n6856)
         );
  INV_X1 U8580 ( .A(n6856), .ZN(n6857) );
  OAI21_X1 U8581 ( .B1(n6858), .B2(n9557), .A(n6857), .ZN(P1_U3462) );
  INV_X1 U8582 ( .A(n7272), .ZN(n7165) );
  AOI211_X1 U8583 ( .C1(n6862), .C2(n6957), .A(n9410), .B(n6861), .ZN(n6911)
         );
  INV_X1 U8584 ( .A(n7093), .ZN(n7270) );
  INV_X1 U8585 ( .A(n6863), .ZN(n6864) );
  AOI21_X1 U8586 ( .B1(n6866), .B2(n6865), .A(n9854), .ZN(n6867) );
  AOI211_X1 U8587 ( .C1(n7270), .C2(n6900), .A(n6868), .B(n6867), .ZN(n6907)
         );
  INV_X1 U8588 ( .A(n6907), .ZN(n6869) );
  AOI211_X1 U8589 ( .C1(n7165), .C2(n6900), .A(n6911), .B(n6869), .ZN(n6959)
         );
  INV_X1 U8590 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6870) );
  OAI22_X1 U8591 ( .A1(n9551), .A2(n8942), .B1(n9927), .B2(n6870), .ZN(n6871)
         );
  INV_X1 U8592 ( .A(n6871), .ZN(n6872) );
  OAI21_X1 U8593 ( .B1(n6959), .B2(n9557), .A(n6872), .ZN(P1_U3456) );
  INV_X1 U8594 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6873) );
  OAI22_X1 U8595 ( .A1(n9551), .A2(n6874), .B1(n9927), .B2(n6873), .ZN(n6875)
         );
  AOI21_X1 U8596 ( .B1(n6876), .B2(n9927), .A(n6875), .ZN(n6877) );
  INV_X1 U8597 ( .A(n6877), .ZN(P1_U3459) );
  OR2_X1 U8598 ( .A1(n6878), .A2(n10048), .ZN(n6879) );
  NAND2_X1 U8599 ( .A1(n6880), .A2(n6879), .ZN(n6925) );
  OR2_X1 U8600 ( .A1(n9033), .A2(n6884), .ZN(n8834) );
  NAND2_X1 U8601 ( .A1(n9033), .A2(n6884), .ZN(n8836) );
  NAND2_X1 U8602 ( .A1(n6925), .A2(n8796), .ZN(n6924) );
  NAND2_X1 U8603 ( .A1(n6924), .A2(n6881), .ZN(n6883) );
  INV_X1 U8604 ( .A(n9032), .ZN(n6882) );
  NAND2_X1 U8605 ( .A1(n6882), .A2(n9715), .ZN(n8838) );
  NAND2_X1 U8606 ( .A1(n9032), .A2(n9887), .ZN(n8951) );
  NAND2_X1 U8607 ( .A1(n6883), .A2(n8797), .ZN(n7081) );
  OAI21_X1 U8608 ( .B1(n6883), .B2(n8797), .A(n7081), .ZN(n9889) );
  AOI211_X1 U8609 ( .C1(n9715), .C2(n6927), .A(n9410), .B(n7105), .ZN(n9882)
         );
  INV_X1 U8610 ( .A(n8796), .ZN(n6885) );
  NAND2_X1 U8611 ( .A1(n6886), .A2(n6885), .ZN(n6931) );
  NAND2_X1 U8612 ( .A1(n6931), .A2(n8834), .ZN(n7086) );
  INV_X1 U8613 ( .A(n8797), .ZN(n7085) );
  XNOR2_X1 U8614 ( .A(n7086), .B(n7085), .ZN(n6888) );
  INV_X1 U8615 ( .A(n9031), .ZN(n7082) );
  OAI22_X1 U8616 ( .A1(n6887), .A2(n9669), .B1(n7082), .B2(n9667), .ZN(n9714)
         );
  AOI21_X1 U8617 ( .B1(n6888), .B2(n9402), .A(n9714), .ZN(n9891) );
  INV_X1 U8618 ( .A(n9891), .ZN(n6889) );
  AOI211_X1 U8619 ( .C1(n9924), .C2(n9889), .A(n9882), .B(n6889), .ZN(n6895)
         );
  INV_X1 U8620 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6890) );
  OAI22_X1 U8621 ( .A1(n9551), .A2(n9887), .B1(n9927), .B2(n6890), .ZN(n6891)
         );
  INV_X1 U8622 ( .A(n6891), .ZN(n6892) );
  OAI21_X1 U8623 ( .B1(n6895), .B2(n9557), .A(n6892), .ZN(P1_U3468) );
  OAI22_X1 U8624 ( .A1(n9491), .A2(n9887), .B1(n9932), .B2(n6443), .ZN(n6893)
         );
  INV_X1 U8625 ( .A(n6893), .ZN(n6894) );
  OAI21_X1 U8626 ( .B1(n6895), .B2(n9929), .A(n6894), .ZN(P1_U3527) );
  INV_X1 U8627 ( .A(n6896), .ZN(n6898) );
  INV_X1 U8628 ( .A(n9831), .ZN(n9122) );
  OAI222_X1 U8629 ( .A1(n9572), .A2(n6897), .B1(n9571), .B2(n6898), .C1(
        P1_U3086), .C2(n9122), .ZN(P1_U3338) );
  INV_X1 U8630 ( .A(n8231), .ZN(n8209) );
  OAI222_X1 U8631 ( .A1(n4406), .A2(n6899), .B1(n8588), .B2(n6898), .C1(
        P2_U3151), .C2(n8209), .ZN(P2_U3278) );
  INV_X1 U8632 ( .A(n6900), .ZN(n6914) );
  INV_X1 U8633 ( .A(n6901), .ZN(n6902) );
  OR3_X1 U8634 ( .A1(n6904), .A2(n6903), .A3(n6902), .ZN(n6905) );
  OR2_X1 U8635 ( .A1(n9904), .A2(n6906), .ZN(n9874) );
  INV_X2 U8636 ( .A(n9421), .ZN(n9416) );
  MUX2_X1 U8637 ( .A(n6414), .B(n6907), .S(n9416), .Z(n6913) );
  INV_X2 U8638 ( .A(n9345), .ZN(n9380) );
  OAI22_X1 U8639 ( .A1(n9897), .A2(n8942), .B1(n9413), .B2(n6909), .ZN(n6910)
         );
  AOI21_X1 U8640 ( .B1(n6911), .B2(n9380), .A(n6910), .ZN(n6912) );
  OAI211_X1 U8641 ( .C1(n6914), .C2(n9874), .A(n6913), .B(n6912), .ZN(P1_U3292) );
  AOI21_X1 U8642 ( .B1(n9380), .B2(n9864), .A(n9872), .ZN(n6923) );
  OAI21_X1 U8643 ( .B1(n5784), .B2(n9413), .A(n6915), .ZN(n6916) );
  AOI21_X1 U8644 ( .B1(n6918), .B2(n6917), .A(n6916), .ZN(n6919) );
  MUX2_X1 U8645 ( .A(n6920), .B(n6919), .S(n9416), .Z(n6921) );
  OAI21_X1 U8646 ( .B1(n6923), .B2(n6922), .A(n6921), .ZN(P1_U3293) );
  OAI21_X1 U8647 ( .B1(n6925), .B2(n8796), .A(n6924), .ZN(n7125) );
  INV_X1 U8648 ( .A(n6926), .ZN(n6929) );
  INV_X1 U8649 ( .A(n6927), .ZN(n6928) );
  AOI211_X1 U8650 ( .C1(n7119), .C2(n6929), .A(n9410), .B(n6928), .ZN(n7117)
         );
  NAND3_X1 U8651 ( .A1(n8835), .A2(n8796), .A3(n8833), .ZN(n6930) );
  AOI21_X1 U8652 ( .B1(n6931), .B2(n6930), .A(n9854), .ZN(n6933) );
  OR2_X1 U8653 ( .A1(n6933), .A2(n6932), .ZN(n7122) );
  AOI211_X1 U8654 ( .C1(n9924), .C2(n7125), .A(n7117), .B(n7122), .ZN(n6971)
         );
  INV_X1 U8655 ( .A(n9551), .ZN(n9554) );
  AOI22_X1 U8656 ( .A1(n9554), .A2(n7119), .B1(n9557), .B2(
        P1_REG0_REG_4__SCAN_IN), .ZN(n6934) );
  OAI21_X1 U8657 ( .B1(n6971), .B2(n9557), .A(n6934), .ZN(P1_U3465) );
  XNOR2_X1 U8658 ( .A(n8109), .B(n6939), .ZN(n7889) );
  XOR2_X1 U8659 ( .A(n6935), .B(n7889), .Z(n9950) );
  XNOR2_X1 U8660 ( .A(n6936), .B(n7889), .ZN(n6937) );
  AOI222_X1 U8661 ( .A1(n8391), .A2(n6937), .B1(n8108), .B2(n8386), .C1(n8110), 
        .C2(n8388), .ZN(n9948) );
  MUX2_X1 U8662 ( .A(n6764), .B(n9948), .S(n9645), .Z(n6941) );
  AOI22_X1 U8663 ( .A1(n8444), .A2(n6939), .B1(n8443), .B2(n6938), .ZN(n6940)
         );
  OAI211_X1 U8664 ( .C1(n8448), .C2(n9950), .A(n6941), .B(n6940), .ZN(P2_U3228) );
  NAND2_X1 U8665 ( .A1(n7946), .A2(n7939), .ZN(n7887) );
  XNOR2_X1 U8666 ( .A(n6943), .B(n7887), .ZN(n9942) );
  INV_X1 U8667 ( .A(n7887), .ZN(n7936) );
  INV_X1 U8668 ( .A(n6944), .ZN(n6945) );
  NOR2_X1 U8669 ( .A1(n6946), .A2(n6945), .ZN(n6947) );
  AOI211_X1 U8670 ( .C1(n7936), .C2(n6948), .A(n9637), .B(n6947), .ZN(n6951)
         );
  OAI22_X1 U8671 ( .A1(n7829), .A2(n9642), .B1(n6949), .B2(n9640), .ZN(n6950)
         );
  NOR2_X1 U8672 ( .A1(n6951), .A2(n6950), .ZN(n9943) );
  MUX2_X1 U8673 ( .A(n6952), .B(n9943), .S(n9645), .Z(n6956) );
  AOI22_X1 U8674 ( .A1(n8444), .A2(n6954), .B1(n8443), .B2(n6953), .ZN(n6955)
         );
  OAI211_X1 U8675 ( .C1(n8448), .C2(n9942), .A(n6956), .B(n6955), .ZN(P2_U3229) );
  AOI22_X1 U8676 ( .A1(n9503), .A2(n6957), .B1(n9929), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6958) );
  OAI21_X1 U8677 ( .B1(n6959), .B2(n9929), .A(n6958), .ZN(P1_U3523) );
  NAND2_X1 U8678 ( .A1(n6961), .A2(n6960), .ZN(n6965) );
  XNOR2_X1 U8679 ( .A(n6963), .B(n6962), .ZN(n6964) );
  XNOR2_X1 U8680 ( .A(n6965), .B(n6964), .ZN(n6969) );
  INV_X1 U8681 ( .A(n9029), .ZN(n7178) );
  OAI22_X1 U8682 ( .A1(n7082), .A2(n9669), .B1(n7178), .B2(n9667), .ZN(n7084)
         );
  AOI22_X1 U8683 ( .A1(n7084), .A2(n9713), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n6966) );
  OAI21_X1 U8684 ( .B1(n7094), .B2(n9719), .A(n6966), .ZN(n6967) );
  AOI21_X1 U8685 ( .B1(n7181), .B2(n9716), .A(n6967), .ZN(n6968) );
  OAI21_X1 U8686 ( .B1(n6969), .B2(n9660), .A(n6968), .ZN(P1_U3213) );
  AOI22_X1 U8687 ( .A1(n9503), .A2(n7119), .B1(n9929), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6970) );
  OAI21_X1 U8688 ( .B1(n6971), .B2(n9929), .A(n6970), .ZN(P1_U3526) );
  INV_X1 U8689 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U8690 ( .A1(n6980), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6972) );
  INV_X1 U8691 ( .A(n7030), .ZN(n6974) );
  AOI21_X1 U8692 ( .B1(n10002), .B2(n6975), .A(n6974), .ZN(n6990) );
  OAI21_X1 U8693 ( .B1(n6977), .B2(n6980), .A(n6976), .ZN(n7027) );
  MUX2_X1 U8694 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8253), .Z(n7023) );
  XNOR2_X1 U8695 ( .A(n7023), .B(n7025), .ZN(n7026) );
  XNOR2_X1 U8696 ( .A(n7027), .B(n7026), .ZN(n6978) );
  NAND2_X1 U8697 ( .A1(n6978), .A2(n8226), .ZN(n6989) );
  INV_X1 U8698 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10372) );
  AND2_X1 U8699 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7008) );
  INV_X1 U8700 ( .A(n7008), .ZN(n6979) );
  OAI21_X1 U8701 ( .B1(n8259), .B2(n10372), .A(n6979), .ZN(n6987) );
  NAND2_X1 U8702 ( .A1(n6980), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6981) );
  INV_X1 U8703 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7065) );
  NAND2_X1 U8704 ( .A1(n6984), .A2(n7065), .ZN(n6985) );
  AOI21_X1 U8705 ( .B1(n7036), .B2(n6985), .A(n8270), .ZN(n6986) );
  AOI211_X1 U8706 ( .C1(n8261), .C2(n7025), .A(n6987), .B(n6986), .ZN(n6988)
         );
  OAI211_X1 U8707 ( .C1(n6990), .C2(n8237), .A(n6989), .B(n6988), .ZN(P2_U3189) );
  INV_X1 U8708 ( .A(n9123), .ZN(n9847) );
  INV_X1 U8709 ( .A(n6991), .ZN(n7020) );
  OAI222_X1 U8710 ( .A1(P1_U3086), .A2(n9847), .B1(n9571), .B2(n7020), .C1(
        n6992), .C2(n9572), .ZN(P1_U3337) );
  XNOR2_X1 U8711 ( .A(n7067), .B(n7735), .ZN(n7205) );
  XNOR2_X1 U8712 ( .A(n7205), .B(n7204), .ZN(n7004) );
  INV_X1 U8713 ( .A(n6993), .ZN(n6994) );
  NOR2_X1 U8714 ( .A1(n6994), .A2(n8109), .ZN(n6995) );
  XNOR2_X1 U8715 ( .A(n9955), .B(n7705), .ZN(n6998) );
  XNOR2_X1 U8716 ( .A(n6998), .B(n8108), .ZN(n7824) );
  INV_X1 U8717 ( .A(n6998), .ZN(n6999) );
  NAND2_X1 U8718 ( .A1(n6999), .A2(n8108), .ZN(n7000) );
  INV_X1 U8719 ( .A(n7207), .ZN(n7002) );
  AOI21_X1 U8720 ( .B1(n7004), .B2(n7003), .A(n7002), .ZN(n7012) );
  INV_X1 U8721 ( .A(n7005), .ZN(n7064) );
  INV_X1 U8722 ( .A(n7851), .ZN(n7714) );
  NOR2_X1 U8723 ( .A1(n7841), .A2(n7006), .ZN(n7007) );
  AOI211_X1 U8724 ( .C1(n7826), .C2(n8106), .A(n7008), .B(n7007), .ZN(n7009)
         );
  OAI21_X1 U8725 ( .B1(n7064), .B2(n7714), .A(n7009), .ZN(n7010) );
  AOI21_X1 U8726 ( .B1(n7067), .B2(n7861), .A(n7010), .ZN(n7011) );
  OAI21_X1 U8727 ( .B1(n7012), .B2(n7856), .A(n7011), .ZN(P2_U3153) );
  NAND2_X1 U8728 ( .A1(n7013), .A2(n7014), .ZN(n7015) );
  AND2_X1 U8729 ( .A1(n7949), .A2(n7941), .ZN(n7890) );
  XNOR2_X1 U8730 ( .A(n7015), .B(n7890), .ZN(n9956) );
  XNOR2_X1 U8731 ( .A(n7016), .B(n7890), .ZN(n7017) );
  AOI222_X1 U8732 ( .A1(n8391), .A2(n7017), .B1(n8107), .B2(n8386), .C1(n8109), 
        .C2(n8388), .ZN(n9954) );
  MUX2_X1 U8733 ( .A(n10327), .B(n9954), .S(n9645), .Z(n7019) );
  AOI22_X1 U8734 ( .A1(n8444), .A2(n7831), .B1(n8443), .B2(n7832), .ZN(n7018)
         );
  OAI211_X1 U8735 ( .C1(n9956), .C2(n8448), .A(n7019), .B(n7018), .ZN(P2_U3227) );
  INV_X1 U8736 ( .A(n8251), .ZN(n8234) );
  OAI222_X1 U8737 ( .A1(n4406), .A2(n7021), .B1(n8234), .B2(P2_U3151), .C1(
        n8588), .C2(n7020), .ZN(P2_U3277) );
  NAND2_X1 U8738 ( .A1(n8225), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7022) );
  OAI21_X1 U8739 ( .B1(n7879), .B2(n8225), .A(n7022), .ZN(P2_U3521) );
  MUX2_X1 U8740 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8253), .Z(n7144) );
  XOR2_X1 U8741 ( .A(n7151), .B(n7144), .Z(n7145) );
  INV_X1 U8742 ( .A(n7023), .ZN(n7024) );
  AOI22_X1 U8743 ( .A1(n7027), .A2(n7026), .B1(n7025), .B2(n7024), .ZN(n7146)
         );
  XOR2_X1 U8744 ( .A(n7145), .B(n7146), .Z(n7045) );
  INV_X1 U8745 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U8746 ( .A(n10004), .B(P2_REG1_REG_8__SCAN_IN), .S(n7151), .Z(n7028)
         );
  NAND3_X1 U8747 ( .A1(n7030), .A2(n4513), .A3(n7029), .ZN(n7031) );
  AOI21_X1 U8748 ( .B1(n7152), .B2(n7031), .A(n8237), .ZN(n7043) );
  INV_X1 U8749 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7134) );
  MUX2_X1 U8750 ( .A(n7134), .B(P2_REG2_REG_8__SCAN_IN), .S(n7151), .Z(n7033)
         );
  NAND2_X1 U8751 ( .A1(n7032), .A2(n7033), .ZN(n7140) );
  INV_X1 U8752 ( .A(n7033), .ZN(n7035) );
  NAND3_X1 U8753 ( .A1(n7036), .A2(n7035), .A3(n7034), .ZN(n7037) );
  AOI21_X1 U8754 ( .B1(n7140), .B2(n7037), .A(n8270), .ZN(n7042) );
  INV_X1 U8755 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U8756 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10296), .ZN(n7208) );
  INV_X1 U8757 ( .A(n7208), .ZN(n7040) );
  NAND2_X1 U8758 ( .A1(n7038), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n7039) );
  OAI211_X1 U8759 ( .C1(n8224), .C2(n7143), .A(n7040), .B(n7039), .ZN(n7041)
         );
  NOR3_X1 U8760 ( .A1(n7043), .A2(n7042), .A3(n7041), .ZN(n7044) );
  OAI21_X1 U8761 ( .B1(n7045), .B2(n8264), .A(n7044), .ZN(P2_U3190) );
  NAND2_X1 U8762 ( .A1(n9416), .A2(n7270), .ZN(n7046) );
  INV_X1 U8763 ( .A(n9413), .ZN(n9894) );
  AOI22_X1 U8764 ( .A1(n9904), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9894), .ZN(n7049) );
  NAND2_X1 U8765 ( .A1(n9872), .A2(n7047), .ZN(n7048) );
  OAI211_X1 U8766 ( .C1(n9345), .C2(n7050), .A(n7049), .B(n7048), .ZN(n7051)
         );
  AOI21_X1 U8767 ( .B1(n7052), .B2(n9901), .A(n7051), .ZN(n7053) );
  OAI21_X1 U8768 ( .B1(n7054), .B2(n9421), .A(n7053), .ZN(P1_U3291) );
  NAND2_X1 U8769 ( .A1(n7057), .A2(n7957), .ZN(n7058) );
  NAND2_X1 U8770 ( .A1(n7059), .A2(n7058), .ZN(n9960) );
  XNOR2_X1 U8771 ( .A(n7060), .B(n7957), .ZN(n7061) );
  NAND2_X1 U8772 ( .A1(n7061), .A2(n8391), .ZN(n7063) );
  AOI22_X1 U8773 ( .A1(n8388), .A2(n8108), .B1(n8106), .B2(n8386), .ZN(n7062)
         );
  OAI211_X1 U8774 ( .C1(n9960), .C2(n7365), .A(n7063), .B(n7062), .ZN(n9962)
         );
  NAND2_X1 U8775 ( .A1(n9962), .A2(n9645), .ZN(n7069) );
  OAI22_X1 U8776 ( .A1(n9645), .A2(n7065), .B1(n7064), .B2(n9632), .ZN(n7066)
         );
  AOI21_X1 U8777 ( .B1(n8444), .B2(n7067), .A(n7066), .ZN(n7068) );
  OAI211_X1 U8778 ( .C1(n9960), .C2(n7371), .A(n7069), .B(n7068), .ZN(P2_U3226) );
  INV_X1 U8779 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10064) );
  INV_X1 U8780 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U8781 ( .A1(n7070), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n7073) );
  NAND2_X1 U8782 ( .A1(n7071), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7072) );
  OAI211_X1 U8783 ( .C1(n7074), .C2(n10286), .A(n7073), .B(n7072), .ZN(n7075)
         );
  INV_X1 U8784 ( .A(n7075), .ZN(n7076) );
  INV_X1 U8785 ( .A(n8272), .ZN(n7078) );
  NAND2_X1 U8786 ( .A1(n7078), .A2(P2_U3893), .ZN(n7079) );
  OAI21_X1 U8787 ( .B1(P2_U3893), .B2(n10064), .A(n7079), .ZN(P2_U3522) );
  NAND2_X1 U8788 ( .A1(n6882), .A2(n9887), .ZN(n7080) );
  NAND2_X1 U8789 ( .A1(n7081), .A2(n7080), .ZN(n7103) );
  INV_X1 U8790 ( .A(n7108), .ZN(n9908) );
  NAND2_X1 U8791 ( .A1(n9908), .A2(n9031), .ZN(n8840) );
  NAND2_X1 U8792 ( .A1(n7082), .A2(n7108), .ZN(n8955) );
  NAND2_X1 U8793 ( .A1(n8840), .A2(n8955), .ZN(n7110) );
  NAND2_X1 U8794 ( .A1(n7103), .A2(n7110), .ZN(n7102) );
  INV_X1 U8795 ( .A(n9030), .ZN(n7262) );
  OR2_X1 U8796 ( .A1(n7181), .A2(n7262), .ZN(n7295) );
  NAND2_X1 U8797 ( .A1(n7181), .A2(n7262), .ZN(n7264) );
  NAND2_X1 U8798 ( .A1(n7295), .A2(n7264), .ZN(n7088) );
  NAND2_X1 U8799 ( .A1(n7083), .A2(n7088), .ZN(n7183) );
  OAI21_X1 U8800 ( .B1(n7083), .B2(n7088), .A(n7183), .ZN(n7164) );
  INV_X1 U8801 ( .A(n7164), .ZN(n7101) );
  INV_X1 U8802 ( .A(n7084), .ZN(n7092) );
  NAND2_X1 U8803 ( .A1(n7086), .A2(n7085), .ZN(n7087) );
  NAND2_X1 U8804 ( .A1(n7087), .A2(n8838), .ZN(n7111) );
  INV_X1 U8805 ( .A(n8955), .ZN(n8798) );
  INV_X1 U8806 ( .A(n7088), .ZN(n8844) );
  NAND3_X1 U8807 ( .A1(n7293), .A2(n8844), .A3(n8840), .ZN(n7265) );
  INV_X1 U8808 ( .A(n7265), .ZN(n7090) );
  AOI21_X1 U8809 ( .B1(n7293), .B2(n8840), .A(n8844), .ZN(n7089) );
  OAI21_X1 U8810 ( .B1(n7090), .B2(n7089), .A(n9402), .ZN(n7091) );
  OAI211_X1 U8811 ( .C1(n7101), .C2(n7093), .A(n7092), .B(n7091), .ZN(n7162)
         );
  NAND2_X1 U8812 ( .A1(n7162), .A2(n9416), .ZN(n7100) );
  NAND2_X1 U8813 ( .A1(n7105), .A2(n9908), .ZN(n7104) );
  NOR2_X1 U8814 ( .A1(n7104), .A2(n7181), .ZN(n7271) );
  AOI211_X1 U8815 ( .C1(n7181), .C2(n7104), .A(n9410), .B(n7271), .ZN(n7163)
         );
  INV_X1 U8816 ( .A(n7181), .ZN(n7097) );
  INV_X1 U8817 ( .A(n7094), .ZN(n7095) );
  AOI22_X1 U8818 ( .A1(n9904), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7095), .B2(
        n9894), .ZN(n7096) );
  OAI21_X1 U8819 ( .B1(n7097), .B2(n9897), .A(n7096), .ZN(n7098) );
  AOI21_X1 U8820 ( .B1(n7163), .B2(n9380), .A(n7098), .ZN(n7099) );
  OAI211_X1 U8821 ( .C1(n7101), .C2(n9874), .A(n7100), .B(n7099), .ZN(P1_U3286) );
  OAI21_X1 U8822 ( .B1(n7103), .B2(n7110), .A(n7102), .ZN(n9911) );
  OAI211_X1 U8823 ( .C1(n7105), .C2(n9908), .A(n7104), .B(n9864), .ZN(n9907)
         );
  INV_X1 U8824 ( .A(n7106), .ZN(n7107) );
  AOI22_X1 U8825 ( .A1(n9872), .A2(n7108), .B1(n7107), .B2(n9894), .ZN(n7109)
         );
  OAI21_X1 U8826 ( .B1(n9907), .B2(n9345), .A(n7109), .ZN(n7115) );
  XNOR2_X1 U8827 ( .A(n7111), .B(n7110), .ZN(n7113) );
  OAI21_X1 U8828 ( .B1(n7113), .B2(n9854), .A(n7112), .ZN(n9909) );
  MUX2_X1 U8829 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n9909), .S(n9416), .Z(n7114)
         );
  AOI211_X1 U8830 ( .C1(n9901), .C2(n9911), .A(n7115), .B(n7114), .ZN(n7116)
         );
  INV_X1 U8831 ( .A(n7116), .ZN(P1_U3287) );
  INV_X1 U8832 ( .A(n7117), .ZN(n7121) );
  AOI22_X1 U8833 ( .A1(n9872), .A2(n7119), .B1(n7118), .B2(n9894), .ZN(n7120)
         );
  OAI21_X1 U8834 ( .B1(n7121), .B2(n9345), .A(n7120), .ZN(n7124) );
  MUX2_X1 U8835 ( .A(n7122), .B(P1_REG2_REG_4__SCAN_IN), .S(n9904), .Z(n7123)
         );
  AOI211_X1 U8836 ( .C1(n9901), .C2(n7125), .A(n7124), .B(n7123), .ZN(n7126)
         );
  INV_X1 U8837 ( .A(n7126), .ZN(P1_U3289) );
  AOI21_X1 U8838 ( .B1(n7128), .B2(n7127), .A(n9637), .ZN(n7131) );
  OAI22_X1 U8839 ( .A1(n7204), .A2(n9640), .B1(n7361), .B2(n9642), .ZN(n7129)
         );
  AOI21_X1 U8840 ( .B1(n7131), .B2(n7130), .A(n7129), .ZN(n9964) );
  XNOR2_X1 U8841 ( .A(n7132), .B(n7892), .ZN(n9967) );
  NOR2_X1 U8842 ( .A1(n9965), .A2(n8277), .ZN(n7136) );
  INV_X1 U8843 ( .A(n7210), .ZN(n7133) );
  OAI22_X1 U8844 ( .A1(n9645), .A2(n7134), .B1(n7133), .B2(n9632), .ZN(n7135)
         );
  AOI211_X1 U8845 ( .C1(n9967), .C2(n7137), .A(n7136), .B(n7135), .ZN(n7138)
         );
  OAI21_X1 U8846 ( .B1(n9964), .B2(n9648), .A(n7138), .ZN(P2_U3225) );
  INV_X1 U8847 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7323) );
  OR2_X1 U8848 ( .A1(n7151), .A2(n7134), .ZN(n7139) );
  NAND2_X1 U8849 ( .A1(n7140), .A2(n7139), .ZN(n7141) );
  AOI21_X1 U8850 ( .B1(n7323), .B2(n7142), .A(n7235), .ZN(n7161) );
  OAI22_X1 U8851 ( .A1(n7146), .A2(n7145), .B1(n7144), .B2(n7143), .ZN(n7148)
         );
  MUX2_X1 U8852 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8253), .Z(n7250) );
  XNOR2_X1 U8853 ( .A(n7250), .B(n7158), .ZN(n7147) );
  NAND2_X1 U8854 ( .A1(n7147), .A2(n7148), .ZN(n7251) );
  OAI21_X1 U8855 ( .B1(n7148), .B2(n7147), .A(n7251), .ZN(n7149) );
  NAND2_X1 U8856 ( .A1(n7149), .A2(n8226), .ZN(n7160) );
  INV_X1 U8857 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10370) );
  NOR2_X1 U8858 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10288), .ZN(n7283) );
  INV_X1 U8859 ( .A(n7283), .ZN(n7150) );
  OAI21_X1 U8860 ( .B1(n8259), .B2(n10370), .A(n7150), .ZN(n7157) );
  INV_X1 U8861 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10287) );
  AOI21_X1 U8862 ( .B1(n7154), .B2(n10287), .A(n7238), .ZN(n7155) );
  NOR2_X1 U8863 ( .A1(n7155), .A2(n8237), .ZN(n7156) );
  AOI211_X1 U8864 ( .C1(n8261), .C2(n7158), .A(n7157), .B(n7156), .ZN(n7159)
         );
  OAI211_X1 U8865 ( .C1(n7161), .C2(n8270), .A(n7160), .B(n7159), .ZN(P2_U3191) );
  AOI211_X1 U8866 ( .C1(n7165), .C2(n7164), .A(n7163), .B(n7162), .ZN(n7171)
         );
  INV_X1 U8867 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7166) );
  NOR2_X1 U8868 ( .A1(n9927), .A2(n7166), .ZN(n7167) );
  AOI21_X1 U8869 ( .B1(n9554), .B2(n7181), .A(n7167), .ZN(n7168) );
  OAI21_X1 U8870 ( .B1(n7171), .B2(n9557), .A(n7168), .ZN(P1_U3474) );
  NOR2_X1 U8871 ( .A1(n9932), .A2(n6446), .ZN(n7169) );
  AOI21_X1 U8872 ( .B1(n9503), .B2(n7181), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8873 ( .B1(n7171), .B2(n9929), .A(n7170), .ZN(P1_U3529) );
  INV_X1 U8874 ( .A(n7172), .ZN(n7174) );
  OAI222_X1 U8875 ( .A1(n4406), .A2(n7173), .B1(n8588), .B2(n7174), .C1(
        P2_U3151), .C2(n8247), .ZN(P2_U3276) );
  OAI222_X1 U8876 ( .A1(n9572), .A2(n7175), .B1(n9571), .B2(n7174), .C1(
        P1_U3086), .C2(n9014), .ZN(P1_U3336) );
  NAND2_X1 U8877 ( .A1(n9873), .A2(n7178), .ZN(n8848) );
  AND2_X1 U8878 ( .A1(n8848), .A2(n7264), .ZN(n8847) );
  OR2_X1 U8879 ( .A1(n9873), .A2(n7178), .ZN(n7296) );
  INV_X1 U8880 ( .A(n7296), .ZN(n7176) );
  AOI21_X1 U8881 ( .B1(n7265), .B2(n8847), .A(n7176), .ZN(n7177) );
  INV_X1 U8882 ( .A(n9028), .ZN(n7263) );
  OR2_X1 U8883 ( .A1(n7306), .A2(n7263), .ZN(n8857) );
  NAND2_X1 U8884 ( .A1(n7306), .A2(n7263), .ZN(n8852) );
  NAND2_X1 U8885 ( .A1(n8857), .A2(n8852), .ZN(n7185) );
  XNOR2_X1 U8886 ( .A(n7177), .B(n7185), .ZN(n7180) );
  NOR2_X1 U8887 ( .A1(n7178), .A2(n9669), .ZN(n7227) );
  INV_X1 U8888 ( .A(n7227), .ZN(n7179) );
  OAI21_X1 U8889 ( .B1(n7180), .B2(n9854), .A(n7179), .ZN(n7196) );
  INV_X1 U8890 ( .A(n7196), .ZN(n7195) );
  NAND2_X1 U8891 ( .A1(n7183), .A2(n7182), .ZN(n7261) );
  NAND2_X1 U8892 ( .A1(n7296), .A2(n8848), .ZN(n7266) );
  NAND2_X1 U8893 ( .A1(n7261), .A2(n7266), .ZN(n7260) );
  OR2_X1 U8894 ( .A1(n9873), .A2(n9029), .ZN(n7184) );
  NAND2_X1 U8895 ( .A1(n7260), .A2(n7184), .ZN(n7186) );
  NAND2_X1 U8896 ( .A1(n7186), .A2(n7185), .ZN(n7304) );
  OAI21_X1 U8897 ( .B1(n7186), .B2(n7185), .A(n7304), .ZN(n7198) );
  NAND2_X1 U8898 ( .A1(n7198), .A2(n9901), .ZN(n7194) );
  INV_X1 U8899 ( .A(n9873), .ZN(n9704) );
  XNOR2_X1 U8900 ( .A(n7307), .B(n7306), .ZN(n7188) );
  NOR2_X1 U8901 ( .A1(n7413), .A2(n9667), .ZN(n7226) );
  INV_X1 U8902 ( .A(n7226), .ZN(n7187) );
  OAI21_X1 U8903 ( .B1(n7188), .B2(n9410), .A(n7187), .ZN(n7197) );
  INV_X1 U8904 ( .A(n7306), .ZN(n7189) );
  NOR2_X1 U8905 ( .A1(n7189), .A2(n9897), .ZN(n7192) );
  INV_X1 U8906 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7190) );
  OAI22_X1 U8907 ( .A1(n9416), .A2(n7190), .B1(n7230), .B2(n9413), .ZN(n7191)
         );
  AOI211_X1 U8908 ( .C1(n7197), .C2(n9380), .A(n7192), .B(n7191), .ZN(n7193)
         );
  OAI211_X1 U8909 ( .C1(n9421), .C2(n7195), .A(n7194), .B(n7193), .ZN(P1_U3284) );
  AOI211_X1 U8910 ( .C1(n7198), .C2(n9924), .A(n7197), .B(n7196), .ZN(n7203)
         );
  AOI22_X1 U8911 ( .A1(n7306), .A2(n9503), .B1(n9929), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7199) );
  OAI21_X1 U8912 ( .B1(n7203), .B2(n9929), .A(n7199), .ZN(P1_U3531) );
  INV_X1 U8913 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7200) );
  NOR2_X1 U8914 ( .A1(n9927), .A2(n7200), .ZN(n7201) );
  AOI21_X1 U8915 ( .B1(n7306), .B2(n9554), .A(n7201), .ZN(n7202) );
  OAI21_X1 U8916 ( .B1(n7203), .B2(n9557), .A(n7202), .ZN(P1_U3480) );
  NAND2_X1 U8917 ( .A1(n7205), .A2(n7204), .ZN(n7206) );
  AND2_X2 U8918 ( .A1(n7207), .A2(n7206), .ZN(n7349) );
  XNOR2_X1 U8919 ( .A(n9965), .B(n7735), .ZN(n7342) );
  XNOR2_X1 U8920 ( .A(n7349), .B(n7342), .ZN(n7280) );
  XNOR2_X1 U8921 ( .A(n7280), .B(n8106), .ZN(n7216) );
  AOI21_X1 U8922 ( .B1(n7850), .B2(n8107), .A(n7208), .ZN(n7214) );
  NAND2_X1 U8923 ( .A1(n7209), .A2(n7861), .ZN(n7213) );
  NAND2_X1 U8924 ( .A1(n7851), .A2(n7210), .ZN(n7212) );
  NAND2_X1 U8925 ( .A1(n7826), .A2(n8105), .ZN(n7211) );
  NAND4_X1 U8926 ( .A1(n7214), .A2(n7213), .A3(n7212), .A4(n7211), .ZN(n7215)
         );
  AOI21_X1 U8927 ( .B1(n7216), .B2(n7839), .A(n7215), .ZN(n7217) );
  INV_X1 U8928 ( .A(n7217), .ZN(P2_U3161) );
  INV_X1 U8929 ( .A(n7218), .ZN(n7219) );
  NOR2_X1 U8930 ( .A1(n7220), .A2(n7219), .ZN(n7222) );
  AOI21_X1 U8931 ( .B1(n7220), .B2(n7219), .A(n7222), .ZN(n9697) );
  NAND2_X1 U8932 ( .A1(n9697), .A2(n9698), .ZN(n9696) );
  NOR2_X1 U8933 ( .A1(n7222), .A2(n7221), .ZN(n7225) );
  INV_X1 U8934 ( .A(n7223), .ZN(n7224) );
  AOI21_X1 U8935 ( .B1(n9696), .B2(n7225), .A(n7224), .ZN(n7233) );
  OAI21_X1 U8936 ( .B1(n7227), .B2(n7226), .A(n9713), .ZN(n7229) );
  OAI211_X1 U8937 ( .C1(n9719), .C2(n7230), .A(n7229), .B(n7228), .ZN(n7231)
         );
  AOI21_X1 U8938 ( .B1(n7306), .B2(n9716), .A(n7231), .ZN(n7232) );
  OAI21_X1 U8939 ( .B1(n7233), .B2(n9660), .A(n7232), .ZN(P1_U3231) );
  INV_X1 U8940 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7234) );
  MUX2_X1 U8941 ( .A(n7234), .B(P2_REG2_REG_10__SCAN_IN), .S(n7248), .Z(n7237)
         );
  OAI21_X1 U8942 ( .B1(n7237), .B2(n7236), .A(n7440), .ZN(n7247) );
  NAND2_X1 U8943 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7351) );
  INV_X1 U8944 ( .A(n7351), .ZN(n7246) );
  INV_X1 U8945 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7240) );
  MUX2_X1 U8946 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n7240), .S(n7248), .Z(n7241)
         );
  AOI21_X1 U8947 ( .B1(n7242), .B2(n7241), .A(n7437), .ZN(n7244) );
  INV_X1 U8948 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7243) );
  OAI22_X1 U8949 ( .A1(n8237), .A2(n7244), .B1(n8259), .B2(n7243), .ZN(n7245)
         );
  AOI211_X1 U8950 ( .C1(n4594), .C2(n7247), .A(n7246), .B(n7245), .ZN(n7257)
         );
  MUX2_X1 U8951 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8253), .Z(n7444) );
  XNOR2_X1 U8952 ( .A(n7444), .B(n7248), .ZN(n7254) );
  OR2_X1 U8953 ( .A1(n7250), .A2(n7249), .ZN(n7252) );
  NAND2_X1 U8954 ( .A1(n7252), .A2(n7251), .ZN(n7253) );
  NAND2_X1 U8955 ( .A1(n7254), .A2(n7253), .ZN(n7445) );
  OAI21_X1 U8956 ( .B1(n7254), .B2(n7253), .A(n7445), .ZN(n7255) );
  NAND2_X1 U8957 ( .A1(n7255), .A2(n8226), .ZN(n7256) );
  OAI211_X1 U8958 ( .C1(n8224), .C2(n7443), .A(n7257), .B(n7256), .ZN(P2_U3192) );
  INV_X1 U8959 ( .A(n7258), .ZN(n7291) );
  OAI222_X1 U8960 ( .A1(n8588), .A2(n7291), .B1(n8084), .B2(P2_U3151), .C1(
        n7259), .C2(n4406), .ZN(P2_U3275) );
  OAI21_X1 U8961 ( .B1(n7261), .B2(n7266), .A(n7260), .ZN(n9878) );
  INV_X1 U8962 ( .A(n9878), .ZN(n7273) );
  OAI22_X1 U8963 ( .A1(n7263), .A2(n9667), .B1(n7262), .B2(n9669), .ZN(n9701)
         );
  NAND2_X1 U8964 ( .A1(n7265), .A2(n7264), .ZN(n7267) );
  XNOR2_X1 U8965 ( .A(n7267), .B(n7266), .ZN(n7268) );
  NOR2_X1 U8966 ( .A1(n7268), .A2(n9854), .ZN(n7269) );
  AOI211_X1 U8967 ( .C1(n9878), .C2(n7270), .A(n9701), .B(n7269), .ZN(n9881)
         );
  OAI211_X1 U8968 ( .C1(n7271), .C2(n9704), .A(n7307), .B(n9864), .ZN(n9875)
         );
  OAI211_X1 U8969 ( .C1(n7273), .C2(n7272), .A(n9881), .B(n9875), .ZN(n7278)
         );
  OAI22_X1 U8970 ( .A1(n9704), .A2(n9491), .B1(n9932), .B2(n6448), .ZN(n7274)
         );
  AOI21_X1 U8971 ( .B1(n7278), .B2(n9932), .A(n7274), .ZN(n7275) );
  INV_X1 U8972 ( .A(n7275), .ZN(P1_U3530) );
  INV_X1 U8973 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7276) );
  OAI22_X1 U8974 ( .A1(n9704), .A2(n9551), .B1(n9927), .B2(n7276), .ZN(n7277)
         );
  AOI21_X1 U8975 ( .B1(n7278), .B2(n9927), .A(n7277), .ZN(n7279) );
  INV_X1 U8976 ( .A(n7279), .ZN(P1_U3477) );
  OAI22_X1 U8977 ( .A1(n7280), .A2(n8106), .B1(n7349), .B2(n7342), .ZN(n7282)
         );
  XNOR2_X1 U8978 ( .A(n7325), .B(n7735), .ZN(n7343) );
  XNOR2_X1 U8979 ( .A(n7343), .B(n8105), .ZN(n7281) );
  XNOR2_X1 U8980 ( .A(n7282), .B(n7281), .ZN(n7289) );
  AOI21_X1 U8981 ( .B1(n7850), .B2(n8106), .A(n7283), .ZN(n7287) );
  NAND2_X1 U8982 ( .A1(n7325), .A2(n7861), .ZN(n7286) );
  NAND2_X1 U8983 ( .A1(n7851), .A2(n7321), .ZN(n7285) );
  NAND2_X1 U8984 ( .A1(n7826), .A2(n8104), .ZN(n7284) );
  NAND4_X1 U8985 ( .A1(n7287), .A2(n7286), .A3(n7285), .A4(n7284), .ZN(n7288)
         );
  AOI21_X1 U8986 ( .B1(n7289), .B2(n7839), .A(n7288), .ZN(n7290) );
  INV_X1 U8987 ( .A(n7290), .ZN(P2_U3171) );
  OAI222_X1 U8988 ( .A1(n9572), .A2(n7292), .B1(n9571), .B2(n7291), .C1(n9007), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  OR2_X1 U8989 ( .A1(n9664), .A2(n7413), .ZN(n8958) );
  NAND2_X1 U8990 ( .A1(n9664), .A2(n7413), .ZN(n8858) );
  NAND2_X1 U8991 ( .A1(n8958), .A2(n8858), .ZN(n8803) );
  INV_X1 U8992 ( .A(n8803), .ZN(n7299) );
  NAND2_X1 U8993 ( .A1(n8847), .A2(n8852), .ZN(n8790) );
  NAND2_X1 U8994 ( .A1(n8857), .A2(n7296), .ZN(n8846) );
  NAND2_X1 U8995 ( .A1(n8846), .A2(n8852), .ZN(n7294) );
  NAND2_X1 U8996 ( .A1(n7294), .A2(n8790), .ZN(n8957) );
  AND2_X1 U8997 ( .A1(n7296), .A2(n7295), .ZN(n8850) );
  NAND3_X1 U8998 ( .A1(n8850), .A2(n8857), .A3(n8840), .ZN(n8954) );
  NAND2_X1 U8999 ( .A1(n8957), .A2(n8954), .ZN(n7297) );
  OAI21_X1 U9000 ( .B1(n7299), .B2(n7298), .A(n7460), .ZN(n7300) );
  NAND2_X1 U9001 ( .A1(n7300), .A2(n9402), .ZN(n7303) );
  NAND2_X1 U9002 ( .A1(n9028), .A2(n9003), .ZN(n7302) );
  NAND2_X1 U9003 ( .A1(n9026), .A2(n9140), .ZN(n7301) );
  AND2_X1 U9004 ( .A1(n7302), .A2(n7301), .ZN(n9657) );
  NAND2_X1 U9005 ( .A1(n7303), .A2(n9657), .ZN(n7328) );
  INV_X1 U9006 ( .A(n7328), .ZN(n7313) );
  OAI21_X1 U9007 ( .B1(n9028), .B2(n7306), .A(n7304), .ZN(n7305) );
  NAND2_X1 U9008 ( .A1(n7305), .A2(n8803), .ZN(n7417) );
  OAI21_X1 U9009 ( .B1(n7305), .B2(n8803), .A(n7417), .ZN(n7330) );
  NAND2_X1 U9010 ( .A1(n7330), .A2(n9901), .ZN(n7312) );
  AOI211_X1 U9011 ( .C1(n9664), .C2(n4690), .A(n9410), .B(n4687), .ZN(n7329)
         );
  NOR2_X1 U9012 ( .A1(n7333), .A2(n9897), .ZN(n7310) );
  OAI22_X1 U9013 ( .A1(n9416), .A2(n7308), .B1(n9666), .B2(n9413), .ZN(n7309)
         );
  AOI211_X1 U9014 ( .C1(n7329), .C2(n9380), .A(n7310), .B(n7309), .ZN(n7311)
         );
  OAI211_X1 U9015 ( .C1(n9421), .C2(n7313), .A(n7312), .B(n7311), .ZN(P1_U3283) );
  NAND2_X1 U9016 ( .A1(n7315), .A2(n7891), .ZN(n7316) );
  NAND2_X1 U9017 ( .A1(n7314), .A2(n7316), .ZN(n9971) );
  XOR2_X1 U9018 ( .A(n7317), .B(n7891), .Z(n7318) );
  NAND2_X1 U9019 ( .A1(n7318), .A2(n8391), .ZN(n7320) );
  AOI22_X1 U9020 ( .A1(n8388), .A2(n8106), .B1(n8104), .B2(n8386), .ZN(n7319)
         );
  OAI211_X1 U9021 ( .C1(n7365), .C2(n9971), .A(n7320), .B(n7319), .ZN(n9973)
         );
  NAND2_X1 U9022 ( .A1(n9973), .A2(n9645), .ZN(n7327) );
  INV_X1 U9023 ( .A(n7321), .ZN(n7322) );
  OAI22_X1 U9024 ( .A1(n9645), .A2(n7323), .B1(n7322), .B2(n9632), .ZN(n7324)
         );
  AOI21_X1 U9025 ( .B1(n8444), .B2(n7325), .A(n7324), .ZN(n7326) );
  OAI211_X1 U9026 ( .C1(n9971), .C2(n7371), .A(n7327), .B(n7326), .ZN(P2_U3224) );
  AOI211_X1 U9027 ( .C1(n7330), .C2(n9924), .A(n7329), .B(n7328), .ZN(n7336)
         );
  INV_X1 U9028 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U9029 ( .A1(n9664), .A2(n9503), .B1(n9929), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7331) );
  OAI21_X1 U9030 ( .B1(n7336), .B2(n9929), .A(n7331), .ZN(P1_U3532) );
  INV_X1 U9031 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7332) );
  OAI22_X1 U9032 ( .A1(n7333), .A2(n9551), .B1(n9927), .B2(n7332), .ZN(n7334)
         );
  INV_X1 U9033 ( .A(n7334), .ZN(n7335) );
  OAI21_X1 U9034 ( .B1(n7336), .B2(n9557), .A(n7335), .ZN(P1_U3483) );
  INV_X1 U9035 ( .A(n7337), .ZN(n7339) );
  OAI222_X1 U9036 ( .A1(n8588), .A2(n7339), .B1(n7916), .B2(P2_U3151), .C1(
        n10262), .C2(n4406), .ZN(P2_U3274) );
  OAI222_X1 U9037 ( .A1(P1_U3086), .A2(n4403), .B1(n9571), .B2(n7339), .C1(
        n7338), .C2(n9572), .ZN(P1_U3334) );
  XNOR2_X1 U9038 ( .A(n7368), .B(n7735), .ZN(n7382) );
  INV_X1 U9039 ( .A(n7342), .ZN(n7341) );
  AOI22_X1 U9040 ( .A1(n7343), .A2(n7361), .B1(n7341), .B2(n7340), .ZN(n7348)
         );
  NAND2_X1 U9041 ( .A1(n7342), .A2(n8106), .ZN(n7344) );
  AOI21_X1 U9042 ( .B1(n7361), .B2(n7344), .A(n7343), .ZN(n7346) );
  NOR2_X1 U9043 ( .A1(n7344), .A2(n7361), .ZN(n7345) );
  XNOR2_X1 U9044 ( .A(n7380), .B(n8104), .ZN(n7372) );
  XOR2_X1 U9045 ( .A(n7382), .B(n7372), .Z(n7356) );
  INV_X1 U9046 ( .A(n7350), .ZN(n7366) );
  OAI21_X1 U9047 ( .B1(n7841), .B2(n7361), .A(n7351), .ZN(n7352) );
  AOI21_X1 U9048 ( .B1(n7826), .B2(n8103), .A(n7352), .ZN(n7353) );
  OAI21_X1 U9049 ( .B1(n7366), .B2(n7714), .A(n7353), .ZN(n7354) );
  AOI21_X1 U9050 ( .B1(n7368), .B2(n7861), .A(n7354), .ZN(n7355) );
  OAI21_X1 U9051 ( .B1(n7356), .B2(n7856), .A(n7355), .ZN(P2_U3157) );
  AND2_X1 U9052 ( .A1(n7973), .A2(n7974), .ZN(n7896) );
  XNOR2_X1 U9053 ( .A(n7358), .B(n7896), .ZN(n9977) );
  XNOR2_X1 U9054 ( .A(n7360), .B(n7896), .ZN(n7363) );
  OAI22_X1 U9055 ( .A1(n7361), .A2(n9640), .B1(n7564), .B2(n9642), .ZN(n7362)
         );
  AOI21_X1 U9056 ( .B1(n7363), .B2(n8391), .A(n7362), .ZN(n7364) );
  OAI21_X1 U9057 ( .B1(n9977), .B2(n7365), .A(n7364), .ZN(n9979) );
  NAND2_X1 U9058 ( .A1(n9979), .A2(n9645), .ZN(n7370) );
  OAI22_X1 U9059 ( .A1(n9645), .A2(n7234), .B1(n7366), .B2(n9632), .ZN(n7367)
         );
  AOI21_X1 U9060 ( .B1(n7368), .B2(n8444), .A(n7367), .ZN(n7369) );
  OAI211_X1 U9061 ( .C1(n9977), .C2(n7371), .A(n7370), .B(n7369), .ZN(P2_U3223) );
  XNOR2_X1 U9062 ( .A(n7409), .B(n8103), .ZN(n7894) );
  XOR2_X1 U9063 ( .A(n7735), .B(n7894), .Z(n7384) );
  AOI22_X1 U9064 ( .A1(n7372), .A2(n7382), .B1(n7381), .B2(n7380), .ZN(n7373)
         );
  XOR2_X1 U9065 ( .A(n7384), .B(n7373), .Z(n7379) );
  INV_X1 U9066 ( .A(n7374), .ZN(n7407) );
  NOR2_X1 U9067 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10285), .ZN(n7450) );
  NOR2_X1 U9068 ( .A1(n7841), .A2(n7381), .ZN(n7375) );
  AOI211_X1 U9069 ( .C1(n7826), .C2(n8102), .A(n7450), .B(n7375), .ZN(n7376)
         );
  OAI21_X1 U9070 ( .B1(n7714), .B2(n7407), .A(n7376), .ZN(n7377) );
  AOI21_X1 U9071 ( .B1(n7409), .B2(n7861), .A(n7377), .ZN(n7378) );
  OAI21_X1 U9072 ( .B1(n7379), .B2(n7856), .A(n7378), .ZN(P2_U3176) );
  INV_X1 U9073 ( .A(n7380), .ZN(n7392) );
  INV_X1 U9074 ( .A(n7894), .ZN(n7402) );
  NAND2_X1 U9075 ( .A1(n7385), .A2(n7705), .ZN(n7386) );
  OAI211_X1 U9076 ( .C1(n7564), .C2(n7705), .A(n7402), .B(n7386), .ZN(n7390)
         );
  NAND2_X1 U9077 ( .A1(n7387), .A2(n7735), .ZN(n7388) );
  OAI211_X1 U9078 ( .C1(n7564), .C2(n7735), .A(n7894), .B(n7388), .ZN(n7389)
         );
  XOR2_X1 U9079 ( .A(n7735), .B(n9991), .Z(n7513) );
  XNOR2_X1 U9080 ( .A(n7513), .B(n8102), .ZN(n7393) );
  XNOR2_X1 U9081 ( .A(n7514), .B(n7393), .ZN(n7400) );
  INV_X1 U9082 ( .A(n7394), .ZN(n7565) );
  NOR2_X1 U9083 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7395), .ZN(n7532) );
  NOR2_X1 U9084 ( .A1(n7841), .A2(n7564), .ZN(n7396) );
  AOI211_X1 U9085 ( .C1(n7826), .C2(n8101), .A(n7532), .B(n7396), .ZN(n7397)
         );
  OAI21_X1 U9086 ( .B1(n7565), .B2(n7714), .A(n7397), .ZN(n7398) );
  AOI21_X1 U9087 ( .B1(n9991), .B2(n7861), .A(n7398), .ZN(n7399) );
  OAI21_X1 U9088 ( .B1(n7400), .B2(n7856), .A(n7399), .ZN(P2_U3164) );
  XNOR2_X1 U9089 ( .A(n7401), .B(n7402), .ZN(n9982) );
  XNOR2_X1 U9090 ( .A(n7403), .B(n7402), .ZN(n7404) );
  NAND2_X1 U9091 ( .A1(n7404), .A2(n8391), .ZN(n7406) );
  AOI22_X1 U9092 ( .A1(n8386), .A2(n8102), .B1(n8104), .B2(n8388), .ZN(n7405)
         );
  NAND2_X1 U9093 ( .A1(n7406), .A2(n7405), .ZN(n9983) );
  NAND2_X1 U9094 ( .A1(n9983), .A2(n9645), .ZN(n7411) );
  INV_X1 U9095 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7441) );
  OAI22_X1 U9096 ( .A1(n9645), .A2(n7441), .B1(n7407), .B2(n9632), .ZN(n7408)
         );
  AOI21_X1 U9097 ( .B1(n7409), .B2(n8444), .A(n7408), .ZN(n7410) );
  OAI211_X1 U9098 ( .C1(n9982), .C2(n8448), .A(n7411), .B(n7410), .ZN(P2_U3222) );
  INV_X1 U9099 ( .A(n9026), .ZN(n9670) );
  OR2_X1 U9100 ( .A1(n9693), .A2(n9670), .ZN(n8860) );
  NAND2_X1 U9101 ( .A1(n9693), .A2(n9670), .ZN(n8861) );
  AND2_X1 U9102 ( .A1(n8860), .A2(n8861), .ZN(n8806) );
  NAND2_X1 U9103 ( .A1(n7460), .A2(n8858), .ZN(n7412) );
  XOR2_X1 U9104 ( .A(n8806), .B(n7412), .Z(n7415) );
  OAI22_X1 U9105 ( .A1(n7466), .A2(n9667), .B1(n7413), .B2(n9669), .ZN(n9692)
         );
  INV_X1 U9106 ( .A(n9692), .ZN(n7414) );
  OAI21_X1 U9107 ( .B1(n7415), .B2(n9854), .A(n7414), .ZN(n7425) );
  INV_X1 U9108 ( .A(n7425), .ZN(n7424) );
  NAND2_X1 U9109 ( .A1(n7417), .A2(n7416), .ZN(n7463) );
  XOR2_X1 U9110 ( .A(n7463), .B(n8806), .Z(n7427) );
  NAND2_X1 U9111 ( .A1(n7427), .A2(n9901), .ZN(n7423) );
  AOI211_X1 U9112 ( .C1(n9693), .C2(n7418), .A(n9410), .B(n9866), .ZN(n7426)
         );
  NOR2_X1 U9113 ( .A1(n4689), .A2(n9897), .ZN(n7421) );
  OAI22_X1 U9114 ( .A1(n9416), .A2(n7419), .B1(n9695), .B2(n9413), .ZN(n7420)
         );
  AOI211_X1 U9115 ( .C1(n7426), .C2(n9380), .A(n7421), .B(n7420), .ZN(n7422)
         );
  OAI211_X1 U9116 ( .C1(n9421), .C2(n7424), .A(n7423), .B(n7422), .ZN(P1_U3282) );
  AOI211_X1 U9117 ( .C1(n7427), .C2(n9924), .A(n7426), .B(n7425), .ZN(n7432)
         );
  INV_X1 U9118 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9112) );
  AOI22_X1 U9119 ( .A1(n9693), .A2(n9503), .B1(n9929), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7428) );
  OAI21_X1 U9120 ( .B1(n7432), .B2(n9929), .A(n7428), .ZN(P1_U3533) );
  INV_X1 U9121 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7429) );
  OAI22_X1 U9122 ( .A1(n4689), .A2(n9551), .B1(n9927), .B2(n7429), .ZN(n7430)
         );
  INV_X1 U9123 ( .A(n7430), .ZN(n7431) );
  OAI21_X1 U9124 ( .B1(n7432), .B2(n9557), .A(n7431), .ZN(P1_U3486) );
  INV_X1 U9125 ( .A(n7433), .ZN(n7435) );
  OAI222_X1 U9126 ( .A1(n9572), .A2(n10282), .B1(n9571), .B2(n7435), .C1(
        P1_U3086), .C2(n7434), .ZN(P1_U3333) );
  OAI222_X1 U9127 ( .A1(n4406), .A2(n7436), .B1(n8588), .B2(n7435), .C1(
        P2_U3151), .C2(n7914), .ZN(P2_U3273) );
  INV_X1 U9128 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10008) );
  NOR2_X1 U9129 ( .A1(n10008), .A2(n7438), .ZN(n7491) );
  AOI21_X1 U9130 ( .B1(n10008), .B2(n7438), .A(n7491), .ZN(n7459) );
  NAND2_X1 U9131 ( .A1(n7443), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7439) );
  XNOR2_X1 U9132 ( .A(n7473), .B(n7490), .ZN(n7442) );
  NOR2_X1 U9133 ( .A1(n7441), .A2(n7442), .ZN(n7474) );
  AOI21_X1 U9134 ( .B1(n7442), .B2(n7441), .A(n7474), .ZN(n7456) );
  INV_X1 U9135 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U9136 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8253), .Z(n7480) );
  XNOR2_X1 U9137 ( .A(n7480), .B(n7490), .ZN(n7448) );
  OR2_X1 U9138 ( .A1(n7444), .A2(n7443), .ZN(n7446) );
  NAND2_X1 U9139 ( .A1(n7446), .A2(n7445), .ZN(n7447) );
  NAND2_X1 U9140 ( .A1(n7448), .A2(n7447), .ZN(n7482) );
  OAI21_X1 U9141 ( .B1(n7448), .B2(n7447), .A(n7482), .ZN(n7449) );
  NAND2_X1 U9142 ( .A1(n7449), .A2(n8226), .ZN(n7452) );
  INV_X1 U9143 ( .A(n7450), .ZN(n7451) );
  OAI211_X1 U9144 ( .C1(n8259), .C2(n10261), .A(n7452), .B(n7451), .ZN(n7453)
         );
  INV_X1 U9145 ( .A(n7453), .ZN(n7455) );
  NAND2_X1 U9146 ( .A1(n8261), .A2(n7490), .ZN(n7454) );
  OAI211_X1 U9147 ( .C1(n7456), .C2(n8270), .A(n7455), .B(n7454), .ZN(n7457)
         );
  INV_X1 U9148 ( .A(n7457), .ZN(n7458) );
  OAI21_X1 U9149 ( .B1(n7459), .B2(n8237), .A(n7458), .ZN(P2_U3193) );
  AND2_X1 U9150 ( .A1(n8861), .A2(n8858), .ZN(n8963) );
  NAND2_X1 U9151 ( .A1(n7461), .A2(n8860), .ZN(n9853) );
  NAND2_X1 U9152 ( .A1(n9861), .A2(n7466), .ZN(n8965) );
  NAND2_X1 U9153 ( .A1(n8862), .A2(n8965), .ZN(n9862) );
  INV_X1 U9154 ( .A(n9862), .ZN(n8807) );
  NAND2_X1 U9155 ( .A1(n9853), .A2(n8807), .ZN(n9857) );
  INV_X1 U9156 ( .A(n9024), .ZN(n9668) );
  OR2_X1 U9157 ( .A1(n9683), .A2(n9668), .ZN(n8967) );
  NAND2_X1 U9158 ( .A1(n9683), .A2(n9668), .ZN(n8966) );
  INV_X1 U9159 ( .A(n8808), .ZN(n7545) );
  XNOR2_X1 U9160 ( .A(n7546), .B(n7545), .ZN(n7462) );
  INV_X1 U9161 ( .A(n9023), .ZN(n7604) );
  OAI22_X1 U9162 ( .A1(n7466), .A2(n9669), .B1(n7604), .B2(n9667), .ZN(n9682)
         );
  AOI21_X1 U9163 ( .B1(n7462), .B2(n9402), .A(n9682), .ZN(n9920) );
  NAND2_X1 U9164 ( .A1(n7463), .A2(n4999), .ZN(n7465) );
  XNOR2_X1 U9165 ( .A(n7552), .B(n8808), .ZN(n9925) );
  NAND2_X1 U9166 ( .A1(n9925), .A2(n9901), .ZN(n7472) );
  INV_X1 U9167 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7467) );
  OAI22_X1 U9168 ( .A1(n9416), .A2(n7467), .B1(n9685), .B2(n9413), .ZN(n7470)
         );
  INV_X1 U9169 ( .A(n9683), .ZN(n9922) );
  NAND2_X1 U9170 ( .A1(n9915), .A2(n9866), .ZN(n9865) );
  INV_X1 U9171 ( .A(n9865), .ZN(n7468) );
  INV_X1 U9172 ( .A(n7553), .ZN(n7555) );
  OAI211_X1 U9173 ( .C1(n9922), .C2(n7468), .A(n7555), .B(n9864), .ZN(n9919)
         );
  NOR2_X1 U9174 ( .A1(n9919), .A2(n9345), .ZN(n7469) );
  AOI211_X1 U9175 ( .C1(n9872), .C2(n9683), .A(n7470), .B(n7469), .ZN(n7471)
         );
  OAI211_X1 U9176 ( .C1(n9421), .C2(n9920), .A(n7472), .B(n7471), .ZN(P1_U3280) );
  NOR2_X1 U9177 ( .A1(n7490), .A2(n7473), .ZN(n7475) );
  NAND2_X1 U9178 ( .A1(n7493), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7477) );
  INV_X1 U9179 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9180 ( .A1(n7542), .A2(n7566), .ZN(n7476) );
  NAND2_X1 U9181 ( .A1(n7477), .A2(n7476), .ZN(n7536) );
  INV_X1 U9182 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n9647) );
  AOI21_X1 U9183 ( .B1(n7478), .B2(n9647), .A(n8115), .ZN(n7503) );
  MUX2_X1 U9184 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8253), .Z(n8121) );
  XNOR2_X1 U9185 ( .A(n8132), .B(n8121), .ZN(n7486) );
  MUX2_X1 U9186 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8253), .Z(n7479) );
  OR2_X1 U9187 ( .A1(n7479), .A2(n7493), .ZN(n7484) );
  XNOR2_X1 U9188 ( .A(n7479), .B(n7542), .ZN(n7530) );
  INV_X1 U9189 ( .A(n7480), .ZN(n7481) );
  NAND2_X1 U9190 ( .A1(n7490), .A2(n7481), .ZN(n7483) );
  NAND2_X1 U9191 ( .A1(n7483), .A2(n7482), .ZN(n7529) );
  NAND2_X1 U9192 ( .A1(n7530), .A2(n7529), .ZN(n7528) );
  NAND2_X1 U9193 ( .A1(n7484), .A2(n7528), .ZN(n7485) );
  NAND2_X1 U9194 ( .A1(n7486), .A2(n7485), .ZN(n8123) );
  OAI21_X1 U9195 ( .B1(n7486), .B2(n7485), .A(n8123), .ZN(n7501) );
  INV_X1 U9196 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9197 ( .A1(n8261), .A2(n8132), .ZN(n7487) );
  OR2_X1 U9198 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5278), .ZN(n7518) );
  OAI211_X1 U9199 ( .C1(n8259), .C2(n7488), .A(n7487), .B(n7518), .ZN(n7500)
         );
  INV_X1 U9200 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9653) );
  NOR2_X1 U9201 ( .A1(n7490), .A2(n7489), .ZN(n7492) );
  NOR2_X1 U9202 ( .A1(n7492), .A2(n7491), .ZN(n7527) );
  NAND2_X1 U9203 ( .A1(n7493), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7496) );
  INV_X1 U9204 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9205 ( .A1(n7542), .A2(n7494), .ZN(n7495) );
  NAND2_X1 U9206 ( .A1(n7496), .A2(n7495), .ZN(n7526) );
  AOI21_X1 U9207 ( .B1(n9653), .B2(n7497), .A(n8133), .ZN(n7498) );
  NOR2_X1 U9208 ( .A1(n7498), .A2(n8237), .ZN(n7499) );
  AOI211_X1 U9209 ( .C1(n8226), .C2(n7501), .A(n7500), .B(n7499), .ZN(n7502)
         );
  OAI21_X1 U9210 ( .B1(n7503), .B2(n8270), .A(n7502), .ZN(P2_U3195) );
  NAND2_X1 U9211 ( .A1(n7507), .A2(n7504), .ZN(n7505) );
  OAI211_X1 U9212 ( .C1(n7506), .C2(n9572), .A(n7505), .B(n9010), .ZN(P1_U3332) );
  NAND2_X1 U9213 ( .A1(n7507), .A2(n8579), .ZN(n7510) );
  INV_X1 U9214 ( .A(n7508), .ZN(n7509) );
  NAND2_X1 U9215 ( .A1(n7509), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8093) );
  OAI211_X1 U9216 ( .C1(n7511), .C2(n4406), .A(n7510), .B(n8093), .ZN(P2_U3272) );
  XNOR2_X1 U9217 ( .A(n9631), .B(n7735), .ZN(n7512) );
  NAND2_X1 U9218 ( .A1(n7512), .A2(n7586), .ZN(n7579) );
  OAI21_X1 U9219 ( .B1(n7512), .B2(n7586), .A(n7579), .ZN(n7516) );
  AOI21_X1 U9220 ( .B1(n7516), .B2(n7515), .A(n7582), .ZN(n7523) );
  INV_X1 U9221 ( .A(n7517), .ZN(n9633) );
  OAI21_X1 U9222 ( .B1(n7841), .B2(n9639), .A(n7518), .ZN(n7519) );
  AOI21_X1 U9223 ( .B1(n7826), .B2(n8100), .A(n7519), .ZN(n7520) );
  OAI21_X1 U9224 ( .B1(n9633), .B2(n7714), .A(n7520), .ZN(n7521) );
  AOI21_X1 U9225 ( .B1(n9631), .B2(n7861), .A(n7521), .ZN(n7522) );
  OAI21_X1 U9226 ( .B1(n7523), .B2(n7856), .A(n7522), .ZN(P2_U3174) );
  INV_X1 U9227 ( .A(n7524), .ZN(n7525) );
  AOI21_X1 U9228 ( .B1(n7527), .B2(n7526), .A(n7525), .ZN(n7544) );
  INV_X1 U9229 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7535) );
  OAI21_X1 U9230 ( .B1(n7530), .B2(n7529), .A(n7528), .ZN(n7531) );
  NAND2_X1 U9231 ( .A1(n7531), .A2(n8226), .ZN(n7534) );
  INV_X1 U9232 ( .A(n7532), .ZN(n7533) );
  OAI211_X1 U9233 ( .C1(n8259), .C2(n7535), .A(n7534), .B(n7533), .ZN(n7541)
         );
  NAND2_X1 U9234 ( .A1(n7537), .A2(n7536), .ZN(n7538) );
  AOI21_X1 U9235 ( .B1(n7539), .B2(n7538), .A(n8270), .ZN(n7540) );
  AOI211_X1 U9236 ( .C1(n8261), .C2(n7542), .A(n7541), .B(n7540), .ZN(n7543)
         );
  OAI21_X1 U9237 ( .B1(n7544), .B2(n8237), .A(n7543), .ZN(P2_U3194) );
  OR2_X1 U9238 ( .A1(n7605), .A2(n7604), .ZN(n8968) );
  NAND2_X1 U9239 ( .A1(n7605), .A2(n7604), .ZN(n8875) );
  NAND2_X1 U9240 ( .A1(n8968), .A2(n8875), .ZN(n8810) );
  INV_X1 U9241 ( .A(n8966), .ZN(n8873) );
  NOR2_X1 U9242 ( .A1(n8810), .A2(n8873), .ZN(n8867) );
  INV_X1 U9243 ( .A(n8810), .ZN(n8872) );
  AOI21_X1 U9244 ( .B1(n7547), .B2(n8966), .A(n8872), .ZN(n7548) );
  NOR3_X1 U9245 ( .A1(n4466), .A2(n7548), .A3(n9854), .ZN(n7551) );
  NAND2_X1 U9246 ( .A1(n9171), .A2(n9140), .ZN(n7550) );
  NAND2_X1 U9247 ( .A1(n9024), .A2(n9003), .ZN(n7549) );
  NAND2_X1 U9248 ( .A1(n7550), .A2(n7549), .ZN(n8597) );
  OR2_X1 U9249 ( .A1(n7551), .A2(n8597), .ZN(n7573) );
  INV_X1 U9250 ( .A(n7573), .ZN(n7561) );
  XNOR2_X1 U9251 ( .A(n7603), .B(n8810), .ZN(n7575) );
  NAND2_X1 U9252 ( .A1(n7575), .A2(n9901), .ZN(n7560) );
  INV_X1 U9253 ( .A(n7605), .ZN(n8600) );
  INV_X1 U9254 ( .A(n7613), .ZN(n7554) );
  AOI211_X1 U9255 ( .C1(n7605), .C2(n7555), .A(n9410), .B(n7554), .ZN(n7574)
         );
  NOR2_X1 U9256 ( .A1(n8600), .A2(n9897), .ZN(n7558) );
  OAI22_X1 U9257 ( .A1(n9416), .A2(n7556), .B1(n8594), .B2(n9413), .ZN(n7557)
         );
  AOI211_X1 U9258 ( .C1(n7574), .C2(n9380), .A(n7558), .B(n7557), .ZN(n7559)
         );
  OAI211_X1 U9259 ( .C1(n9421), .C2(n7561), .A(n7560), .B(n7559), .ZN(P1_U3279) );
  INV_X1 U9260 ( .A(n7979), .ZN(n7898) );
  XNOR2_X1 U9261 ( .A(n7562), .B(n7898), .ZN(n7563) );
  OAI222_X1 U9262 ( .A1(n9642), .A2(n7586), .B1(n9640), .B2(n7564), .C1(n9637), 
        .C2(n7563), .ZN(n9989) );
  INV_X1 U9263 ( .A(n9989), .ZN(n7572) );
  OAI22_X1 U9264 ( .A1(n9645), .A2(n7566), .B1(n7565), .B2(n9632), .ZN(n7570)
         );
  NOR2_X1 U9265 ( .A1(n7567), .A2(n7979), .ZN(n9988) );
  INV_X1 U9266 ( .A(n7568), .ZN(n9987) );
  NOR3_X1 U9267 ( .A1(n9988), .A2(n9987), .A3(n8448), .ZN(n7569) );
  AOI211_X1 U9268 ( .C1(n8444), .C2(n9991), .A(n7570), .B(n7569), .ZN(n7571)
         );
  OAI21_X1 U9269 ( .B1(n9648), .B2(n7572), .A(n7571), .ZN(P2_U3221) );
  AOI211_X1 U9270 ( .C1(n7575), .C2(n9924), .A(n7574), .B(n7573), .ZN(n7578)
         );
  AOI22_X1 U9271 ( .A1(n7605), .A2(n9503), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9929), .ZN(n7576) );
  OAI21_X1 U9272 ( .B1(n7578), .B2(n9929), .A(n7576), .ZN(P1_U3536) );
  AOI22_X1 U9273 ( .A1(n7605), .A2(n9554), .B1(P1_REG0_REG_14__SCAN_IN), .B2(
        n9557), .ZN(n7577) );
  OAI21_X1 U9274 ( .B1(n7578), .B2(n9557), .A(n7577), .ZN(P1_U3495) );
  INV_X1 U9275 ( .A(n7627), .ZN(n7633) );
  INV_X1 U9276 ( .A(n7579), .ZN(n7581) );
  XNOR2_X1 U9277 ( .A(n7627), .B(n7735), .ZN(n7671) );
  XNOR2_X1 U9278 ( .A(n7671), .B(n8100), .ZN(n7580) );
  OAI21_X2 U9279 ( .B1(n7582), .B2(n7581), .A(n7580), .ZN(n7673) );
  INV_X1 U9280 ( .A(n7673), .ZN(n7584) );
  NOR3_X1 U9281 ( .A1(n7582), .A2(n7581), .A3(n7580), .ZN(n7583) );
  OAI21_X1 U9282 ( .B1(n7584), .B2(n7583), .A(n7839), .ZN(n7589) );
  NOR2_X1 U9283 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10192), .ZN(n8127) );
  AOI21_X1 U9284 ( .B1(n7826), .B2(n8099), .A(n8127), .ZN(n7585) );
  OAI21_X1 U9285 ( .B1(n7586), .B2(n7841), .A(n7585), .ZN(n7587) );
  AOI21_X1 U9286 ( .B1(n7631), .B2(n7851), .A(n7587), .ZN(n7588) );
  OAI211_X1 U9287 ( .C1(n7633), .C2(n7848), .A(n7589), .B(n7588), .ZN(P2_U3155) );
  INV_X1 U9288 ( .A(n7590), .ZN(n7594) );
  INV_X1 U9289 ( .A(n7591), .ZN(n7592) );
  OAI222_X1 U9290 ( .A1(n8588), .A2(n7594), .B1(P2_U3151), .B2(n7592), .C1(
        n10061), .C2(n4406), .ZN(P2_U3271) );
  OAI222_X1 U9291 ( .A1(n7595), .A2(P1_U3086), .B1(n9571), .B2(n7594), .C1(
        n7593), .C2(n9572), .ZN(P1_U3331) );
  INV_X1 U9292 ( .A(n7596), .ZN(n7601) );
  INV_X1 U9293 ( .A(n7597), .ZN(n7599) );
  OAI222_X1 U9294 ( .A1(n8588), .A2(n7601), .B1(P2_U3151), .B2(n7599), .C1(
        n7598), .C2(n4406), .ZN(P2_U3270) );
  OAI222_X1 U9295 ( .A1(n7602), .A2(P1_U3086), .B1(n9575), .B2(n7601), .C1(
        n7600), .C2(n9572), .ZN(P1_U3330) );
  INV_X1 U9296 ( .A(n9171), .ZN(n9167) );
  OR2_X1 U9297 ( .A1(n9555), .A2(n9167), .ZN(n8971) );
  NAND2_X1 U9298 ( .A1(n9555), .A2(n9167), .ZN(n8876) );
  NAND2_X1 U9299 ( .A1(n8971), .A2(n8876), .ZN(n8789) );
  XNOR2_X1 U9300 ( .A(n9169), .B(n8789), .ZN(n9502) );
  INV_X1 U9301 ( .A(n9502), .ZN(n7619) );
  INV_X1 U9302 ( .A(n9901), .ZN(n9398) );
  INV_X1 U9303 ( .A(n8968), .ZN(n7607) );
  OAI21_X1 U9304 ( .B1(n4466), .B2(n7607), .A(n8789), .ZN(n7609) );
  NOR2_X1 U9305 ( .A1(n8789), .A2(n7607), .ZN(n7608) );
  AOI21_X1 U9306 ( .B1(n7609), .B2(n8769), .A(n9854), .ZN(n7612) );
  NAND2_X1 U9307 ( .A1(n9172), .A2(n9140), .ZN(n7611) );
  NAND2_X1 U9308 ( .A1(n9023), .A2(n9003), .ZN(n7610) );
  NAND2_X1 U9309 ( .A1(n7611), .A2(n7610), .ZN(n8749) );
  OR2_X1 U9310 ( .A1(n7612), .A2(n8749), .ZN(n9500) );
  INV_X1 U9311 ( .A(n9555), .ZN(n9168) );
  AOI211_X1 U9312 ( .C1(n9555), .C2(n7613), .A(n9410), .B(n9407), .ZN(n9501)
         );
  NAND2_X1 U9313 ( .A1(n9501), .A2(n9380), .ZN(n7616) );
  INV_X1 U9314 ( .A(n8746), .ZN(n7614) );
  AOI22_X1 U9315 ( .A1(n9904), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n7614), .B2(
        n9894), .ZN(n7615) );
  OAI211_X1 U9316 ( .C1(n9168), .C2(n9897), .A(n7616), .B(n7615), .ZN(n7617)
         );
  AOI21_X1 U9317 ( .B1(n9416), .B2(n9500), .A(n7617), .ZN(n7618) );
  OAI21_X1 U9318 ( .B1(n7619), .B2(n9398), .A(n7618), .ZN(P1_U3278) );
  XNOR2_X1 U9319 ( .A(n7621), .B(n7991), .ZN(n7638) );
  INV_X1 U9320 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7624) );
  XNOR2_X1 U9321 ( .A(n7622), .B(n4652), .ZN(n7623) );
  AOI222_X1 U9322 ( .A1(n8391), .A2(n7623), .B1(n8099), .B2(n8386), .C1(n8101), 
        .C2(n8388), .ZN(n7630) );
  MUX2_X1 U9323 ( .A(n7624), .B(n7630), .S(n9993), .Z(n7626) );
  NAND2_X1 U9324 ( .A1(n7627), .A2(n8568), .ZN(n7625) );
  OAI211_X1 U9325 ( .C1(n7638), .C2(n8572), .A(n7626), .B(n7625), .ZN(P2_U3432) );
  NAND2_X1 U9326 ( .A1(n10012), .A2(n9968), .ZN(n8500) );
  INV_X1 U9327 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8135) );
  MUX2_X1 U9328 ( .A(n8135), .B(n7630), .S(n10012), .Z(n7629) );
  INV_X1 U9329 ( .A(n8460), .ZN(n8497) );
  NAND2_X1 U9330 ( .A1(n7627), .A2(n8497), .ZN(n7628) );
  OAI211_X1 U9331 ( .C1(n7638), .C2(n8500), .A(n7629), .B(n7628), .ZN(P2_U3473) );
  INV_X1 U9332 ( .A(n7630), .ZN(n7635) );
  INV_X1 U9333 ( .A(n7631), .ZN(n7632) );
  OAI22_X1 U9334 ( .A1(n7633), .A2(n8331), .B1(n7632), .B2(n9632), .ZN(n7634)
         );
  OAI21_X1 U9335 ( .B1(n7635), .B2(n7634), .A(n9645), .ZN(n7637) );
  NAND2_X1 U9336 ( .A1(n9648), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7636) );
  OAI211_X1 U9337 ( .C1(n7638), .C2(n8448), .A(n7637), .B(n7636), .ZN(P2_U3219) );
  INV_X1 U9338 ( .A(n7639), .ZN(n9574) );
  INV_X1 U9339 ( .A(n7640), .ZN(n7642) );
  OAI222_X1 U9340 ( .A1(n8588), .A2(n9574), .B1(P2_U3151), .B2(n7642), .C1(
        n7641), .C2(n4406), .ZN(P2_U3269) );
  NAND2_X1 U9341 ( .A1(n7643), .A2(n7992), .ZN(n7644) );
  NAND3_X1 U9342 ( .A1(n7645), .A2(n8391), .A3(n7644), .ZN(n7648) );
  OAI22_X1 U9343 ( .A1(n9641), .A2(n9640), .B1(n8418), .B2(n9642), .ZN(n7646)
         );
  INV_X1 U9344 ( .A(n7646), .ZN(n7647) );
  NAND2_X1 U9345 ( .A1(n7648), .A2(n7647), .ZN(n8440) );
  MUX2_X1 U9346 ( .A(n8440), .B(P2_REG1_REG_15__SCAN_IN), .S(n10010), .Z(n7652) );
  XNOR2_X1 U9347 ( .A(n7650), .B(n7992), .ZN(n8449) );
  INV_X1 U9348 ( .A(n8445), .ZN(n7653) );
  OAI22_X1 U9349 ( .A1(n8449), .A2(n8500), .B1(n7653), .B2(n8460), .ZN(n7651)
         );
  OR2_X1 U9350 ( .A1(n7652), .A2(n7651), .ZN(P2_U3474) );
  MUX2_X1 U9351 ( .A(n8440), .B(P2_REG0_REG_15__SCAN_IN), .S(n9994), .Z(n7655)
         );
  OAI22_X1 U9352 ( .A1(n8449), .A2(n8572), .B1(n7653), .B2(n8516), .ZN(n7654)
         );
  OR2_X1 U9353 ( .A1(n7655), .A2(n7654), .ZN(P2_U3435) );
  INV_X1 U9354 ( .A(n8761), .ZN(n9569) );
  OAI222_X1 U9355 ( .A1(n8588), .A2(n9569), .B1(n7657), .B2(P2_U3151), .C1(
        n7656), .C2(n4406), .ZN(P2_U3266) );
  INV_X1 U9356 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8622) );
  INV_X1 U9357 ( .A(n8621), .ZN(n8583) );
  OAI222_X1 U9358 ( .A1(n9572), .A2(n8622), .B1(n9575), .B2(n8583), .C1(n5801), 
        .C2(P1_U3086), .ZN(P1_U3327) );
  INV_X1 U9359 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7863) );
  NAND2_X1 U9360 ( .A1(n7658), .A2(SI_29_), .ZN(n7663) );
  INV_X1 U9361 ( .A(n7659), .ZN(n7661) );
  NAND2_X1 U9362 ( .A1(n7661), .A2(n7660), .ZN(n7662) );
  INV_X1 U9363 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10221) );
  MUX2_X1 U9364 ( .A(n7863), .B(n10221), .S(n7868), .Z(n7665) );
  INV_X1 U9365 ( .A(SI_30_), .ZN(n7664) );
  NAND2_X1 U9366 ( .A1(n7665), .A2(n7664), .ZN(n7865) );
  INV_X1 U9367 ( .A(n7665), .ZN(n7666) );
  NAND2_X1 U9368 ( .A1(n7666), .A2(SI_30_), .ZN(n7667) );
  NAND2_X1 U9369 ( .A1(n7865), .A2(n7667), .ZN(n7866) );
  INV_X1 U9370 ( .A(n8752), .ZN(n7670) );
  OAI222_X1 U9371 ( .A1(n4406), .A2(n7863), .B1(n8588), .B2(n7670), .C1(
        P2_U3151), .C2(n7668), .ZN(P2_U3265) );
  OAI222_X1 U9372 ( .A1(n9572), .A2(n10221), .B1(n9575), .B2(n7670), .C1(
        P1_U3086), .C2(n7669), .ZN(P1_U3325) );
  INV_X1 U9373 ( .A(n8299), .ZN(n8517) );
  XNOR2_X1 U9374 ( .A(n8467), .B(n7735), .ZN(n7703) );
  XNOR2_X1 U9375 ( .A(n8490), .B(n7735), .ZN(n7681) );
  NAND2_X1 U9376 ( .A1(n7671), .A2(n9641), .ZN(n7672) );
  XNOR2_X1 U9377 ( .A(n8445), .B(n7735), .ZN(n7674) );
  XNOR2_X1 U9378 ( .A(n7674), .B(n8432), .ZN(n7858) );
  INV_X1 U9379 ( .A(n7674), .ZN(n7675) );
  XNOR2_X1 U9380 ( .A(n8569), .B(n7735), .ZN(n7676) );
  NAND2_X1 U9381 ( .A1(n7676), .A2(n8418), .ZN(n7677) );
  OAI21_X1 U9382 ( .B1(n7676), .B2(n8418), .A(n7677), .ZN(n7765) );
  INV_X1 U9383 ( .A(n7677), .ZN(n7775) );
  XNOR2_X1 U9384 ( .A(n8562), .B(n7735), .ZN(n7678) );
  NAND2_X1 U9385 ( .A1(n7678), .A2(n8433), .ZN(n7813) );
  INV_X1 U9386 ( .A(n7678), .ZN(n7679) );
  NAND2_X1 U9387 ( .A1(n7679), .A2(n8097), .ZN(n7680) );
  AND2_X1 U9388 ( .A1(n7813), .A2(n7680), .ZN(n7774) );
  XNOR2_X1 U9389 ( .A(n7681), .B(n8419), .ZN(n7814) );
  XNOR2_X1 U9390 ( .A(n8485), .B(n7735), .ZN(n7683) );
  XNOR2_X1 U9391 ( .A(n7683), .B(n8379), .ZN(n7725) );
  XNOR2_X1 U9392 ( .A(n8553), .B(n7705), .ZN(n7682) );
  NOR2_X1 U9393 ( .A1(n7682), .A2(n8387), .ZN(n7744) );
  AOI21_X1 U9394 ( .B1(n7682), .B2(n8387), .A(n7744), .ZN(n7793) );
  INV_X1 U9395 ( .A(n7683), .ZN(n7684) );
  NAND2_X1 U9396 ( .A1(n7684), .A2(n8379), .ZN(n7794) );
  INV_X1 U9397 ( .A(n7744), .ZN(n7685) );
  XNOR2_X1 U9398 ( .A(n8548), .B(n7735), .ZN(n7687) );
  NAND2_X1 U9399 ( .A1(n7687), .A2(n7686), .ZN(n7691) );
  INV_X1 U9400 ( .A(n7687), .ZN(n7688) );
  NAND2_X1 U9401 ( .A1(n7688), .A2(n8378), .ZN(n7689) );
  AND2_X1 U9402 ( .A1(n7691), .A2(n7689), .ZN(n7743) );
  NAND2_X1 U9403 ( .A1(n7690), .A2(n7743), .ZN(n7745) );
  NAND2_X1 U9404 ( .A1(n7745), .A2(n7691), .ZN(n7804) );
  XNOR2_X1 U9405 ( .A(n7812), .B(n7735), .ZN(n7692) );
  XNOR2_X1 U9406 ( .A(n7692), .B(n8342), .ZN(n7805) );
  NAND2_X1 U9407 ( .A1(n7804), .A2(n7805), .ZN(n7803) );
  INV_X1 U9408 ( .A(n7692), .ZN(n7693) );
  NAND2_X1 U9409 ( .A1(n7693), .A2(n8342), .ZN(n7694) );
  NAND2_X1 U9410 ( .A1(n7803), .A2(n7694), .ZN(n7698) );
  INV_X1 U9411 ( .A(n7698), .ZN(n7696) );
  XNOR2_X1 U9412 ( .A(n8474), .B(n7735), .ZN(n7697) );
  INV_X1 U9413 ( .A(n7697), .ZN(n7695) );
  NAND2_X1 U9414 ( .A1(n7718), .A2(n7783), .ZN(n7702) );
  XNOR2_X1 U9415 ( .A(n8532), .B(n7735), .ZN(n7699) );
  NAND2_X1 U9416 ( .A1(n7699), .A2(n8343), .ZN(n7755) );
  INV_X1 U9417 ( .A(n7699), .ZN(n7700) );
  NAND2_X1 U9418 ( .A1(n7700), .A2(n8096), .ZN(n7701) );
  NAND2_X1 U9419 ( .A1(n7702), .A2(n7784), .ZN(n7754) );
  NAND2_X1 U9420 ( .A1(n7754), .A2(n7755), .ZN(n7704) );
  XNOR2_X1 U9421 ( .A(n7703), .B(n8329), .ZN(n7756) );
  XNOR2_X1 U9422 ( .A(n8523), .B(n7705), .ZN(n7706) );
  INV_X1 U9423 ( .A(n7706), .ZN(n7707) );
  NAND2_X1 U9424 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  XNOR2_X1 U9425 ( .A(n8299), .B(n7735), .ZN(n7732) );
  XNOR2_X1 U9426 ( .A(n7732), .B(n7843), .ZN(n7710) );
  AOI21_X1 U9427 ( .B1(n7711), .B2(n7710), .A(n7856), .ZN(n7712) );
  INV_X1 U9428 ( .A(n8298), .ZN(n7715) );
  AOI22_X1 U9429 ( .A1(n8095), .A2(n7850), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7713) );
  OAI21_X1 U9430 ( .B1(n7715), .B2(n7714), .A(n7713), .ZN(n7716) );
  AOI21_X1 U9431 ( .B1(n7826), .B2(n8295), .A(n7716), .ZN(n7717) );
  INV_X1 U9432 ( .A(n7718), .ZN(n7786) );
  AOI21_X1 U9433 ( .B1(n8356), .B2(n7719), .A(n7786), .ZN(n7724) );
  AOI22_X1 U9434 ( .A1(n8367), .A2(n7850), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7721) );
  NAND2_X1 U9435 ( .A1(n8344), .A2(n7851), .ZN(n7720) );
  OAI211_X1 U9436 ( .C1(n8343), .C2(n7854), .A(n7721), .B(n7720), .ZN(n7722)
         );
  AOI21_X1 U9437 ( .B1(n8474), .B2(n7861), .A(n7722), .ZN(n7723) );
  OAI21_X1 U9438 ( .B1(n7724), .B2(n7856), .A(n7723), .ZN(P2_U3156) );
  INV_X1 U9439 ( .A(n8485), .ZN(n7731) );
  OAI211_X1 U9440 ( .C1(n7726), .C2(n7725), .A(n7795), .B(n7839), .ZN(n7730)
         );
  NAND2_X1 U9441 ( .A1(n7826), .A2(n8387), .ZN(n7727) );
  NAND2_X1 U9442 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8258) );
  OAI211_X1 U9443 ( .C1(n8419), .C2(n7841), .A(n7727), .B(n8258), .ZN(n7728)
         );
  AOI21_X1 U9444 ( .B1(n8396), .B2(n7851), .A(n7728), .ZN(n7729) );
  OAI211_X1 U9445 ( .C1(n7731), .C2(n7848), .A(n7730), .B(n7729), .ZN(P2_U3159) );
  INV_X1 U9446 ( .A(n7732), .ZN(n7733) );
  XNOR2_X1 U9447 ( .A(n8279), .B(n7735), .ZN(n7736) );
  NAND2_X1 U9448 ( .A1(n8282), .A2(n7826), .ZN(n7738) );
  AOI22_X1 U9449 ( .A1(n8287), .A2(n7851), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7737) );
  OAI211_X1 U9450 ( .C1(n7843), .C2(n7841), .A(n7738), .B(n7737), .ZN(n7739)
         );
  AOI21_X1 U9451 ( .B1(n8511), .B2(n7861), .A(n7739), .ZN(n7740) );
  OAI21_X1 U9452 ( .B1(n7741), .B2(n7856), .A(n7740), .ZN(P2_U3160) );
  INV_X1 U9453 ( .A(n8548), .ZN(n7753) );
  INV_X1 U9454 ( .A(n7742), .ZN(n7797) );
  NOR3_X1 U9455 ( .A1(n7797), .A2(n7744), .A3(n7743), .ZN(n7747) );
  INV_X1 U9456 ( .A(n7745), .ZN(n7746) );
  OAI21_X1 U9457 ( .B1(n7747), .B2(n7746), .A(n7839), .ZN(n7752) );
  AOI22_X1 U9458 ( .A1(n8367), .A2(n7826), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7748) );
  OAI21_X1 U9459 ( .B1(n7749), .B2(n7841), .A(n7748), .ZN(n7750) );
  AOI21_X1 U9460 ( .B1(n8370), .B2(n7851), .A(n7750), .ZN(n7751) );
  OAI211_X1 U9461 ( .C1(n7753), .C2(n7848), .A(n7752), .B(n7751), .ZN(P2_U3163) );
  INV_X1 U9462 ( .A(n8467), .ZN(n8319) );
  INV_X1 U9463 ( .A(n7754), .ZN(n7787) );
  INV_X1 U9464 ( .A(n7755), .ZN(n7757) );
  NOR3_X1 U9465 ( .A1(n7787), .A2(n7757), .A3(n7756), .ZN(n7760) );
  INV_X1 U9466 ( .A(n7758), .ZN(n7759) );
  OAI21_X1 U9467 ( .B1(n7760), .B2(n7759), .A(n7839), .ZN(n7764) );
  AOI22_X1 U9468 ( .A1(n8096), .A2(n7850), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7761) );
  OAI21_X1 U9469 ( .B1(n8316), .B2(n7854), .A(n7761), .ZN(n7762) );
  AOI21_X1 U9470 ( .B1(n8317), .B2(n7851), .A(n7762), .ZN(n7763) );
  OAI211_X1 U9471 ( .C1(n8319), .C2(n7848), .A(n7764), .B(n7763), .ZN(P2_U3165) );
  INV_X1 U9472 ( .A(n8569), .ZN(n7773) );
  OAI21_X1 U9473 ( .B1(n7855), .B2(n7766), .A(n7765), .ZN(n7767) );
  INV_X1 U9474 ( .A(n7767), .ZN(n7768) );
  OAI21_X1 U9475 ( .B1(n4468), .B2(n7768), .A(n7839), .ZN(n7772) );
  NAND2_X1 U9476 ( .A1(n7826), .A2(n8097), .ZN(n7769) );
  NAND2_X1 U9477 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8181) );
  OAI211_X1 U9478 ( .C1(n8432), .C2(n7841), .A(n7769), .B(n8181), .ZN(n7770)
         );
  AOI21_X1 U9479 ( .B1(n8437), .B2(n7851), .A(n7770), .ZN(n7771) );
  OAI211_X1 U9480 ( .C1(n7773), .C2(n7848), .A(n7772), .B(n7771), .ZN(P2_U3166) );
  INV_X1 U9481 ( .A(n8562), .ZN(n7782) );
  INV_X1 U9482 ( .A(n7815), .ZN(n7777) );
  NOR3_X1 U9483 ( .A1(n4468), .A2(n7775), .A3(n7774), .ZN(n7776) );
  OAI21_X1 U9484 ( .B1(n7777), .B2(n7776), .A(n7839), .ZN(n7781) );
  NAND2_X1 U9485 ( .A1(n7826), .A2(n8389), .ZN(n7778) );
  NAND2_X1 U9486 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8207) );
  OAI211_X1 U9487 ( .C1(n8418), .C2(n7841), .A(n7778), .B(n8207), .ZN(n7779)
         );
  AOI21_X1 U9488 ( .B1(n8424), .B2(n7851), .A(n7779), .ZN(n7780) );
  OAI211_X1 U9489 ( .C1(n7782), .C2(n7848), .A(n7781), .B(n7780), .ZN(P2_U3168) );
  INV_X1 U9490 ( .A(n8532), .ZN(n8332) );
  INV_X1 U9491 ( .A(n7783), .ZN(n7785) );
  NOR3_X1 U9492 ( .A1(n7786), .A2(n7785), .A3(n7784), .ZN(n7788) );
  OAI21_X1 U9493 ( .B1(n7788), .B2(n7787), .A(n7839), .ZN(n7792) );
  AOI22_X1 U9494 ( .A1(n8329), .A2(n7826), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7789) );
  OAI21_X1 U9495 ( .B1(n7808), .B2(n7841), .A(n7789), .ZN(n7790) );
  AOI21_X1 U9496 ( .B1(n8334), .B2(n7851), .A(n7790), .ZN(n7791) );
  OAI211_X1 U9497 ( .C1(n8332), .C2(n7848), .A(n7792), .B(n7791), .ZN(P2_U3169) );
  INV_X1 U9498 ( .A(n8553), .ZN(n7802) );
  AOI21_X1 U9499 ( .B1(n7795), .B2(n7794), .A(n7793), .ZN(n7796) );
  OAI21_X1 U9500 ( .B1(n7797), .B2(n7796), .A(n7839), .ZN(n7801) );
  AOI22_X1 U9501 ( .A1(n8378), .A2(n7826), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7798) );
  OAI21_X1 U9502 ( .B1(n8403), .B2(n7841), .A(n7798), .ZN(n7799) );
  AOI21_X1 U9503 ( .B1(n8382), .B2(n7851), .A(n7799), .ZN(n7800) );
  OAI211_X1 U9504 ( .C1(n7802), .C2(n7848), .A(n7801), .B(n7800), .ZN(P2_U3173) );
  OAI21_X1 U9505 ( .B1(n7805), .B2(n7804), .A(n7803), .ZN(n7806) );
  NAND2_X1 U9506 ( .A1(n7806), .A2(n7839), .ZN(n7811) );
  AOI22_X1 U9507 ( .A1(n8378), .A2(n7850), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7807) );
  OAI21_X1 U9508 ( .B1(n7808), .B2(n7854), .A(n7807), .ZN(n7809) );
  AOI21_X1 U9509 ( .B1(n8359), .B2(n7851), .A(n7809), .ZN(n7810) );
  OAI211_X1 U9510 ( .C1(n7812), .C2(n7848), .A(n7811), .B(n7810), .ZN(P2_U3175) );
  INV_X1 U9511 ( .A(n8490), .ZN(n7822) );
  AND3_X1 U9512 ( .A1(n7815), .A2(n7814), .A3(n7813), .ZN(n7816) );
  OAI21_X1 U9513 ( .B1(n7817), .B2(n7816), .A(n7839), .ZN(n7821) );
  NAND2_X1 U9514 ( .A1(n7826), .A2(n8379), .ZN(n7818) );
  NAND2_X1 U9515 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8228) );
  OAI211_X1 U9516 ( .C1(n8433), .C2(n7841), .A(n7818), .B(n8228), .ZN(n7819)
         );
  AOI21_X1 U9517 ( .B1(n8408), .B2(n7851), .A(n7819), .ZN(n7820) );
  OAI211_X1 U9518 ( .C1(n7822), .C2(n7848), .A(n7821), .B(n7820), .ZN(P2_U3178) );
  OAI211_X1 U9519 ( .C1(n7825), .C2(n7824), .A(n7823), .B(n7839), .ZN(n7836)
         );
  NAND2_X1 U9520 ( .A1(n7826), .A2(n8107), .ZN(n7828) );
  OAI211_X1 U9521 ( .C1(n7829), .C2(n7841), .A(n7828), .B(n7827), .ZN(n7830)
         );
  INV_X1 U9522 ( .A(n7830), .ZN(n7835) );
  NAND2_X1 U9523 ( .A1(n7861), .A2(n7831), .ZN(n7834) );
  NAND2_X1 U9524 ( .A1(n7851), .A2(n7832), .ZN(n7833) );
  NAND4_X1 U9525 ( .A1(n7836), .A2(n7835), .A3(n7834), .A4(n7833), .ZN(
        P2_U3179) );
  INV_X1 U9526 ( .A(n8523), .ZN(n7849) );
  OAI21_X1 U9527 ( .B1(n8316), .B2(n7838), .A(n7837), .ZN(n7840) );
  NAND2_X1 U9528 ( .A1(n7840), .A2(n7839), .ZN(n7847) );
  OAI22_X1 U9529 ( .A1(n7842), .A2(n7841), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10055), .ZN(n7845) );
  NOR2_X1 U9530 ( .A1(n7843), .A2(n7854), .ZN(n7844) );
  AOI211_X1 U9531 ( .C1(n8307), .C2(n7851), .A(n7845), .B(n7844), .ZN(n7846)
         );
  OAI211_X1 U9532 ( .C1(n7849), .C2(n7848), .A(n7847), .B(n7846), .ZN(P2_U3180) );
  INV_X1 U9533 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10269) );
  NOR2_X1 U9534 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10269), .ZN(n8153) );
  AOI21_X1 U9535 ( .B1(n7850), .B2(n8100), .A(n8153), .ZN(n7853) );
  NAND2_X1 U9536 ( .A1(n7851), .A2(n8442), .ZN(n7852) );
  OAI211_X1 U9537 ( .C1(n7854), .C2(n8418), .A(n7853), .B(n7852), .ZN(n7860)
         );
  AOI211_X1 U9538 ( .C1(n7858), .C2(n7857), .A(n7856), .B(n7855), .ZN(n7859)
         );
  AOI211_X1 U9539 ( .C1(n8445), .C2(n7861), .A(n7860), .B(n7859), .ZN(n7862)
         );
  INV_X1 U9540 ( .A(n7862), .ZN(P2_U3181) );
  NOR2_X1 U9541 ( .A1(n7873), .A2(n7863), .ZN(n7864) );
  INV_X1 U9542 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8575) );
  MUX2_X1 U9543 ( .A(n8575), .B(n10064), .S(n7868), .Z(n7869) );
  XNOR2_X1 U9544 ( .A(n7869), .B(SI_31_), .ZN(n7870) );
  NAND2_X1 U9545 ( .A1(n9559), .A2(n7872), .ZN(n7875) );
  OR2_X1 U9546 ( .A1(n7873), .A2(n8575), .ZN(n7874) );
  OAI22_X1 U9547 ( .A1(n7877), .A2(n7876), .B1(n8454), .B2(n8501), .ZN(n7880)
         );
  INV_X1 U9548 ( .A(n8454), .ZN(n8506) );
  NAND2_X1 U9549 ( .A1(n8506), .A2(n7879), .ZN(n8067) );
  AND2_X1 U9550 ( .A1(n8067), .A2(n7878), .ZN(n8075) );
  NAND2_X1 U9551 ( .A1(n8071), .A2(n8075), .ZN(n7881) );
  OR2_X1 U9552 ( .A1(n8506), .A2(n7879), .ZN(n8068) );
  INV_X1 U9553 ( .A(n7881), .ZN(n7907) );
  AND2_X1 U9554 ( .A1(n8068), .A2(n8057), .ZN(n8058) );
  INV_X1 U9555 ( .A(n8037), .ZN(n8029) );
  INV_X1 U9556 ( .A(n8030), .ZN(n7882) );
  NAND2_X1 U9557 ( .A1(n7884), .A2(n7883), .ZN(n9635) );
  NOR4_X1 U9558 ( .A1(n7887), .A2(n7913), .A3(n7886), .A4(n7885), .ZN(n7888)
         );
  NAND4_X1 U9559 ( .A1(n7890), .A2(n7926), .A3(n7889), .A4(n7888), .ZN(n7893)
         );
  NOR4_X1 U9560 ( .A1(n7893), .A2(n7957), .A3(n7892), .A4(n7891), .ZN(n7895)
         );
  NAND4_X1 U9561 ( .A1(n9635), .A2(n7896), .A3(n7895), .A4(n7894), .ZN(n7897)
         );
  NOR4_X1 U9562 ( .A1(n7899), .A2(n7898), .A3(n4652), .A4(n7897), .ZN(n7900)
         );
  NAND4_X1 U9563 ( .A1(n5653), .A2(n8416), .A3(n8430), .A4(n7900), .ZN(n7901)
         );
  NOR4_X1 U9564 ( .A1(n8363), .A2(n7902), .A3(n8376), .A4(n7901), .ZN(n7903)
         );
  NAND4_X1 U9565 ( .A1(n8339), .A2(n8354), .A3(n8328), .A4(n7903), .ZN(n7904)
         );
  NOR4_X1 U9566 ( .A1(n8291), .A2(n7905), .A3(n8302), .A4(n7904), .ZN(n7906)
         );
  NAND4_X1 U9567 ( .A1(n7907), .A2(n8058), .A3(n7906), .A4(n8279), .ZN(n7908)
         );
  NAND2_X1 U9568 ( .A1(n7908), .A2(n7916), .ZN(n7909) );
  INV_X1 U9569 ( .A(n7915), .ZN(n7912) );
  NAND2_X1 U9570 ( .A1(n7923), .A2(n8070), .ZN(n7921) );
  OAI21_X1 U9571 ( .B1(n7913), .B2(n7912), .A(n7921), .ZN(n7920) );
  NAND2_X1 U9572 ( .A1(n7915), .A2(n7914), .ZN(n7918) );
  MUX2_X1 U9573 ( .A(n7918), .B(n7917), .S(n7916), .Z(n7919) );
  NAND2_X1 U9574 ( .A1(n7920), .A2(n7919), .ZN(n7928) );
  INV_X1 U9575 ( .A(n7921), .ZN(n7925) );
  INV_X1 U9576 ( .A(n7922), .ZN(n7924) );
  AOI22_X1 U9577 ( .A1(n7925), .A2(n7924), .B1(n8066), .B2(n4802), .ZN(n7927)
         );
  NAND3_X1 U9578 ( .A1(n7928), .A2(n7927), .A3(n7926), .ZN(n7935) );
  NAND2_X1 U9579 ( .A1(n8112), .A2(n5071), .ZN(n7929) );
  NAND2_X1 U9580 ( .A1(n7944), .A2(n7929), .ZN(n7932) );
  NAND2_X1 U9581 ( .A1(n7938), .A2(n7930), .ZN(n7931) );
  MUX2_X1 U9582 ( .A(n7932), .B(n7931), .S(n8070), .Z(n7933) );
  INV_X1 U9583 ( .A(n7933), .ZN(n7934) );
  NAND2_X1 U9584 ( .A1(n7935), .A2(n7934), .ZN(n7937) );
  NAND2_X1 U9585 ( .A1(n7937), .A2(n7936), .ZN(n7948) );
  INV_X1 U9586 ( .A(n7938), .ZN(n7940) );
  OAI211_X1 U9587 ( .C1(n7948), .C2(n7940), .A(n7951), .B(n7939), .ZN(n7943)
         );
  NAND2_X1 U9588 ( .A1(n7945), .A2(n7941), .ZN(n7942) );
  NAND3_X1 U9589 ( .A1(n7943), .A2(n7949), .A3(n7942), .ZN(n7954) );
  INV_X1 U9590 ( .A(n7944), .ZN(n7947) );
  OAI211_X1 U9591 ( .C1(n7948), .C2(n7947), .A(n5642), .B(n7946), .ZN(n7952)
         );
  INV_X1 U9592 ( .A(n7949), .ZN(n7950) );
  AOI21_X1 U9593 ( .B1(n7952), .B2(n7951), .A(n7950), .ZN(n7953) );
  MUX2_X1 U9594 ( .A(n7954), .B(n7953), .S(n8070), .Z(n7972) );
  NAND2_X1 U9595 ( .A1(n7964), .A2(n7963), .ZN(n7956) );
  NAND2_X1 U9596 ( .A1(n7960), .A2(n7959), .ZN(n7955) );
  MUX2_X1 U9597 ( .A(n7956), .B(n7955), .S(n8070), .Z(n7967) );
  NOR2_X1 U9598 ( .A1(n7967), .A2(n7957), .ZN(n7971) );
  AND2_X1 U9599 ( .A1(n7959), .A2(n7958), .ZN(n7961) );
  OAI211_X1 U9600 ( .C1(n7967), .C2(n7961), .A(n7974), .B(n7960), .ZN(n7969)
         );
  AND2_X1 U9601 ( .A1(n7963), .A2(n7962), .ZN(n7966) );
  AND2_X1 U9602 ( .A1(n7973), .A2(n7964), .ZN(n7965) );
  OAI21_X1 U9603 ( .B1(n7967), .B2(n7966), .A(n7965), .ZN(n7968) );
  MUX2_X1 U9604 ( .A(n7969), .B(n7968), .S(n8070), .Z(n7970) );
  AOI21_X1 U9605 ( .B1(n7972), .B2(n7971), .A(n7970), .ZN(n7981) );
  NAND2_X1 U9606 ( .A1(n7977), .A2(n7973), .ZN(n7976) );
  NAND2_X1 U9607 ( .A1(n4997), .A2(n7974), .ZN(n7975) );
  MUX2_X1 U9608 ( .A(n7976), .B(n7975), .S(n8070), .Z(n7980) );
  MUX2_X1 U9609 ( .A(n7977), .B(n4997), .S(n8066), .Z(n7978) );
  OAI211_X1 U9610 ( .C1(n7981), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7987)
         );
  AND2_X1 U9611 ( .A1(n9991), .A2(n9639), .ZN(n7984) );
  INV_X1 U9612 ( .A(n7982), .ZN(n7983) );
  MUX2_X1 U9613 ( .A(n7984), .B(n7983), .S(n8066), .Z(n7985) );
  INV_X1 U9614 ( .A(n7985), .ZN(n7986) );
  MUX2_X1 U9615 ( .A(n7989), .B(n7988), .S(n8066), .Z(n7990) );
  NAND2_X1 U9616 ( .A1(n7993), .A2(n7992), .ZN(n8000) );
  INV_X1 U9617 ( .A(n7994), .ZN(n7996) );
  OAI21_X1 U9618 ( .B1(n8000), .B2(n7996), .A(n7995), .ZN(n8002) );
  INV_X1 U9619 ( .A(n7997), .ZN(n7999) );
  OAI211_X1 U9620 ( .C1(n8000), .C2(n7999), .A(n8006), .B(n7998), .ZN(n8001)
         );
  MUX2_X1 U9621 ( .A(n8002), .B(n8001), .S(n8066), .Z(n8004) );
  INV_X1 U9622 ( .A(n8003), .ZN(n8005) );
  INV_X1 U9623 ( .A(n8006), .ZN(n8007) );
  NAND2_X1 U9624 ( .A1(n8013), .A2(n8008), .ZN(n8010) );
  OAI211_X1 U9625 ( .C1(n8015), .C2(n8010), .A(n8009), .B(n8016), .ZN(n8011)
         );
  NAND3_X1 U9626 ( .A1(n8011), .A2(n8014), .A3(n8018), .ZN(n8012) );
  NAND3_X1 U9627 ( .A1(n8015), .A2(n8014), .A3(n8013), .ZN(n8017) );
  NAND3_X1 U9628 ( .A1(n8017), .A2(n8374), .A3(n8016), .ZN(n8019) );
  NAND3_X1 U9629 ( .A1(n8019), .A2(n8018), .A3(n8022), .ZN(n8020) );
  MUX2_X1 U9630 ( .A(n8022), .B(n8021), .S(n8070), .Z(n8023) );
  NAND2_X1 U9631 ( .A1(n8323), .A2(n8024), .ZN(n8025) );
  MUX2_X1 U9632 ( .A(n8026), .B(n8025), .S(n8070), .Z(n8027) );
  INV_X1 U9633 ( .A(n8027), .ZN(n8028) );
  NAND2_X1 U9634 ( .A1(n8036), .A2(n8032), .ZN(n8031) );
  AOI21_X1 U9635 ( .B1(n8031), .B2(n8030), .A(n8029), .ZN(n8040) );
  INV_X1 U9636 ( .A(n8032), .ZN(n8035) );
  INV_X1 U9637 ( .A(n8033), .ZN(n8034) );
  OAI21_X1 U9638 ( .B1(n8036), .B2(n8035), .A(n8034), .ZN(n8038) );
  NAND2_X1 U9639 ( .A1(n8038), .A2(n8037), .ZN(n8039) );
  MUX2_X1 U9640 ( .A(n8040), .B(n8039), .S(n8066), .Z(n8041) );
  MUX2_X1 U9641 ( .A(n4819), .B(n8043), .S(n8066), .Z(n8044) );
  NOR2_X1 U9642 ( .A1(n8302), .A2(n8044), .ZN(n8045) );
  INV_X1 U9643 ( .A(n8046), .ZN(n8047) );
  MUX2_X1 U9644 ( .A(n8048), .B(n8047), .S(n8070), .Z(n8049) );
  INV_X1 U9645 ( .A(n8050), .ZN(n8052) );
  MUX2_X1 U9646 ( .A(n8052), .B(n8051), .S(n8066), .Z(n8053) );
  MUX2_X1 U9647 ( .A(n8077), .B(n8060), .S(n8070), .Z(n8064) );
  NAND2_X1 U9648 ( .A1(n8054), .A2(n8066), .ZN(n8056) );
  AND2_X1 U9649 ( .A1(n8282), .A2(n8066), .ZN(n8055) );
  AOI21_X1 U9650 ( .B1(n8057), .B2(n8056), .A(n8055), .ZN(n8063) );
  INV_X1 U9651 ( .A(n8058), .ZN(n8059) );
  AOI21_X1 U9652 ( .B1(n8078), .B2(n8060), .A(n8059), .ZN(n8062) );
  INV_X1 U9653 ( .A(n8071), .ZN(n8061) );
  INV_X1 U9654 ( .A(n8064), .ZN(n8065) );
  NAND3_X1 U9655 ( .A1(n4662), .A2(n4444), .A3(n8065), .ZN(n8074) );
  NAND2_X1 U9656 ( .A1(n8067), .A2(n8066), .ZN(n8069) );
  NAND2_X1 U9657 ( .A1(n8069), .A2(n8068), .ZN(n8079) );
  NAND2_X1 U9658 ( .A1(n8071), .A2(n8079), .ZN(n8073) );
  NAND3_X1 U9659 ( .A1(n8074), .A2(n8071), .A3(n8070), .ZN(n8072) );
  OAI211_X1 U9660 ( .C1(n8074), .C2(n8073), .A(n8072), .B(n5005), .ZN(n8083)
         );
  INV_X1 U9661 ( .A(n8075), .ZN(n8076) );
  AOI21_X1 U9662 ( .B1(n8078), .B2(n8077), .A(n8076), .ZN(n8082) );
  INV_X1 U9663 ( .A(n8079), .ZN(n8080) );
  NAND2_X1 U9664 ( .A1(n8080), .A2(n5005), .ZN(n8081) );
  XNOR2_X1 U9665 ( .A(n8086), .B(n8247), .ZN(n8094) );
  INV_X1 U9666 ( .A(n8087), .ZN(n8088) );
  NAND3_X1 U9667 ( .A1(n8089), .A2(n8088), .A3(n8253), .ZN(n8090) );
  OAI211_X1 U9668 ( .C1(n8091), .C2(n8093), .A(n8090), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8092) );
  OAI21_X1 U9669 ( .B1(n8094), .B2(n8093), .A(n8092), .ZN(P2_U3296) );
  MUX2_X1 U9670 ( .A(n8282), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8225), .Z(
        P2_U3520) );
  MUX2_X1 U9671 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8295), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9672 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8304), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9673 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8095), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9674 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8329), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9675 ( .A(n8096), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8225), .Z(
        P2_U3515) );
  MUX2_X1 U9676 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8356), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9677 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8367), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9678 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8378), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9679 ( .A(n8387), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8225), .Z(
        P2_U3511) );
  MUX2_X1 U9680 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8379), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9681 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8389), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U9682 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8097), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9683 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8098), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9684 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8099), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9685 ( .A(n8100), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8225), .Z(
        P2_U3505) );
  MUX2_X1 U9686 ( .A(n8101), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8225), .Z(
        P2_U3504) );
  MUX2_X1 U9687 ( .A(n8102), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8225), .Z(
        P2_U3503) );
  MUX2_X1 U9688 ( .A(n8103), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8225), .Z(
        P2_U3502) );
  MUX2_X1 U9689 ( .A(n8104), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8225), .Z(
        P2_U3501) );
  MUX2_X1 U9690 ( .A(n8105), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8225), .Z(
        P2_U3500) );
  MUX2_X1 U9691 ( .A(n8106), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8225), .Z(
        P2_U3499) );
  MUX2_X1 U9692 ( .A(n8107), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8225), .Z(
        P2_U3498) );
  MUX2_X1 U9693 ( .A(n8108), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8225), .Z(
        P2_U3497) );
  MUX2_X1 U9694 ( .A(n8109), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8225), .Z(
        P2_U3496) );
  MUX2_X1 U9695 ( .A(n8110), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8225), .Z(
        P2_U3495) );
  MUX2_X1 U9696 ( .A(n8111), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8225), .Z(
        P2_U3494) );
  MUX2_X1 U9697 ( .A(n8112), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8225), .Z(
        P2_U3493) );
  MUX2_X1 U9698 ( .A(n8113), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8225), .Z(
        P2_U3492) );
  NOR2_X1 U9699 ( .A1(n8132), .A2(n8114), .ZN(n8116) );
  INV_X1 U9700 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8117) );
  MUX2_X1 U9701 ( .A(n8117), .B(P2_REG2_REG_14__SCAN_IN), .S(n8136), .Z(n8118)
         );
  INV_X1 U9702 ( .A(n8118), .ZN(n8119) );
  NOR2_X1 U9703 ( .A1(n8120), .A2(n8119), .ZN(n8157) );
  AOI21_X1 U9704 ( .B1(n8120), .B2(n8119), .A(n8157), .ZN(n8144) );
  MUX2_X1 U9705 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8253), .Z(n8148) );
  XNOR2_X1 U9706 ( .A(n8136), .B(n8148), .ZN(n8126) );
  INV_X1 U9707 ( .A(n8121), .ZN(n8122) );
  NAND2_X1 U9708 ( .A1(n8132), .A2(n8122), .ZN(n8124) );
  NAND2_X1 U9709 ( .A1(n8124), .A2(n8123), .ZN(n8125) );
  NAND2_X1 U9710 ( .A1(n8126), .A2(n8125), .ZN(n8149) );
  OAI21_X1 U9711 ( .B1(n8126), .B2(n8125), .A(n8149), .ZN(n8142) );
  INV_X1 U9712 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8130) );
  NAND2_X1 U9713 ( .A1(n8261), .A2(n8136), .ZN(n8129) );
  INV_X1 U9714 ( .A(n8127), .ZN(n8128) );
  OAI211_X1 U9715 ( .C1(n8130), .C2(n8259), .A(n8129), .B(n8128), .ZN(n8141)
         );
  NOR2_X1 U9716 ( .A1(n8132), .A2(n8131), .ZN(n8134) );
  AOI22_X1 U9717 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8136), .B1(n8158), .B2(
        n8135), .ZN(n8137) );
  AOI21_X1 U9718 ( .B1(n8138), .B2(n8137), .A(n8145), .ZN(n8139) );
  NOR2_X1 U9719 ( .A1(n8139), .A2(n8237), .ZN(n8140) );
  AOI211_X1 U9720 ( .C1(n8226), .C2(n8142), .A(n8141), .B(n8140), .ZN(n8143)
         );
  OAI21_X1 U9721 ( .B1(n8144), .B2(n8270), .A(n8143), .ZN(P2_U3196) );
  INV_X1 U9722 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8147) );
  AOI21_X1 U9723 ( .B1(n8147), .B2(n8146), .A(n8186), .ZN(n8166) );
  MUX2_X1 U9724 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8253), .Z(n8175) );
  XNOR2_X1 U9725 ( .A(n8185), .B(n8175), .ZN(n8152) );
  OR2_X1 U9726 ( .A1(n8148), .A2(n8158), .ZN(n8150) );
  NAND2_X1 U9727 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U9728 ( .A1(n8152), .A2(n8151), .ZN(n8176) );
  OAI21_X1 U9729 ( .B1(n8152), .B2(n8151), .A(n8176), .ZN(n8164) );
  INV_X1 U9730 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U9731 ( .A1(n8261), .A2(n8185), .ZN(n8155) );
  INV_X1 U9732 ( .A(n8153), .ZN(n8154) );
  OAI211_X1 U9733 ( .C1(n8156), .C2(n8259), .A(n8155), .B(n8154), .ZN(n8163)
         );
  AOI21_X1 U9734 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n8158), .A(n8157), .ZN(
        n8167) );
  XNOR2_X1 U9735 ( .A(n8185), .B(n8167), .ZN(n8160) );
  INV_X1 U9736 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8159) );
  AOI21_X1 U9737 ( .B1(n8160), .B2(n8159), .A(n8168), .ZN(n8161) );
  NOR2_X1 U9738 ( .A1(n8161), .A2(n8270), .ZN(n8162) );
  AOI211_X1 U9739 ( .C1(n8226), .C2(n8164), .A(n8163), .B(n8162), .ZN(n8165)
         );
  OAI21_X1 U9740 ( .B1(n8166), .B2(n8237), .A(n8165), .ZN(P2_U3197) );
  NOR2_X1 U9741 ( .A1(n8185), .A2(n8167), .ZN(n8169) );
  INV_X1 U9742 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8171) );
  NOR2_X1 U9743 ( .A1(n8204), .A2(n8171), .ZN(n8170) );
  AOI21_X1 U9744 ( .B1(n8171), .B2(n8204), .A(n8170), .ZN(n8172) );
  AOI21_X1 U9745 ( .B1(n8173), .B2(n8172), .A(n8203), .ZN(n8195) );
  INV_X1 U9746 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8183) );
  MUX2_X1 U9747 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8253), .Z(n8198) );
  XNOR2_X1 U9748 ( .A(n8198), .B(n8193), .ZN(n8179) );
  OR2_X1 U9749 ( .A1(n8175), .A2(n8174), .ZN(n8177) );
  NAND2_X1 U9750 ( .A1(n8177), .A2(n8176), .ZN(n8178) );
  NAND2_X1 U9751 ( .A1(n8179), .A2(n8178), .ZN(n8199) );
  OAI21_X1 U9752 ( .B1(n8179), .B2(n8178), .A(n8199), .ZN(n8180) );
  NAND2_X1 U9753 ( .A1(n8180), .A2(n8226), .ZN(n8182) );
  OAI211_X1 U9754 ( .C1(n8259), .C2(n8183), .A(n8182), .B(n8181), .ZN(n8192)
         );
  NOR2_X1 U9755 ( .A1(n8185), .A2(n8184), .ZN(n8187) );
  INV_X1 U9756 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8496) );
  AOI22_X1 U9757 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8193), .B1(n8204), .B2(
        n8496), .ZN(n8188) );
  AOI21_X1 U9758 ( .B1(n8189), .B2(n8188), .A(n8196), .ZN(n8190) );
  NOR2_X1 U9759 ( .A1(n8190), .A2(n8237), .ZN(n8191) );
  AOI211_X1 U9760 ( .C1(n8261), .C2(n8193), .A(n8192), .B(n8191), .ZN(n8194)
         );
  OAI21_X1 U9761 ( .B1(n8195), .B2(n8270), .A(n8194), .ZN(P2_U3198) );
  INV_X1 U9762 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8493) );
  XNOR2_X1 U9763 ( .A(n8231), .B(n8230), .ZN(n8197) );
  NOR2_X1 U9764 ( .A1(n8493), .A2(n8197), .ZN(n8232) );
  AOI21_X1 U9765 ( .B1(n8493), .B2(n8197), .A(n8232), .ZN(n8212) );
  INV_X1 U9766 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8423) );
  MUX2_X1 U9767 ( .A(n8423), .B(n8493), .S(n8253), .Z(n8220) );
  XNOR2_X1 U9768 ( .A(n8220), .B(n8209), .ZN(n8202) );
  OR2_X1 U9769 ( .A1(n8198), .A2(n8204), .ZN(n8200) );
  NAND2_X1 U9770 ( .A1(n8200), .A2(n8199), .ZN(n8201) );
  NAND2_X1 U9771 ( .A1(n8202), .A2(n8201), .ZN(n8218) );
  OAI21_X1 U9772 ( .B1(n8202), .B2(n8201), .A(n8218), .ZN(n8211) );
  INV_X1 U9773 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8208) );
  NOR2_X1 U9774 ( .A1(n8423), .A2(n8205), .ZN(n8214) );
  AOI21_X1 U9775 ( .B1(n8205), .B2(n8423), .A(n8214), .ZN(n8206) );
  NOR2_X1 U9776 ( .A1(n8224), .A2(n8209), .ZN(n8210) );
  NOR2_X1 U9777 ( .A1(n8231), .A2(n8213), .ZN(n8215) );
  NOR2_X1 U9778 ( .A1(n8215), .A2(n8214), .ZN(n8217) );
  NAND2_X1 U9779 ( .A1(n8234), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8241) );
  OAI21_X1 U9780 ( .B1(n8234), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8241), .ZN(
        n8216) );
  AOI21_X1 U9781 ( .B1(n8217), .B2(n8216), .A(n8243), .ZN(n8240) );
  INV_X1 U9782 ( .A(n8218), .ZN(n8219) );
  AOI21_X1 U9783 ( .B1(n8220), .B2(n8231), .A(n8219), .ZN(n8222) );
  MUX2_X1 U9784 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8253), .Z(n8221) );
  NOR2_X1 U9785 ( .A1(n8222), .A2(n8221), .ZN(n8249) );
  INV_X1 U9786 ( .A(n8249), .ZN(n8223) );
  NAND2_X1 U9787 ( .A1(n8222), .A2(n8221), .ZN(n8250) );
  NAND2_X1 U9788 ( .A1(n8223), .A2(n8250), .ZN(n8227) );
  OAI21_X1 U9789 ( .B1(n8227), .B2(n8225), .A(n8224), .ZN(n8239) );
  INV_X1 U9790 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10023) );
  NAND3_X1 U9791 ( .A1(n8227), .A2(n8226), .A3(n8234), .ZN(n8229) );
  OAI211_X1 U9792 ( .C1(n10023), .C2(n8259), .A(n8229), .B(n8228), .ZN(n8238)
         );
  NOR2_X1 U9793 ( .A1(n8231), .A2(n8230), .ZN(n8233) );
  NOR2_X1 U9794 ( .A1(n8233), .A2(n8232), .ZN(n8236) );
  NAND2_X1 U9795 ( .A1(n8234), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8244) );
  OAI21_X1 U9796 ( .B1(n8234), .B2(P2_REG1_REG_18__SCAN_IN), .A(n8244), .ZN(
        n8235) );
  NOR2_X1 U9797 ( .A1(n8236), .A2(n8235), .ZN(n8246) );
  INV_X1 U9798 ( .A(n8241), .ZN(n8242) );
  INV_X1 U9799 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10244) );
  MUX2_X1 U9800 ( .A(n10244), .B(P2_REG2_REG_19__SCAN_IN), .S(n8262), .Z(n8255) );
  INV_X1 U9801 ( .A(n8244), .ZN(n8245) );
  NOR2_X1 U9802 ( .A1(n8246), .A2(n8245), .ZN(n8248) );
  XNOR2_X1 U9803 ( .A(n8247), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8252) );
  XNOR2_X1 U9804 ( .A(n8248), .B(n8252), .ZN(n8268) );
  AOI21_X1 U9805 ( .B1(n8251), .B2(n8250), .A(n8249), .ZN(n8257) );
  INV_X1 U9806 ( .A(n8252), .ZN(n8254) );
  MUX2_X1 U9807 ( .A(n8255), .B(n8254), .S(n8253), .Z(n8256) );
  XNOR2_X1 U9808 ( .A(n8257), .B(n8256), .ZN(n8265) );
  OAI21_X1 U9809 ( .B1(n8259), .B2(n4629), .A(n8258), .ZN(n8260) );
  AOI21_X1 U9810 ( .B1(n8262), .B2(n8261), .A(n8260), .ZN(n8263) );
  OAI21_X1 U9811 ( .B1(n8265), .B2(n8264), .A(n8263), .ZN(n8266) );
  AOI21_X1 U9812 ( .B1(n8268), .B2(n8267), .A(n8266), .ZN(n8269) );
  OAI21_X1 U9813 ( .B1(n9648), .B2(n8502), .A(n8273), .ZN(n8275) );
  AOI21_X1 U9814 ( .B1(n9648), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8275), .ZN(
        n8274) );
  OAI21_X1 U9815 ( .B1(n8451), .B2(n8277), .A(n8274), .ZN(P2_U3202) );
  AOI21_X1 U9816 ( .B1(n9648), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8275), .ZN(
        n8276) );
  OAI21_X1 U9817 ( .B1(n8454), .B2(n8277), .A(n8276), .ZN(P2_U3203) );
  XNOR2_X1 U9818 ( .A(n8281), .B(n8280), .ZN(n8286) );
  NAND2_X1 U9819 ( .A1(n8282), .A2(n8386), .ZN(n8284) );
  AOI21_X1 U9820 ( .B1(n8286), .B2(n8391), .A(n8285), .ZN(n8510) );
  MUX2_X1 U9821 ( .A(n10340), .B(n8510), .S(n9645), .Z(n8289) );
  AOI22_X1 U9822 ( .A1(n8511), .A2(n8444), .B1(n8443), .B2(n8287), .ZN(n8288)
         );
  XOR2_X1 U9823 ( .A(n8290), .B(n8291), .Z(n8518) );
  NOR2_X1 U9824 ( .A1(n8316), .A2(n9640), .ZN(n8294) );
  AOI21_X1 U9825 ( .B1(n8295), .B2(n8386), .A(n8294), .ZN(n8296) );
  AOI22_X1 U9826 ( .A1(n8299), .A2(n8444), .B1(n8443), .B2(n8298), .ZN(n8300)
         );
  XNOR2_X1 U9827 ( .A(n8301), .B(n8302), .ZN(n8526) );
  XNOR2_X1 U9828 ( .A(n8303), .B(n8302), .ZN(n8305) );
  AOI222_X1 U9829 ( .A1(n8391), .A2(n8305), .B1(n8329), .B2(n8388), .C1(n8304), 
        .C2(n8386), .ZN(n8521) );
  MUX2_X1 U9830 ( .A(n8306), .B(n8521), .S(n9645), .Z(n8309) );
  AOI22_X1 U9831 ( .A1(n8523), .A2(n8444), .B1(n8443), .B2(n8307), .ZN(n8308)
         );
  OAI211_X1 U9832 ( .C1(n8526), .C2(n8448), .A(n8309), .B(n8308), .ZN(P2_U3207) );
  XNOR2_X1 U9833 ( .A(n8310), .B(n8314), .ZN(n8530) );
  INV_X1 U9834 ( .A(n8311), .ZN(n8312) );
  AOI21_X1 U9835 ( .B1(n8314), .B2(n8313), .A(n8312), .ZN(n8315) );
  OAI222_X1 U9836 ( .A1(n9640), .A2(n8343), .B1(n9642), .B2(n8316), .C1(n9637), 
        .C2(n8315), .ZN(n8466) );
  INV_X1 U9837 ( .A(n8317), .ZN(n8318) );
  OAI22_X1 U9838 ( .A1(n8319), .A2(n8331), .B1(n8318), .B2(n9632), .ZN(n8320)
         );
  OAI21_X1 U9839 ( .B1(n8466), .B2(n8320), .A(n9645), .ZN(n8322) );
  NAND2_X1 U9840 ( .A1(n9648), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8321) );
  OAI211_X1 U9841 ( .C1(n8530), .C2(n8448), .A(n8322), .B(n8321), .ZN(P2_U3208) );
  INV_X1 U9842 ( .A(n8323), .ZN(n8324) );
  NOR2_X1 U9843 ( .A1(n8325), .A2(n8324), .ZN(n8326) );
  XNOR2_X1 U9844 ( .A(n8326), .B(n8328), .ZN(n8535) );
  XOR2_X1 U9845 ( .A(n8328), .B(n8327), .Z(n8330) );
  AOI222_X1 U9846 ( .A1(n8391), .A2(n8330), .B1(n8356), .B2(n8388), .C1(n8329), 
        .C2(n8386), .ZN(n8531) );
  OAI21_X1 U9847 ( .B1(n8332), .B2(n8331), .A(n8531), .ZN(n8333) );
  NAND2_X1 U9848 ( .A1(n8333), .A2(n9645), .ZN(n8336) );
  AOI22_X1 U9849 ( .A1(n8334), .A2(n8443), .B1(n9648), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8335) );
  OAI211_X1 U9850 ( .C1(n8535), .C2(n8448), .A(n8336), .B(n8335), .ZN(P2_U3209) );
  INV_X1 U9851 ( .A(n8339), .ZN(n8337) );
  XNOR2_X1 U9852 ( .A(n8338), .B(n8337), .ZN(n8539) );
  XNOR2_X1 U9853 ( .A(n8340), .B(n8339), .ZN(n8341) );
  OAI222_X1 U9854 ( .A1(n9642), .A2(n8343), .B1(n9640), .B2(n8342), .C1(n9637), 
        .C2(n8341), .ZN(n8473) );
  NAND2_X1 U9855 ( .A1(n8473), .A2(n9645), .ZN(n8349) );
  INV_X1 U9856 ( .A(n8344), .ZN(n8346) );
  INV_X1 U9857 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8345) );
  OAI22_X1 U9858 ( .A1(n8346), .A2(n9632), .B1(n9645), .B2(n8345), .ZN(n8347)
         );
  AOI21_X1 U9859 ( .B1(n8474), .B2(n8444), .A(n8347), .ZN(n8348) );
  OAI211_X1 U9860 ( .C1(n8539), .C2(n8448), .A(n8349), .B(n8348), .ZN(P2_U3210) );
  XNOR2_X1 U9861 ( .A(n8350), .B(n8354), .ZN(n8545) );
  NAND3_X1 U9862 ( .A1(n8352), .A2(n8354), .A3(n8353), .ZN(n8355) );
  NAND2_X1 U9863 ( .A1(n8351), .A2(n8355), .ZN(n8357) );
  AOI222_X1 U9864 ( .A1(n8391), .A2(n8357), .B1(n8356), .B2(n8386), .C1(n8378), 
        .C2(n8388), .ZN(n8540) );
  MUX2_X1 U9865 ( .A(n8358), .B(n8540), .S(n9645), .Z(n8361) );
  AOI22_X1 U9866 ( .A1(n8542), .A2(n8444), .B1(n8443), .B2(n8359), .ZN(n8360)
         );
  OAI211_X1 U9867 ( .C1(n8545), .C2(n8448), .A(n8361), .B(n8360), .ZN(P2_U3211) );
  XNOR2_X1 U9868 ( .A(n8362), .B(n8363), .ZN(n8551) );
  INV_X1 U9869 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8369) );
  INV_X1 U9870 ( .A(n8363), .ZN(n8365) );
  NAND3_X1 U9871 ( .A1(n8375), .A2(n8365), .A3(n8364), .ZN(n8366) );
  NAND2_X1 U9872 ( .A1(n8352), .A2(n8366), .ZN(n8368) );
  AOI222_X1 U9873 ( .A1(n8391), .A2(n8368), .B1(n8387), .B2(n8388), .C1(n8367), 
        .C2(n8386), .ZN(n8546) );
  MUX2_X1 U9874 ( .A(n8369), .B(n8546), .S(n9645), .Z(n8372) );
  AOI22_X1 U9875 ( .A1(n8548), .A2(n8444), .B1(n8443), .B2(n8370), .ZN(n8371)
         );
  OAI211_X1 U9876 ( .C1(n8551), .C2(n8448), .A(n8372), .B(n8371), .ZN(P2_U3212) );
  XNOR2_X1 U9877 ( .A(n8373), .B(n8374), .ZN(n8556) );
  INV_X1 U9878 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8381) );
  OAI21_X1 U9879 ( .B1(n8377), .B2(n8376), .A(n8375), .ZN(n8380) );
  AOI222_X1 U9880 ( .A1(n8391), .A2(n8380), .B1(n8379), .B2(n8388), .C1(n8378), 
        .C2(n8386), .ZN(n8552) );
  MUX2_X1 U9881 ( .A(n8381), .B(n8552), .S(n9645), .Z(n8384) );
  AOI22_X1 U9882 ( .A1(n8553), .A2(n8444), .B1(n8443), .B2(n8382), .ZN(n8383)
         );
  OAI211_X1 U9883 ( .C1(n8556), .C2(n8448), .A(n8384), .B(n8383), .ZN(P2_U3213) );
  XNOR2_X1 U9884 ( .A(n8385), .B(n8392), .ZN(n8390) );
  AOI222_X1 U9885 ( .A1(n8391), .A2(n8390), .B1(n8389), .B2(n8388), .C1(n8387), 
        .C2(n8386), .ZN(n8487) );
  OR2_X1 U9886 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  NAND2_X1 U9887 ( .A1(n8395), .A2(n8394), .ZN(n8488) );
  AOI22_X1 U9888 ( .A1(n9648), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8443), .B2(
        n8396), .ZN(n8398) );
  NAND2_X1 U9889 ( .A1(n8485), .A2(n8444), .ZN(n8397) );
  OAI211_X1 U9890 ( .C1(n8488), .C2(n8448), .A(n8398), .B(n8397), .ZN(n8399)
         );
  INV_X1 U9891 ( .A(n8399), .ZN(n8400) );
  OAI21_X1 U9892 ( .B1(n8487), .B2(n9648), .A(n8400), .ZN(P2_U3214) );
  XNOR2_X1 U9893 ( .A(n8401), .B(n8406), .ZN(n8402) );
  OAI222_X1 U9894 ( .A1(n9640), .A2(n8433), .B1(n9642), .B2(n8403), .C1(n8402), 
        .C2(n9637), .ZN(n8489) );
  NAND2_X1 U9895 ( .A1(n8405), .A2(n8406), .ZN(n8407) );
  NAND2_X1 U9896 ( .A1(n8404), .A2(n8407), .ZN(n8560) );
  AOI22_X1 U9897 ( .A1(n9648), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8443), .B2(
        n8408), .ZN(n8410) );
  NAND2_X1 U9898 ( .A1(n8490), .A2(n8444), .ZN(n8409) );
  OAI211_X1 U9899 ( .C1(n8560), .C2(n8448), .A(n8410), .B(n8409), .ZN(n8411)
         );
  AOI21_X1 U9900 ( .B1(n8489), .B2(n9645), .A(n8411), .ZN(n8412) );
  INV_X1 U9901 ( .A(n8412), .ZN(P2_U3215) );
  XNOR2_X1 U9902 ( .A(n8414), .B(n8416), .ZN(n8565) );
  INV_X1 U9903 ( .A(n8415), .ZN(n8417) );
  AOI21_X1 U9904 ( .B1(n8417), .B2(n8416), .A(n9637), .ZN(n8422) );
  OAI22_X1 U9905 ( .A1(n8419), .A2(n9642), .B1(n8418), .B2(n9640), .ZN(n8420)
         );
  AOI21_X1 U9906 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8561) );
  MUX2_X1 U9907 ( .A(n8423), .B(n8561), .S(n9645), .Z(n8426) );
  AOI22_X1 U9908 ( .A1(n8562), .A2(n8444), .B1(n8443), .B2(n8424), .ZN(n8425)
         );
  OAI211_X1 U9909 ( .C1(n8565), .C2(n8448), .A(n8426), .B(n8425), .ZN(P2_U3216) );
  XNOR2_X1 U9910 ( .A(n8427), .B(n8430), .ZN(n8573) );
  INV_X1 U9911 ( .A(n8429), .ZN(n8431) );
  AOI21_X1 U9912 ( .B1(n8431), .B2(n8430), .A(n9637), .ZN(n8436) );
  OAI22_X1 U9913 ( .A1(n8433), .A2(n9642), .B1(n8432), .B2(n9640), .ZN(n8434)
         );
  AOI21_X1 U9914 ( .B1(n8436), .B2(n8435), .A(n8434), .ZN(n8566) );
  MUX2_X1 U9915 ( .A(n8171), .B(n8566), .S(n9645), .Z(n8439) );
  AOI22_X1 U9916 ( .A1(n8569), .A2(n8444), .B1(n8443), .B2(n8437), .ZN(n8438)
         );
  OAI211_X1 U9917 ( .C1(n8573), .C2(n8448), .A(n8439), .B(n8438), .ZN(P2_U3217) );
  MUX2_X1 U9918 ( .A(n8440), .B(P2_REG2_REG_15__SCAN_IN), .S(n9648), .Z(n8441)
         );
  INV_X1 U9919 ( .A(n8441), .ZN(n8447) );
  AOI22_X1 U9920 ( .A1(n8445), .A2(n8444), .B1(n8443), .B2(n8442), .ZN(n8446)
         );
  OAI211_X1 U9921 ( .C1(n8449), .C2(n8448), .A(n8447), .B(n8446), .ZN(P2_U3218) );
  NOR2_X1 U9922 ( .A1(n8502), .A2(n10010), .ZN(n8452) );
  AOI21_X1 U9923 ( .B1(P2_REG1_REG_31__SCAN_IN), .B2(n10010), .A(n8452), .ZN(
        n8450) );
  OAI21_X1 U9924 ( .B1(n8451), .B2(n8460), .A(n8450), .ZN(P2_U3490) );
  AOI21_X1 U9925 ( .B1(P2_REG1_REG_30__SCAN_IN), .B2(n10010), .A(n8452), .ZN(
        n8453) );
  OAI21_X1 U9926 ( .B1(n8454), .B2(n8460), .A(n8453), .ZN(P2_U3489) );
  NAND2_X1 U9927 ( .A1(n8510), .A2(n10012), .ZN(n8457) );
  INV_X1 U9928 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8455) );
  NAND2_X1 U9929 ( .A1(n10010), .A2(n8455), .ZN(n8456) );
  NAND2_X1 U9930 ( .A1(n8511), .A2(n8497), .ZN(n8458) );
  OAI211_X1 U9931 ( .C1(n8514), .C2(n8500), .A(n8459), .B(n8458), .ZN(P2_U3487) );
  MUX2_X1 U9932 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8515), .S(n10012), .Z(n8462) );
  OAI22_X1 U9933 ( .A1(n8518), .A2(n8500), .B1(n8517), .B2(n8460), .ZN(n8461)
         );
  INV_X1 U9934 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8463) );
  MUX2_X1 U9935 ( .A(n8463), .B(n8521), .S(n10012), .Z(n8465) );
  NAND2_X1 U9936 ( .A1(n8523), .A2(n8497), .ZN(n8464) );
  OAI211_X1 U9937 ( .C1(n8500), .C2(n8526), .A(n8465), .B(n8464), .ZN(P2_U3485) );
  AOI21_X1 U9938 ( .B1(n9992), .B2(n8467), .A(n8466), .ZN(n8527) );
  MUX2_X1 U9939 ( .A(n8468), .B(n8527), .S(n10012), .Z(n8469) );
  OAI21_X1 U9940 ( .B1(n8530), .B2(n8500), .A(n8469), .ZN(P2_U3484) );
  INV_X1 U9941 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8470) );
  MUX2_X1 U9942 ( .A(n8470), .B(n8531), .S(n10012), .Z(n8472) );
  NAND2_X1 U9943 ( .A1(n8532), .A2(n8497), .ZN(n8471) );
  OAI211_X1 U9944 ( .C1(n8500), .C2(n8535), .A(n8472), .B(n8471), .ZN(P2_U3483) );
  AOI21_X1 U9945 ( .B1(n9992), .B2(n8474), .A(n8473), .ZN(n8536) );
  MUX2_X1 U9946 ( .A(n10283), .B(n8536), .S(n10012), .Z(n8475) );
  OAI21_X1 U9947 ( .B1(n8539), .B2(n8500), .A(n8475), .ZN(P2_U3482) );
  INV_X1 U9948 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8476) );
  MUX2_X1 U9949 ( .A(n8476), .B(n8540), .S(n10012), .Z(n8478) );
  NAND2_X1 U9950 ( .A1(n8542), .A2(n8497), .ZN(n8477) );
  OAI211_X1 U9951 ( .C1(n8545), .C2(n8500), .A(n8478), .B(n8477), .ZN(P2_U3481) );
  INV_X1 U9952 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8479) );
  MUX2_X1 U9953 ( .A(n8479), .B(n8546), .S(n10012), .Z(n8481) );
  NAND2_X1 U9954 ( .A1(n8548), .A2(n8497), .ZN(n8480) );
  OAI211_X1 U9955 ( .C1(n8500), .C2(n8551), .A(n8481), .B(n8480), .ZN(P2_U3480) );
  INV_X1 U9956 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8482) );
  MUX2_X1 U9957 ( .A(n8482), .B(n8552), .S(n10012), .Z(n8484) );
  NAND2_X1 U9958 ( .A1(n8553), .A2(n8497), .ZN(n8483) );
  OAI211_X1 U9959 ( .C1(n8556), .C2(n8500), .A(n8484), .B(n8483), .ZN(P2_U3479) );
  NAND2_X1 U9960 ( .A1(n8485), .A2(n9992), .ZN(n8486) );
  OAI211_X1 U9961 ( .C1(n9986), .C2(n8488), .A(n8487), .B(n8486), .ZN(n8557)
         );
  MUX2_X1 U9962 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8557), .S(n10012), .Z(
        P2_U3478) );
  INV_X1 U9963 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8491) );
  AOI21_X1 U9964 ( .B1(n9992), .B2(n8490), .A(n8489), .ZN(n8558) );
  MUX2_X1 U9965 ( .A(n8491), .B(n8558), .S(n10012), .Z(n8492) );
  OAI21_X1 U9966 ( .B1(n8500), .B2(n8560), .A(n8492), .ZN(P2_U3477) );
  MUX2_X1 U9967 ( .A(n8493), .B(n8561), .S(n10012), .Z(n8495) );
  NAND2_X1 U9968 ( .A1(n8562), .A2(n8497), .ZN(n8494) );
  OAI211_X1 U9969 ( .C1(n8565), .C2(n8500), .A(n8495), .B(n8494), .ZN(P2_U3476) );
  MUX2_X1 U9970 ( .A(n8496), .B(n8566), .S(n10012), .Z(n8499) );
  NAND2_X1 U9971 ( .A1(n8569), .A2(n8497), .ZN(n8498) );
  OAI211_X1 U9972 ( .C1(n8573), .C2(n8500), .A(n8499), .B(n8498), .ZN(P2_U3475) );
  INV_X1 U9973 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U9974 ( .A1(n8501), .A2(n8568), .ZN(n8504) );
  INV_X1 U9975 ( .A(n8502), .ZN(n8503) );
  NAND2_X1 U9976 ( .A1(n8503), .A2(n9993), .ZN(n8507) );
  OAI211_X1 U9977 ( .C1(n8505), .C2(n9993), .A(n8504), .B(n8507), .ZN(P2_U3458) );
  INV_X1 U9978 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U9979 ( .A1(n8506), .A2(n8568), .ZN(n8508) );
  OAI211_X1 U9980 ( .C1(n8509), .C2(n9993), .A(n8508), .B(n8507), .ZN(P2_U3457) );
  INV_X1 U9981 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10293) );
  MUX2_X1 U9982 ( .A(n10293), .B(n8510), .S(n9993), .Z(n8513) );
  NAND2_X1 U9983 ( .A1(n8511), .A2(n8568), .ZN(n8512) );
  OAI211_X1 U9984 ( .C1(n8514), .C2(n8572), .A(n8513), .B(n8512), .ZN(P2_U3455) );
  MUX2_X1 U9985 ( .A(n8515), .B(P2_REG0_REG_27__SCAN_IN), .S(n9994), .Z(n8520)
         );
  OAI22_X1 U9986 ( .A1(n8518), .A2(n8572), .B1(n8517), .B2(n8516), .ZN(n8519)
         );
  INV_X1 U9987 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8522) );
  MUX2_X1 U9988 ( .A(n8522), .B(n8521), .S(n9993), .Z(n8525) );
  NAND2_X1 U9989 ( .A1(n8523), .A2(n8568), .ZN(n8524) );
  OAI211_X1 U9990 ( .C1(n8526), .C2(n8572), .A(n8525), .B(n8524), .ZN(P2_U3453) );
  INV_X1 U9991 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8528) );
  MUX2_X1 U9992 ( .A(n8528), .B(n8527), .S(n9993), .Z(n8529) );
  OAI21_X1 U9993 ( .B1(n8530), .B2(n8572), .A(n8529), .ZN(P2_U3452) );
  MUX2_X1 U9994 ( .A(n10190), .B(n8531), .S(n9993), .Z(n8534) );
  NAND2_X1 U9995 ( .A1(n8532), .A2(n8568), .ZN(n8533) );
  OAI211_X1 U9996 ( .C1(n8535), .C2(n8572), .A(n8534), .B(n8533), .ZN(P2_U3451) );
  INV_X1 U9997 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8537) );
  MUX2_X1 U9998 ( .A(n8537), .B(n8536), .S(n9993), .Z(n8538) );
  OAI21_X1 U9999 ( .B1(n8539), .B2(n8572), .A(n8538), .ZN(P2_U3450) );
  INV_X1 U10000 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8541) );
  MUX2_X1 U10001 ( .A(n8541), .B(n8540), .S(n9993), .Z(n8544) );
  NAND2_X1 U10002 ( .A1(n8542), .A2(n8568), .ZN(n8543) );
  OAI211_X1 U10003 ( .C1(n8545), .C2(n8572), .A(n8544), .B(n8543), .ZN(
        P2_U3449) );
  INV_X1 U10004 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8547) );
  MUX2_X1 U10005 ( .A(n8547), .B(n8546), .S(n9993), .Z(n8550) );
  NAND2_X1 U10006 ( .A1(n8548), .A2(n8568), .ZN(n8549) );
  OAI211_X1 U10007 ( .C1(n8551), .C2(n8572), .A(n8550), .B(n8549), .ZN(
        P2_U3448) );
  INV_X1 U10008 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n10125) );
  MUX2_X1 U10009 ( .A(n10125), .B(n8552), .S(n9993), .Z(n8555) );
  NAND2_X1 U10010 ( .A1(n8553), .A2(n8568), .ZN(n8554) );
  OAI211_X1 U10011 ( .C1(n8556), .C2(n8572), .A(n8555), .B(n8554), .ZN(
        P2_U3447) );
  MUX2_X1 U10012 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8557), .S(n9993), .Z(
        P2_U3446) );
  INV_X1 U10013 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n10343) );
  MUX2_X1 U10014 ( .A(n10343), .B(n8558), .S(n9993), .Z(n8559) );
  OAI21_X1 U10015 ( .B1(n8560), .B2(n8572), .A(n8559), .ZN(P2_U3444) );
  INV_X1 U10016 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n10344) );
  MUX2_X1 U10017 ( .A(n10344), .B(n8561), .S(n9993), .Z(n8564) );
  NAND2_X1 U10018 ( .A1(n8562), .A2(n8568), .ZN(n8563) );
  OAI211_X1 U10019 ( .C1(n8565), .C2(n8572), .A(n8564), .B(n8563), .ZN(
        P2_U3441) );
  INV_X1 U10020 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8567) );
  MUX2_X1 U10021 ( .A(n8567), .B(n8566), .S(n9993), .Z(n8571) );
  NAND2_X1 U10022 ( .A1(n8569), .A2(n8568), .ZN(n8570) );
  OAI211_X1 U10023 ( .C1(n8573), .C2(n8572), .A(n8571), .B(n8570), .ZN(
        P2_U3438) );
  NAND3_X1 U10024 ( .A1(n8574), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n8576) );
  OAI22_X1 U10025 ( .A1(n8577), .A2(n8576), .B1(n8575), .B2(n4406), .ZN(n8578)
         );
  AOI21_X1 U10026 ( .B1(n9559), .B2(n8579), .A(n8578), .ZN(n8580) );
  INV_X1 U10027 ( .A(n8580), .ZN(P2_U3264) );
  AOI21_X1 U10028 ( .B1(n8586), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n8581), .ZN(
        n8582) );
  OAI21_X1 U10029 ( .B1(n8583), .B2(n8588), .A(n8582), .ZN(P2_U3267) );
  INV_X1 U10030 ( .A(n8584), .ZN(n9570) );
  AOI21_X1 U10031 ( .B1(n8586), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8585), .ZN(
        n8587) );
  OAI21_X1 U10032 ( .B1(n9570), .B2(n8588), .A(n8587), .ZN(P2_U3268) );
  MUX2_X1 U10033 ( .A(n8589), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  OAI21_X1 U10034 ( .B1(n8592), .B2(n8591), .A(n8590), .ZN(n8593) );
  NAND2_X1 U10035 ( .A1(n8593), .A2(n6298), .ZN(n8599) );
  NAND2_X1 U10036 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9795) );
  INV_X1 U10037 ( .A(n9795), .ZN(n8596) );
  NOR2_X1 U10038 ( .A1(n9719), .A2(n8594), .ZN(n8595) );
  AOI211_X1 U10039 ( .C1(n9713), .C2(n8597), .A(n8596), .B(n8595), .ZN(n8598)
         );
  OAI211_X1 U10040 ( .C1(n8600), .C2(n9703), .A(n8599), .B(n8598), .ZN(
        P1_U3215) );
  NAND2_X1 U10041 ( .A1(n8603), .A2(n8602), .ZN(n8604) );
  XNOR2_X1 U10042 ( .A(n8601), .B(n8604), .ZN(n8610) );
  AND2_X1 U10043 ( .A1(n9189), .A2(n9003), .ZN(n8605) );
  AOI21_X1 U10044 ( .B1(n9194), .B2(n9140), .A(n8605), .ZN(n9293) );
  NOR2_X1 U10045 ( .A1(n9293), .A2(n9656), .ZN(n8608) );
  OAI22_X1 U10046 ( .A1(n9297), .A2(n9719), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8606), .ZN(n8607) );
  AOI211_X1 U10047 ( .C1(n9296), .C2(n9716), .A(n8608), .B(n8607), .ZN(n8609)
         );
  OAI21_X1 U10048 ( .B1(n8610), .B2(n9660), .A(n8609), .ZN(P1_U3216) );
  OAI21_X1 U10049 ( .B1(n8614), .B2(n8611), .A(n8613), .ZN(n8615) );
  NAND2_X1 U10050 ( .A1(n8615), .A2(n6298), .ZN(n8620) );
  NAND2_X1 U10051 ( .A1(n9183), .A2(n9140), .ZN(n8617) );
  NAND2_X1 U10052 ( .A1(n9177), .A2(n9003), .ZN(n8616) );
  NAND2_X1 U10053 ( .A1(n8617), .A2(n8616), .ZN(n9351) );
  NOR2_X1 U10054 ( .A1(n10178), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9134) );
  NOR2_X1 U10055 ( .A1(n9719), .A2(n9358), .ZN(n8618) );
  AOI211_X1 U10056 ( .C1(n9351), .C2(n9713), .A(n9134), .B(n8618), .ZN(n8619)
         );
  OAI211_X1 U10057 ( .C1(n9545), .C2(n9703), .A(n8620), .B(n8619), .ZN(
        P1_U3219) );
  NAND2_X1 U10058 ( .A1(n8621), .A2(n8781), .ZN(n8624) );
  OR2_X1 U10059 ( .A1(n8782), .A2(n8622), .ZN(n8623) );
  NAND2_X1 U10060 ( .A1(n9226), .A2(n8625), .ZN(n8628) );
  NAND2_X1 U10061 ( .A1(n9021), .A2(n8626), .ZN(n8627) );
  NAND2_X1 U10062 ( .A1(n8628), .A2(n8627), .ZN(n8630) );
  XNOR2_X1 U10063 ( .A(n8630), .B(n8629), .ZN(n8633) );
  AOI22_X1 U10064 ( .A1(n9226), .A2(n8631), .B1(n6194), .B2(n9021), .ZN(n8632)
         );
  XNOR2_X1 U10065 ( .A(n8633), .B(n8632), .ZN(n8644) );
  INV_X1 U10066 ( .A(n8644), .ZN(n8634) );
  NAND2_X1 U10067 ( .A1(n8634), .A2(n6298), .ZN(n8650) );
  NAND4_X1 U10068 ( .A1(n8649), .A2(n6298), .A3(n8643), .A4(n8644), .ZN(n8648)
         );
  NAND2_X1 U10069 ( .A1(n8757), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U10070 ( .A1(n8755), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U10071 ( .A1(n8756), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8637) );
  OR2_X1 U10072 ( .A1(n8635), .A2(n9205), .ZN(n8636) );
  NAND4_X1 U10073 ( .A1(n8639), .A2(n8638), .A3(n8637), .A4(n8636), .ZN(n9020)
         );
  NAND2_X1 U10074 ( .A1(n9020), .A2(n9140), .ZN(n8641) );
  NAND2_X1 U10075 ( .A1(n9201), .A2(n9003), .ZN(n8640) );
  NAND2_X1 U10076 ( .A1(n8641), .A2(n8640), .ZN(n9214) );
  AOI22_X1 U10077 ( .A1(n9214), .A2(n9713), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8642) );
  OAI21_X1 U10078 ( .B1(n9221), .B2(n9719), .A(n8642), .ZN(n8646) );
  NOR3_X1 U10079 ( .A1(n8644), .A2(n9660), .A3(n8643), .ZN(n8645) );
  AOI211_X1 U10080 ( .C1(n9226), .C2(n9716), .A(n8646), .B(n8645), .ZN(n8647)
         );
  OAI211_X1 U10081 ( .C1(n8650), .C2(n8649), .A(n8648), .B(n8647), .ZN(
        P1_U3220) );
  OAI21_X1 U10082 ( .B1(n8653), .B2(n8651), .A(n8652), .ZN(n8654) );
  NAND2_X1 U10083 ( .A1(n8654), .A2(n6298), .ZN(n8660) );
  INV_X1 U10084 ( .A(n8655), .ZN(n9327) );
  AND2_X1 U10085 ( .A1(n9183), .A2(n9003), .ZN(n8656) );
  AOI21_X1 U10086 ( .B1(n9189), .B2(n9140), .A(n8656), .ZN(n9323) );
  OAI22_X1 U10087 ( .A1(n9323), .A2(n9656), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8657), .ZN(n8658) );
  AOI21_X1 U10088 ( .B1(n9327), .B2(n8737), .A(n8658), .ZN(n8659) );
  OAI211_X1 U10089 ( .C1(n9537), .C2(n9703), .A(n8660), .B(n8659), .ZN(
        P1_U3223) );
  OAI21_X1 U10090 ( .B1(n8663), .B2(n8662), .A(n8661), .ZN(n8664) );
  NAND2_X1 U10091 ( .A1(n8664), .A2(n6298), .ZN(n8669) );
  NAND2_X1 U10092 ( .A1(n9022), .A2(n9140), .ZN(n8666) );
  NAND2_X1 U10093 ( .A1(n9194), .A2(n9003), .ZN(n8665) );
  NAND2_X1 U10094 ( .A1(n8666), .A2(n8665), .ZN(n9264) );
  INV_X1 U10095 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n10298) );
  OAI22_X1 U10096 ( .A1(n9267), .A2(n9719), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10298), .ZN(n8667) );
  AOI21_X1 U10097 ( .B1(n9264), .B2(n9713), .A(n8667), .ZN(n8668) );
  OAI211_X1 U10098 ( .C1(n9259), .C2(n9703), .A(n8669), .B(n8668), .ZN(
        P1_U3225) );
  INV_X1 U10099 ( .A(n9494), .ZN(n9412) );
  OAI21_X1 U10100 ( .B1(n8672), .B2(n8670), .A(n8671), .ZN(n8673) );
  NAND2_X1 U10101 ( .A1(n8673), .A2(n6298), .ZN(n8679) );
  NAND2_X1 U10102 ( .A1(n9171), .A2(n9003), .ZN(n8675) );
  NAND2_X1 U10103 ( .A1(n9173), .A2(n9140), .ZN(n8674) );
  NAND2_X1 U10104 ( .A1(n8675), .A2(n8674), .ZN(n9401) );
  NAND2_X1 U10105 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9822) );
  INV_X1 U10106 ( .A(n9822), .ZN(n8677) );
  NOR2_X1 U10107 ( .A1(n9719), .A2(n9414), .ZN(n8676) );
  AOI211_X1 U10108 ( .C1(n9713), .C2(n9401), .A(n8677), .B(n8676), .ZN(n8678)
         );
  OAI211_X1 U10109 ( .C1(n9412), .C2(n9703), .A(n8679), .B(n8678), .ZN(
        P1_U3226) );
  INV_X1 U10110 ( .A(n9392), .ZN(n9552) );
  OAI21_X1 U10111 ( .B1(n8683), .B2(n8680), .A(n8682), .ZN(n8684) );
  NAND2_X1 U10112 ( .A1(n8684), .A2(n6298), .ZN(n8689) );
  NAND2_X1 U10113 ( .A1(n9177), .A2(n9140), .ZN(n8686) );
  NAND2_X1 U10114 ( .A1(n9172), .A2(n9003), .ZN(n8685) );
  AND2_X1 U10115 ( .A1(n8686), .A2(n8685), .ZN(n9389) );
  NAND2_X1 U10116 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9834) );
  OAI21_X1 U10117 ( .B1(n9389), .B2(n9656), .A(n9834), .ZN(n8687) );
  AOI21_X1 U10118 ( .B1(n9393), .B2(n8737), .A(n8687), .ZN(n8688) );
  OAI211_X1 U10119 ( .C1(n9552), .C2(n9703), .A(n8689), .B(n8688), .ZN(
        P1_U3228) );
  OAI21_X1 U10120 ( .B1(n8693), .B2(n8692), .A(n8691), .ZN(n8694) );
  NAND2_X1 U10121 ( .A1(n8694), .A2(n6298), .ZN(n8700) );
  NAND2_X1 U10122 ( .A1(n9196), .A2(n9140), .ZN(n8696) );
  NAND2_X1 U10123 ( .A1(n9191), .A2(n9003), .ZN(n8695) );
  NAND2_X1 U10124 ( .A1(n8696), .A2(n8695), .ZN(n9275) );
  OAI22_X1 U10125 ( .A1(n9282), .A2(n9719), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8697), .ZN(n8698) );
  AOI21_X1 U10126 ( .B1(n9275), .B2(n9713), .A(n8698), .ZN(n8699) );
  OAI211_X1 U10127 ( .C1(n9526), .C2(n9703), .A(n8700), .B(n8699), .ZN(
        P1_U3229) );
  INV_X1 U10128 ( .A(n8702), .ZN(n8704) );
  NOR2_X1 U10129 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  XNOR2_X1 U10130 ( .A(n8701), .B(n8705), .ZN(n8711) );
  NAND2_X1 U10131 ( .A1(n9185), .A2(n9140), .ZN(n8707) );
  NAND2_X1 U10132 ( .A1(n9179), .A2(n9003), .ZN(n8706) );
  NAND2_X1 U10133 ( .A1(n8707), .A2(n8706), .ZN(n9336) );
  AOI22_X1 U10134 ( .A1(n9336), .A2(n9713), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n8708) );
  OAI21_X1 U10135 ( .B1(n9340), .B2(n9719), .A(n8708), .ZN(n8709) );
  AOI21_X1 U10136 ( .B1(n9342), .B2(n9716), .A(n8709), .ZN(n8710) );
  OAI21_X1 U10137 ( .B1(n8711), .B2(n9660), .A(n8710), .ZN(P1_U3233) );
  XNOR2_X1 U10138 ( .A(n8714), .B(n8713), .ZN(n8715) );
  XNOR2_X1 U10139 ( .A(n8712), .B(n8715), .ZN(n8720) );
  AND2_X1 U10140 ( .A1(n9185), .A2(n9003), .ZN(n8716) );
  AOI21_X1 U10141 ( .B1(n9191), .B2(n9140), .A(n8716), .ZN(n9306) );
  AOI22_X1 U10142 ( .A1(n9312), .A2(n8737), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n8717) );
  OAI21_X1 U10143 ( .B1(n9306), .B2(n9656), .A(n8717), .ZN(n8718) );
  AOI21_X1 U10144 ( .B1(n9311), .B2(n9716), .A(n8718), .ZN(n8719) );
  OAI21_X1 U10145 ( .B1(n8720), .B2(n9660), .A(n8719), .ZN(P1_U3235) );
  INV_X1 U10146 ( .A(n8722), .ZN(n8723) );
  AOI21_X1 U10147 ( .B1(n8724), .B2(n8721), .A(n8723), .ZN(n8728) );
  NOR2_X1 U10148 ( .A1(n9719), .A2(n9365), .ZN(n8726) );
  AOI22_X1 U10149 ( .A1(n9179), .A2(n9140), .B1(n9003), .B2(n9173), .ZN(n9369)
         );
  NAND2_X1 U10150 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9850) );
  OAI21_X1 U10151 ( .B1(n9369), .B2(n9656), .A(n9850), .ZN(n8725) );
  AOI211_X1 U10152 ( .C1(n9377), .C2(n9716), .A(n8726), .B(n8725), .ZN(n8727)
         );
  OAI21_X1 U10153 ( .B1(n8728), .B2(n9660), .A(n8727), .ZN(P1_U3238) );
  INV_X1 U10154 ( .A(n8729), .ZN(n8732) );
  INV_X1 U10155 ( .A(n8730), .ZN(n8731) );
  INV_X1 U10156 ( .A(n8733), .ZN(n8735) );
  NAND3_X1 U10157 ( .A1(n8735), .A2(n6298), .A3(n8734), .ZN(n8741) );
  AND2_X1 U10158 ( .A1(n9201), .A2(n9140), .ZN(n8736) );
  AOI21_X1 U10159 ( .B1(n9196), .B2(n9003), .A(n8736), .ZN(n9247) );
  AOI22_X1 U10160 ( .A1(n9251), .A2(n8737), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n8738) );
  OAI21_X1 U10161 ( .B1(n9247), .B2(n9656), .A(n8738), .ZN(n8739) );
  AOI21_X1 U10162 ( .B1(n9445), .B2(n9716), .A(n8739), .ZN(n8740) );
  NAND2_X1 U10163 ( .A1(n8741), .A2(n8740), .ZN(P1_U3240) );
  OAI21_X1 U10164 ( .B1(n8742), .B2(n8744), .A(n8743), .ZN(n8745) );
  NAND2_X1 U10165 ( .A1(n8745), .A2(n6298), .ZN(n8751) );
  NAND2_X1 U10166 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9807) );
  INV_X1 U10167 ( .A(n9807), .ZN(n8748) );
  NOR2_X1 U10168 ( .A1(n9719), .A2(n8746), .ZN(n8747) );
  AOI211_X1 U10169 ( .C1(n9713), .C2(n8749), .A(n8748), .B(n8747), .ZN(n8750)
         );
  OAI211_X1 U10170 ( .C1(n9168), .C2(n9703), .A(n8751), .B(n8750), .ZN(
        P1_U3241) );
  NAND2_X1 U10171 ( .A1(n8752), .A2(n8781), .ZN(n8754) );
  OR2_X1 U10172 ( .A1(n8782), .A2(n10221), .ZN(n8753) );
  INV_X1 U10173 ( .A(n9142), .ZN(n8822) );
  NAND2_X1 U10174 ( .A1(n8755), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8760) );
  NAND2_X1 U10175 ( .A1(n8756), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8759) );
  NAND2_X1 U10176 ( .A1(n8757), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8758) );
  AND3_X1 U10177 ( .A1(n8760), .A2(n8759), .A3(n8758), .ZN(n9165) );
  NOR2_X1 U10178 ( .A1(n8822), .A2(n9165), .ZN(n8923) );
  NAND2_X1 U10179 ( .A1(n9148), .A2(n9165), .ZN(n8819) );
  NAND2_X1 U10180 ( .A1(n8761), .A2(n8781), .ZN(n8763) );
  INV_X1 U10181 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10337) );
  OR2_X1 U10182 ( .A1(n8782), .A2(n10337), .ZN(n8762) );
  INV_X1 U10183 ( .A(n9020), .ZN(n8776) );
  NAND2_X1 U10184 ( .A1(n9430), .A2(n8776), .ZN(n8921) );
  NAND2_X1 U10185 ( .A1(n8819), .A2(n8921), .ZN(n8991) );
  NAND2_X1 U10186 ( .A1(n9226), .A2(n9202), .ZN(n8787) );
  INV_X1 U10187 ( .A(n9201), .ZN(n8774) );
  NAND2_X1 U10188 ( .A1(n8787), .A2(n9160), .ZN(n8988) );
  INV_X1 U10189 ( .A(n8988), .ZN(n8778) );
  INV_X1 U10190 ( .A(n9196), .ZN(n9197) );
  OR2_X1 U10191 ( .A1(n9281), .A2(n9193), .ZN(n9157) );
  INV_X1 U10192 ( .A(n9191), .ZN(n9192) );
  OR2_X1 U10193 ( .A1(n9296), .A2(n9192), .ZN(n8825) );
  INV_X1 U10194 ( .A(n9189), .ZN(n9188) );
  OR2_X1 U10195 ( .A1(n9311), .A2(n9188), .ZN(n9290) );
  NAND2_X1 U10196 ( .A1(n8825), .A2(n9290), .ZN(n8764) );
  NAND2_X1 U10197 ( .A1(n9296), .A2(n9192), .ZN(n9155) );
  NAND2_X1 U10198 ( .A1(n8764), .A2(n9155), .ZN(n8827) );
  NAND2_X1 U10199 ( .A1(n9157), .A2(n8827), .ZN(n8765) );
  NAND2_X1 U10200 ( .A1(n9281), .A2(n9193), .ZN(n8905) );
  NAND2_X1 U10201 ( .A1(n8765), .A2(n8905), .ZN(n8766) );
  NAND2_X1 U10202 ( .A1(n9158), .A2(n8766), .ZN(n8987) );
  NAND2_X1 U10203 ( .A1(n9311), .A2(n9188), .ZN(n8788) );
  NAND2_X1 U10204 ( .A1(n9155), .A2(n8788), .ZN(n8826) );
  INV_X1 U10205 ( .A(n8826), .ZN(n8767) );
  INV_X1 U10206 ( .A(n9185), .ZN(n9186) );
  NAND2_X1 U10207 ( .A1(n9326), .A2(n9186), .ZN(n8899) );
  INV_X1 U10208 ( .A(n9183), .ZN(n9182) );
  NAND2_X1 U10209 ( .A1(n9342), .A2(n9182), .ZN(n8882) );
  NAND2_X1 U10210 ( .A1(n8899), .A2(n8882), .ZN(n8894) );
  OR2_X1 U10211 ( .A1(n9326), .A2(n9186), .ZN(n8982) );
  NAND2_X1 U10212 ( .A1(n8894), .A2(n8982), .ZN(n9153) );
  AND3_X1 U10213 ( .A1(n8905), .A2(n8767), .A3(n9153), .ZN(n8768) );
  NAND2_X1 U10214 ( .A1(n9450), .A2(n9197), .ZN(n8907) );
  OAI21_X1 U10215 ( .B1(n8987), .B2(n8768), .A(n8907), .ZN(n8984) );
  NAND2_X1 U10216 ( .A1(n8769), .A2(n8876), .ZN(n9400) );
  INV_X1 U10217 ( .A(n9172), .ZN(n8770) );
  OR2_X1 U10218 ( .A1(n9494), .A2(n8770), .ZN(n8879) );
  NAND2_X1 U10219 ( .A1(n9494), .A2(n8770), .ZN(n8880) );
  NAND2_X1 U10220 ( .A1(n9400), .A2(n9406), .ZN(n8771) );
  NAND2_X1 U10221 ( .A1(n8771), .A2(n8880), .ZN(n9387) );
  INV_X1 U10222 ( .A(n9173), .ZN(n9174) );
  OR2_X1 U10223 ( .A1(n9392), .A2(n9174), .ZN(n8976) );
  NAND2_X1 U10224 ( .A1(n9387), .A2(n8976), .ZN(n8772) );
  NAND2_X1 U10225 ( .A1(n9392), .A2(n9174), .ZN(n8881) );
  NAND2_X1 U10226 ( .A1(n8772), .A2(n8881), .ZN(n9367) );
  OR2_X1 U10227 ( .A1(n9377), .A2(n9176), .ZN(n8886) );
  NAND2_X1 U10228 ( .A1(n9377), .A2(n9176), .ZN(n8888) );
  NAND2_X1 U10229 ( .A1(n9367), .A2(n9372), .ZN(n9366) );
  NAND2_X1 U10230 ( .A1(n9366), .A2(n8888), .ZN(n9349) );
  INV_X1 U10231 ( .A(n9179), .ZN(n9180) );
  OR2_X1 U10232 ( .A1(n9357), .A2(n9180), .ZN(n8892) );
  NAND2_X1 U10233 ( .A1(n9357), .A2(n9180), .ZN(n8939) );
  NAND2_X1 U10234 ( .A1(n9349), .A2(n9355), .ZN(n8773) );
  OR2_X1 U10235 ( .A1(n9342), .A2(n9182), .ZN(n9319) );
  OAI21_X1 U10236 ( .B1(n8987), .B2(n9154), .A(n9159), .ZN(n8775) );
  NAND2_X1 U10237 ( .A1(n8915), .A2(n8916), .ZN(n8909) );
  INV_X1 U10238 ( .A(n8909), .ZN(n8990) );
  OAI21_X1 U10239 ( .B1(n8984), .B2(n8775), .A(n8990), .ZN(n8777) );
  NAND2_X1 U10240 ( .A1(n8920), .A2(n9162), .ZN(n8993) );
  AOI21_X1 U10241 ( .B1(n8778), .B2(n8777), .A(n8993), .ZN(n8779) );
  AOI211_X1 U10242 ( .C1(n8822), .C2(n9148), .A(n8991), .B(n8779), .ZN(n8780)
         );
  AOI21_X1 U10243 ( .B1(n9512), .B2(n8923), .A(n8780), .ZN(n8786) );
  NAND2_X1 U10244 ( .A1(n9559), .A2(n8781), .ZN(n8784) );
  OR2_X1 U10245 ( .A1(n8782), .A2(n10064), .ZN(n8783) );
  OAI21_X1 U10246 ( .B1(n8786), .B2(n8995), .A(n8785), .ZN(n8824) );
  OR2_X1 U10247 ( .A1(n9148), .A2(n9165), .ZN(n8936) );
  INV_X1 U10248 ( .A(n9243), .ZN(n9245) );
  AND2_X1 U10249 ( .A1(n9291), .A2(n4457), .ZN(n8901) );
  XNOR2_X1 U10250 ( .A(n9326), .B(n9186), .ZN(n9320) );
  NAND2_X1 U10251 ( .A1(n9319), .A2(n8882), .ZN(n9334) );
  NAND2_X1 U10252 ( .A1(n8976), .A2(n8881), .ZN(n9385) );
  INV_X1 U10253 ( .A(n8789), .ZN(n8812) );
  INV_X1 U10254 ( .A(n8954), .ZN(n8802) );
  INV_X1 U10255 ( .A(n8790), .ZN(n8801) );
  INV_X1 U10256 ( .A(n8792), .ZN(n8794) );
  NAND4_X1 U10257 ( .A1(n8795), .A2(n8794), .A3(n8793), .A4(n4403), .ZN(n8799)
         );
  NOR4_X1 U10258 ( .A1(n8799), .A2(n8798), .A3(n8797), .A4(n8796), .ZN(n8800)
         );
  NAND3_X1 U10259 ( .A1(n8802), .A2(n8801), .A3(n8800), .ZN(n8804) );
  NOR2_X1 U10260 ( .A1(n8804), .A2(n8803), .ZN(n8805) );
  NAND4_X1 U10261 ( .A1(n8808), .A2(n8807), .A3(n8806), .A4(n8805), .ZN(n8809)
         );
  NOR2_X1 U10262 ( .A1(n8810), .A2(n8809), .ZN(n8811) );
  NAND3_X1 U10263 ( .A1(n9406), .A2(n8812), .A3(n8811), .ZN(n8813) );
  NOR2_X1 U10264 ( .A1(n9385), .A2(n8813), .ZN(n8814) );
  NAND3_X1 U10265 ( .A1(n9355), .A2(n9372), .A3(n8814), .ZN(n8815) );
  OR3_X1 U10266 ( .A1(n9320), .A2(n9334), .A3(n8815), .ZN(n8816) );
  NOR2_X1 U10267 ( .A1(n4537), .A2(n8816), .ZN(n8817) );
  AND4_X1 U10268 ( .A1(n9233), .A2(n9262), .A3(n9274), .A4(n8817), .ZN(n8818)
         );
  AND3_X1 U10269 ( .A1(n9217), .A2(n9245), .A3(n8818), .ZN(n8820) );
  AND4_X1 U10270 ( .A1(n9203), .A2(n8936), .A3(n8820), .A4(n8819), .ZN(n8821)
         );
  INV_X1 U10271 ( .A(n8995), .ZN(n9013) );
  AND2_X1 U10272 ( .A1(n8821), .A2(n9013), .ZN(n8932) );
  INV_X1 U10273 ( .A(n8932), .ZN(n8823) );
  AOI21_X1 U10274 ( .B1(n8824), .B2(n8823), .A(n8938), .ZN(n8933) );
  INV_X1 U10275 ( .A(n9162), .ZN(n8919) );
  NAND2_X1 U10276 ( .A1(n8826), .A2(n8825), .ZN(n8828) );
  MUX2_X1 U10277 ( .A(n8828), .B(n8827), .S(n8934), .Z(n8904) );
  NAND2_X1 U10278 ( .A1(n8829), .A2(n8833), .ZN(n8940) );
  AND2_X1 U10279 ( .A1(n8836), .A2(n8830), .ZN(n8947) );
  NAND2_X1 U10280 ( .A1(n8838), .A2(n8834), .ZN(n8952) );
  AOI21_X1 U10281 ( .B1(n8940), .B2(n8947), .A(n8952), .ZN(n8832) );
  NAND2_X1 U10282 ( .A1(n8840), .A2(n8951), .ZN(n8831) );
  OAI21_X1 U10283 ( .B1(n8832), .B2(n8831), .A(n8955), .ZN(n8843) );
  NAND3_X1 U10284 ( .A1(n8835), .A2(n8834), .A3(n8833), .ZN(n8837) );
  NAND3_X1 U10285 ( .A1(n8837), .A2(n8951), .A3(n8836), .ZN(n8839) );
  NAND3_X1 U10286 ( .A1(n8839), .A2(n8955), .A3(n8838), .ZN(n8841) );
  NAND2_X1 U10287 ( .A1(n8841), .A2(n8840), .ZN(n8842) );
  MUX2_X1 U10288 ( .A(n8843), .B(n8842), .S(n8934), .Z(n8845) );
  NAND2_X1 U10289 ( .A1(n8845), .A2(n8844), .ZN(n8851) );
  NAND2_X1 U10290 ( .A1(n8852), .A2(n8848), .ZN(n8849) );
  INV_X1 U10291 ( .A(n8852), .ZN(n8853) );
  OAI21_X1 U10292 ( .B1(n8859), .B2(n8853), .A(n8958), .ZN(n8854) );
  NAND2_X1 U10293 ( .A1(n8854), .A2(n8963), .ZN(n8856) );
  AND2_X1 U10294 ( .A1(n8862), .A2(n8860), .ZN(n8961) );
  INV_X1 U10295 ( .A(n8965), .ZN(n8855) );
  AOI21_X1 U10296 ( .B1(n8856), .B2(n8961), .A(n8855), .ZN(n8866) );
  AND2_X1 U10297 ( .A1(n8965), .A2(n8861), .ZN(n8863) );
  AOI21_X1 U10298 ( .B1(n8864), .B2(n8863), .A(n4867), .ZN(n8865) );
  MUX2_X1 U10299 ( .A(n8866), .B(n8865), .S(n8934), .Z(n8874) );
  INV_X1 U10300 ( .A(n8967), .ZN(n8868) );
  OAI21_X1 U10301 ( .B1(n8874), .B2(n8868), .A(n8867), .ZN(n8869) );
  NAND3_X1 U10302 ( .A1(n8869), .A2(n8971), .A3(n8968), .ZN(n8870) );
  NAND2_X1 U10303 ( .A1(n8870), .A2(n8876), .ZN(n8871) );
  INV_X1 U10304 ( .A(n8880), .ZN(n8977) );
  OAI211_X1 U10305 ( .C1(n8874), .C2(n8873), .A(n8872), .B(n8967), .ZN(n8877)
         );
  AND2_X1 U10306 ( .A1(n8876), .A2(n8875), .ZN(n8975) );
  NAND2_X1 U10307 ( .A1(n8877), .A2(n8975), .ZN(n8878) );
  INV_X1 U10308 ( .A(n8879), .ZN(n8972) );
  NAND2_X1 U10309 ( .A1(n8892), .A2(n8886), .ZN(n8979) );
  INV_X1 U10310 ( .A(n8979), .ZN(n8884) );
  AND2_X1 U10311 ( .A1(n8888), .A2(n8881), .ZN(n8981) );
  OAI211_X1 U10312 ( .C1(n8981), .C2(n8979), .A(n8882), .B(n8939), .ZN(n8883)
         );
  AOI21_X1 U10313 ( .B1(n8885), .B2(n8884), .A(n8883), .ZN(n8891) );
  NAND3_X1 U10314 ( .A1(n8887), .A2(n8886), .A3(n8976), .ZN(n8889) );
  NAND3_X1 U10315 ( .A1(n8889), .A2(n8939), .A3(n8888), .ZN(n8890) );
  MUX2_X1 U10316 ( .A(n8891), .B(n8890), .S(n8934), .Z(n8898) );
  NAND2_X1 U10317 ( .A1(n9319), .A2(n8892), .ZN(n8893) );
  NAND2_X1 U10318 ( .A1(n8893), .A2(n8934), .ZN(n8897) );
  NAND2_X1 U10319 ( .A1(n8982), .A2(n9319), .ZN(n8895) );
  MUX2_X1 U10320 ( .A(n8895), .B(n8894), .S(n8934), .Z(n8896) );
  AOI21_X1 U10321 ( .B1(n8898), .B2(n8897), .A(n8896), .ZN(n8903) );
  MUX2_X1 U10322 ( .A(n8899), .B(n8982), .S(n8934), .Z(n8900) );
  INV_X1 U10323 ( .A(n8900), .ZN(n8902) );
  MUX2_X1 U10324 ( .A(n8905), .B(n9157), .S(n8934), .Z(n8906) );
  NAND2_X1 U10325 ( .A1(n9159), .A2(n8907), .ZN(n8911) );
  AOI21_X1 U10326 ( .B1(n8914), .B2(n9158), .A(n8911), .ZN(n8910) );
  NOR2_X1 U10327 ( .A1(n8988), .A2(n8934), .ZN(n8908) );
  INV_X1 U10328 ( .A(n9158), .ZN(n8913) );
  INV_X1 U10329 ( .A(n8911), .ZN(n8912) );
  OAI21_X1 U10330 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8917) );
  NAND2_X1 U10331 ( .A1(n8988), .A2(n8934), .ZN(n8918) );
  INV_X1 U10332 ( .A(n9203), .ZN(n9163) );
  MUX2_X1 U10333 ( .A(n8921), .B(n8920), .S(n8934), .Z(n8922) );
  MUX2_X1 U10334 ( .A(n8926), .B(n4549), .S(n9148), .Z(n8930) );
  NAND2_X1 U10335 ( .A1(n9013), .A2(n8924), .ZN(n8929) );
  INV_X1 U10336 ( .A(n9165), .ZN(n9019) );
  NAND2_X1 U10337 ( .A1(n9148), .A2(n9019), .ZN(n8925) );
  OAI22_X1 U10338 ( .A1(n8926), .A2(n8925), .B1(n8934), .B2(n8936), .ZN(n8927)
         );
  INV_X1 U10339 ( .A(n8938), .ZN(n9006) );
  NAND2_X1 U10340 ( .A1(n8934), .A2(n8943), .ZN(n8935) );
  INV_X1 U10341 ( .A(n8936), .ZN(n8937) );
  NOR2_X1 U10342 ( .A1(n8938), .A2(n8937), .ZN(n8997) );
  INV_X1 U10343 ( .A(n8940), .ZN(n8950) );
  INV_X1 U10344 ( .A(n8941), .ZN(n8945) );
  NAND2_X1 U10345 ( .A1(n5813), .A2(n8942), .ZN(n8944) );
  NAND4_X1 U10346 ( .A1(n8946), .A2(n8945), .A3(n8944), .A4(n8943), .ZN(n8949)
         );
  INV_X1 U10347 ( .A(n8947), .ZN(n8948) );
  AOI21_X1 U10348 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8953) );
  OAI21_X1 U10349 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8956) );
  AOI21_X1 U10350 ( .B1(n8956), .B2(n8955), .A(n8954), .ZN(n8960) );
  INV_X1 U10351 ( .A(n8957), .ZN(n8959) );
  OAI21_X1 U10352 ( .B1(n8960), .B2(n8959), .A(n8958), .ZN(n8964) );
  INV_X1 U10353 ( .A(n8961), .ZN(n8962) );
  AOI21_X1 U10354 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8970) );
  NAND2_X1 U10355 ( .A1(n8966), .A2(n8965), .ZN(n8969) );
  OAI211_X1 U10356 ( .C1(n8970), .C2(n8969), .A(n8968), .B(n8967), .ZN(n8974)
         );
  INV_X1 U10357 ( .A(n8971), .ZN(n8973) );
  AOI211_X1 U10358 ( .C1(n8975), .C2(n8974), .A(n8973), .B(n8972), .ZN(n8978)
         );
  OAI21_X1 U10359 ( .B1(n8978), .B2(n8977), .A(n8976), .ZN(n8980) );
  AOI21_X1 U10360 ( .B1(n8981), .B2(n8980), .A(n8979), .ZN(n8983) );
  OAI211_X1 U10361 ( .C1(n4861), .C2(n8983), .A(n8982), .B(n9319), .ZN(n8986)
         );
  INV_X1 U10362 ( .A(n8984), .ZN(n8985) );
  OAI211_X1 U10363 ( .C1(n8987), .C2(n8986), .A(n8985), .B(n9159), .ZN(n8989)
         );
  AOI21_X1 U10364 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8994) );
  INV_X1 U10365 ( .A(n8991), .ZN(n8992) );
  OAI21_X1 U10366 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(n8996) );
  AOI21_X1 U10367 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n9001) );
  NAND2_X1 U10368 ( .A1(n9001), .A2(n9002), .ZN(n8999) );
  INV_X1 U10369 ( .A(n9010), .ZN(n8998) );
  OAI211_X1 U10370 ( .C1(n9001), .C2(n9000), .A(n8999), .B(n8998), .ZN(n9017)
         );
  NAND4_X1 U10371 ( .A1(n9004), .A2(n9003), .A3(n9138), .A4(n9002), .ZN(n9005)
         );
  OAI211_X1 U10372 ( .C1(n9009), .C2(n9010), .A(n9005), .B(P1_B_REG_SCAN_IN), 
        .ZN(n9016) );
  OAI21_X1 U10373 ( .B1(n4549), .B2(n9006), .A(n8931), .ZN(n9012) );
  NOR4_X1 U10374 ( .A1(n9010), .A2(n9009), .A3(n4403), .A4(n9007), .ZN(n9011)
         );
  OAI211_X1 U10375 ( .C1(n9014), .C2(n9013), .A(n9012), .B(n9011), .ZN(n9015)
         );
  OAI211_X1 U10376 ( .C1(n9018), .C2(n9017), .A(n9016), .B(n9015), .ZN(
        P1_U3242) );
  MUX2_X1 U10377 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9019), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10378 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9020), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10379 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9021), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10380 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9201), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9022), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9196), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9191), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9189), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9185), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9183), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9179), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9177), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9173), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9172), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9171), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9023), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9024), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9025), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9026), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9027), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9028), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9029), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9030), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9031), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9032), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9033), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9034), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n5813), .S(P1_U3973), .Z(
        P1_U3555) );
  INV_X1 U10406 ( .A(n9812), .ZN(n9841) );
  OAI211_X1 U10407 ( .C1(n9037), .C2(n9036), .A(n9841), .B(n9035), .ZN(n9044)
         );
  INV_X1 U10408 ( .A(n9816), .ZN(n9837) );
  OAI211_X1 U10409 ( .C1(n9040), .C2(n9039), .A(n9837), .B(n9038), .ZN(n9043)
         );
  NAND2_X1 U10410 ( .A1(n9830), .A2(n5804), .ZN(n9042) );
  AOI22_X1 U10411 ( .A1(n9728), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9041) );
  NAND4_X1 U10412 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(
        P1_U3244) );
  INV_X1 U10413 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9046) );
  NAND2_X1 U10414 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9045) );
  OAI21_X1 U10415 ( .B1(n9852), .B2(n9046), .A(n9045), .ZN(n9047) );
  AOI21_X1 U10416 ( .B1(n9048), .B2(n9830), .A(n9047), .ZN(n9057) );
  OAI211_X1 U10417 ( .C1(n9051), .C2(n9050), .A(n9837), .B(n9049), .ZN(n9056)
         );
  OAI211_X1 U10418 ( .C1(n9054), .C2(n9053), .A(n9841), .B(n9052), .ZN(n9055)
         );
  NAND3_X1 U10419 ( .A1(n9057), .A2(n9056), .A3(n9055), .ZN(P1_U3246) );
  INV_X1 U10420 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9614) );
  NAND2_X1 U10421 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9717) );
  OAI21_X1 U10422 ( .B1(n9852), .B2(n9614), .A(n9717), .ZN(n9058) );
  AOI21_X1 U10423 ( .B1(n9059), .B2(n9830), .A(n9058), .ZN(n9068) );
  OAI211_X1 U10424 ( .C1(n9062), .C2(n9061), .A(n9837), .B(n9060), .ZN(n9067)
         );
  OAI211_X1 U10425 ( .C1(n9065), .C2(n9064), .A(n9841), .B(n9063), .ZN(n9066)
         );
  NAND3_X1 U10426 ( .A1(n9068), .A2(n9067), .A3(n9066), .ZN(P1_U3248) );
  INV_X1 U10427 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9615) );
  NAND2_X1 U10428 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9069) );
  OAI21_X1 U10429 ( .B1(n9852), .B2(n9615), .A(n9069), .ZN(n9070) );
  AOI21_X1 U10430 ( .B1(n9071), .B2(n9830), .A(n9070), .ZN(n9080) );
  OAI211_X1 U10431 ( .C1(n9074), .C2(n9073), .A(n9841), .B(n9072), .ZN(n9079)
         );
  OAI211_X1 U10432 ( .C1(n9077), .C2(n9076), .A(n9837), .B(n9075), .ZN(n9078)
         );
  NAND3_X1 U10433 ( .A1(n9080), .A2(n9079), .A3(n9078), .ZN(P1_U3249) );
  INV_X1 U10434 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U10435 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9081) );
  OAI21_X1 U10436 ( .B1(n9852), .B2(n10232), .A(n9081), .ZN(n9082) );
  AOI21_X1 U10437 ( .B1(n9083), .B2(n9830), .A(n9082), .ZN(n9092) );
  OAI211_X1 U10438 ( .C1(n9086), .C2(n9085), .A(n9841), .B(n9084), .ZN(n9091)
         );
  OAI211_X1 U10439 ( .C1(n9089), .C2(n9088), .A(n9837), .B(n9087), .ZN(n9090)
         );
  NAND3_X1 U10440 ( .A1(n9092), .A2(n9091), .A3(n9090), .ZN(P1_U3250) );
  XNOR2_X1 U10441 ( .A(n9781), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n9777) );
  NOR2_X1 U10442 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9113), .ZN(n9093) );
  AOI21_X1 U10443 ( .B1(n9113), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9093), .ZN(
        n9763) );
  OR2_X1 U10444 ( .A1(n9107), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9094) );
  NAND2_X1 U10445 ( .A1(n9095), .A2(n9094), .ZN(n9579) );
  NAND2_X1 U10446 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n9111), .ZN(n9096) );
  OAI21_X1 U10447 ( .B1(n9111), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9096), .ZN(
        n9578) );
  NOR2_X1 U10448 ( .A1(n9579), .A2(n9578), .ZN(n9581) );
  AOI21_X1 U10449 ( .B1(n9111), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9581), .ZN(
        n9748) );
  NAND2_X1 U10450 ( .A1(n9754), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9097) );
  OAI21_X1 U10451 ( .B1(n9754), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9097), .ZN(
        n9747) );
  NOR2_X1 U10452 ( .A1(n9748), .A2(n9747), .ZN(n9746) );
  AOI21_X1 U10453 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9754), .A(n9746), .ZN(
        n9762) );
  NAND2_X1 U10454 ( .A1(n9763), .A2(n9762), .ZN(n9761) );
  OAI21_X1 U10455 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9113), .A(n9761), .ZN(
        n9778) );
  NOR2_X1 U10456 ( .A1(n9777), .A2(n9778), .ZN(n9776) );
  AOI21_X1 U10457 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n9781), .A(n9776), .ZN(
        n9791) );
  NAND2_X1 U10458 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9794), .ZN(n9098) );
  OAI21_X1 U10459 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9794), .A(n9098), .ZN(
        n9790) );
  NOR2_X1 U10460 ( .A1(n9791), .A2(n9790), .ZN(n9789) );
  AOI21_X1 U10461 ( .B1(n9794), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9789), .ZN(
        n9099) );
  NOR2_X1 U10462 ( .A1(n9099), .A2(n9119), .ZN(n9100) );
  INV_X1 U10463 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9802) );
  XOR2_X1 U10464 ( .A(n9806), .B(n9099), .Z(n9803) );
  NOR2_X1 U10465 ( .A1(n9802), .A2(n9803), .ZN(n9801) );
  NOR2_X1 U10466 ( .A1(n9100), .A2(n9801), .ZN(n9818) );
  XNOR2_X1 U10467 ( .A(n9821), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9817) );
  OR2_X1 U10468 ( .A1(n9818), .A2(n9817), .ZN(n9814) );
  NAND2_X1 U10469 ( .A1(n9821), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9101) );
  AND2_X1 U10470 ( .A1(n9814), .A2(n9101), .ZN(n9826) );
  INV_X1 U10471 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U10472 ( .A(n9831), .B(n9102), .ZN(n9827) );
  NAND2_X1 U10473 ( .A1(n9826), .A2(n9827), .ZN(n9825) );
  OR2_X1 U10474 ( .A1(n9831), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9103) );
  AND2_X1 U10475 ( .A1(n9825), .A2(n9103), .ZN(n9840) );
  NAND2_X1 U10476 ( .A1(n9123), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9105) );
  OR2_X1 U10477 ( .A1(n9123), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9104) );
  AND2_X1 U10478 ( .A1(n9105), .A2(n9104), .ZN(n9839) );
  NAND2_X1 U10479 ( .A1(n9840), .A2(n9839), .ZN(n9838) );
  NAND2_X1 U10480 ( .A1(n9838), .A2(n9105), .ZN(n9106) );
  XNOR2_X1 U10481 ( .A(n9106), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9130) );
  INV_X1 U10482 ( .A(n9130), .ZN(n9127) );
  INV_X1 U10483 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10264) );
  MUX2_X1 U10484 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n10264), .S(n9781), .Z(
        n9774) );
  OR2_X1 U10485 ( .A1(n9113), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9115) );
  OR2_X1 U10486 ( .A1(n9107), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9108) );
  NAND2_X1 U10487 ( .A1(n9109), .A2(n9108), .ZN(n9583) );
  MUX2_X1 U10488 ( .A(n9110), .B(P1_REG1_REG_10__SCAN_IN), .S(n9111), .Z(n9582) );
  NOR2_X1 U10489 ( .A1(n9583), .A2(n9582), .ZN(n9585) );
  AOI21_X1 U10490 ( .B1(n9111), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9585), .ZN(
        n9751) );
  MUX2_X1 U10491 ( .A(n9112), .B(P1_REG1_REG_11__SCAN_IN), .S(n9754), .Z(n9750) );
  NOR2_X1 U10492 ( .A1(n9751), .A2(n9750), .ZN(n9749) );
  AOI21_X1 U10493 ( .B1(n9754), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9749), .ZN(
        n9758) );
  INV_X1 U10494 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U10495 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9114), .S(n9113), .Z(n9759) );
  NAND2_X1 U10496 ( .A1(n9758), .A2(n9759), .ZN(n9757) );
  AND2_X1 U10497 ( .A1(n9115), .A2(n9757), .ZN(n9773) );
  NAND2_X1 U10498 ( .A1(n9774), .A2(n9773), .ZN(n9772) );
  NAND2_X1 U10499 ( .A1(n9781), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9116) );
  NAND2_X1 U10500 ( .A1(n9772), .A2(n9116), .ZN(n9786) );
  INV_X1 U10501 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9117) );
  XNOR2_X1 U10502 ( .A(n9794), .B(n9117), .ZN(n9785) );
  AND2_X1 U10503 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  AOI21_X1 U10504 ( .B1(n9794), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9787), .ZN(
        n9118) );
  NOR2_X1 U10505 ( .A1(n9118), .A2(n9119), .ZN(n9120) );
  XNOR2_X1 U10506 ( .A(n9119), .B(n9118), .ZN(n9800) );
  NOR2_X1 U10507 ( .A1(n9799), .A2(n9800), .ZN(n9798) );
  NOR2_X1 U10508 ( .A1(n9120), .A2(n9798), .ZN(n9811) );
  INV_X1 U10509 ( .A(n9811), .ZN(n9121) );
  XNOR2_X1 U10510 ( .A(n9821), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9810) );
  OAI22_X1 U10511 ( .A1(n9121), .A2(n9810), .B1(P1_REG1_REG_16__SCAN_IN), .B2(
        n9821), .ZN(n9829) );
  INV_X1 U10512 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9489) );
  XNOR2_X1 U10513 ( .A(n9831), .B(n9489), .ZN(n9828) );
  AOI22_X1 U10514 ( .A1(n9829), .A2(n9828), .B1(n9489), .B2(n9122), .ZN(n9844)
         );
  INV_X1 U10515 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9484) );
  AND2_X1 U10516 ( .A1(n9123), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9124) );
  AOI21_X1 U10517 ( .B1(n9484), .B2(n9847), .A(n9124), .ZN(n9843) );
  NAND2_X1 U10518 ( .A1(n9844), .A2(n9843), .ZN(n9842) );
  INV_X1 U10519 ( .A(n9124), .ZN(n9125) );
  NAND2_X1 U10520 ( .A1(n9842), .A2(n9125), .ZN(n9126) );
  XNOR2_X1 U10521 ( .A(n9126), .B(n10323), .ZN(n9128) );
  AOI22_X1 U10522 ( .A1(n9127), .A2(n9837), .B1(n9128), .B2(n9841), .ZN(n9133)
         );
  OAI21_X1 U10523 ( .B1(n9128), .B2(n9812), .A(n9848), .ZN(n9129) );
  AOI21_X1 U10524 ( .B1(n9130), .B2(n9837), .A(n9129), .ZN(n9132) );
  MUX2_X1 U10525 ( .A(n9133), .B(n9132), .S(n9131), .Z(n9136) );
  INV_X1 U10526 ( .A(n9134), .ZN(n9135) );
  OAI211_X1 U10527 ( .C1(n4628), .C2(n9852), .A(n9136), .B(n9135), .ZN(
        P1_U3262) );
  NOR2_X1 U10528 ( .A1(n9408), .A2(n9392), .ZN(n9391) );
  NAND2_X1 U10529 ( .A1(n9548), .A2(n9391), .ZN(n9374) );
  NOR2_X1 U10530 ( .A1(n9308), .A2(n9296), .ZN(n9295) );
  NAND2_X1 U10531 ( .A1(n9517), .A2(n9235), .ZN(n9223) );
  NAND2_X1 U10532 ( .A1(n9422), .A2(n9380), .ZN(n9144) );
  NAND2_X1 U10533 ( .A1(n9138), .A2(P1_B_REG_SCAN_IN), .ZN(n9139) );
  NAND2_X1 U10534 ( .A1(n9140), .A2(n9139), .ZN(n9166) );
  INV_X1 U10535 ( .A(n9166), .ZN(n9141) );
  AND2_X1 U10536 ( .A1(n9142), .A2(n9141), .ZN(n9425) );
  AND2_X1 U10537 ( .A1(n9416), .A2(n9425), .ZN(n9150) );
  AOI21_X1 U10538 ( .B1(n9421), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9150), .ZN(
        n9143) );
  OAI211_X1 U10539 ( .C1(n9508), .C2(n9897), .A(n9144), .B(n9143), .ZN(
        P1_U3263) );
  INV_X1 U10540 ( .A(n9204), .ZN(n9147) );
  INV_X1 U10541 ( .A(n9145), .ZN(n9146) );
  AOI211_X1 U10542 ( .C1(n9148), .C2(n9147), .A(n9410), .B(n9146), .ZN(n9426)
         );
  NAND2_X1 U10543 ( .A1(n9426), .A2(n9380), .ZN(n9152) );
  AND2_X1 U10544 ( .A1(n9904), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9149) );
  NOR2_X1 U10545 ( .A1(n9150), .A2(n9149), .ZN(n9151) );
  OAI211_X1 U10546 ( .C1(n9512), .C2(n9897), .A(n9152), .B(n9151), .ZN(
        P1_U3264) );
  NAND3_X1 U10547 ( .A1(n9291), .A2(n9290), .A3(n9305), .ZN(n9156) );
  NAND2_X1 U10548 ( .A1(n9274), .A2(n9273), .ZN(n9272) );
  NAND2_X1 U10549 ( .A1(n9272), .A2(n9157), .ZN(n9263) );
  NAND2_X1 U10550 ( .A1(n9263), .A2(n9262), .ZN(n9261) );
  INV_X1 U10551 ( .A(n9160), .ZN(n9161) );
  NAND2_X1 U10552 ( .A1(n9213), .A2(n9217), .ZN(n9212) );
  NAND2_X1 U10553 ( .A1(n9212), .A2(n9162), .ZN(n9164) );
  NAND2_X1 U10554 ( .A1(n9169), .A2(n5000), .ZN(n9170) );
  NOR2_X1 U10555 ( .A1(n9392), .A2(n9173), .ZN(n9175) );
  NOR2_X1 U10556 ( .A1(n9548), .A2(n9176), .ZN(n9178) );
  NOR2_X1 U10557 ( .A1(n9357), .A2(n9179), .ZN(n9181) );
  NOR2_X1 U10558 ( .A1(n9541), .A2(n9182), .ZN(n9184) );
  OAI22_X2 U10559 ( .A1(n9333), .A2(n9184), .B1(n9183), .B2(n9342), .ZN(n9318)
         );
  NOR2_X1 U10560 ( .A1(n9326), .A2(n9185), .ZN(n9187) );
  NOR2_X1 U10561 ( .A1(n9450), .A2(n9196), .ZN(n9198) );
  NAND2_X1 U10562 ( .A1(n9244), .A2(n9243), .ZN(n9199) );
  OAI21_X1 U10563 ( .B1(n9200), .B2(n9254), .A(n9199), .ZN(n9234) );
  NAND2_X1 U10564 ( .A1(n9428), .A2(n9901), .ZN(n9211) );
  AOI211_X1 U10565 ( .C1(n9430), .C2(n9223), .A(n9410), .B(n9204), .ZN(n9429)
         );
  INV_X1 U10566 ( .A(n9430), .ZN(n9208) );
  INV_X1 U10567 ( .A(n9205), .ZN(n9206) );
  AOI22_X1 U10568 ( .A1(n9421), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n9206), .B2(
        n9894), .ZN(n9207) );
  OAI21_X1 U10569 ( .B1(n9208), .B2(n9897), .A(n9207), .ZN(n9209) );
  AOI21_X1 U10570 ( .B1(n9429), .B2(n9380), .A(n9209), .ZN(n9210) );
  OAI211_X1 U10571 ( .C1(n4460), .C2(n9421), .A(n9211), .B(n9210), .ZN(
        P1_U3356) );
  OAI211_X1 U10572 ( .C1(n9213), .C2(n9217), .A(n9212), .B(n9402), .ZN(n9216)
         );
  INV_X1 U10573 ( .A(n9214), .ZN(n9215) );
  NAND2_X1 U10574 ( .A1(n9218), .A2(n9217), .ZN(n9219) );
  NAND2_X1 U10575 ( .A1(n9435), .A2(n9901), .ZN(n9228) );
  INV_X1 U10576 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9222) );
  OAI22_X1 U10577 ( .A1(n9416), .A2(n9222), .B1(n9221), .B2(n9413), .ZN(n9225)
         );
  OAI211_X1 U10578 ( .C1(n9517), .C2(n9235), .A(n9864), .B(n9223), .ZN(n9432)
         );
  NOR2_X1 U10579 ( .A1(n9432), .A2(n9345), .ZN(n9224) );
  AOI211_X1 U10580 ( .C1(n9872), .C2(n9226), .A(n9225), .B(n9224), .ZN(n9227)
         );
  OAI211_X1 U10581 ( .C1(n9421), .C2(n9433), .A(n9228), .B(n9227), .ZN(
        P1_U3265) );
  XNOR2_X1 U10582 ( .A(n9229), .B(n9233), .ZN(n9230) );
  NAND2_X1 U10583 ( .A1(n9230), .A2(n9402), .ZN(n9232) );
  NAND2_X1 U10584 ( .A1(n9232), .A2(n9231), .ZN(n9438) );
  INV_X1 U10585 ( .A(n9438), .ZN(n9242) );
  XNOR2_X1 U10586 ( .A(n9234), .B(n9233), .ZN(n9440) );
  NAND2_X1 U10587 ( .A1(n9440), .A2(n9901), .ZN(n9241) );
  AOI211_X1 U10588 ( .C1(n9236), .C2(n9249), .A(n9410), .B(n9235), .ZN(n9439)
         );
  AOI22_X1 U10589 ( .A1(n9421), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9894), .B2(
        n9237), .ZN(n9238) );
  OAI21_X1 U10590 ( .B1(n4680), .B2(n9897), .A(n9238), .ZN(n9239) );
  AOI21_X1 U10591 ( .B1(n9439), .B2(n9380), .A(n9239), .ZN(n9240) );
  OAI211_X1 U10592 ( .C1(n9242), .C2(n9421), .A(n9241), .B(n9240), .ZN(
        P1_U3266) );
  XNOR2_X1 U10593 ( .A(n9244), .B(n9243), .ZN(n9447) );
  XNOR2_X1 U10594 ( .A(n9246), .B(n9245), .ZN(n9248) );
  OAI21_X1 U10595 ( .B1(n9248), .B2(n9854), .A(n9247), .ZN(n9444) );
  INV_X1 U10596 ( .A(n9249), .ZN(n9250) );
  AOI211_X1 U10597 ( .C1(n9445), .C2(n4683), .A(n9410), .B(n9250), .ZN(n9443)
         );
  NAND2_X1 U10598 ( .A1(n9443), .A2(n9380), .ZN(n9253) );
  AOI22_X1 U10599 ( .A1(n9251), .A2(n9894), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9421), .ZN(n9252) );
  OAI211_X1 U10600 ( .C1(n9254), .C2(n9897), .A(n9253), .B(n9252), .ZN(n9255)
         );
  AOI21_X1 U10601 ( .B1(n9416), .B2(n9444), .A(n9255), .ZN(n9256) );
  OAI21_X1 U10602 ( .B1(n9447), .B2(n9398), .A(n9256), .ZN(P1_U3267) );
  XNOR2_X1 U10603 ( .A(n9257), .B(n9262), .ZN(n9452) );
  AOI211_X1 U10604 ( .C1(n9450), .C2(n9278), .A(n9410), .B(n9258), .ZN(n9448)
         );
  OAI22_X1 U10605 ( .A1(n9259), .A2(n9897), .B1(n10181), .B2(n9416), .ZN(n9260) );
  AOI21_X1 U10606 ( .B1(n9448), .B2(n9380), .A(n9260), .ZN(n9270) );
  OAI211_X1 U10607 ( .C1(n9263), .C2(n9262), .A(n9261), .B(n9402), .ZN(n9266)
         );
  INV_X1 U10608 ( .A(n9264), .ZN(n9265) );
  NAND2_X1 U10609 ( .A1(n9266), .A2(n9265), .ZN(n9449) );
  NOR2_X1 U10610 ( .A1(n9267), .A2(n9413), .ZN(n9268) );
  OAI21_X1 U10611 ( .B1(n9449), .B2(n9268), .A(n9416), .ZN(n9269) );
  OAI211_X1 U10612 ( .C1(n9452), .C2(n9398), .A(n9270), .B(n9269), .ZN(
        P1_U3268) );
  XNOR2_X1 U10613 ( .A(n9271), .B(n9274), .ZN(n9455) );
  INV_X1 U10614 ( .A(n9455), .ZN(n9288) );
  OAI211_X1 U10615 ( .C1(n9274), .C2(n9273), .A(n9272), .B(n9402), .ZN(n9277)
         );
  INV_X1 U10616 ( .A(n9275), .ZN(n9276) );
  NAND2_X1 U10617 ( .A1(n9277), .A2(n9276), .ZN(n9453) );
  INV_X1 U10618 ( .A(n9295), .ZN(n9280) );
  INV_X1 U10619 ( .A(n9278), .ZN(n9279) );
  AOI211_X1 U10620 ( .C1(n9281), .C2(n9280), .A(n9410), .B(n9279), .ZN(n9454)
         );
  NAND2_X1 U10621 ( .A1(n9454), .A2(n9380), .ZN(n9285) );
  INV_X1 U10622 ( .A(n9282), .ZN(n9283) );
  AOI22_X1 U10623 ( .A1(n9283), .A2(n9894), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9421), .ZN(n9284) );
  OAI211_X1 U10624 ( .C1(n9526), .C2(n9897), .A(n9285), .B(n9284), .ZN(n9286)
         );
  AOI21_X1 U10625 ( .B1(n9416), .B2(n9453), .A(n9286), .ZN(n9287) );
  OAI21_X1 U10626 ( .B1(n9288), .B2(n9398), .A(n9287), .ZN(P1_U3269) );
  XOR2_X1 U10627 ( .A(n9291), .B(n9289), .Z(n9460) );
  INV_X1 U10628 ( .A(n9460), .ZN(n9303) );
  NAND2_X1 U10629 ( .A1(n9305), .A2(n9290), .ZN(n9292) );
  XNOR2_X1 U10630 ( .A(n9292), .B(n9291), .ZN(n9294) );
  OAI21_X1 U10631 ( .B1(n9294), .B2(n9854), .A(n9293), .ZN(n9458) );
  AOI211_X1 U10632 ( .C1(n9296), .C2(n9308), .A(n9410), .B(n9295), .ZN(n9459)
         );
  NAND2_X1 U10633 ( .A1(n9459), .A2(n9380), .ZN(n9300) );
  INV_X1 U10634 ( .A(n9297), .ZN(n9298) );
  AOI22_X1 U10635 ( .A1(n9298), .A2(n9894), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9421), .ZN(n9299) );
  OAI211_X1 U10636 ( .C1(n9530), .C2(n9897), .A(n9300), .B(n9299), .ZN(n9301)
         );
  AOI21_X1 U10637 ( .B1(n9416), .B2(n9458), .A(n9301), .ZN(n9302) );
  OAI21_X1 U10638 ( .B1(n9303), .B2(n9398), .A(n9302), .ZN(P1_U3270) );
  XNOR2_X1 U10639 ( .A(n9304), .B(n4457), .ZN(n9465) );
  INV_X1 U10640 ( .A(n9465), .ZN(n9317) );
  OAI211_X1 U10641 ( .C1(n4445), .C2(n4457), .A(n9305), .B(n9402), .ZN(n9307)
         );
  NAND2_X1 U10642 ( .A1(n9307), .A2(n9306), .ZN(n9463) );
  INV_X1 U10643 ( .A(n9325), .ZN(n9310) );
  INV_X1 U10644 ( .A(n9308), .ZN(n9309) );
  AOI211_X1 U10645 ( .C1(n9311), .C2(n9310), .A(n9410), .B(n9309), .ZN(n9464)
         );
  NAND2_X1 U10646 ( .A1(n9464), .A2(n9380), .ZN(n9314) );
  AOI22_X1 U10647 ( .A1(n9312), .A2(n9894), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9421), .ZN(n9313) );
  OAI211_X1 U10648 ( .C1(n9534), .C2(n9897), .A(n9314), .B(n9313), .ZN(n9315)
         );
  AOI21_X1 U10649 ( .B1(n9416), .B2(n9463), .A(n9315), .ZN(n9316) );
  OAI21_X1 U10650 ( .B1(n9317), .B2(n9398), .A(n9316), .ZN(P1_U3271) );
  XNOR2_X1 U10651 ( .A(n9318), .B(n9320), .ZN(n9470) );
  INV_X1 U10652 ( .A(n9470), .ZN(n9332) );
  OR2_X1 U10653 ( .A1(n9335), .A2(n9334), .ZN(n9337) );
  NAND2_X1 U10654 ( .A1(n9337), .A2(n9319), .ZN(n9321) );
  XNOR2_X1 U10655 ( .A(n9321), .B(n9320), .ZN(n9322) );
  NAND2_X1 U10656 ( .A1(n9322), .A2(n9402), .ZN(n9324) );
  NAND2_X1 U10657 ( .A1(n9324), .A2(n9323), .ZN(n9468) );
  AOI211_X1 U10658 ( .C1(n9326), .C2(n9339), .A(n9410), .B(n9325), .ZN(n9469)
         );
  NAND2_X1 U10659 ( .A1(n9469), .A2(n9380), .ZN(n9329) );
  AOI22_X1 U10660 ( .A1(n9327), .A2(n9894), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9904), .ZN(n9328) );
  OAI211_X1 U10661 ( .C1(n9537), .C2(n9897), .A(n9329), .B(n9328), .ZN(n9330)
         );
  AOI21_X1 U10662 ( .B1(n9416), .B2(n9468), .A(n9330), .ZN(n9331) );
  OAI21_X1 U10663 ( .B1(n9332), .B2(n9398), .A(n9331), .ZN(P1_U3272) );
  XNOR2_X1 U10664 ( .A(n9333), .B(n9334), .ZN(n9474) );
  AOI21_X1 U10665 ( .B1(n9335), .B2(n9334), .A(n9854), .ZN(n9338) );
  AOI21_X1 U10666 ( .B1(n9338), .B2(n9337), .A(n9336), .ZN(n9473) );
  INV_X1 U10667 ( .A(n9473), .ZN(n9347) );
  OAI211_X1 U10668 ( .C1(n9356), .C2(n9541), .A(n9864), .B(n9339), .ZN(n9472)
         );
  INV_X1 U10669 ( .A(n9340), .ZN(n9341) );
  AOI22_X1 U10670 ( .A1(P1_REG2_REG_20__SCAN_IN), .A2(n9421), .B1(n9341), .B2(
        n9894), .ZN(n9344) );
  NAND2_X1 U10671 ( .A1(n9342), .A2(n9872), .ZN(n9343) );
  OAI211_X1 U10672 ( .C1(n9472), .C2(n9345), .A(n9344), .B(n9343), .ZN(n9346)
         );
  AOI21_X1 U10673 ( .B1(n9347), .B2(n9416), .A(n9346), .ZN(n9348) );
  OAI21_X1 U10674 ( .B1(n9474), .B2(n9398), .A(n9348), .ZN(P1_U3273) );
  XNOR2_X1 U10675 ( .A(n9349), .B(n9355), .ZN(n9350) );
  NAND2_X1 U10676 ( .A1(n9350), .A2(n9402), .ZN(n9353) );
  INV_X1 U10677 ( .A(n9351), .ZN(n9352) );
  NAND2_X1 U10678 ( .A1(n9353), .A2(n9352), .ZN(n9477) );
  INV_X1 U10679 ( .A(n9477), .ZN(n9364) );
  XOR2_X1 U10680 ( .A(n9355), .B(n9354), .Z(n9479) );
  NAND2_X1 U10681 ( .A1(n9479), .A2(n9901), .ZN(n9363) );
  AOI211_X1 U10682 ( .C1(n9357), .C2(n9374), .A(n9410), .B(n9356), .ZN(n9478)
         );
  NOR2_X1 U10683 ( .A1(n9545), .A2(n9897), .ZN(n9361) );
  OAI22_X1 U10684 ( .A1(n9416), .A2(n9359), .B1(n9358), .B2(n9413), .ZN(n9360)
         );
  AOI211_X1 U10685 ( .C1(n9478), .C2(n9380), .A(n9361), .B(n9360), .ZN(n9362)
         );
  OAI211_X1 U10686 ( .C1(n9421), .C2(n9364), .A(n9363), .B(n9362), .ZN(
        P1_U3274) );
  INV_X1 U10687 ( .A(n9365), .ZN(n9371) );
  OAI21_X1 U10688 ( .B1(n9372), .B2(n9367), .A(n9366), .ZN(n9368) );
  NAND2_X1 U10689 ( .A1(n9368), .A2(n9402), .ZN(n9370) );
  NAND2_X1 U10690 ( .A1(n9370), .A2(n9369), .ZN(n9481) );
  AOI21_X1 U10691 ( .B1(n9371), .B2(n9894), .A(n9481), .ZN(n9383) );
  XNOR2_X1 U10692 ( .A(n9373), .B(n9372), .ZN(n9483) );
  NAND2_X1 U10693 ( .A1(n9483), .A2(n9901), .ZN(n9382) );
  INV_X1 U10694 ( .A(n9391), .ZN(n9376) );
  INV_X1 U10695 ( .A(n9374), .ZN(n9375) );
  AOI211_X1 U10696 ( .C1(n9377), .C2(n9376), .A(n9410), .B(n9375), .ZN(n9482)
         );
  INV_X1 U10697 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9378) );
  OAI22_X1 U10698 ( .A1(n9548), .A2(n9897), .B1(n9378), .B2(n9416), .ZN(n9379)
         );
  AOI21_X1 U10699 ( .B1(n9482), .B2(n9380), .A(n9379), .ZN(n9381) );
  OAI211_X1 U10700 ( .C1(n9421), .C2(n9383), .A(n9382), .B(n9381), .ZN(
        P1_U3275) );
  XNOR2_X1 U10701 ( .A(n9384), .B(n9385), .ZN(n9488) );
  INV_X1 U10702 ( .A(n9488), .ZN(n9399) );
  INV_X1 U10703 ( .A(n9385), .ZN(n9386) );
  XNOR2_X1 U10704 ( .A(n9387), .B(n9386), .ZN(n9388) );
  NAND2_X1 U10705 ( .A1(n9388), .A2(n9402), .ZN(n9390) );
  NAND2_X1 U10706 ( .A1(n9390), .A2(n9389), .ZN(n9486) );
  AOI211_X1 U10707 ( .C1(n9392), .C2(n9408), .A(n9410), .B(n9391), .ZN(n9487)
         );
  NAND2_X1 U10708 ( .A1(n9487), .A2(n9380), .ZN(n9395) );
  AOI22_X1 U10709 ( .A1(n9421), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9393), .B2(
        n9894), .ZN(n9394) );
  OAI211_X1 U10710 ( .C1(n9552), .C2(n9897), .A(n9395), .B(n9394), .ZN(n9396)
         );
  AOI21_X1 U10711 ( .B1(n9416), .B2(n9486), .A(n9396), .ZN(n9397) );
  OAI21_X1 U10712 ( .B1(n9399), .B2(n9398), .A(n9397), .ZN(P1_U3276) );
  XNOR2_X1 U10713 ( .A(n9400), .B(n9406), .ZN(n9403) );
  AOI21_X1 U10714 ( .B1(n9403), .B2(n9402), .A(n9401), .ZN(n9497) );
  AOI21_X1 U10715 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9492) );
  NAND2_X1 U10716 ( .A1(n9492), .A2(n9901), .ZN(n9420) );
  INV_X1 U10717 ( .A(n9407), .ZN(n9411) );
  INV_X1 U10718 ( .A(n9408), .ZN(n9409) );
  AOI211_X1 U10719 ( .C1(n9494), .C2(n9411), .A(n9410), .B(n9409), .ZN(n9493)
         );
  NOR2_X1 U10720 ( .A1(n9412), .A2(n9897), .ZN(n9418) );
  INV_X1 U10721 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9415) );
  OAI22_X1 U10722 ( .A1(n9416), .A2(n9415), .B1(n9414), .B2(n9413), .ZN(n9417)
         );
  AOI211_X1 U10723 ( .C1(n9493), .C2(n9380), .A(n9418), .B(n9417), .ZN(n9419)
         );
  OAI211_X1 U10724 ( .C1(n9421), .C2(n9497), .A(n9420), .B(n9419), .ZN(
        P1_U3277) );
  INV_X1 U10725 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9423) );
  NOR2_X1 U10726 ( .A1(n9422), .A2(n9425), .ZN(n9505) );
  MUX2_X1 U10727 ( .A(n9423), .B(n9505), .S(n9932), .Z(n9424) );
  OAI21_X1 U10728 ( .B1(n9508), .B2(n9491), .A(n9424), .ZN(P1_U3553) );
  INV_X1 U10729 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U10730 ( .A1(n9426), .A2(n9425), .ZN(n9509) );
  MUX2_X1 U10731 ( .A(n10230), .B(n9509), .S(n9932), .Z(n9427) );
  OAI21_X1 U10732 ( .B1(n9512), .B2(n9491), .A(n9427), .ZN(P1_U3552) );
  NAND2_X1 U10733 ( .A1(n9428), .A2(n9924), .ZN(n9431) );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9513), .S(n9932), .Z(
        P1_U3551) );
  INV_X1 U10735 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9436) );
  NAND2_X1 U10736 ( .A1(n9433), .A2(n9432), .ZN(n9434) );
  OAI21_X1 U10737 ( .B1(n9517), .B2(n9491), .A(n9437), .ZN(P1_U3550) );
  INV_X1 U10738 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9441) );
  MUX2_X1 U10739 ( .A(n9441), .B(n9518), .S(n9932), .Z(n9442) );
  OAI21_X1 U10740 ( .B1(n4680), .B2(n9491), .A(n9442), .ZN(P1_U3549) );
  AOI211_X1 U10741 ( .C1(n9495), .C2(n9445), .A(n9444), .B(n9443), .ZN(n9446)
         );
  OAI21_X1 U10742 ( .B1(n9447), .B2(n9498), .A(n9446), .ZN(n9521) );
  MUX2_X1 U10743 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9521), .S(n9932), .Z(
        P1_U3548) );
  AOI211_X1 U10744 ( .C1(n9495), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9451)
         );
  OAI21_X1 U10745 ( .B1(n9452), .B2(n9498), .A(n9451), .ZN(n9522) );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9522), .S(n9932), .Z(
        P1_U3547) );
  AOI211_X1 U10747 ( .C1(n9455), .C2(n9924), .A(n9454), .B(n9453), .ZN(n9523)
         );
  MUX2_X1 U10748 ( .A(n9456), .B(n9523), .S(n9932), .Z(n9457) );
  OAI21_X1 U10749 ( .B1(n9526), .B2(n9491), .A(n9457), .ZN(P1_U3546) );
  AOI211_X1 U10750 ( .C1(n9460), .C2(n9924), .A(n9459), .B(n9458), .ZN(n9527)
         );
  MUX2_X1 U10751 ( .A(n9461), .B(n9527), .S(n9932), .Z(n9462) );
  OAI21_X1 U10752 ( .B1(n9530), .B2(n9491), .A(n9462), .ZN(P1_U3545) );
  AOI211_X1 U10753 ( .C1(n9465), .C2(n9924), .A(n9464), .B(n9463), .ZN(n9531)
         );
  MUX2_X1 U10754 ( .A(n9466), .B(n9531), .S(n9932), .Z(n9467) );
  OAI21_X1 U10755 ( .B1(n9534), .B2(n9491), .A(n9467), .ZN(P1_U3544) );
  INV_X1 U10756 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n10312) );
  AOI211_X1 U10757 ( .C1(n9470), .C2(n9924), .A(n9469), .B(n9468), .ZN(n9535)
         );
  MUX2_X1 U10758 ( .A(n10312), .B(n9535), .S(n9932), .Z(n9471) );
  OAI21_X1 U10759 ( .B1(n9537), .B2(n9491), .A(n9471), .ZN(P1_U3543) );
  OAI211_X1 U10760 ( .C1(n9474), .C2(n9498), .A(n9473), .B(n9472), .ZN(n9538)
         );
  MUX2_X1 U10761 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9538), .S(n9932), .Z(n9475) );
  INV_X1 U10762 ( .A(n9475), .ZN(n9476) );
  OAI21_X1 U10763 ( .B1(n9541), .B2(n9491), .A(n9476), .ZN(P1_U3542) );
  AOI211_X1 U10764 ( .C1(n9479), .C2(n9924), .A(n9478), .B(n9477), .ZN(n9542)
         );
  MUX2_X1 U10765 ( .A(n10323), .B(n9542), .S(n9932), .Z(n9480) );
  OAI21_X1 U10766 ( .B1(n9545), .B2(n9491), .A(n9480), .ZN(P1_U3541) );
  AOI211_X1 U10767 ( .C1(n9483), .C2(n9924), .A(n9482), .B(n9481), .ZN(n9546)
         );
  MUX2_X1 U10768 ( .A(n9484), .B(n9546), .S(n9932), .Z(n9485) );
  OAI21_X1 U10769 ( .B1(n9548), .B2(n9491), .A(n9485), .ZN(P1_U3540) );
  AOI211_X1 U10770 ( .C1(n9488), .C2(n9924), .A(n9487), .B(n9486), .ZN(n9549)
         );
  MUX2_X1 U10771 ( .A(n9489), .B(n9549), .S(n9932), .Z(n9490) );
  OAI21_X1 U10772 ( .B1(n9552), .B2(n9491), .A(n9490), .ZN(P1_U3539) );
  INV_X1 U10773 ( .A(n9492), .ZN(n9499) );
  AOI21_X1 U10774 ( .B1(n9495), .B2(n9494), .A(n9493), .ZN(n9496) );
  OAI211_X1 U10775 ( .C1(n9499), .C2(n9498), .A(n9497), .B(n9496), .ZN(n9553)
         );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9553), .S(n9932), .Z(
        P1_U3538) );
  AOI211_X1 U10777 ( .C1(n9502), .C2(n9924), .A(n9501), .B(n9500), .ZN(n9558)
         );
  AOI22_X1 U10778 ( .A1(n9555), .A2(n9503), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9929), .ZN(n9504) );
  OAI21_X1 U10779 ( .B1(n9558), .B2(n9929), .A(n9504), .ZN(P1_U3537) );
  INV_X1 U10780 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9506) );
  MUX2_X1 U10781 ( .A(n9506), .B(n9505), .S(n9927), .Z(n9507) );
  OAI21_X1 U10782 ( .B1(n9508), .B2(n9551), .A(n9507), .ZN(P1_U3521) );
  INV_X1 U10783 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9510) );
  MUX2_X1 U10784 ( .A(n9510), .B(n9509), .S(n9927), .Z(n9511) );
  OAI21_X1 U10785 ( .B1(n9512), .B2(n9551), .A(n9511), .ZN(P1_U3520) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9513), .S(n9927), .Z(
        P1_U3519) );
  INV_X1 U10787 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9515) );
  OAI21_X1 U10788 ( .B1(n9517), .B2(n9551), .A(n9516), .ZN(P1_U3518) );
  INV_X1 U10789 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9519) );
  MUX2_X1 U10790 ( .A(n9519), .B(n9518), .S(n9927), .Z(n9520) );
  OAI21_X1 U10791 ( .B1(n4680), .B2(n9551), .A(n9520), .ZN(P1_U3517) );
  MUX2_X1 U10792 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9521), .S(n9927), .Z(
        P1_U3516) );
  MUX2_X1 U10793 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9522), .S(n9927), .Z(
        P1_U3515) );
  INV_X1 U10794 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9524) );
  MUX2_X1 U10795 ( .A(n9524), .B(n9523), .S(n9927), .Z(n9525) );
  OAI21_X1 U10796 ( .B1(n9526), .B2(n9551), .A(n9525), .ZN(P1_U3514) );
  INV_X1 U10797 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9528) );
  MUX2_X1 U10798 ( .A(n9528), .B(n9527), .S(n9927), .Z(n9529) );
  OAI21_X1 U10799 ( .B1(n9530), .B2(n9551), .A(n9529), .ZN(P1_U3513) );
  INV_X1 U10800 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9532) );
  MUX2_X1 U10801 ( .A(n9532), .B(n9531), .S(n9927), .Z(n9533) );
  OAI21_X1 U10802 ( .B1(n9534), .B2(n9551), .A(n9533), .ZN(P1_U3512) );
  INV_X1 U10803 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10271) );
  MUX2_X1 U10804 ( .A(n10271), .B(n9535), .S(n9927), .Z(n9536) );
  OAI21_X1 U10805 ( .B1(n9537), .B2(n9551), .A(n9536), .ZN(P1_U3511) );
  MUX2_X1 U10806 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9538), .S(n9927), .Z(n9539) );
  INV_X1 U10807 ( .A(n9539), .ZN(n9540) );
  OAI21_X1 U10808 ( .B1(n9541), .B2(n9551), .A(n9540), .ZN(P1_U3510) );
  INV_X1 U10809 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9543) );
  MUX2_X1 U10810 ( .A(n9543), .B(n9542), .S(n9927), .Z(n9544) );
  OAI21_X1 U10811 ( .B1(n9545), .B2(n9551), .A(n9544), .ZN(P1_U3509) );
  MUX2_X1 U10812 ( .A(n10315), .B(n9546), .S(n9927), .Z(n9547) );
  OAI21_X1 U10813 ( .B1(n9548), .B2(n9551), .A(n9547), .ZN(P1_U3507) );
  MUX2_X1 U10814 ( .A(n10051), .B(n9549), .S(n9927), .Z(n9550) );
  OAI21_X1 U10815 ( .B1(n9552), .B2(n9551), .A(n9550), .ZN(P1_U3504) );
  MUX2_X1 U10816 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9553), .S(n9927), .Z(
        P1_U3501) );
  AOI22_X1 U10817 ( .A1(n9555), .A2(n9554), .B1(P1_REG0_REG_15__SCAN_IN), .B2(
        n9557), .ZN(n9556) );
  OAI21_X1 U10818 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(P1_U3498) );
  INV_X1 U10819 ( .A(n9559), .ZN(n9567) );
  INV_X1 U10820 ( .A(n9560), .ZN(n9563) );
  NOR4_X1 U10821 ( .A1(n9563), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9562), .A4(
        P1_U3086), .ZN(n9564) );
  AOI21_X1 U10822 ( .B1(n9565), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9564), .ZN(
        n9566) );
  OAI21_X1 U10823 ( .B1(n9567), .B2(n9575), .A(n9566), .ZN(P1_U3324) );
  OAI222_X1 U10824 ( .A1(n9572), .A2(n10337), .B1(n9575), .B2(n9569), .C1(
        n9568), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U10825 ( .A1(n9572), .A2(n10324), .B1(n9571), .B2(n9570), .C1(
        P1_U3086), .C2(n9721), .ZN(P1_U3328) );
  OAI222_X1 U10826 ( .A1(n9576), .A2(P1_U3086), .B1(n9575), .B2(n9574), .C1(
        n9573), .C2(n9572), .ZN(P1_U3329) );
  MUX2_X1 U10827 ( .A(n9577), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10828 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9592) );
  AND2_X1 U10829 ( .A1(n9579), .A2(n9578), .ZN(n9580) );
  OR3_X1 U10830 ( .A1(n9581), .A2(n9580), .A3(n9816), .ZN(n9587) );
  AND2_X1 U10831 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  OR3_X1 U10832 ( .A1(n9585), .A2(n9584), .A3(n9812), .ZN(n9586) );
  OAI211_X1 U10833 ( .C1(n9848), .C2(n9588), .A(n9587), .B(n9586), .ZN(n9589)
         );
  INV_X1 U10834 ( .A(n9589), .ZN(n9591) );
  OR2_X1 U10835 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9590), .ZN(n9655) );
  OAI211_X1 U10836 ( .C1(n9592), .C2(n9852), .A(n9591), .B(n9655), .ZN(
        P1_U3253) );
  INV_X1 U10837 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n10347) );
  OAI211_X1 U10838 ( .C1(n9595), .C2(n9594), .A(n9841), .B(n9593), .ZN(n9600)
         );
  OAI211_X1 U10839 ( .C1(n9598), .C2(n9597), .A(n9837), .B(n9596), .ZN(n9599)
         );
  OAI211_X1 U10840 ( .C1(n9848), .C2(n9601), .A(n9600), .B(n9599), .ZN(n9602)
         );
  INV_X1 U10841 ( .A(n9602), .ZN(n9603) );
  NAND2_X1 U10842 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9699) );
  OAI211_X1 U10843 ( .C1(n10347), .C2(n9852), .A(n9603), .B(n9699), .ZN(
        P1_U3251) );
  INV_X1 U10844 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10280) );
  NOR2_X1 U10845 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9604) );
  AOI21_X1 U10846 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9604), .ZN(n10026) );
  NOR2_X1 U10847 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9605) );
  AOI21_X1 U10848 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9605), .ZN(n10029) );
  NOR2_X1 U10849 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9606) );
  AOI21_X1 U10850 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9606), .ZN(n10032) );
  NOR2_X1 U10851 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9607) );
  AOI21_X1 U10852 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9607), .ZN(n10035) );
  NOR2_X1 U10853 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9608) );
  AOI21_X1 U10854 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9608), .ZN(n10038) );
  NOR2_X1 U10855 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9609) );
  AOI21_X1 U10856 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9609), .ZN(n10041) );
  NOR2_X1 U10857 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9610) );
  AOI21_X1 U10858 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n9610), .ZN(n10385) );
  NAND2_X1 U10859 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n10015) );
  INV_X1 U10860 ( .A(n10015), .ZN(n10017) );
  NAND2_X1 U10861 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  AOI22_X1 U10862 ( .A1(n10017), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P2_ADDR_REG_1__SCAN_IN), .B2(n10013), .ZN(n10379) );
  NAND2_X1 U10863 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9611) );
  OAI21_X1 U10864 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n9611), .ZN(n10378) );
  NOR2_X1 U10865 ( .A1(n10379), .A2(n10378), .ZN(n10377) );
  AOI21_X1 U10866 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10377), .ZN(n10382) );
  NAND2_X1 U10867 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9612) );
  OAI21_X1 U10868 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n9612), .ZN(n10381) );
  NOR2_X1 U10869 ( .A1(n10382), .A2(n10381), .ZN(n10380) );
  AOI21_X1 U10870 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10380), .ZN(n10384) );
  NAND2_X1 U10871 ( .A1(n10385), .A2(n10384), .ZN(n10383) );
  OAI21_X1 U10872 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10383), .ZN(n9613) );
  NAND2_X1 U10873 ( .A1(n9614), .A2(n9613), .ZN(n10365) );
  INV_X1 U10874 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n10367) );
  OR2_X1 U10875 ( .A1(n9614), .A2(n9613), .ZN(n10366) );
  NAND2_X1 U10876 ( .A1(n10367), .A2(n10366), .ZN(n10363) );
  NAND2_X1 U10877 ( .A1(n10365), .A2(n10363), .ZN(n9616) );
  NOR2_X1 U10878 ( .A1(n9616), .A2(n9615), .ZN(n9617) );
  XNOR2_X1 U10879 ( .A(n9616), .B(n9615), .ZN(n10362) );
  NOR2_X1 U10880 ( .A1(n9618), .A2(n10232), .ZN(n9619) );
  XNOR2_X1 U10881 ( .A(n10232), .B(n9618), .ZN(n10373) );
  NOR2_X1 U10882 ( .A1(n9620), .A2(n10347), .ZN(n9621) );
  INV_X1 U10883 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10376) );
  XNOR2_X1 U10884 ( .A(n10347), .B(n9620), .ZN(n10375) );
  NOR2_X1 U10885 ( .A1(n9622), .A2(n10335), .ZN(n9623) );
  XNOR2_X1 U10886 ( .A(n10335), .B(n9622), .ZN(n10369) );
  NAND2_X1 U10887 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9624) );
  OAI21_X1 U10888 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9624), .ZN(n10046) );
  INV_X1 U10889 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10112) );
  AOI22_X1 U10890 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(n10112), .B1(
        P1_ADDR_REG_11__SCAN_IN), .B2(n10261), .ZN(n10043) );
  AOI21_X1 U10891 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10042), .ZN(n10040) );
  NAND2_X1 U10892 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  OAI21_X1 U10893 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10039), .ZN(n10037) );
  NAND2_X1 U10894 ( .A1(n10038), .A2(n10037), .ZN(n10036) );
  OAI21_X1 U10895 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10036), .ZN(n10034) );
  NAND2_X1 U10896 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  OAI21_X1 U10897 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10033), .ZN(n10031) );
  NAND2_X1 U10898 ( .A1(n10032), .A2(n10031), .ZN(n10030) );
  OAI21_X1 U10899 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10030), .ZN(n10028) );
  NAND2_X1 U10900 ( .A1(n10029), .A2(n10028), .ZN(n10027) );
  OAI21_X1 U10901 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10027), .ZN(n10025) );
  NAND2_X1 U10902 ( .A1(n10026), .A2(n10025), .ZN(n10024) );
  OAI21_X1 U10903 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10024), .ZN(n9625) );
  OR2_X1 U10904 ( .A1(n10280), .A2(n9625), .ZN(n10022) );
  NAND2_X1 U10905 ( .A1(n10023), .A2(n10022), .ZN(n10019) );
  NAND2_X1 U10906 ( .A1(n10280), .A2(n9625), .ZN(n10021) );
  NAND2_X1 U10907 ( .A1(n10019), .A2(n10021), .ZN(n9627) );
  XOR2_X1 U10908 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9626) );
  XNOR2_X1 U10909 ( .A(n9627), .B(n9626), .ZN(ADD_1068_U4) );
  XOR2_X1 U10910 ( .A(n9629), .B(n9635), .Z(n9652) );
  INV_X1 U10911 ( .A(n9630), .ZN(n9644) );
  NAND2_X1 U10912 ( .A1(n9631), .A2(n9992), .ZN(n9649) );
  OAI22_X1 U10913 ( .A1(n9649), .A2(n9634), .B1(n9633), .B2(n9632), .ZN(n9643)
         );
  XNOR2_X1 U10914 ( .A(n9636), .B(n9635), .ZN(n9638) );
  OAI222_X1 U10915 ( .A1(n9642), .A2(n9641), .B1(n9640), .B2(n9639), .C1(n9638), .C2(n9637), .ZN(n9650) );
  AOI211_X1 U10916 ( .C1(n9652), .C2(n9644), .A(n9643), .B(n9650), .ZN(n9646)
         );
  AOI22_X1 U10917 ( .A1(n9648), .A2(n9647), .B1(n9646), .B2(n9645), .ZN(
        P2_U3220) );
  INV_X1 U10918 ( .A(n9649), .ZN(n9651) );
  AOI211_X1 U10919 ( .C1(n9652), .C2(n9968), .A(n9651), .B(n9650), .ZN(n9654)
         );
  AOI22_X1 U10920 ( .A1(n10012), .A2(n9654), .B1(n9653), .B2(n10010), .ZN(
        P2_U3472) );
  INV_X1 U10921 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U10922 ( .A1(n9994), .A2(n10088), .B1(n9654), .B2(n9993), .ZN(
        P2_U3429) );
  OAI21_X1 U10923 ( .B1(n9657), .B2(n9656), .A(n9655), .ZN(n9663) );
  AOI21_X1 U10924 ( .B1(n9659), .B2(n9658), .A(n9688), .ZN(n9661) );
  NOR2_X1 U10925 ( .A1(n9661), .A2(n9660), .ZN(n9662) );
  AOI211_X1 U10926 ( .C1(n9664), .C2(n9716), .A(n9663), .B(n9662), .ZN(n9665)
         );
  OAI21_X1 U10927 ( .B1(n9666), .B2(n9719), .A(n9665), .ZN(P1_U3217) );
  OAI22_X1 U10928 ( .A1(n9670), .A2(n9669), .B1(n9668), .B2(n9667), .ZN(n9856)
         );
  INV_X1 U10929 ( .A(n9671), .ZN(n9675) );
  NAND3_X1 U10930 ( .A1(n9690), .A2(n9673), .A3(n9672), .ZN(n9674) );
  NAND2_X1 U10931 ( .A1(n9675), .A2(n9674), .ZN(n9676) );
  AOI222_X1 U10932 ( .A1(n9716), .A2(n9861), .B1(n9856), .B2(n9713), .C1(n9676), .C2(n6298), .ZN(n9677) );
  NAND2_X1 U10933 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9769) );
  OAI211_X1 U10934 ( .C1(n9719), .C2(n9859), .A(n9677), .B(n9769), .ZN(
        P1_U3224) );
  AOI21_X1 U10935 ( .B1(n9679), .B2(n9678), .A(n4470), .ZN(n9680) );
  INV_X1 U10936 ( .A(n9680), .ZN(n9681) );
  AOI222_X1 U10937 ( .A1(n9716), .A2(n9683), .B1(n9682), .B2(n9713), .C1(n9681), .C2(n6298), .ZN(n9684) );
  NAND2_X1 U10938 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9782) );
  OAI211_X1 U10939 ( .C1(n9719), .C2(n9685), .A(n9684), .B(n9782), .ZN(
        P1_U3234) );
  OR3_X1 U10940 ( .A1(n9688), .A2(n9687), .A3(n9686), .ZN(n9689) );
  NAND2_X1 U10941 ( .A1(n9690), .A2(n9689), .ZN(n9691) );
  AOI222_X1 U10942 ( .A1(n9716), .A2(n9693), .B1(n9692), .B2(n9713), .C1(n9691), .C2(n6298), .ZN(n9694) );
  NAND2_X1 U10943 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9755) );
  OAI211_X1 U10944 ( .C1(n9719), .C2(n9695), .A(n9694), .B(n9755), .ZN(
        P1_U3236) );
  XNOR2_X1 U10945 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10946 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10947 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9706) );
  INV_X1 U10948 ( .A(n9699), .ZN(n9700) );
  AOI21_X1 U10949 ( .B1(n9701), .B2(n9713), .A(n9700), .ZN(n9702) );
  OAI21_X1 U10950 ( .B1(n9704), .B2(n9703), .A(n9702), .ZN(n9705) );
  AOI21_X1 U10951 ( .B1(n9706), .B2(n6298), .A(n9705), .ZN(n9707) );
  OAI21_X1 U10952 ( .B1(n9870), .B2(n9719), .A(n9707), .ZN(P1_U3221) );
  NAND2_X1 U10953 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  XOR2_X1 U10954 ( .A(n9711), .B(n9710), .Z(n9712) );
  AOI222_X1 U10955 ( .A1(n9716), .A2(n9715), .B1(n9714), .B2(n9713), .C1(n9712), .C2(n6298), .ZN(n9718) );
  OAI211_X1 U10956 ( .C1(n9719), .C2(n9883), .A(n9718), .B(n9717), .ZN(
        P1_U3227) );
  INV_X1 U10957 ( .A(n9720), .ZN(n9722) );
  NAND2_X1 U10958 ( .A1(n9721), .A2(n10073), .ZN(n9724) );
  NAND2_X1 U10959 ( .A1(n9722), .A2(n9724), .ZN(n9725) );
  MUX2_X1 U10960 ( .A(n9725), .B(n9724), .S(n9723), .Z(n9727) );
  NAND2_X1 U10961 ( .A1(n9727), .A2(n9726), .ZN(n9730) );
  AOI22_X1 U10962 ( .A1(n9728), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n9729) );
  OAI21_X1 U10963 ( .B1(n9731), .B2(n9730), .A(n9729), .ZN(P1_U3243) );
  INV_X1 U10964 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9745) );
  OAI211_X1 U10965 ( .C1(n9734), .C2(n9733), .A(n9841), .B(n9732), .ZN(n9739)
         );
  OAI211_X1 U10966 ( .C1(n9737), .C2(n9736), .A(n9837), .B(n9735), .ZN(n9738)
         );
  OAI211_X1 U10967 ( .C1(n9848), .C2(n9740), .A(n9739), .B(n9738), .ZN(n9741)
         );
  NOR2_X1 U10968 ( .A1(n9742), .A2(n9741), .ZN(n9744) );
  OAI211_X1 U10969 ( .C1(n9852), .C2(n9745), .A(n9744), .B(n9743), .ZN(
        P1_U3247) );
  AOI211_X1 U10970 ( .C1(n9748), .C2(n9747), .A(n9746), .B(n9816), .ZN(n9753)
         );
  AOI211_X1 U10971 ( .C1(n9751), .C2(n9750), .A(n9749), .B(n9812), .ZN(n9752)
         );
  AOI211_X1 U10972 ( .C1(n9830), .C2(n9754), .A(n9753), .B(n9752), .ZN(n9756)
         );
  OAI211_X1 U10973 ( .C1(n10112), .C2(n9852), .A(n9756), .B(n9755), .ZN(
        P1_U3254) );
  INV_X1 U10974 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9771) );
  OAI21_X1 U10975 ( .B1(n9759), .B2(n9758), .A(n9757), .ZN(n9760) );
  NAND2_X1 U10976 ( .A1(n9841), .A2(n9760), .ZN(n9766) );
  OAI21_X1 U10977 ( .B1(n9763), .B2(n9762), .A(n9761), .ZN(n9764) );
  NAND2_X1 U10978 ( .A1(n9837), .A2(n9764), .ZN(n9765) );
  OAI211_X1 U10979 ( .C1(n9848), .C2(n9767), .A(n9766), .B(n9765), .ZN(n9768)
         );
  INV_X1 U10980 ( .A(n9768), .ZN(n9770) );
  OAI211_X1 U10981 ( .C1(n9771), .C2(n9852), .A(n9770), .B(n9769), .ZN(
        P1_U3255) );
  INV_X1 U10982 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9784) );
  OAI211_X1 U10983 ( .C1(n9774), .C2(n9773), .A(n9841), .B(n9772), .ZN(n9775)
         );
  INV_X1 U10984 ( .A(n9775), .ZN(n9780) );
  AOI211_X1 U10985 ( .C1(n9778), .C2(n9777), .A(n9776), .B(n9816), .ZN(n9779)
         );
  AOI211_X1 U10986 ( .C1(n9830), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9783)
         );
  OAI211_X1 U10987 ( .C1(n9784), .C2(n9852), .A(n9783), .B(n9782), .ZN(
        P1_U3256) );
  INV_X1 U10988 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9797) );
  OAI21_X1 U10989 ( .B1(n9786), .B2(n9785), .A(n9841), .ZN(n9788) );
  NOR2_X1 U10990 ( .A1(n9788), .A2(n9787), .ZN(n9793) );
  AOI211_X1 U10991 ( .C1(n9791), .C2(n9790), .A(n9789), .B(n9816), .ZN(n9792)
         );
  AOI211_X1 U10992 ( .C1(n9830), .C2(n9794), .A(n9793), .B(n9792), .ZN(n9796)
         );
  OAI211_X1 U10993 ( .C1(n9797), .C2(n9852), .A(n9796), .B(n9795), .ZN(
        P1_U3257) );
  INV_X1 U10994 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9809) );
  AOI211_X1 U10995 ( .C1(n9800), .C2(n9799), .A(n9798), .B(n9812), .ZN(n9805)
         );
  AOI211_X1 U10996 ( .C1(n9803), .C2(n9802), .A(n9801), .B(n9816), .ZN(n9804)
         );
  AOI211_X1 U10997 ( .C1(n9830), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9808)
         );
  OAI211_X1 U10998 ( .C1(n9809), .C2(n9852), .A(n9808), .B(n9807), .ZN(
        P1_U3258) );
  INV_X1 U10999 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9824) );
  XNOR2_X1 U11000 ( .A(n9811), .B(n9810), .ZN(n9813) );
  NOR2_X1 U11001 ( .A1(n9813), .A2(n9812), .ZN(n9820) );
  INV_X1 U11002 ( .A(n9814), .ZN(n9815) );
  AOI211_X1 U11003 ( .C1(n9818), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9819)
         );
  AOI211_X1 U11004 ( .C1(n9830), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9823)
         );
  OAI211_X1 U11005 ( .C1(n9824), .C2(n9852), .A(n9823), .B(n9822), .ZN(
        P1_U3259) );
  INV_X1 U11006 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9836) );
  OAI21_X1 U11007 ( .B1(n9827), .B2(n9826), .A(n9825), .ZN(n9833) );
  XNOR2_X1 U11008 ( .A(n9829), .B(n9828), .ZN(n9832) );
  AOI222_X1 U11009 ( .A1(n9833), .A2(n9837), .B1(n9841), .B2(n9832), .C1(n9831), .C2(n9830), .ZN(n9835) );
  OAI211_X1 U11010 ( .C1(n9836), .C2(n9852), .A(n9835), .B(n9834), .ZN(
        P1_U3260) );
  OAI211_X1 U11011 ( .C1(n9840), .C2(n9839), .A(n9838), .B(n9837), .ZN(n9846)
         );
  OAI211_X1 U11012 ( .C1(n9844), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9845)
         );
  OAI211_X1 U11013 ( .C1(n9848), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9849)
         );
  INV_X1 U11014 ( .A(n9849), .ZN(n9851) );
  OAI211_X1 U11015 ( .C1(n10280), .C2(n9852), .A(n9851), .B(n9850), .ZN(
        P1_U3261) );
  INV_X1 U11016 ( .A(n9853), .ZN(n9855) );
  AOI21_X1 U11017 ( .B1(n9855), .B2(n9862), .A(n9854), .ZN(n9858) );
  AOI21_X1 U11018 ( .B1(n9858), .B2(n9857), .A(n9856), .ZN(n9914) );
  INV_X1 U11019 ( .A(n9859), .ZN(n9860) );
  AOI222_X1 U11020 ( .A1(n9861), .A2(n9872), .B1(n9860), .B2(n9894), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(n9421), .ZN(n9869) );
  XNOR2_X1 U11021 ( .A(n9863), .B(n9862), .ZN(n9917) );
  OAI211_X1 U11022 ( .C1(n9866), .C2(n9915), .A(n9865), .B(n9864), .ZN(n9913)
         );
  INV_X1 U11023 ( .A(n9913), .ZN(n9867) );
  AOI22_X1 U11024 ( .A1(n9917), .A2(n9901), .B1(n9867), .B2(n9380), .ZN(n9868)
         );
  OAI211_X1 U11025 ( .C1(n9904), .C2(n9914), .A(n9869), .B(n9868), .ZN(
        P1_U3281) );
  INV_X1 U11026 ( .A(n9870), .ZN(n9871) );
  AOI222_X1 U11027 ( .A1(n9873), .A2(n9872), .B1(n9871), .B2(n9894), .C1(
        P1_REG2_REG_8__SCAN_IN), .C2(n9421), .ZN(n9880) );
  INV_X1 U11028 ( .A(n9874), .ZN(n9877) );
  INV_X1 U11029 ( .A(n9875), .ZN(n9876) );
  AOI22_X1 U11030 ( .A1(n9878), .A2(n9877), .B1(n9380), .B2(n9876), .ZN(n9879)
         );
  OAI211_X1 U11031 ( .C1(n9904), .C2(n9881), .A(n9880), .B(n9879), .ZN(
        P1_U3285) );
  NAND2_X1 U11032 ( .A1(n9882), .A2(n9380), .ZN(n9886) );
  INV_X1 U11033 ( .A(n9883), .ZN(n9884) );
  AOI22_X1 U11034 ( .A1(n9904), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n9884), .B2(
        n9894), .ZN(n9885) );
  OAI211_X1 U11035 ( .C1(n9887), .C2(n9897), .A(n9886), .B(n9885), .ZN(n9888)
         );
  AOI21_X1 U11036 ( .B1(n9889), .B2(n9901), .A(n9888), .ZN(n9890) );
  OAI21_X1 U11037 ( .B1(n9904), .B2(n9891), .A(n9890), .ZN(P1_U3288) );
  NAND2_X1 U11038 ( .A1(n9892), .A2(n9380), .ZN(n9896) );
  INV_X1 U11039 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9893) );
  AOI22_X1 U11040 ( .A1(n9904), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9894), .B2(
        n9893), .ZN(n9895) );
  OAI211_X1 U11041 ( .C1(n9898), .C2(n9897), .A(n9896), .B(n9895), .ZN(n9899)
         );
  AOI21_X1 U11042 ( .B1(n9901), .B2(n9900), .A(n9899), .ZN(n9902) );
  OAI21_X1 U11043 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(P1_U3290) );
  AND2_X1 U11044 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9906), .ZN(P1_U3294) );
  AND2_X1 U11045 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9906), .ZN(P1_U3295) );
  AND2_X1 U11046 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9906), .ZN(P1_U3296) );
  AND2_X1 U11047 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9906), .ZN(P1_U3297) );
  AND2_X1 U11048 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9906), .ZN(P1_U3298) );
  INV_X1 U11049 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10063) );
  NOR2_X1 U11050 ( .A1(n9905), .A2(n10063), .ZN(P1_U3299) );
  AND2_X1 U11051 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9906), .ZN(P1_U3300) );
  AND2_X1 U11052 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9906), .ZN(P1_U3301) );
  AND2_X1 U11053 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9906), .ZN(P1_U3302) );
  AND2_X1 U11054 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9906), .ZN(P1_U3303) );
  AND2_X1 U11055 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9906), .ZN(P1_U3304) );
  AND2_X1 U11056 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9906), .ZN(P1_U3305) );
  AND2_X1 U11057 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9906), .ZN(P1_U3306) );
  INV_X1 U11058 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10239) );
  NOR2_X1 U11059 ( .A1(n9905), .A2(n10239), .ZN(P1_U3307) );
  AND2_X1 U11060 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9906), .ZN(P1_U3308) );
  INV_X1 U11061 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10164) );
  NOR2_X1 U11062 ( .A1(n9905), .A2(n10164), .ZN(P1_U3309) );
  AND2_X1 U11063 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9906), .ZN(P1_U3310) );
  AND2_X1 U11064 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9906), .ZN(P1_U3311) );
  INV_X1 U11065 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10076) );
  NOR2_X1 U11066 ( .A1(n9905), .A2(n10076), .ZN(P1_U3312) );
  INV_X1 U11067 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10085) );
  NOR2_X1 U11068 ( .A1(n9905), .A2(n10085), .ZN(P1_U3313) );
  INV_X1 U11069 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U11070 ( .A1(n9905), .A2(n10215), .ZN(P1_U3314) );
  AND2_X1 U11071 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9906), .ZN(P1_U3315) );
  AND2_X1 U11072 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9906), .ZN(P1_U3316) );
  AND2_X1 U11073 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9906), .ZN(P1_U3317) );
  AND2_X1 U11074 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9906), .ZN(P1_U3318) );
  INV_X1 U11075 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10166) );
  NOR2_X1 U11076 ( .A1(n9905), .A2(n10166), .ZN(P1_U3319) );
  INV_X1 U11077 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10101) );
  NOR2_X1 U11078 ( .A1(n9905), .A2(n10101), .ZN(P1_U3320) );
  INV_X1 U11079 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10176) );
  NOR2_X1 U11080 ( .A1(n9905), .A2(n10176), .ZN(P1_U3321) );
  AND2_X1 U11081 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9906), .ZN(P1_U3322) );
  AND2_X1 U11082 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9906), .ZN(P1_U3323) );
  OAI21_X1 U11083 ( .B1(n9908), .B2(n9921), .A(n9907), .ZN(n9910) );
  AOI211_X1 U11084 ( .C1(n9924), .C2(n9911), .A(n9910), .B(n9909), .ZN(n9928)
         );
  INV_X1 U11085 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9912) );
  AOI22_X1 U11086 ( .A1(n9927), .A2(n9928), .B1(n9912), .B2(n9557), .ZN(
        P1_U3471) );
  OAI211_X1 U11087 ( .C1(n9915), .C2(n9921), .A(n9914), .B(n9913), .ZN(n9916)
         );
  AOI21_X1 U11088 ( .B1(n9917), .B2(n9924), .A(n9916), .ZN(n9930) );
  INV_X1 U11089 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U11090 ( .A1(n9927), .A2(n9930), .B1(n9918), .B2(n9557), .ZN(
        P1_U3489) );
  OAI211_X1 U11091 ( .C1(n9922), .C2(n9921), .A(n9920), .B(n9919), .ZN(n9923)
         );
  AOI21_X1 U11092 ( .B1(n9925), .B2(n9924), .A(n9923), .ZN(n9931) );
  INV_X1 U11093 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U11094 ( .A1(n9927), .A2(n9931), .B1(n9926), .B2(n9557), .ZN(
        P1_U3492) );
  AOI22_X1 U11095 ( .A1(n9932), .A2(n9928), .B1(n10284), .B2(n9929), .ZN(
        P1_U3528) );
  AOI22_X1 U11096 ( .A1(n9932), .A2(n9930), .B1(n9114), .B2(n9929), .ZN(
        P1_U3534) );
  AOI22_X1 U11097 ( .A1(n9932), .A2(n9931), .B1(n10264), .B2(n9929), .ZN(
        P1_U3535) );
  INV_X1 U11098 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n9936) );
  OAI22_X1 U11099 ( .A1(n9933), .A2(n9976), .B1(n5071), .B2(n9980), .ZN(n9934)
         );
  NOR2_X1 U11100 ( .A1(n9935), .A2(n9934), .ZN(n9996) );
  AOI22_X1 U11101 ( .A1(n9994), .A2(n9936), .B1(n9996), .B2(n9993), .ZN(
        P2_U3396) );
  INV_X1 U11102 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U11103 ( .A1(n9938), .A2(n9968), .B1(n9992), .B2(n9937), .ZN(n9939)
         );
  AND2_X1 U11104 ( .A1(n9940), .A2(n9939), .ZN(n9997) );
  AOI22_X1 U11105 ( .A1(n9994), .A2(n9941), .B1(n9997), .B2(n9993), .ZN(
        P2_U3399) );
  INV_X1 U11106 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9947) );
  INV_X1 U11107 ( .A(n9942), .ZN(n9946) );
  OAI21_X1 U11108 ( .B1(n9944), .B2(n9980), .A(n9943), .ZN(n9945) );
  AOI21_X1 U11109 ( .B1(n9946), .B2(n9968), .A(n9945), .ZN(n9998) );
  AOI22_X1 U11110 ( .A1(n9994), .A2(n9947), .B1(n9998), .B2(n9993), .ZN(
        P2_U3402) );
  INV_X1 U11111 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9953) );
  INV_X1 U11112 ( .A(n9948), .ZN(n9952) );
  OAI22_X1 U11113 ( .A1(n9950), .A2(n9986), .B1(n9949), .B2(n9980), .ZN(n9951)
         );
  NOR2_X1 U11114 ( .A1(n9952), .A2(n9951), .ZN(n9999) );
  AOI22_X1 U11115 ( .A1(n9994), .A2(n9953), .B1(n9999), .B2(n9993), .ZN(
        P2_U3405) );
  INV_X1 U11116 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10124) );
  INV_X1 U11117 ( .A(n9954), .ZN(n9958) );
  OAI22_X1 U11118 ( .A1(n9956), .A2(n9986), .B1(n9955), .B2(n9980), .ZN(n9957)
         );
  NOR2_X1 U11119 ( .A1(n9958), .A2(n9957), .ZN(n10001) );
  AOI22_X1 U11120 ( .A1(n9994), .A2(n10124), .B1(n10001), .B2(n9993), .ZN(
        P2_U3408) );
  INV_X1 U11121 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9963) );
  OAI22_X1 U11122 ( .A1(n9960), .A2(n9976), .B1(n9959), .B2(n9980), .ZN(n9961)
         );
  NOR2_X1 U11123 ( .A1(n9962), .A2(n9961), .ZN(n10003) );
  AOI22_X1 U11124 ( .A1(n9994), .A2(n9963), .B1(n10003), .B2(n9993), .ZN(
        P2_U3411) );
  INV_X1 U11125 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9969) );
  OAI21_X1 U11126 ( .B1(n9965), .B2(n9980), .A(n9964), .ZN(n9966) );
  AOI21_X1 U11127 ( .B1(n9968), .B2(n9967), .A(n9966), .ZN(n10005) );
  AOI22_X1 U11128 ( .A1(n9994), .A2(n9969), .B1(n10005), .B2(n9993), .ZN(
        P2_U3414) );
  INV_X1 U11129 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9974) );
  OAI22_X1 U11130 ( .A1(n9971), .A2(n9976), .B1(n9970), .B2(n9980), .ZN(n9972)
         );
  NOR2_X1 U11131 ( .A1(n9973), .A2(n9972), .ZN(n10006) );
  AOI22_X1 U11132 ( .A1(n9994), .A2(n9974), .B1(n10006), .B2(n9993), .ZN(
        P2_U3417) );
  INV_X1 U11133 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10155) );
  OAI22_X1 U11134 ( .A1(n9977), .A2(n9976), .B1(n9975), .B2(n9980), .ZN(n9978)
         );
  NOR2_X1 U11135 ( .A1(n9979), .A2(n9978), .ZN(n10007) );
  AOI22_X1 U11136 ( .A1(n9994), .A2(n10155), .B1(n10007), .B2(n9993), .ZN(
        P2_U3420) );
  INV_X1 U11137 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9985) );
  OAI22_X1 U11138 ( .A1(n9982), .A2(n9986), .B1(n9981), .B2(n9980), .ZN(n9984)
         );
  NOR2_X1 U11139 ( .A1(n9984), .A2(n9983), .ZN(n10009) );
  AOI22_X1 U11140 ( .A1(n9994), .A2(n9985), .B1(n10009), .B2(n9993), .ZN(
        P2_U3423) );
  INV_X1 U11141 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10152) );
  NOR3_X1 U11142 ( .A1(n9988), .A2(n9987), .A3(n9986), .ZN(n9990) );
  AOI211_X1 U11143 ( .C1(n9992), .C2(n9991), .A(n9990), .B(n9989), .ZN(n10011)
         );
  AOI22_X1 U11144 ( .A1(n9994), .A2(n10152), .B1(n10011), .B2(n9993), .ZN(
        P2_U3426) );
  AOI22_X1 U11145 ( .A1(n10012), .A2(n9996), .B1(n9995), .B2(n10010), .ZN(
        P2_U3461) );
  AOI22_X1 U11146 ( .A1(n10012), .A2(n9997), .B1(n10128), .B2(n10010), .ZN(
        P2_U3462) );
  AOI22_X1 U11147 ( .A1(n10012), .A2(n9998), .B1(n6352), .B2(n10010), .ZN(
        P2_U3463) );
  AOI22_X1 U11148 ( .A1(n10012), .A2(n9999), .B1(n10279), .B2(n10010), .ZN(
        P2_U3464) );
  AOI22_X1 U11149 ( .A1(n10012), .A2(n10001), .B1(n10000), .B2(n10010), .ZN(
        P2_U3465) );
  AOI22_X1 U11150 ( .A1(n10012), .A2(n10003), .B1(n10002), .B2(n10010), .ZN(
        P2_U3466) );
  AOI22_X1 U11151 ( .A1(n10012), .A2(n10005), .B1(n10004), .B2(n10010), .ZN(
        P2_U3467) );
  AOI22_X1 U11152 ( .A1(n10012), .A2(n10006), .B1(n10287), .B2(n10010), .ZN(
        P2_U3468) );
  AOI22_X1 U11153 ( .A1(n10012), .A2(n10007), .B1(n7240), .B2(n10010), .ZN(
        P2_U3469) );
  AOI22_X1 U11154 ( .A1(n10012), .A2(n10009), .B1(n10008), .B2(n10010), .ZN(
        P2_U3470) );
  AOI22_X1 U11155 ( .A1(n10012), .A2(n10011), .B1(n7494), .B2(n10010), .ZN(
        P2_U3471) );
  OAI21_X1 U11156 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(n10016) );
  XNOR2_X1 U11157 ( .A(n10016), .B(P2_ADDR_REG_1__SCAN_IN), .ZN(ADD_1068_U5)
         );
  INV_X1 U11158 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10018) );
  INV_X1 U11159 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10229) );
  AOI21_X1 U11160 ( .B1(n10018), .B2(n10229), .A(n10017), .ZN(ADD_1068_U46) );
  INV_X1 U11161 ( .A(n10021), .ZN(n10020) );
  OAI222_X1 U11162 ( .A1(n10023), .A2(n10022), .B1(n10023), .B2(n10021), .C1(
        n10020), .C2(n10019), .ZN(ADD_1068_U55) );
  OAI21_X1 U11163 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(ADD_1068_U56) );
  OAI21_X1 U11164 ( .B1(n10029), .B2(n10028), .A(n10027), .ZN(ADD_1068_U57) );
  OAI21_X1 U11165 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(ADD_1068_U58) );
  OAI21_X1 U11166 ( .B1(n10035), .B2(n10034), .A(n10033), .ZN(ADD_1068_U59) );
  OAI21_X1 U11167 ( .B1(n10038), .B2(n10037), .A(n10036), .ZN(ADD_1068_U60) );
  OAI21_X1 U11168 ( .B1(n10041), .B2(n10040), .A(n10039), .ZN(ADD_1068_U61) );
  AOI21_X1 U11169 ( .B1(n10044), .B2(n10043), .A(n10042), .ZN(ADD_1068_U62) );
  AOI21_X1 U11170 ( .B1(n10047), .B2(n10046), .A(n10045), .ZN(ADD_1068_U63) );
  MUX2_X1 U11171 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10048), .S(P1_U3973), .Z(
        n10258) );
  AOI22_X1 U11172 ( .A1(n10051), .A2(keyinput111), .B1(keyinput4), .B2(n10050), 
        .ZN(n10049) );
  OAI221_X1 U11173 ( .B1(n10051), .B2(keyinput111), .C1(n10050), .C2(keyinput4), .A(n10049), .ZN(n10059) );
  AOI22_X1 U11174 ( .A1(n9415), .A2(keyinput103), .B1(keyinput55), .B2(n5278), 
        .ZN(n10052) );
  OAI221_X1 U11175 ( .B1(n9415), .B2(keyinput103), .C1(n5278), .C2(keyinput55), 
        .A(n10052), .ZN(n10058) );
  AOI22_X1 U11176 ( .A1(n5768), .A2(keyinput81), .B1(keyinput33), .B2(n10312), 
        .ZN(n10053) );
  OAI221_X1 U11177 ( .B1(n5768), .B2(keyinput81), .C1(n10312), .C2(keyinput33), 
        .A(n10053), .ZN(n10057) );
  AOI22_X1 U11178 ( .A1(n4978), .A2(keyinput3), .B1(keyinput87), .B2(n10055), 
        .ZN(n10054) );
  OAI221_X1 U11179 ( .B1(n4978), .B2(keyinput3), .C1(n10055), .C2(keyinput87), 
        .A(n10054), .ZN(n10056) );
  NOR4_X1 U11180 ( .A1(n10059), .A2(n10058), .A3(n10057), .A4(n10056), .ZN(
        n10098) );
  AOI22_X1 U11181 ( .A1(n10061), .A2(keyinput57), .B1(keyinput64), .B2(n6631), 
        .ZN(n10060) );
  OAI221_X1 U11182 ( .B1(n10061), .B2(keyinput57), .C1(n6631), .C2(keyinput64), 
        .A(n10060), .ZN(n10071) );
  AOI22_X1 U11183 ( .A1(n10063), .A2(keyinput122), .B1(keyinput105), .B2(
        n10316), .ZN(n10062) );
  OAI221_X1 U11184 ( .B1(n10063), .B2(keyinput122), .C1(n10316), .C2(
        keyinput105), .A(n10062), .ZN(n10070) );
  XOR2_X1 U11185 ( .A(n10064), .B(keyinput72), .Z(n10068) );
  XNOR2_X1 U11186 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(keyinput13), .ZN(n10067)
         );
  XNOR2_X1 U11187 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput88), .ZN(n10066)
         );
  XNOR2_X1 U11188 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput114), .ZN(n10065) );
  NAND4_X1 U11189 ( .A1(n10068), .A2(n10067), .A3(n10066), .A4(n10065), .ZN(
        n10069) );
  NOR3_X1 U11190 ( .A1(n10071), .A2(n10070), .A3(n10069), .ZN(n10097) );
  AOI22_X1 U11191 ( .A1(n10073), .A2(keyinput112), .B1(n10262), .B2(
        keyinput113), .ZN(n10072) );
  OAI221_X1 U11192 ( .B1(n10073), .B2(keyinput112), .C1(n10262), .C2(
        keyinput113), .A(n10072), .ZN(n10082) );
  AOI22_X1 U11193 ( .A1(n10279), .A2(keyinput35), .B1(n5779), .B2(keyinput75), 
        .ZN(n10074) );
  OAI221_X1 U11194 ( .B1(n10279), .B2(keyinput35), .C1(n5779), .C2(keyinput75), 
        .A(n10074), .ZN(n10081) );
  AOI22_X1 U11195 ( .A1(n10076), .A2(keyinput34), .B1(keyinput107), .B2(n10259), .ZN(n10075) );
  OAI221_X1 U11196 ( .B1(n10076), .B2(keyinput34), .C1(n10259), .C2(
        keyinput107), .A(n10075), .ZN(n10080) );
  XNOR2_X1 U11197 ( .A(SI_0_), .B(keyinput101), .ZN(n10078) );
  XNOR2_X1 U11198 ( .A(SI_28_), .B(keyinput49), .ZN(n10077) );
  NAND2_X1 U11199 ( .A1(n10078), .A2(n10077), .ZN(n10079) );
  NOR4_X1 U11200 ( .A1(n10082), .A2(n10081), .A3(n10080), .A4(n10079), .ZN(
        n10096) );
  AOI22_X1 U11201 ( .A1(n5253), .A2(keyinput102), .B1(keyinput47), .B2(n10261), 
        .ZN(n10083) );
  OAI221_X1 U11202 ( .B1(n5253), .B2(keyinput102), .C1(n10261), .C2(keyinput47), .A(n10083), .ZN(n10094) );
  AOI22_X1 U11203 ( .A1(n5578), .A2(keyinput28), .B1(n10085), .B2(keyinput79), 
        .ZN(n10084) );
  OAI221_X1 U11204 ( .B1(n5578), .B2(keyinput28), .C1(n10085), .C2(keyinput79), 
        .A(n10084), .ZN(n10093) );
  AOI22_X1 U11205 ( .A1(n10088), .A2(keyinput98), .B1(n10087), .B2(keyinput83), 
        .ZN(n10086) );
  OAI221_X1 U11206 ( .B1(n10088), .B2(keyinput98), .C1(n10087), .C2(keyinput83), .A(n10086), .ZN(n10092) );
  XOR2_X1 U11207 ( .A(n7243), .B(keyinput115), .Z(n10090) );
  XNOR2_X1 U11208 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput61), .ZN(n10089) );
  NAND2_X1 U11209 ( .A1(n10090), .A2(n10089), .ZN(n10091) );
  NOR4_X1 U11210 ( .A1(n10094), .A2(n10093), .A3(n10092), .A4(n10091), .ZN(
        n10095) );
  NAND4_X1 U11211 ( .A1(n10098), .A2(n10097), .A3(n10096), .A4(n10095), .ZN(
        n10256) );
  AOI22_X1 U11212 ( .A1(n9359), .A2(keyinput31), .B1(keyinput69), .B2(n6952), 
        .ZN(n10099) );
  OAI221_X1 U11213 ( .B1(n9359), .B2(keyinput31), .C1(n6952), .C2(keyinput69), 
        .A(n10099), .ZN(n10109) );
  AOI22_X1 U11214 ( .A1(n10101), .A2(keyinput66), .B1(keyinput10), .B2(n10266), 
        .ZN(n10100) );
  OAI221_X1 U11215 ( .B1(n10101), .B2(keyinput66), .C1(n10266), .C2(keyinput10), .A(n10100), .ZN(n10104) );
  XNOR2_X1 U11216 ( .A(n10335), .B(keyinput116), .ZN(n10103) );
  XNOR2_X1 U11217 ( .A(n10267), .B(keyinput42), .ZN(n10102) );
  OR3_X1 U11218 ( .A1(n10104), .A2(n10103), .A3(n10102), .ZN(n10108) );
  AOI22_X1 U11219 ( .A1(n10106), .A2(keyinput5), .B1(keyinput53), .B2(n7308), 
        .ZN(n10105) );
  OAI221_X1 U11220 ( .B1(n10106), .B2(keyinput5), .C1(n7308), .C2(keyinput53), 
        .A(n10105), .ZN(n10107) );
  NOR3_X1 U11221 ( .A1(n10109), .A2(n10108), .A3(n10107), .ZN(n10149) );
  INV_X1 U11222 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10270) );
  AOI22_X1 U11223 ( .A1(n10270), .A2(keyinput17), .B1(keyinput30), .B2(n10269), 
        .ZN(n10110) );
  OAI221_X1 U11224 ( .B1(n10270), .B2(keyinput17), .C1(n10269), .C2(keyinput30), .A(n10110), .ZN(n10121) );
  AOI22_X1 U11225 ( .A1(n5741), .A2(keyinput37), .B1(keyinput78), .B2(n10271), 
        .ZN(n10111) );
  OAI221_X1 U11226 ( .B1(n5741), .B2(keyinput37), .C1(n10271), .C2(keyinput78), 
        .A(n10111), .ZN(n10116) );
  XNOR2_X1 U11227 ( .A(n10112), .B(keyinput60), .ZN(n10115) );
  XNOR2_X1 U11228 ( .A(n10113), .B(keyinput92), .ZN(n10114) );
  OR3_X1 U11229 ( .A1(n10116), .A2(n10115), .A3(n10114), .ZN(n10120) );
  AOI22_X1 U11230 ( .A1(n10118), .A2(keyinput2), .B1(keyinput7), .B2(n6481), 
        .ZN(n10117) );
  OAI221_X1 U11231 ( .B1(n10118), .B2(keyinput2), .C1(n6481), .C2(keyinput7), 
        .A(n10117), .ZN(n10119) );
  NOR3_X1 U11232 ( .A1(n10121), .A2(n10120), .A3(n10119), .ZN(n10148) );
  AOI22_X1 U11233 ( .A1(n10343), .A2(keyinput25), .B1(keyinput106), .B2(n8423), 
        .ZN(n10122) );
  OAI221_X1 U11234 ( .B1(n10343), .B2(keyinput25), .C1(n8423), .C2(keyinput106), .A(n10122), .ZN(n10134) );
  AOI22_X1 U11235 ( .A1(n10125), .A2(keyinput9), .B1(keyinput124), .B2(n10124), 
        .ZN(n10123) );
  OAI221_X1 U11236 ( .B1(n10125), .B2(keyinput9), .C1(n10124), .C2(keyinput124), .A(n10123), .ZN(n10133) );
  INV_X1 U11237 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U11238 ( .A1(n10264), .A2(keyinput0), .B1(n10127), .B2(keyinput117), 
        .ZN(n10126) );
  OAI221_X1 U11239 ( .B1(n10264), .B2(keyinput0), .C1(n10127), .C2(keyinput117), .A(n10126), .ZN(n10132) );
  XOR2_X1 U11240 ( .A(n10128), .B(keyinput89), .Z(n10130) );
  XNOR2_X1 U11241 ( .A(P2_IR_REG_28__SCAN_IN), .B(keyinput38), .ZN(n10129) );
  NAND2_X1 U11242 ( .A1(n10130), .A2(n10129), .ZN(n10131) );
  NOR4_X1 U11243 ( .A1(n10134), .A2(n10133), .A3(n10132), .A4(n10131), .ZN(
        n10147) );
  INV_X1 U11244 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U11245 ( .A1(n10344), .A2(keyinput16), .B1(n10136), .B2(keyinput100), .ZN(n10135) );
  OAI221_X1 U11246 ( .B1(n10344), .B2(keyinput16), .C1(n10136), .C2(
        keyinput100), .A(n10135), .ZN(n10145) );
  AOI22_X1 U11247 ( .A1(n10337), .A2(keyinput6), .B1(n10138), .B2(keyinput119), 
        .ZN(n10137) );
  OAI221_X1 U11248 ( .B1(n10337), .B2(keyinput6), .C1(n10138), .C2(keyinput119), .A(n10137), .ZN(n10144) );
  XNOR2_X1 U11249 ( .A(P1_REG2_REG_2__SCAN_IN), .B(keyinput86), .ZN(n10142) );
  XNOR2_X1 U11250 ( .A(P2_IR_REG_22__SCAN_IN), .B(keyinput73), .ZN(n10141) );
  XNOR2_X1 U11251 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput46), .ZN(n10140)
         );
  XNOR2_X1 U11252 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput70), .ZN(n10139) );
  NAND4_X1 U11253 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10143) );
  NOR3_X1 U11254 ( .A1(n10145), .A2(n10144), .A3(n10143), .ZN(n10146) );
  NAND4_X1 U11255 ( .A1(n10149), .A2(n10148), .A3(n10147), .A4(n10146), .ZN(
        n10255) );
  AOI22_X1 U11256 ( .A1(n10152), .A2(keyinput59), .B1(n10151), .B2(keyinput23), 
        .ZN(n10150) );
  OAI221_X1 U11257 ( .B1(n10152), .B2(keyinput59), .C1(n10151), .C2(keyinput23), .A(n10150), .ZN(n10162) );
  INV_X1 U11258 ( .A(SI_21_), .ZN(n10311) );
  AOI22_X1 U11259 ( .A1(n10311), .A2(keyinput84), .B1(keyinput125), .B2(n10154), .ZN(n10153) );
  OAI221_X1 U11260 ( .B1(n10311), .B2(keyinput84), .C1(n10154), .C2(
        keyinput125), .A(n10153), .ZN(n10161) );
  XOR2_X1 U11261 ( .A(n10155), .B(keyinput45), .Z(n10159) );
  XNOR2_X1 U11262 ( .A(P1_REG3_REG_10__SCAN_IN), .B(keyinput74), .ZN(n10158)
         );
  XNOR2_X1 U11263 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput14), .ZN(n10157) );
  XNOR2_X1 U11264 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput11), .ZN(n10156) );
  NAND4_X1 U11265 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  NOR3_X1 U11266 ( .A1(n10162), .A2(n10161), .A3(n10160), .ZN(n10203) );
  AOI22_X1 U11267 ( .A1(n10164), .A2(keyinput65), .B1(keyinput126), .B2(n10327), .ZN(n10163) );
  OAI221_X1 U11268 ( .B1(n10164), .B2(keyinput65), .C1(n10327), .C2(
        keyinput126), .A(n10163), .ZN(n10173) );
  AOI22_X1 U11269 ( .A1(n10336), .A2(keyinput91), .B1(n10166), .B2(keyinput58), 
        .ZN(n10165) );
  OAI221_X1 U11270 ( .B1(n10336), .B2(keyinput91), .C1(n10166), .C2(keyinput58), .A(n10165), .ZN(n10172) );
  AOI22_X1 U11271 ( .A1(n10168), .A2(keyinput121), .B1(keyinput15), .B2(n5293), 
        .ZN(n10167) );
  OAI221_X1 U11272 ( .B1(n10168), .B2(keyinput121), .C1(n5293), .C2(keyinput15), .A(n10167), .ZN(n10171) );
  AOI22_X1 U11273 ( .A1(n10347), .A2(keyinput118), .B1(n10323), .B2(keyinput94), .ZN(n10169) );
  OAI221_X1 U11274 ( .B1(n10347), .B2(keyinput118), .C1(n10323), .C2(
        keyinput94), .A(n10169), .ZN(n10170) );
  NOR4_X1 U11275 ( .A1(n10173), .A2(n10172), .A3(n10171), .A4(n10170), .ZN(
        n10202) );
  AOI22_X1 U11276 ( .A1(n10176), .A2(keyinput21), .B1(keyinput67), .B2(n10175), 
        .ZN(n10174) );
  OAI221_X1 U11277 ( .B1(n10176), .B2(keyinput21), .C1(n10175), .C2(keyinput67), .A(n10174), .ZN(n10187) );
  AOI22_X1 U11278 ( .A1(n10179), .A2(keyinput51), .B1(n10178), .B2(keyinput48), 
        .ZN(n10177) );
  OAI221_X1 U11279 ( .B1(n10179), .B2(keyinput51), .C1(n10178), .C2(keyinput48), .A(n10177), .ZN(n10186) );
  AOI22_X1 U11280 ( .A1(n10340), .A2(keyinput44), .B1(n10181), .B2(keyinput85), 
        .ZN(n10180) );
  OAI221_X1 U11281 ( .B1(n10340), .B2(keyinput44), .C1(n10181), .C2(keyinput85), .A(n10180), .ZN(n10185) );
  XNOR2_X1 U11282 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(keyinput18), .ZN(n10183)
         );
  XNOR2_X1 U11283 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput68), .ZN(n10182)
         );
  NAND2_X1 U11284 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  NOR4_X1 U11285 ( .A1(n10187), .A2(n10186), .A3(n10185), .A4(n10184), .ZN(
        n10201) );
  AOI22_X1 U11286 ( .A1(n10190), .A2(keyinput120), .B1(n10189), .B2(keyinput1), 
        .ZN(n10188) );
  OAI221_X1 U11287 ( .B1(n10190), .B2(keyinput120), .C1(n10189), .C2(keyinput1), .A(n10188), .ZN(n10199) );
  AOI22_X1 U11288 ( .A1(n10308), .A2(keyinput29), .B1(n10192), .B2(keyinput93), 
        .ZN(n10191) );
  OAI221_X1 U11289 ( .B1(n10308), .B2(keyinput29), .C1(n10192), .C2(keyinput93), .A(n10191), .ZN(n10198) );
  AOI22_X1 U11290 ( .A1(n6243), .A2(keyinput27), .B1(n10295), .B2(keyinput110), 
        .ZN(n10193) );
  OAI221_X1 U11291 ( .B1(n6243), .B2(keyinput27), .C1(n10295), .C2(keyinput110), .A(n10193), .ZN(n10197) );
  XNOR2_X1 U11292 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput95), .ZN(n10195)
         );
  XNOR2_X1 U11293 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput32), .ZN(n10194)
         );
  NAND2_X1 U11294 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  NOR4_X1 U11295 ( .A1(n10199), .A2(n10198), .A3(n10197), .A4(n10196), .ZN(
        n10200) );
  NAND4_X1 U11296 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10254) );
  INV_X1 U11297 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U11298 ( .A1(n10298), .A2(keyinput36), .B1(keyinput96), .B2(n10205), 
        .ZN(n10204) );
  OAI221_X1 U11299 ( .B1(n10298), .B2(keyinput36), .C1(n10205), .C2(keyinput96), .A(n10204), .ZN(n10213) );
  AOI22_X1 U11300 ( .A1(n5948), .A2(keyinput41), .B1(n10294), .B2(keyinput99), 
        .ZN(n10206) );
  OAI221_X1 U11301 ( .B1(n5948), .B2(keyinput41), .C1(n10294), .C2(keyinput99), 
        .A(n10206), .ZN(n10212) );
  AOI22_X1 U11302 ( .A1(n10299), .A2(keyinput104), .B1(n10300), .B2(keyinput20), .ZN(n10207) );
  OAI221_X1 U11303 ( .B1(n10299), .B2(keyinput104), .C1(n10300), .C2(
        keyinput20), .A(n10207), .ZN(n10211) );
  XNOR2_X1 U11304 ( .A(P2_REG1_REG_25__SCAN_IN), .B(keyinput56), .ZN(n10209)
         );
  XNOR2_X1 U11305 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput90), .ZN(n10208) );
  NAND2_X1 U11306 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  NOR4_X1 U11307 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10252) );
  AOI22_X1 U11308 ( .A1(n10284), .A2(keyinput54), .B1(keyinput123), .B2(n10283), .ZN(n10214) );
  OAI221_X1 U11309 ( .B1(n10284), .B2(keyinput54), .C1(n10283), .C2(
        keyinput123), .A(n10214), .ZN(n10219) );
  XNOR2_X1 U11310 ( .A(n10215), .B(keyinput82), .ZN(n10218) );
  XNOR2_X1 U11311 ( .A(n10216), .B(keyinput62), .ZN(n10217) );
  OR3_X1 U11312 ( .A1(n10219), .A2(n10218), .A3(n10217), .ZN(n10225) );
  AOI22_X1 U11313 ( .A1(n10221), .A2(keyinput77), .B1(n5900), .B2(keyinput40), 
        .ZN(n10220) );
  OAI221_X1 U11314 ( .B1(n10221), .B2(keyinput77), .C1(n5900), .C2(keyinput40), 
        .A(n10220), .ZN(n10224) );
  INV_X1 U11315 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11316 ( .A1(n10296), .A2(keyinput22), .B1(n10297), .B2(keyinput71), 
        .ZN(n10222) );
  OAI221_X1 U11317 ( .B1(n10296), .B2(keyinput22), .C1(n10297), .C2(keyinput71), .A(n10222), .ZN(n10223) );
  NOR3_X1 U11318 ( .A1(n10225), .A2(n10224), .A3(n10223), .ZN(n10251) );
  AOI22_X1 U11319 ( .A1(n10285), .A2(keyinput63), .B1(n10282), .B2(keyinput43), 
        .ZN(n10226) );
  OAI221_X1 U11320 ( .B1(n10285), .B2(keyinput63), .C1(n10282), .C2(keyinput43), .A(n10226), .ZN(n10236) );
  AOI22_X1 U11321 ( .A1(n10280), .A2(keyinput26), .B1(n10281), .B2(keyinput80), 
        .ZN(n10227) );
  OAI221_X1 U11322 ( .B1(n10280), .B2(keyinput26), .C1(n10281), .C2(keyinput80), .A(n10227), .ZN(n10235) );
  AOI22_X1 U11323 ( .A1(n10230), .A2(keyinput76), .B1(keyinput50), .B2(n10229), 
        .ZN(n10228) );
  OAI221_X1 U11324 ( .B1(n10230), .B2(keyinput76), .C1(n10229), .C2(keyinput50), .A(n10228), .ZN(n10234) );
  AOI22_X1 U11325 ( .A1(n10288), .A2(keyinput109), .B1(keyinput12), .B2(n10232), .ZN(n10231) );
  OAI221_X1 U11326 ( .B1(n10288), .B2(keyinput109), .C1(n10232), .C2(
        keyinput12), .A(n10231), .ZN(n10233) );
  NOR4_X1 U11327 ( .A1(n10236), .A2(n10235), .A3(n10234), .A4(n10233), .ZN(
        n10250) );
  AOI22_X1 U11328 ( .A1(n10287), .A2(keyinput127), .B1(n5621), .B2(keyinput39), 
        .ZN(n10237) );
  OAI221_X1 U11329 ( .B1(n10287), .B2(keyinput127), .C1(n5621), .C2(keyinput39), .A(n10237), .ZN(n10248) );
  AOI22_X1 U11330 ( .A1(n10286), .A2(keyinput8), .B1(n10239), .B2(keyinput19), 
        .ZN(n10238) );
  OAI221_X1 U11331 ( .B1(n10286), .B2(keyinput8), .C1(n10239), .C2(keyinput19), 
        .A(n10238), .ZN(n10247) );
  AOI22_X1 U11332 ( .A1(n10242), .A2(keyinput97), .B1(keyinput52), .B2(n10241), 
        .ZN(n10240) );
  OAI221_X1 U11333 ( .B1(n10242), .B2(keyinput97), .C1(n10241), .C2(keyinput52), .A(n10240), .ZN(n10246) );
  INV_X1 U11334 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n10325) );
  AOI22_X1 U11335 ( .A1(n10325), .A2(keyinput108), .B1(keyinput24), .B2(n10244), .ZN(n10243) );
  OAI221_X1 U11336 ( .B1(n10325), .B2(keyinput108), .C1(n10244), .C2(
        keyinput24), .A(n10243), .ZN(n10245) );
  NOR4_X1 U11337 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10249) );
  NAND4_X1 U11338 ( .A1(n10252), .A2(n10251), .A3(n10250), .A4(n10249), .ZN(
        n10253) );
  NOR4_X1 U11339 ( .A1(n10256), .A2(n10255), .A3(n10254), .A4(n10253), .ZN(
        n10257) );
  XOR2_X1 U11340 ( .A(n10258), .B(n10257), .Z(n10360) );
  NOR4_X1 U11341 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(SI_0_), .A3(SI_28_), 
        .A4(P1_REG3_REG_2__SCAN_IN), .ZN(n10260) );
  NAND3_X1 U11342 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(n10260), .A3(n10259), 
        .ZN(n10278) );
  NAND4_X1 U11343 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .A3(n10262), .A4(n10261), .ZN(n10263) );
  NOR3_X1 U11344 ( .A1(SI_12_), .A2(P1_REG3_REG_12__SCAN_IN), .A3(n10263), 
        .ZN(n10276) );
  NAND4_X1 U11345 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P2_REG0_REG_20__SCAN_IN), 
        .A3(P2_REG0_REG_6__SCAN_IN), .A4(n10264), .ZN(n10265) );
  NOR3_X1 U11346 ( .A1(n10266), .A2(n10265), .A3(P2_REG2_REG_4__SCAN_IN), .ZN(
        n10268) );
  NAND3_X1 U11347 ( .A1(n10268), .A2(P1_REG2_REG_19__SCAN_IN), .A3(n10267), 
        .ZN(n10274) );
  NAND4_X1 U11348 ( .A1(SI_17_), .A2(P1_REG2_REG_10__SCAN_IN), .A3(n10270), 
        .A4(n10269), .ZN(n10273) );
  NAND4_X1 U11349 ( .A1(SI_3_), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P1_ADDR_REG_11__SCAN_IN), .A4(n10271), .ZN(n10272) );
  NOR3_X1 U11350 ( .A1(n10274), .A2(n10273), .A3(n10272), .ZN(n10275) );
  NAND4_X1 U11351 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10276), .A3(n10275), .A4(
        n5578), .ZN(n10277) );
  NOR4_X1 U11352 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10279), .A3(n10278), .A4(
        n10277), .ZN(n10358) );
  NAND4_X1 U11353 ( .A1(P1_REG1_REG_30__SCAN_IN), .A2(n10282), .A3(n10281), 
        .A4(n10280), .ZN(n10292) );
  NAND4_X1 U11354 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(n10285), .A3(n10284), 
        .A4(n10283), .ZN(n10291) );
  NAND4_X1 U11355 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_DATAO_REG_15__SCAN_IN), 
        .A3(P2_DATAO_REG_12__SCAN_IN), .A4(P2_REG2_REG_19__SCAN_IN), .ZN(
        n10290) );
  NAND4_X1 U11356 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(n10288), .A3(n10287), .A4(
        n10286), .ZN(n10289) );
  NOR4_X1 U11357 ( .A1(n10292), .A2(n10291), .A3(n10290), .A4(n10289), .ZN(
        n10357) );
  NAND4_X1 U11358 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(P1_REG1_REG_9__SCAN_IN), 
        .A3(n10294), .A4(n10293), .ZN(n10304) );
  NAND4_X1 U11359 ( .A1(P1_REG2_REG_26__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .A3(P2_REG0_REG_24__SCAN_IN), .A4(n10295), .ZN(n10303) );
  NAND4_X1 U11360 ( .A1(P2_REG1_REG_25__SCAN_IN), .A2(P2_DATAO_REG_30__SCAN_IN), .A3(n10297), .A4(n10296), .ZN(n10302) );
  NAND4_X1 U11361 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(n10300), .A3(n10299), .A4(
        n10298), .ZN(n10301) );
  NOR4_X1 U11362 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10356) );
  INV_X1 U11363 ( .A(n10305), .ZN(n10354) );
  INV_X1 U11364 ( .A(n10306), .ZN(n10353) );
  INV_X1 U11365 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10307) );
  NAND4_X1 U11366 ( .A1(n10307), .A2(P1_REG2_REG_25__SCAN_IN), .A3(
        P1_REG3_REG_10__SCAN_IN), .A4(P2_DATAO_REG_6__SCAN_IN), .ZN(n10334) );
  NOR2_X1 U11367 ( .A1(P1_REG0_REG_4__SCAN_IN), .A2(n10308), .ZN(n10322) );
  INV_X1 U11368 ( .A(n10309), .ZN(n10310) );
  AND2_X1 U11369 ( .A1(n10310), .A2(n4978), .ZN(n10321) );
  NAND4_X1 U11370 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(SI_11_), .A3(
        P2_REG0_REG_12__SCAN_IN), .A4(n10311), .ZN(n10314) );
  NAND4_X1 U11371 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(P2_REG3_REG_26__SCAN_IN), 
        .A3(P2_REG3_REG_13__SCAN_IN), .A4(n10312), .ZN(n10313) );
  NOR2_X1 U11372 ( .A1(n10314), .A2(n10313), .ZN(n10320) );
  NAND4_X1 U11373 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_DATAO_REG_31__SCAN_IN), 
        .A3(n10316), .A4(n10315), .ZN(n10318) );
  NAND4_X1 U11374 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), 
        .A3(P1_IR_REG_30__SCAN_IN), .A4(P1_REG0_REG_17__SCAN_IN), .ZN(n10317)
         );
  NOR2_X1 U11375 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NAND4_X1 U11376 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10330) );
  NOR4_X1 U11377 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .A3(n10324), .A4(n10323), .ZN(n10326) );
  AND2_X1 U11378 ( .A1(n10326), .A2(n10325), .ZN(n10328) );
  NAND4_X1 U11379 ( .A1(n10328), .A2(n8423), .A3(n10327), .A4(n5779), .ZN(
        n10329) );
  NOR2_X1 U11380 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  NAND3_X1 U11381 ( .A1(n10332), .A2(P1_D_REG_16__SCAN_IN), .A3(n10331), .ZN(
        n10333) );
  NOR3_X1 U11382 ( .A1(n10335), .A2(n10334), .A3(n10333), .ZN(n10351) );
  NAND4_X1 U11383 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_REG0_REG_15__SCAN_IN), 
        .A3(P2_IR_REG_13__SCAN_IN), .A4(n10336), .ZN(n10339) );
  NAND4_X1 U11384 ( .A1(n10337), .A2(n5043), .A3(P2_REG1_REG_3__SCAN_IN), .A4(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n10338) );
  NOR2_X1 U11385 ( .A1(n10339), .A2(n10338), .ZN(n10350) );
  NAND4_X1 U11386 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(
        P2_IR_REG_22__SCAN_IN), .ZN(n10346) );
  NAND4_X1 U11387 ( .A1(n10344), .A2(n10343), .A3(P2_REG0_REG_10__SCAN_IN), 
        .A4(P2_REG1_REG_24__SCAN_IN), .ZN(n10345) );
  NOR2_X1 U11388 ( .A1(n10346), .A2(n10345), .ZN(n10349) );
  AND4_X1 U11389 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_1__SCAN_IN), 
        .A3(P1_ADDR_REG_7__SCAN_IN), .A4(n10347), .ZN(n10348) );
  NAND4_X1 U11390 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NOR3_X1 U11391 ( .A1(n10354), .A2(n10353), .A3(n10352), .ZN(n10355) );
  NAND4_X1 U11392 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  XNOR2_X1 U11393 ( .A(n10360), .B(n10359), .ZN(P1_U3557) );
  AOI21_X1 U11394 ( .B1(n10362), .B2(n6365), .A(n10361), .ZN(ADD_1068_U50) );
  INV_X1 U11395 ( .A(n10365), .ZN(n10364) );
  OAI222_X1 U11396 ( .A1(n10367), .A2(n10366), .B1(n10367), .B2(n10365), .C1(
        n10364), .C2(n10363), .ZN(ADD_1068_U51) );
  AOI21_X1 U11397 ( .B1(n10370), .B2(n10369), .A(n10368), .ZN(ADD_1068_U47) );
  AOI21_X1 U11398 ( .B1(n10373), .B2(n10372), .A(n10371), .ZN(ADD_1068_U49) );
  AOI21_X1 U11399 ( .B1(n10376), .B2(n10375), .A(n10374), .ZN(ADD_1068_U48) );
  AOI21_X1 U11400 ( .B1(n10379), .B2(n10378), .A(n10377), .ZN(ADD_1068_U54) );
  AOI21_X1 U11401 ( .B1(n10382), .B2(n10381), .A(n10380), .ZN(ADD_1068_U53) );
  OAI21_X1 U11402 ( .B1(n10385), .B2(n10384), .A(n10383), .ZN(ADD_1068_U52) );
  CLKBUF_X2 U4914 ( .A(n5080), .Z(n5100) );
  CLKBUF_X3 U4930 ( .A(n5834), .Z(n8755) );
  CLKBUF_X1 U4940 ( .A(n5837), .Z(n8635) );
  CLKBUF_X1 U4941 ( .A(n9008), .Z(n4403) );
endmodule

